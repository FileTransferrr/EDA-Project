// ****** Basic Gate Module Defination ******
module or2(out, in1, in2);
  output out;
  input in1, in2;
  wire in1, in2, out;
  assign out = in1 || in2;
endmodule

module and2(out, in1, in2);
  output out;
  input in1, in2;
  wire in1, in2, out;
  assign out = in1 && in2;
endmodule

module not1(out, in);
  output out;
  input in;
  wire in,out;
  assign out = ~in;
endmodule

module nand2(out, in1, in2);
  output out;
  input in1, in2;
  wire in1, in2, out;
  assign out = ~(in1 && in2);
endmodule
// ****** Basic Gate Module Defination End ******

// ****** Combined Logic Module Defination ******
module combLogic( w_000_000, w_000_001, w_000_002, w_000_003, w_000_004, w_000_005, w_000_006, w_000_007, w_000_008, w_000_009, w_000_010, w_000_011, w_000_012, w_000_013, w_000_014, w_000_015, w_000_016, w_000_017, w_000_018, w_000_019, w_000_020, w_000_021, w_000_022, w_000_023, w_000_024, w_000_025, w_000_026, w_000_027, w_000_028, w_000_029, w_000_030, w_000_031, w_000_032, w_000_033, w_000_034, w_000_035, w_000_036, w_000_037, w_000_038, w_000_039, w_000_040, w_000_041, w_000_042, w_000_043, w_000_044, w_000_045, w_000_046, w_000_047, w_000_048, w_000_049, w_000_050, w_000_051, w_000_052, w_000_053, w_000_054, w_000_055, w_000_056, w_000_057, w_000_058, w_000_059, w_000_060, w_000_061, w_000_062, w_000_063, w_000_064, w_000_065, w_000_066, w_000_067, w_000_068, w_000_069, w_000_070, w_000_071, w_000_072, w_000_073, w_000_074, w_000_075, w_000_076, w_000_077, w_000_078, w_000_079, w_000_080, w_000_081, w_000_082, w_000_083, w_000_084, w_000_085, w_000_086, w_000_087, w_000_088, w_000_089, w_000_090, w_000_091, w_000_092, w_000_093, w_000_094, w_000_095, w_000_096, w_000_097, w_000_098, w_000_099, w_000_100, w_000_101, w_000_102, w_000_103, w_000_104, w_000_105, w_000_106, w_000_107, w_000_108, w_000_109, w_000_110, w_000_111, w_000_112, w_000_113, w_000_114, w_000_115, w_000_116, w_000_117, w_000_118, w_000_119, w_000_120, w_000_121, w_000_122, w_000_123, w_000_124, w_000_125, w_000_126, w_000_127, w_000_128, w_000_129, w_000_130, w_000_131, w_000_132, w_000_133, w_000_134, w_000_135, w_000_136, w_000_137, w_000_138, w_000_139, w_000_140, w_000_141, w_000_142, w_000_143, w_000_144, w_000_145, w_000_146, w_000_147, w_000_148, w_000_149, w_000_150, w_000_151, w_000_152, w_000_153, w_000_154, w_000_155, w_000_156, w_000_157, w_000_158, w_000_159, w_000_160, w_000_161, w_000_162, w_000_163, w_000_164, w_000_165, w_000_166, w_000_167, w_000_168, w_000_169, w_000_170, w_000_171, w_000_172, w_000_173, w_000_174, w_000_175, w_000_176, w_000_177, w_000_178, w_000_179, w_000_180, w_000_181, w_000_182, w_000_183, w_000_184, w_000_185, w_000_186, w_000_187, w_000_188, w_000_189, w_000_190, w_000_191, w_000_192, w_000_193, w_000_194, w_000_195, w_000_196, w_000_197, w_000_198, w_000_199, w_000_200, w_000_201, w_000_202, w_000_203, w_000_204, w_000_205, w_000_206, w_000_207, w_000_208, w_000_209, w_000_210, w_000_211, w_000_212, w_000_213, w_000_214, w_000_215, w_000_216, w_000_217, w_000_218, w_000_219, w_000_220, w_000_221, w_000_222, w_000_223, w_000_224, w_000_225, w_000_226, w_000_227, w_000_228, w_000_229, w_000_230, w_000_231, w_000_232, w_000_233, w_000_234, w_000_235, w_000_236, w_000_237, w_000_238, w_000_239, w_000_240, w_000_241, w_000_242, w_000_243, w_000_244, w_000_245, w_000_246, w_000_247, w_000_248, w_000_249, w_000_250, w_000_251, w_000_252, w_000_253, w_000_254, w_000_255, w_000_256, w_000_257, w_000_258, w_000_259, w_000_260, w_000_261, w_000_262, w_000_263, w_000_264, w_000_265, w_000_266, w_000_267, w_000_268, w_000_269, w_000_270, w_000_271, w_000_272, w_000_273, w_000_274, w_000_275, w_000_276, w_000_277, w_000_278, w_000_279, w_000_280, w_000_281, w_000_282, w_000_283, w_000_284, w_000_285, w_000_286, w_000_287, w_000_288, w_000_289, w_000_290, w_000_291, w_000_292, w_000_293, w_000_294, w_000_295, w_000_296, w_000_297, w_000_298, w_000_299, w_000_300, w_000_301, w_000_302, w_000_303, w_000_304, w_000_305, w_000_306, w_000_307, w_000_308, w_000_309, w_000_310, w_000_311, w_000_312, w_000_313, w_000_314, w_000_315, w_000_316, w_000_317, w_000_318, w_000_319, w_000_320, w_000_321, w_000_322, w_000_323, w_000_324, w_000_325, w_000_326, w_000_327, w_000_328, w_000_329, w_000_330, w_000_331, w_000_332, w_000_333, w_000_334, w_000_335, w_000_336, w_000_337, w_000_338, w_000_339, w_000_340, w_000_341, w_000_342, w_000_343, w_000_344, w_000_345, w_000_346, w_000_347, w_000_348, w_000_349, w_000_350, w_000_351, w_000_352, w_000_353, w_000_354, w_000_355, w_000_356, w_000_357, w_000_358, w_000_359, w_000_360, w_000_361, w_000_362, w_000_363, w_000_364, w_000_365, w_000_366, w_000_367, w_000_368, w_000_369, w_000_370, w_000_371, w_000_372, w_000_373, w_000_374, w_000_375, w_000_376, w_000_377, w_000_378, w_000_379, w_000_380, w_000_381, w_000_382, w_000_383, w_000_384, w_000_385, w_000_386, w_000_387, w_000_388, w_000_389, w_000_390, w_000_391, w_000_392, w_000_393, w_000_394, w_000_395, w_000_396, w_000_397, w_000_398, w_000_399, w_000_400, w_000_401, w_000_402, w_000_403, w_000_404, w_000_405, w_000_406, w_000_407, w_000_408, w_000_409, w_000_410, w_000_411, w_000_412, w_000_413, w_000_414, w_000_415, w_000_416, w_000_417, w_000_418, w_000_419, w_000_420, w_000_421, w_000_422, w_000_423, w_000_424, w_000_425, w_000_426, w_000_427, w_000_428, w_000_429, w_000_430, w_000_431, w_000_432, w_000_433, w_000_434, w_000_435, w_000_436, w_000_437, w_000_438, w_000_439, w_000_440, w_000_441, w_000_442, w_000_443, w_000_444, w_000_445, w_000_446, w_000_447, w_000_448, w_000_449, w_000_450, w_000_451, w_000_452, w_000_453, w_000_454, w_000_455, w_000_456, w_000_457, w_000_458, w_000_459, w_000_460, w_000_461, w_000_462, w_000_463, w_000_464, w_000_465, w_000_466, w_000_467, w_000_468, w_000_469, w_000_470, w_000_471, w_000_472, w_000_473, w_000_474, w_000_475, w_000_476, w_000_477, w_000_478, w_000_479, w_000_480, w_000_481, w_000_482, w_000_483, w_000_484, w_000_485, w_000_486, w_000_487, w_000_488, w_000_489, w_000_490, w_000_491, w_000_492, w_000_493, w_000_494, w_000_495, w_000_496, w_000_497, w_000_498, w_000_499, w_000_500, w_000_501, w_000_502, w_000_503, w_000_504, w_000_505, w_000_506, w_000_507, w_000_508, w_000_509, w_000_510, w_000_511, w_000_512, w_000_513, w_000_514, w_000_515, w_000_516, w_000_517, w_000_518, w_000_519, w_000_520, w_000_521, w_000_522, w_000_523, w_000_524, w_000_525, w_000_526, w_000_527, w_000_528, w_000_529, w_000_530, w_000_531, w_000_532, w_000_533, w_000_534, w_000_535, w_000_536, w_000_537, w_000_538, w_000_539, w_000_540, w_000_541, w_000_542, w_000_543, w_000_544, w_000_545, w_000_546, w_000_547, w_000_548, w_000_549, w_000_550, w_000_551, w_000_552, w_000_553, w_000_554, w_000_555, w_000_556, w_000_557, w_000_558, w_000_559, w_000_560, w_000_561, w_000_562, w_000_563, w_000_564, w_000_565, w_000_566, w_000_567, w_000_568, w_000_569, w_000_570, w_000_571, w_000_572, w_000_573, w_000_574, w_000_575, w_000_576, w_000_577, w_000_578, w_000_579, w_000_580, w_000_581, w_000_582, w_000_583, w_000_584, w_000_585, w_000_586, w_000_587, w_000_588, w_000_589, w_000_590, w_000_591, w_000_592, w_000_593, w_000_594, w_000_595, w_000_596, w_000_597, w_000_598, w_000_599, w_000_600, w_000_601, w_000_602, w_000_603, w_000_604, w_000_605, w_000_606, w_000_607, w_000_608, w_000_609, w_000_610, w_000_611, w_000_612, w_000_613, w_000_614, w_000_615, w_000_616, w_000_617, w_000_618, w_000_619, w_000_620, w_000_621, w_000_622, w_000_623, w_000_624, w_000_625, w_000_626, w_000_627, w_000_628, w_000_629, w_000_630, w_000_631, w_000_632, w_000_633, w_000_634, w_000_635, w_000_636, w_000_637, w_000_638, w_000_639, w_000_640, w_000_641, w_000_642, w_000_643, w_000_644, w_000_645, w_000_646, w_000_647, w_000_648, w_000_649, w_000_650, w_000_651, w_000_652, w_000_653, w_000_654, w_000_655, w_000_656, w_000_657, w_000_658, w_000_659, w_000_660, w_000_661, w_000_662, w_000_663, w_000_664, w_000_665, w_000_666, w_000_667, w_000_668, w_000_669, w_000_670, w_000_671, w_000_672, w_000_673, w_000_674, w_000_675, w_000_676, w_000_677, w_000_678, w_000_679, w_000_680, w_000_681, w_000_682, w_000_683, w_000_684, w_000_685, w_000_686, w_000_687, w_000_688, w_000_689, w_000_690, w_000_691, w_000_692, w_000_693, w_000_694, w_000_695, w_000_696, w_000_697, w_000_698, w_000_699, w_000_700, w_000_701, w_000_702, w_000_703, w_000_704, w_000_705, w_000_706, w_000_707, w_000_708, w_000_709, w_000_710, w_000_711, w_000_712, w_000_713, w_000_714, w_000_715, w_000_716, w_000_717, w_000_718, w_000_719, w_000_720, w_000_721, w_000_722, w_000_723, w_000_724, w_000_725, w_000_726, w_000_727, w_000_728, w_000_729, w_000_730, w_000_731, w_000_732, w_000_733, w_000_734, w_000_735, w_000_736, w_000_737, w_000_738, w_000_739, w_000_740, w_000_741, w_000_742, w_000_743, w_000_744, w_000_745, w_000_746, w_000_747, w_000_748, w_000_749, w_000_750, w_000_751, w_000_752, w_000_753, w_000_754, w_000_755, w_000_756, w_000_757, w_000_758, w_000_759, w_000_760, w_000_761, w_000_762, w_000_763, w_000_764, w_000_765, w_000_766, w_000_767, w_000_768, w_000_769, w_000_770, w_000_771, w_000_772, w_000_773, w_000_774, w_000_775, w_000_776, w_000_777, w_000_778, w_000_779, w_000_780, w_000_781, w_000_782, w_000_783, w_000_784, w_000_785, w_000_786, w_000_787, w_000_788, w_000_789, w_000_790, w_000_791, w_000_792, w_000_793, w_000_794, w_000_795, w_000_796, w_000_797, w_000_798, w_000_799, w_000_800, w_000_801, w_000_802, w_000_803, w_000_804, w_000_805, w_000_806, w_000_807, w_000_808, w_000_809, w_000_810, w_000_811, w_000_812, w_000_813, w_000_814, w_000_815, w_000_816, w_000_817, w_000_818, w_000_819, w_000_820, w_000_821, w_000_822, w_000_823, w_000_824, w_000_825, w_000_826, w_000_827, w_000_828, w_000_829, w_000_830, w_000_831, w_000_832, w_000_833, w_000_834, w_000_835, w_000_836, w_000_837, w_000_838, w_000_839, w_000_840, w_000_841, w_000_842, w_000_843, w_000_844, w_000_845, w_000_846, w_000_847, w_000_848, w_000_849, w_000_850, w_000_851, w_000_852, w_000_853, w_000_854, w_000_855, w_000_856, w_000_857, w_000_858, w_000_859, w_000_860, w_000_861, w_000_862, w_000_863, w_000_864, w_000_865, w_000_866, w_000_867, w_000_868, w_000_869, w_000_870, w_000_871, w_000_872, w_000_873, w_000_874, w_000_875, w_000_876, w_000_877, w_000_878, w_000_879, w_000_880, w_000_881, w_000_882, w_000_883, w_000_884, w_000_885, w_000_886, w_000_887, w_000_888, w_000_889, w_000_890, w_000_891, w_000_892, w_000_893, w_000_894, w_000_895, w_000_896, w_000_897, w_000_898, w_000_899, w_000_900, w_000_901, w_000_902, w_000_903, w_000_904, w_000_905, w_000_906, w_000_907, w_000_908, w_000_909, w_000_910, w_000_911, w_000_912, w_000_913, w_000_914, w_000_915, w_000_916, w_000_917, w_000_918, w_000_919, w_000_920, w_000_921, w_000_922, w_000_923, w_000_924, w_000_925, w_000_926, w_000_927, w_000_928, w_000_929, w_000_930, w_000_931, w_000_932, w_000_933, w_000_934, w_000_935, w_000_936, w_000_937, w_000_938, w_000_939, w_000_940, w_000_941, w_000_942, w_000_943, w_000_944, w_000_945, w_000_946, w_000_947, w_000_948, w_000_949, w_000_950, w_000_951, w_000_952, w_000_953, w_000_954, w_000_955, w_000_956, w_000_957, w_000_958, w_000_959, w_000_960, w_000_961, w_000_962, w_000_963, w_000_964, w_000_965, w_000_966, w_000_967, w_000_968, w_000_969, w_000_970, w_000_971, w_000_972, w_000_973, w_000_974, w_000_975, w_000_976, w_000_977, w_000_978, w_000_979, w_000_980, w_000_981, w_000_982, w_000_983, w_000_984, w_000_985, w_000_986, w_000_987, w_000_988, w_000_989, w_000_990, w_000_991, w_000_992, w_000_993, w_000_994, w_000_995, w_000_996, w_000_997, w_000_998, w_000_999, w_000_1000, w_000_1001, w_000_1002, w_000_1003, w_000_1004, w_000_1005, w_000_1006, w_000_1007, w_000_1008, w_000_1009, w_000_1010, w_000_1011, w_000_1012, w_000_1013, w_000_1014, w_000_1015, w_000_1016, w_000_1017, w_000_1018, w_000_1019, w_000_1020, w_000_1021, w_000_1022, w_000_1023, w_000_1024, w_000_1025, w_000_1026, w_000_1027, w_000_1028, w_000_1029, w_000_1030, w_000_1031, w_000_1032, w_000_1033, w_000_1034, w_000_1035, w_000_1036, w_000_1037, w_000_1038, w_000_1039, w_000_1040, w_000_1041, w_000_1042, w_000_1043, w_000_1044, w_000_1045, w_000_1046, w_000_1047, w_000_1048, w_000_1049, w_000_1050, w_000_1051, w_000_1052, w_000_1053, w_000_1054, w_000_1055, w_000_1056, w_000_1057, w_000_1058, w_000_1059, w_000_1060, w_000_1061, w_000_1062, w_000_1063, w_000_1064, w_000_1065, w_000_1066, w_000_1067, w_000_1068, w_000_1069, w_000_1070, w_000_1071, w_000_1072, w_000_1073, w_000_1074, w_000_1075, w_000_1076, w_000_1077, w_000_1078, w_000_1079, w_000_1080, w_000_1081, w_000_1082, w_000_1083, w_000_1084, w_000_1085, w_000_1086, w_000_1087, w_000_1088, w_000_1089, w_000_1090, w_000_1091, w_000_1092, w_000_1093, w_000_1094, w_000_1095, w_000_1096, w_000_1097, w_000_1098, w_000_1099, w_000_1100, w_000_1101, w_000_1102, w_000_1103, w_000_1104, w_000_1105, w_000_1106, w_000_1107, w_000_1108, w_000_1109, w_000_1110, w_000_1111, w_000_1112, w_000_1113, w_000_1114, w_000_1115, w_000_1116, w_000_1117, w_000_1118, w_000_1119, w_000_1120, w_000_1121, w_000_1122, w_000_1123, w_000_1124, w_000_1125, w_000_1126, w_000_1127, w_000_1128, w_000_1129, w_000_1130, w_000_1131, w_000_1132, w_000_1133, w_000_1134, w_000_1135, w_000_1136, w_000_1137, w_000_1138, w_000_1139, w_000_1140, w_000_1141, w_000_1142, w_000_1143, w_000_1144, w_000_1145, w_000_1146, w_000_1147, w_000_1148, w_000_1149, w_000_1150, w_000_1151, w_000_1152, w_000_1153, w_000_1154, w_000_1155, w_000_1156, w_000_1157, w_000_1158, w_000_1159, w_000_1160, w_000_1161, w_000_1162, w_000_1163, w_000_1164, w_000_1165, w_000_1166, w_000_1167, w_000_1168, w_000_1169, w_000_1170, w_000_1171, w_000_1172, w_000_1173, w_000_1174, w_000_1175, w_000_1176, w_000_1177, w_000_1178, w_000_1179, w_000_1180, w_000_1181, w_000_1182, w_000_1183, w_000_1184, w_000_1185, w_000_1186, w_000_1187, w_000_1188, w_000_1189, w_000_1190, w_000_1191, w_000_1192, w_000_1193, w_000_1194, w_000_1195, w_000_1196, w_000_1197, w_000_1198, w_000_1199, w_000_1200, w_000_1201, w_000_1202, w_000_1203, w_000_1204, w_000_1205, w_000_1206, w_000_1207, w_000_1208, w_000_1209, w_000_1210, w_000_1211, w_000_1212, w_000_1213, w_000_1214, w_000_1215, w_000_1216, w_000_1217, w_000_1218, w_000_1219, w_000_1220, w_000_1221, w_000_1222, w_000_1223, w_000_1224, w_000_1225, w_000_1226, w_000_1227, w_000_1228, w_000_1229, w_000_1230, w_000_1231, w_000_1232, w_000_1233, w_000_1234, w_000_1235, w_000_1236, w_000_1237, w_000_1238, w_000_1239, w_000_1240, w_000_1241, w_000_1242, w_000_1243, w_000_1244, w_000_1245, w_000_1246, w_000_1247, w_000_1248, w_000_1249, w_000_1250, w_000_1251, w_000_1252, w_000_1253, w_000_1254, w_000_1255, w_000_1256, w_000_1257, w_000_1258, w_000_1259, w_000_1260, w_000_1261, w_000_1262, w_000_1263, w_000_1264, w_000_1265, w_000_1266, w_000_1267, w_000_1268, w_000_1269, w_000_1270, w_000_1271, w_000_1272, w_000_1273, w_000_1274, w_000_1275, w_000_1276, w_000_1277, w_000_1278, w_000_1279, w_000_1280, w_000_1281, w_000_1282, w_000_1283, w_000_1284, w_000_1285, w_000_1286, w_000_1287, w_000_1288, w_000_1289, w_000_1290, w_000_1291, w_000_1292, w_000_1293, w_000_1294, w_000_1295, w_000_1296, w_000_1297, w_000_1298, w_000_1299, w_000_1300, w_000_1301, w_000_1302, w_000_1303, w_000_1304, w_000_1305, w_000_1306, w_000_1307, w_000_1308, w_000_1309, w_000_1310, w_000_1311, w_000_1312, w_000_1313, w_000_1314, w_000_1315, w_000_1316, w_000_1317, w_000_1318, w_000_1319, w_000_1320, w_000_1321, w_000_1322, w_000_1323, w_000_1324, w_000_1325, w_000_1326, w_000_1327, w_000_1328, w_000_1329, w_000_1330, w_000_1331, w_000_1332, w_000_1333, w_000_1334, w_000_1335, w_000_1336, w_000_1337, w_000_1338, w_000_1339, w_000_1340, w_000_1341, w_000_1342, w_000_1343, w_000_1344, w_000_1345, w_000_1346, w_000_1347, w_000_1348, w_000_1349, w_000_1350, w_000_1351, w_000_1352, w_000_1353, w_000_1354, w_000_1355, w_000_1356, w_000_1357, w_000_1358, w_000_1359, w_000_1360, w_000_1361, w_000_1362, w_000_1363, w_000_1364, w_000_1365, w_000_1366, w_000_1367, w_000_1368, w_000_1369, w_000_1370, w_000_1371, w_000_1372, w_000_1373, w_000_1374, w_000_1375, w_000_1376, w_000_1377, w_000_1378, w_000_1379, w_000_1380, w_000_1381, w_000_1382, w_000_1383, w_000_1384, w_000_1385, w_000_1386, w_000_1387, w_000_1388, w_000_1389, w_000_1390, w_000_1391, w_000_1392, w_000_1393, w_000_1394, w_000_1395, w_000_1396, w_000_1397, w_000_1398, w_000_1399, w_000_1400, w_000_1401, w_000_1402, w_000_1403, w_000_1404, w_000_1405, w_000_1406, w_000_1407, w_000_1408, w_000_1409, w_000_1410, w_000_1411, w_000_1412, w_000_1413, w_000_1414, w_000_1415, w_000_1416, w_000_1417, w_000_1418, w_000_1419, w_000_1420, w_000_1421, w_000_1422, w_000_1423, w_000_1424, w_000_1425, w_000_1426, w_000_1427, w_000_1428, w_000_1429, w_000_1430, w_000_1431, w_000_1432, w_000_1433, w_000_1434, w_000_1435, w_000_1436, w_000_1437, w_000_1438, w_000_1439, w_000_1440, w_000_1441, w_000_1442, w_000_1443, w_000_1444, w_000_1445, w_000_1446, w_000_1447, w_000_1448, w_000_1449, w_000_1450, w_000_1451, w_000_1452, w_000_1453, w_000_1454, w_000_1455, w_000_1456, w_000_1457, w_000_1458, w_000_1459, w_000_1460, w_000_1461, w_000_1462, w_000_1463, w_000_1464, w_000_1465, w_000_1466, w_000_1467, w_000_1468, w_000_1469, w_000_1470, w_000_1471, w_000_1472, w_000_1473, w_000_1474, w_000_1475, w_000_1476, w_000_1477, w_000_1478, w_000_1479, w_000_1480, w_000_1481, w_000_1482, w_000_1483, w_000_1484, w_000_1485, w_000_1486, w_000_1487, w_000_1488, w_000_1489, w_000_1490, w_000_1491, w_000_1492, w_000_1493, w_000_1494, w_000_1495, w_000_1496, w_000_1497, w_000_1498, w_000_1499, w_000_1500, w_000_1501, w_000_1502, w_000_1503, w_000_1504, w_000_1505, w_000_1506, w_000_1507, w_000_1508, w_000_1509, w_000_1510, w_000_1511, w_000_1512, w_000_1513, w_000_1514, w_000_1515, w_000_1516, w_000_1517, w_000_1518, w_000_1519, w_000_1520, w_000_1521, w_000_1522, w_000_1523, w_000_1524, w_000_1525, w_000_1526, w_000_1527, w_000_1528, w_000_1529, w_000_1530, w_000_1531, w_000_1532, w_000_1533, w_000_1534, w_000_1535, w_000_1536, w_000_1537, w_000_1538, w_000_1539, w_000_1540, w_000_1541, w_000_1542, w_000_1543, w_000_1544, w_000_1545, w_000_1546, w_000_1547, w_000_1548, w_000_1549, w_000_1550, w_000_1551, w_000_1552, w_000_1553, w_000_1554, w_000_1555, w_000_1556, w_000_1557, w_000_1558, w_000_1559, w_000_1560, w_000_1561, w_000_1562, w_000_1563, w_000_1564, w_000_1565, w_000_1566, w_000_1567, w_000_1568, w_000_1569, w_000_1570, w_000_1571, w_000_1572, w_000_1573, w_000_1574, w_000_1575, w_000_1576, w_000_1577, w_000_1578, w_000_1579, w_000_1580, w_000_1581, w_000_1582, w_000_1583, w_000_1584, w_000_1585, w_000_1586, w_000_1587, w_000_1588, w_000_1589, w_000_1590, w_000_1591, w_000_1592, w_000_1593, w_000_1594, w_000_1595, w_000_1596, w_000_1597, w_000_1598, w_000_1599, w_000_1600, w_000_1601, w_000_1602, w_000_1603, w_000_1604, w_000_1605, w_000_1606, w_000_1607, w_000_1608, w_000_1609, w_000_1610, w_000_1611, w_000_1612, w_000_1613, w_000_1614, w_000_1615, w_000_1616, w_000_1617, w_000_1618, w_000_1619, w_000_1620, w_000_1621, w_000_1622, w_000_1623, w_000_1624, w_000_1625, w_000_1626, w_000_1627, w_000_1628, w_000_1629, w_000_1630, w_000_1631, w_000_1632, w_000_1633, w_000_1634, w_000_1635, w_000_1636, w_000_1637, w_000_1638, w_000_1639, w_000_1640, w_000_1641, w_000_1642, w_000_1643, w_000_1644, w_000_1645, w_000_1646, w_000_1647, w_000_1648, w_000_1649, w_000_1650, w_000_1651, w_000_1652, w_000_1653, w_000_1654, w_000_1655, w_000_1656, w_000_1657, w_000_1658, w_000_1659, w_000_1660, w_000_1661, w_000_1662, w_000_1663, w_000_1664, w_000_1665, w_000_1666, w_000_1667, w_000_1668, w_000_1669, w_000_1670, w_000_1671, w_000_1672, w_000_1673, w_000_1674, w_000_1675, w_000_1676, w_000_1677, w_000_1678, w_000_1679, w_000_1680, w_000_1681, w_000_1682, w_000_1683, w_000_1684, w_000_1685, w_000_1686, w_000_1687, w_000_1688, w_000_1689, w_000_1690, w_000_1691, w_000_1692, w_000_1693, w_000_1694, w_000_1695, w_000_1696, w_000_1697, w_000_1698, w_000_1699, w_000_1700, w_000_1701, w_000_1702, w_000_1703, w_000_1704, w_000_1705, w_000_1706, w_000_1707, w_000_1708, w_000_1709, w_000_1710, w_000_1711, w_000_1712, w_000_1713, w_000_1714, w_000_1715, w_000_1716, w_000_1717, w_000_1718, w_000_1719, w_000_1720, w_000_1721, w_000_1722, w_000_1723, w_000_1724, w_000_1725, w_000_1726, w_000_1727, w_000_1728, w_000_1729, w_000_1730, w_000_1731, w_000_1732, w_000_1733, w_000_1734, w_000_1735, w_000_1736, w_000_1737, w_000_1738, w_000_1739, w_000_1740, w_000_1741, w_000_1742, w_000_1743, w_000_1744, w_000_1745, w_000_1746, w_000_1747, w_000_1748, w_000_1749, w_000_1750, w_000_1751, w_000_1752, w_000_1753, w_000_1754, w_000_1755, w_000_1756, w_000_1757, w_000_1758, w_000_1759, w_000_1760, w_000_1761, w_000_1762, w_000_1763, w_000_1764, w_000_1765, w_000_1766, w_000_1767, w_000_1768, w_000_1769, w_000_1770, w_000_1771, w_000_1772, w_000_1773, w_000_1774, w_000_1775, w_000_1776, w_000_1777, w_000_1778, w_000_1779, w_000_1780, w_000_1781, w_000_1782, w_000_1783, w_000_1784, w_000_1785, w_000_1786, w_000_1787, w_000_1788, w_000_1789, w_000_1790, w_000_1791, w_000_1792, w_000_1793, w_000_1794, w_000_1795, w_000_1796, w_000_1797, w_000_1798, w_000_1799, w_000_1800, w_000_1801, w_000_1802, w_000_1803, w_000_1804, w_000_1805, w_000_1806, w_000_1807, w_000_1808, w_000_1809, w_000_1810, w_000_1811, w_000_1812, w_000_1813, w_000_1814, w_000_1815, w_000_1816, w_000_1817, w_000_1818, w_000_1819, w_000_1820, w_000_1821, w_000_1822, w_000_1823, w_000_1824, w_000_1825, w_000_1826, w_000_1827, w_000_1828, w_000_1829, w_000_1830, w_000_1831, w_000_1832, w_000_1833, w_000_1834, w_000_1835, w_000_1836, w_000_1837, w_000_1838, w_000_1839, w_000_1840, w_000_1841, w_000_1842, w_000_1843, w_000_1844, w_000_1845, w_000_1846, w_000_1847, w_000_1848, w_000_1849, w_000_1850, w_000_1851, w_000_1852, w_000_1853, w_000_1854, w_000_1855, w_000_1856, w_000_1857, w_000_1858, w_000_1859, w_000_1860, w_000_1861, w_000_1862, w_000_1863, w_000_1864, w_000_1865, w_000_1866, w_000_1867, w_000_1868, w_000_1869, w_000_1870, w_000_1871, w_000_1872, w_000_1873, w_000_1874, w_000_1875, w_000_1876, w_000_1877, w_000_1878, w_000_1879, w_000_1880, w_000_1881, w_000_1882, w_000_1883, w_000_1884, w_000_1885, w_000_1886, w_000_1887, w_000_1888, w_000_1889, w_000_1890, w_000_1891, w_000_1892, w_000_1893, w_000_1894, w_000_1895, w_000_1896, w_000_1897, w_000_1898, w_000_1899, w_000_1900, w_000_1901, w_000_1902, w_000_1903, w_000_1904, w_000_1905, w_000_1906, w_000_1907, w_000_1908, w_000_1909, w_000_1910, w_000_1911, w_000_1912, w_000_1913, w_000_1914, w_000_1915, w_000_1916, w_000_1917, w_000_1918, w_000_1919, w_000_1920, w_000_1921, w_000_1922, w_000_1923, w_000_1924, w_000_1925, w_000_1926, w_000_1927, w_000_1928, w_000_1929, w_000_1930, w_000_1931, w_000_1932, w_000_1933, w_000_1934, w_000_1935, w_000_1936, w_000_1937, w_000_1938, w_000_1939, w_000_1940, w_000_1941, w_000_1942, w_000_1943, w_000_1944, w_000_1945, w_000_1946, w_000_1947, w_000_1948, w_000_1949, w_000_1950, w_000_1951, w_000_1952, w_000_1953, w_000_1954, w_000_1955, w_000_1956, w_000_1957, w_000_1958, w_000_1959, w_000_1960, w_000_1961, w_000_1962, w_000_1963, w_000_1964, w_000_1965, w_000_1966, w_000_1967, w_000_1968, w_000_1969, w_000_1970, w_000_1971, w_000_1972, w_000_1973, w_000_1974, w_000_1975, w_000_1976, w_000_1977, w_000_1978, w_000_1979, w_000_1980, w_000_1981, w_000_1982, w_000_1983, w_000_1984, w_000_1985, w_000_1986, w_000_1987, w_000_1988, w_000_1989, w_000_1990, w_000_1991, w_000_1992, w_000_1993, w_000_1994, w_000_1995, w_000_1996, w_000_1997, w_000_1998, w_000_1999, w_000_2000, w_000_2001, w_000_2002, w_000_2003, w_000_2004, w_000_2005, w_000_2006, w_000_2007, w_000_2008, w_000_2009, w_000_2010, w_000_2011, w_000_2012, w_000_2013, w_000_2014, w_000_2015, w_000_2016, w_000_2017, w_000_2018, w_000_2019, w_000_2020, w_000_2021, w_000_2022, w_000_2023, w_000_2024, w_000_2025, w_000_2026, w_000_2027, w_000_2028, w_000_2029, w_000_2030, w_000_2031, w_000_2032, w_000_2033, w_000_2034, w_000_2035, w_000_2036, w_000_2037, w_000_2038, w_000_2039, w_000_2040, w_000_2041, w_000_2042, w_000_2043, w_000_2044, w_000_2045, w_000_2046, w_000_2047, w_000_2048, w_000_2049, w_000_2050, w_000_2051, w_000_2052, w_000_2053, w_000_2054, w_000_2055, w_000_2056, w_000_2057, w_000_2058, w_000_2059, w_000_2060, w_000_2061, w_000_2062, w_000_2063, w_000_2064, w_000_2065, w_000_2066, w_000_2067, w_000_2068, w_000_2069, w_000_2070, w_000_2071, w_000_2072, w_000_2073, w_000_2074, w_000_2075, w_000_2076, w_000_2077, w_000_2078, w_000_2079, w_000_2080, w_000_2081, w_000_2082, w_000_2083, w_000_2084, w_000_2085, w_000_2086, w_000_2087, w_000_2088, w_000_2089, w_000_2090, w_000_2091, w_000_2092, w_000_2093, w_000_2094, w_000_2095, w_000_2096, w_000_2097, w_000_2098, w_000_2099, w_000_2100, w_000_2101, w_000_2102, w_000_2103, w_000_2104, w_000_2105, w_000_2106, w_000_2107, w_000_2108, w_000_2109, w_000_2110, w_000_2111, w_000_2112, w_000_2113, w_000_2114, w_000_2115, w_000_2116, w_000_2117, w_000_2118, w_000_2119, w_000_2120, w_000_2121, w_000_2122, w_000_2123, w_000_2124, w_000_2125, w_000_2126, w_000_2127, w_000_2128, w_000_2129, w_000_2130, w_000_2131, w_000_2132, w_000_2133, w_000_2134, w_000_2135, w_000_2136, w_000_2137, w_000_2138, w_000_2139, w_000_2140, w_000_2141, w_000_2142, w_000_2143, w_000_2144, w_000_2145, w_000_2146, w_000_2147, w_000_2148, w_000_2149, w_000_2150, w_000_2151, w_000_2152, w_000_2153, w_000_2154, w_000_2155, w_000_2156, w_000_2157, w_000_2158, w_000_2160, w_000_2161, w_000_2162, w_000_2163, w_000_2164, w_000_2165, w_000_2166, w_000_2167, w_000_2168, w_000_2169, w_000_2170, w_000_2171, w_000_2172, w_000_2173, w_000_2174, w_000_2175, w_000_2176, w_000_2177, w_000_2178, w_000_2179, w_000_2180, w_000_2181, w_000_2182, w_000_2183, w_000_2184, w_000_2185, w_000_2186, w_000_2187, w_000_2188, w_000_2189, w_000_2190, w_000_2191, w_000_2192, w_000_2193, w_000_2194, w_000_2195, w_000_2196, w_000_2197, w_000_2198, w_000_2199, w_000_2200, w_000_2201, w_000_2202, w_000_2203, w_000_2204, w_000_2205, w_000_2206, w_000_2207, w_000_2208, w_000_2209, w_000_2210, w_000_2211, w_000_2212, w_000_2213, w_000_2214, w_000_2215, w_000_2216, w_000_2217, w_000_2218, w_000_2219, w_000_2220, w_000_2221, w_000_2222, w_000_2223, w_000_2224, w_000_2225, w_000_2226, w_000_2227, w_000_2228, w_000_2229, w_000_2230, w_000_2231, w_000_2232, w_000_2233, w_000_2234, w_000_2235, w_000_2236, w_000_2237, w_000_2238, w_000_2239, w_000_2240, w_000_2241, w_000_2242, w_000_2243, w_000_2244, w_000_2245, w_000_2246, w_000_2247, w_000_2248, w_000_2249, w_000_2250, w_000_2251, w_000_2252, w_000_2253, w_000_2254, w_000_2255, w_000_2256, w_000_2257, w_000_2258, w_000_2259, w_000_2260, w_000_2261, w_000_2262, w_000_2263, w_000_2264, w_000_2265, w_000_2266, w_000_2267, w_000_2268, w_000_2269, w_000_2270, w_000_2271, w_000_2272, w_000_2273, w_000_2274, w_000_2275, w_000_2276, w_000_2277, w_000_2278, w_000_2279, w_000_2280, w_000_2281, w_000_2282, w_000_2283, w_000_2284, w_000_2285, w_000_2286, w_000_2287, w_000_2288, w_000_2289, w_000_2290, w_000_2291, w_000_2292, w_000_2293, w_000_2294, w_000_2295, w_000_2296, w_000_2297, w_000_2298, w_000_2299, w_000_2300, w_000_2301, w_000_2302, w_000_2303, w_000_2304, w_000_2305, w_000_2306, w_000_2307, w_000_2308, w_000_2309, w_000_2310, w_000_2311, w_000_2312, w_000_2313, w_000_2314, w_000_2315, w_000_2316, w_000_2317, w_000_2318, w_000_2319, w_000_2320, w_000_2321, w_000_2322, w_000_2323, w_000_2324, w_000_2325, w_000_2326, w_000_2327, w_000_2328, w_000_2329, w_000_2330, w_000_2331, w_000_2332, w_000_2333, w_000_2334, w_000_2335, w_000_2336, w_000_2337, w_000_2338, w_000_2339, w_000_2340, w_000_2341, w_000_2342, w_000_2343, w_000_2344, w_000_2345, w_000_2346, w_000_2347, w_000_2348, w_000_2349, w_000_2350, w_000_2351, w_000_2352, w_000_2353, w_000_2354, w_000_2355, w_000_2356, w_000_2357, w_000_2358, w_000_2359, w_000_2360, w_000_2361, w_000_2362, w_000_2363, w_000_2364, w_000_2365, w_000_2366, w_000_2367, w_000_2368, w_000_2369, w_000_2370, w_000_2371, w_000_2372, w_000_2373, w_000_2374, w_000_2375, w_000_2376, w_000_2377, w_000_2378, w_000_2379, w_000_2380, w_000_2381, w_000_2382, w_000_2383, w_000_2384, w_000_2385, w_000_2386, w_000_2387, w_000_2388, w_000_2389, w_000_2390, w_000_2391, w_000_2392, w_000_2393, w_000_2394, w_000_2395, w_000_2396, w_000_2397, w_000_2398, w_000_2399, w_000_2400, w_000_2401, w_000_2402, w_000_2403, w_000_2404, w_000_2405, w_000_2406, w_000_2407, w_000_2408, w_000_2410, w_000_2411, w_000_2412, w_000_2413, w_000_2414, w_000_2415, w_000_2416, w_000_2417, w_000_2418, w_000_2419, w_000_2420, w_000_2421, w_000_2422, w_000_2423, w_000_2424, w_000_2425, w_000_2426, w_000_2427, w_000_2428, w_000_2429, w_000_2430, w_000_2431, w_000_2432, w_000_2433, w_000_2434, w_000_2435, w_000_2436, w_000_2437, w_000_2438, w_000_2439, w_000_2440, w_000_2441, w_000_2442, w_000_2443, w_000_2444, w_000_2445, w_000_2446, w_000_2447, w_000_2448, w_000_2449, w_000_2450, w_000_2451, w_000_2452, w_000_2453, w_000_2454, w_000_2455, w_000_2456, w_000_2457, w_000_2458, w_000_2459, w_000_2460, w_000_2461, w_000_2462, w_000_2463, w_000_2464, w_000_2465, w_000_2466, w_000_2467, w_000_2468, w_000_2469, w_000_2470, w_000_2471, w_000_2472, w_000_2473, w_000_2474, w_000_2475, w_000_2476, w_000_2477, w_000_2478, w_000_2479, w_000_2480, w_000_2481, w_000_2482, w_000_2483, w_000_2484, w_000_2485, w_000_2486, w_000_2487, w_000_2488, w_000_2489, w_000_2490, w_000_2491, w_000_2492, w_000_2493, w_000_2494, w_000_2495, w_000_2496, w_000_2497, w_000_2498, w_000_2499, w_000_2500, w_000_2501, w_000_2502, w_000_2503, w_000_2504, w_000_2505, w_000_2506, w_000_2507, w_000_2508, w_000_2509, w_000_2510, w_000_2511, w_000_2512, w_000_2513, w_000_2514, w_000_2515, w_000_2516, w_000_2517, w_000_2518, w_000_2519, w_000_2520, w_000_2521, w_000_2522, w_000_2523, w_000_2524, w_000_2525, w_000_2526, w_000_2527, w_000_2528, w_000_2529, w_000_2530, w_000_2531, w_000_2532, w_000_2533, w_000_2534, w_000_2535, w_000_2536, w_000_2537, w_000_2538, w_000_2539, w_000_2540, w_000_2541, w_000_2542, w_000_2543, w_000_2544, w_000_2545, w_000_2546, w_000_2547, w_000_2548, w_000_2549, w_000_2550, w_000_2551, w_000_2552, w_000_2553, w_000_2554, w_000_2555, w_000_2556, w_000_2557, w_000_2558, w_000_2559, w_000_2560, w_000_2561, w_000_2562, w_000_2563, w_000_2564, w_000_2565, w_000_2566, w_000_2567, w_000_2568, w_000_2569, w_000_2570, w_000_2571, w_000_2572, w_000_2573, w_000_2574, w_000_2575, w_000_2576, w_000_2577, w_000_2578, w_000_2579, w_000_2580, w_000_2581, w_000_2582, w_000_2583, w_000_2584, w_000_2585, w_000_2586, w_000_2587, w_000_2588, w_000_2589, w_000_2590, w_000_2591, w_000_2592, w_000_2593, w_000_2594, w_000_2595, w_000_2596, w_000_2597, w_000_2598, w_000_2599, w_000_2600, w_000_2601, w_000_2602, w_000_2603, w_000_2604, w_000_2605, w_000_2606, w_000_2607, w_000_2608, w_000_2609, w_000_2610, w_000_2611, w_000_2612, w_000_2613, w_000_2614, w_000_2615, w_000_2616, w_000_2617, w_000_2618, w_000_2619, w_000_2620, w_000_2621, w_000_2622, w_000_2623, w_000_2624, w_000_2625, w_000_2626, w_000_2627, w_000_2628, w_000_2629, w_000_2630, w_000_2631, w_000_2632, w_000_2633, w_000_2634, w_000_2635, w_000_2636, w_000_2637, w_000_2638, w_000_2639, w_000_2640, w_000_2641, w_000_2642, w_000_2643, w_000_2644, w_000_2645, w_000_2646, w_000_2647, w_000_2648, w_000_2649, w_000_2650, w_000_2651, w_000_2652, w_000_2653, w_000_2654, w_000_2655, w_000_2656, w_000_2657, w_000_2658, w_000_2659, w_000_2660, w_000_2661, w_000_2662, w_000_2663, w_000_2664, w_000_2665, w_000_2666, w_000_2667, w_000_2668, w_000_2669, w_000_2670, w_000_2671, w_000_2672, w_000_2673, w_000_2674, w_000_2675, w_000_2676, w_000_2677, w_000_2678, w_000_2679, w_000_2680, w_000_2681, w_000_2682, w_000_2683, w_000_2684, w_000_2685, w_000_2686, w_000_2687, w_000_2688, w_000_2689, w_000_2690, w_000_2691, w_000_2692, w_000_2693, w_000_2694, w_000_2695, w_000_2696, w_000_2697, w_000_2698, w_000_2699, w_000_2700, w_000_2701, w_000_2702, w_000_2703, w_000_2704, w_000_2705, w_000_2706, w_000_2707, w_000_2708, w_000_2709, w_000_2710, w_000_2711, w_000_2712, w_000_2713, w_000_2714, w_000_2715, w_000_2716, w_000_2717, w_000_2718, w_000_2719, w_000_2720, w_000_2721, w_000_2722, w_000_2723, w_000_2724, w_000_2725, w_000_2726, w_000_2727, w_000_2728, w_000_2729, w_000_2730, w_000_2731, w_000_2732, w_000_2733, w_000_2734, w_000_2735, w_000_2736, w_000_2737, w_000_2738, w_000_2739, w_000_2740, w_000_2741, w_000_2742, w_000_2743, w_000_2744, w_000_2745, w_000_2746, w_000_2747, w_000_2748, w_000_2749, w_000_2750, w_000_2751, w_000_2752, w_000_2753, w_000_2754, w_000_2755, w_000_2756, w_000_2757, w_000_2758, w_000_2759, w_000_2760, w_000_2761, w_000_2762, w_000_2763, w_000_2764, w_000_2765, w_000_2766, w_000_2767, w_000_2768, w_000_2769, w_000_2770, w_000_2771, w_000_2772, w_000_2773, w_000_2774, w_000_2775, w_000_2776, w_000_2777, w_000_2778, w_000_2779, w_000_2780, w_000_2781, w_000_2782, w_000_2783, w_000_2784, w_000_2785, w_000_2786, w_000_2787, w_000_2788, w_000_2789, w_000_2790, w_000_2791, w_000_2792, w_000_2793, w_000_2794, w_000_2795, w_000_2796, w_000_2797, w_000_2798, w_000_2799, w_000_2800, w_000_2801, w_000_2802, w_000_2803, w_000_2804, w_000_2805, w_000_2806, w_000_2807, w_000_2808, w_000_2809, w_000_2810, w_000_2811, w_000_2812, w_000_2813, w_000_2814, w_000_2815, w_000_2816, w_000_2817, w_000_2818, w_000_2819, w_000_2820, w_000_2821, w_000_2822, w_000_2823, w_000_2824, w_000_2825, w_000_2826, w_000_2827, w_000_2828, w_000_2829, w_000_2830, w_000_2831, w_000_2832, w_000_2834, w_000_2835, w_000_2836, w_000_2837, w_000_2838, w_000_2839, w_000_2840, w_000_2841, w_000_2842, w_000_2843, w_000_2844, w_000_2845, w_000_2846, w_000_2847, w_000_2848, w_000_2849, w_000_2850, w_000_2851, w_000_2852, w_000_2853, w_000_2854, w_000_2855, w_000_2856, w_000_2857, w_000_2858, w_000_2859, w_000_2860, w_000_2861, w_000_2862, w_000_2863, w_000_2864, w_000_2865, w_000_2866, w_000_2867, w_000_2868, w_000_2869, w_000_2870, w_000_2871, w_000_2872, w_000_2873, w_000_2874, w_000_2875, w_000_2876, w_000_2877, w_000_2878, w_000_2879, w_000_2880, w_000_2881, w_000_2882, w_000_2883, w_000_2884, w_000_2885, w_000_2886, w_000_2887, w_000_2888, w_000_2889, w_000_2890, w_000_2891, w_000_2892, w_000_2893, w_000_2894, w_000_2895, w_000_2896, w_000_2897, w_000_2898, w_000_2899, w_000_2900, w_000_2901, w_000_2902, w_000_2903, w_000_2904, w_000_2905, w_000_2906, w_000_2907, w_000_2908, w_000_2909, w_000_2910, w_000_2911, w_000_2912, w_000_2913, w_000_2914, w_000_2915, w_000_2916, w_000_2917, w_000_2918, w_000_2919, w_000_2920, w_000_2921, w_000_2922, w_000_2923, w_000_2924, w_000_2925, w_000_2926, w_000_2927, w_000_2928, w_000_2929, w_000_2930, w_000_2931, w_000_2932, w_000_2933, w_000_2934, w_000_2935, w_000_2936, w_000_2937, w_000_2938, w_000_2939, w_000_2940, w_000_2941, w_000_2942, w_000_2943, w_000_2944, w_000_2945, w_000_2946, w_000_2947, w_000_2948, w_000_2949, w_000_2950, w_000_2951, w_000_2952, w_000_2953, w_000_2954, w_000_2955, w_000_2956, w_000_2957, w_000_2958, w_000_2959, w_000_2960, w_000_2961, w_000_2962, w_000_2963, w_000_2964, w_000_2965, w_000_2966, w_000_2967, w_000_2968, w_000_2969, w_000_2970, w_000_2971, w_000_2972, w_000_2973, w_000_2974, w_000_2975, w_000_2976, w_000_2977, w_000_2978, w_000_2979, w_000_2980, w_000_2981, w_000_2982, w_000_2983, w_000_2984, w_000_2985, w_000_2986, w_000_2987, w_000_2988, w_000_2989, w_000_2990, w_000_2991, w_000_2992, w_000_2993, w_000_2994, w_000_2995, w_000_2996, w_000_2997, w_000_2998, w_000_2999, w_000_3000, w_000_3001, w_000_3002, w_000_3003, w_000_3004, w_000_3005, w_000_3006, w_000_3007, w_000_3008, w_000_3009, w_000_3010, w_000_3011, w_000_3012, w_000_3013, w_000_3014, w_000_3015, w_000_3016, w_000_3017, w_000_3018, w_000_3019, w_000_3020, w_000_3021, w_000_3022, w_000_3023, w_000_3024, w_000_3025, w_000_3026, w_000_3027, w_000_3028, w_000_3029, w_000_3030, w_000_3031, w_000_3032, w_000_3033, w_000_3034, w_000_3035, w_000_3036, w_000_3037, w_000_3038, w_000_3039, w_000_3040, w_000_3041, w_000_3042, w_000_3043, w_000_3044, w_000_3045, w_000_3046, w_000_3047, w_000_3048, w_000_3049, w_000_3050, w_000_3051, w_000_3052, w_000_3053, w_000_3054, w_000_3055, w_000_3056, w_000_3057, w_000_3058, w_000_3059, w_000_3060, w_000_3061, w_000_3062, w_000_3063, w_000_3064, w_000_3065, w_000_3066, w_000_3067, w_000_3068, w_000_3069, w_000_3070, w_000_3071, w_000_3072, w_000_3073, w_000_3074, w_000_3075, w_000_3076, w_000_3077, w_000_3078, w_000_3079, w_000_3080, w_000_3081, w_000_3082, w_000_3083, w_000_3084, w_000_3085, w_000_3086, w_000_3087, w_000_3088, w_000_3089, w_000_3090, w_000_3091, w_000_3092, w_000_3093, w_000_3094, w_000_3095, w_000_3096, w_000_3097, w_000_3098, w_000_3099, w_000_3100, w_000_3101, w_000_3102, w_000_3103, w_000_3104, w_000_3105, w_000_3106, w_000_3107, w_000_3108, w_000_3109, w_000_3110, w_000_3111, w_000_3112, w_000_3113, w_000_3114, w_000_3115, w_000_3116, w_000_3117, w_000_3118, w_000_3119, w_000_3120, w_000_3121, w_000_3122, w_000_3123, w_000_3124, w_000_3125, w_000_3126, w_000_3127, w_000_3128, w_000_3129, w_000_3130, w_000_3131, w_000_3132, w_000_3133, w_000_3134, w_000_3135, w_000_3136, w_000_3137, w_000_3138, w_000_3139, w_000_3140, w_000_3141, w_000_3142, w_000_3143, w_000_3144, w_000_3145, w_000_3146, w_000_3147, w_000_3148, w_000_3149, w_000_3150, w_000_3151, w_000_3152, w_000_3153, w_000_3154, w_000_3155, w_000_3156, w_000_3157, w_000_3158, w_000_3159, w_000_3160, w_000_3161, w_000_3162, w_000_3163, w_000_3164, w_000_3165, w_000_3166, w_000_3167, w_000_3168, w_000_3169, w_000_3170, w_000_3171, w_000_3172, w_000_3173, w_000_3174, w_000_3175, w_000_3176, w_000_3177, w_000_3178, w_000_3179, w_000_3180, w_000_3181, w_000_3182, w_000_3183, w_000_3184, w_000_3185, w_000_3186, w_000_3187, w_000_3188, w_000_3189, w_000_3190, w_000_3191, w_000_3192, w_000_3193, w_000_3194, w_000_3195, w_000_3196, w_000_3197, w_000_3198, w_000_3199, w_000_3200, w_000_3201, w_000_3202, w_000_3203, w_000_3204, w_000_3205, w_000_3206, w_000_3207, w_000_3208, w_000_3209, w_000_3210, w_000_3211, w_000_3212, w_000_3213, w_000_3214, w_000_3215, w_000_3216, w_000_3217, w_000_3218, w_000_3219, w_000_3220, w_000_3221, w_000_3222, w_000_3223, w_000_3224, w_000_3225, w_000_3226, w_000_3227, w_000_3228, w_000_3229, w_000_3230, w_000_3231, w_000_3232, w_000_3233, w_000_3234, w_000_3235, w_000_3236, w_000_3237, w_000_3238, w_000_3239, w_000_3240, w_000_3241, w_000_3242, w_000_3243, w_000_3244, w_000_3245, w_000_3246, w_000_3247, w_000_3248, w_000_3249, w_000_3250, w_000_3251, w_000_3252, w_000_3253, w_000_3254, w_000_3255, w_000_3256, w_000_3257, w_000_3258, w_000_3259, w_000_3260, w_000_3261, w_000_3262, w_000_3263, w_000_3264, w_000_3265, w_000_3266, w_000_3267, w_000_3268, w_000_3269, w_000_3270, w_000_3271, w_000_3272, w_000_3273, w_000_3274, w_000_3275, w_000_3276, w_000_3277, w_000_3278, w_000_3279, w_000_3280, w_000_3281, w_000_3282, w_000_3283, w_000_3284, w_000_3285, w_000_3286, w_000_3287, w_000_3288, w_000_3289, w_000_3290, w_000_3291, w_000_3292, w_000_3293, w_000_3294, w_000_3295, w_000_3296, w_000_3297, w_000_3298, w_000_3299, w_000_3300, w_000_3301, w_000_3302, w_000_3303, w_000_3304, w_000_3305, w_000_3306, w_000_3307, w_000_3308, w_000_3309, w_000_3310, w_000_3311, w_000_3312, w_000_3313, w_000_3314, w_000_3315, w_000_3316, w_000_3317, w_000_3318, w_000_3319, w_000_3320, w_000_3321, w_000_3322, w_000_3323, w_000_3324, w_000_3325, w_000_3326, w_000_3327, w_000_3328, w_000_3329, w_000_3330, w_000_3331, w_000_3332, w_000_3333, w_000_3334, w_000_3335, w_000_3336, w_000_3337, w_000_3338, w_000_3339, w_000_3340, w_000_3341, w_000_3342, w_000_3343, w_000_3344, w_000_3345, w_000_3346, w_000_3347, w_000_3348, w_000_3349, w_000_3350, w_000_3351, w_000_3352, w_000_3353, w_000_3354, w_000_3355, w_000_3356, w_000_3357, w_000_3358, w_000_3359, w_000_3360, w_000_3361, w_000_3362, w_000_3363, w_000_3364, w_000_3365, w_000_3366, w_000_3367, w_000_3368, w_000_3369, w_000_3370, w_000_3371, w_000_3372, w_000_3373, w_000_3374, w_000_3375, w_000_3376, w_000_3377, w_000_3378, w_000_3379, w_000_3380, w_000_3381, w_000_3382, w_000_3383, w_000_3384, w_000_3385, w_000_3386, w_000_3387, w_000_3388, w_000_3389, w_000_3390, w_000_3391, w_000_3392, w_000_3393, w_000_3394, w_000_3395, w_000_3396, w_000_3397, w_000_3398, w_000_3399, w_000_3400, w_000_3401, w_000_3402, w_000_3403, w_000_3404, w_000_3405, w_000_3406, w_000_3407, w_000_3408, w_000_3409, w_000_3410, w_000_3411, w_000_3412, w_000_3413, w_000_3414, w_000_3415, w_000_3416, w_000_3417, w_000_3418, w_000_3419, w_000_3420, w_000_3421, w_000_3422, w_000_3423, w_000_3424, w_000_3425, w_000_3426, w_000_3427, w_000_3428, w_000_3429, w_000_3430, w_000_3431, w_000_3432, w_000_3433, w_000_3434, w_000_3435, w_000_3436, w_000_3437, w_000_3438, w_000_3439, w_000_3440, w_000_3441, w_000_3442, w_000_3443, w_000_3444, w_000_3445, w_000_3446, w_000_3447, w_000_3448, w_000_3449, w_000_3450, w_000_3451, w_000_3452, w_000_3453, w_000_3454, w_000_3455, w_000_3456, w_000_3457, w_000_3458, w_000_3459, w_000_3460, w_000_3461, w_000_3462, w_000_3463, w_000_3464, w_000_3465, w_000_3466, w_000_3467, w_000_3468, w_000_3469, w_000_3470, w_000_3471, w_000_3472, w_000_3473, w_000_3474, w_000_3475, w_000_3476, w_000_3477, w_000_3478, w_000_3479, w_000_3480, w_000_3481, w_000_3482, w_000_3483, w_000_3484, w_000_3485, w_000_3486, w_000_3487, w_000_3488, w_000_3489, w_000_3490, w_000_3491, w_000_3492, w_000_3493, w_000_3494, w_000_3495, w_000_3496, w_000_3497, w_000_3498, w_000_3499, w_000_3500, w_000_3501, w_000_3502, w_000_3503, w_000_3504, w_000_3505, w_000_3506, w_000_3507, w_000_3508, w_000_3509, w_000_3510, w_000_3511, w_000_3512, w_000_3513, w_000_3514, w_000_3515, w_000_3516, w_000_3517, w_000_3518, w_000_3519, w_000_3520, w_000_3521, w_000_3522, w_000_3523, w_000_3524, w_000_3525, w_000_3526, w_000_3527, w_000_3528, w_000_3529, w_000_3530, w_000_3531, w_000_3532, w_000_3533, w_000_3534, w_000_3535, w_000_3536, w_000_3537, w_000_3538, w_000_3539, w_000_3540, w_000_3541, w_000_3542, w_000_3543, w_000_3544, w_000_3545, w_000_3546, w_000_3547, w_000_3548, w_000_3549, w_000_3550, w_000_3551, w_000_3552, w_000_3553, w_000_3554, w_000_3555, w_000_3556, w_000_3557, w_000_3558, w_000_3559, w_000_3560, w_000_3561, w_000_3562, w_000_3563, w_000_3564, w_000_3565, w_000_3566, w_000_3567, w_000_3568, w_000_3569, w_000_3570, w_000_3571, w_000_3572, w_000_3573, w_000_3574, w_000_3575, w_000_3576, w_000_3577, w_000_3578, w_000_3579, w_000_3580, w_000_3581, w_000_3582, w_000_3583, w_000_3584, w_000_3585, w_000_3586, w_000_3587, w_000_3588, w_000_3589, w_000_3590, w_000_3591, w_000_3592, w_000_3593, w_000_3594, w_000_3595, w_000_3596, w_000_3597, w_000_3598, w_000_3599, w_000_3600, w_000_3601, w_000_3602, w_000_3603, w_000_3604, w_000_3605, w_000_3606, w_000_3607, w_000_3608, w_000_3609, w_000_3610, w_000_3611, w_000_3612, w_000_3613, w_000_3614, w_000_3615, w_000_3616, w_000_3617, w_000_3618, w_000_3619, w_000_3620, w_000_3621, w_000_3622, w_000_3623, w_000_3624, w_000_3625, w_000_3626, w_000_3627, w_000_3628, w_000_3629, w_000_3630, w_000_3631, w_000_3632, w_000_3633, w_000_3634, w_000_3635, w_000_3636, w_000_3637, w_000_3638, w_000_3639, w_000_3640, w_000_3641, w_000_3642, w_000_3643, w_000_3644, w_000_3645, w_000_3646, w_000_3647, w_000_3648, w_000_3649, w_000_3650, w_000_3651, w_000_3652, w_000_3653, w_000_3654, w_000_3655, w_000_3656, w_000_3657, w_000_3658, w_000_3659, w_000_3660, w_000_3661, w_000_3662, w_000_3663, w_000_3664, w_000_3665, w_000_3666, w_000_3667, w_000_3668, w_000_3669, w_000_3670, w_000_3671, w_000_3672, w_000_3673, w_000_3674, w_000_3675, w_000_3676, w_000_3677, w_000_3678, w_000_3679, w_000_3680, w_000_3681, w_000_3682, w_000_3683, w_000_3684, w_000_3685, w_000_3686, w_000_3687, w_000_3688, w_000_3689, w_000_3690, w_000_3691, w_000_3692, w_000_3693, w_000_3694, w_000_3695, w_000_3696, w_000_3697, w_000_3698, w_000_3699, w_000_3700, w_000_3701, w_000_3702, w_000_3703, w_000_3704, w_000_3705, w_000_3706, w_000_3707, w_000_3708, w_000_3709, w_000_3710, w_000_3711, w_000_3712, w_000_3713, w_000_3714, w_000_3715, w_000_3716, w_000_3717, w_000_3718, w_000_3719, w_000_3720, w_000_3721, w_000_3722, w_000_3723, w_000_3724, w_000_3725, w_000_3726, w_000_3727, w_000_3728, w_000_3729, w_000_3730, w_000_3731, w_000_3732, w_000_3733, w_000_3734, w_000_3735, w_000_3736, w_000_3737, w_000_3738, w_000_3739, w_000_3740, w_000_3741, w_000_3742, w_000_3743, w_000_3744, w_000_3745, w_000_3746, w_000_3747, w_000_3748, w_000_3749, w_000_3750, w_000_3751, w_000_3752, w_000_3753, w_000_3754, w_000_3755, w_000_3756, w_000_3757, w_000_3758, w_000_3759, w_000_3760, w_000_3761, w_000_3762, w_000_3763, w_000_3764, w_000_3765, w_000_3766, w_000_3767, w_000_3768, w_000_3769, w_000_3770, w_000_3771, w_000_3772, w_000_3773, w_000_3774, w_000_3775, w_000_3776, w_000_3777, w_000_3778, w_000_3779, w_000_3780, w_000_3781, w_000_3782, w_000_3783, w_000_3784, w_000_3785, w_000_3786, w_000_3787, w_000_3788, w_000_3789, w_000_3790, w_000_3791, w_000_3792, w_000_3793, w_000_3794, w_000_3795, w_000_3796, w_000_3797, w_000_3798, w_000_3799, w_000_3800, w_000_3801, w_000_3802, w_000_3803, w_000_3804, w_000_3805, w_000_3806, w_000_3807, w_000_3808, w_000_3809, w_000_3810, w_000_3811, w_000_3812, w_000_3813, w_000_3814, w_000_3815, w_000_3816, w_000_3817, w_000_3818, w_000_3819, w_000_3820, w_000_3821, w_000_3822, w_000_3823, w_000_3824, w_000_3825, w_000_3826, w_000_3827, w_000_3828, w_000_3829, w_000_3830, w_000_3831, w_000_3832, w_000_3833, w_000_3834, w_000_3835, w_000_3836, w_000_3837, w_000_3838, w_000_3839, w_000_3840, w_000_3841, w_000_3842, w_000_3843, w_000_3844, w_000_3845, w_000_3846, w_000_3847, w_000_3848, w_000_3849, w_000_3850, w_000_3851, w_000_3852, w_000_3853, w_000_3854, w_000_3855, w_000_3856, w_000_3857, w_000_3858, w_000_3859, w_000_3860, w_000_3861, w_000_3862, w_000_3863, w_000_3864, w_000_3865, w_000_3866, w_000_3867, w_000_3868, w_000_3869, w_000_3870, w_000_3871, w_000_3872, w_000_3873, w_000_3874, w_000_3875, w_000_3876, w_000_3877, w_000_3878, w_000_3879, w_000_3880, w_000_3881, w_000_3882, w_000_3883, w_000_3884, w_000_3885, w_000_3886, w_000_3887, w_000_3888, w_000_3889, w_000_3890, w_000_3891, w_000_3892, w_000_3893, w_000_3894, w_000_3895, w_000_3896, w_000_3897, w_000_3898, w_000_3899, w_000_3900, w_000_3901, w_000_3902, w_000_3903, w_000_3904, w_000_3905, w_000_3906, w_000_3907, w_000_3908, w_000_3909, w_000_3910, w_000_3911, w_000_3912, w_000_3913, w_000_3914, w_000_3915, w_000_3916, w_000_3917, w_000_3918, w_000_3919, w_000_3920, w_000_3921, w_000_3922, w_000_3923, w_000_3924, w_000_3925, w_000_3926, w_000_3927, w_000_3928, w_000_3929, w_000_3930, w_000_3931, w_000_3932, w_000_3933, w_000_3934, w_000_3935, w_000_3936, w_000_3937, w_000_3938, w_000_3939, w_000_3940, w_000_3941, w_000_3942, w_000_3943, w_000_3944, w_000_3945, w_000_3946, w_000_3947, w_000_3948, w_000_3949, w_000_3950, w_000_3951, w_000_3952, w_000_3953, w_000_3954, w_000_3955, w_000_3956, w_000_3957, w_000_3958, w_000_3959, w_000_3960, w_000_3961, w_000_3962, w_000_3963, w_000_3964, w_000_3965, w_000_3966, w_000_3967, w_000_3968, w_000_3969, w_000_3970, w_000_3971, w_000_3972, w_000_3973, w_000_3974, w_000_3975, w_000_3976, w_000_3977, w_000_3978, w_000_3979, w_000_3980, w_000_3981, w_000_3982, w_000_3983, w_000_3984, w_000_3985, w_000_3986, w_000_3987, w_000_3988, w_000_3989, w_000_3990, w_000_3991, w_000_3992, w_000_3993, w_000_3994, w_000_3995, w_000_3996, w_000_3997, w_000_3998, w_000_3999, w_000_4000, w_000_4001, w_000_4002, w_000_4003, w_000_4004, w_000_4005, w_000_4006, w_000_4007, w_000_4008, w_000_4009, w_000_4010, w_000_4011, w_000_4012, w_000_4013, w_000_4014, w_000_4015, w_000_4016, w_000_4017, w_000_4018, w_000_4019, w_000_4020, w_000_4022, w_000_4023, w_000_4024, w_000_4025, w_000_4026, w_000_4027, w_000_4028, w_000_4029, w_000_4030, w_000_4031, w_000_4032, w_000_4033, w_000_4034, w_000_4035, w_000_4036, w_000_4037, w_000_4038, w_000_4039, w_000_4040, w_000_4041, w_000_4042, w_000_4043, w_000_4044, w_000_4045, w_000_4046, w_000_4047, w_000_4048, w_000_4049, w_000_4050, w_000_4051, w_000_4052, w_000_4053, w_000_4054, w_000_4055, w_000_4056, w_000_4057, w_000_4058, w_000_4059, w_000_4060, w_000_4061, w_000_4062, w_000_4063, w_000_4064, w_000_4065, w_000_4066, w_000_4067, w_000_4068, w_000_4069, w_000_4070, w_000_4071, w_000_4072, w_000_4073, w_000_4074, w_000_4075, w_000_4076, w_000_4077, w_000_4078, w_000_4079, w_000_4080, w_000_4081, w_000_4082, w_000_4083, w_000_4084, w_000_4085, w_000_4086, w_000_4087, w_000_4088, w_000_4089, w_000_4090, w_000_4091, w_000_4092, w_000_4093, w_000_4094, w_000_4095, w_000_4096, w_000_4097, w_000_4098, w_000_4099, w_000_4100, w_000_4101, w_000_4102, w_000_4103, w_000_4104, w_000_4105, w_000_4106, w_000_4107, w_000_4108, w_000_4109, w_000_4110, w_000_4111, w_000_4112, w_000_4113, w_000_4114, w_000_4115, w_000_4116, w_000_4117, w_000_4118, w_000_4119, w_000_4120, w_000_4121, w_000_4122, w_000_4123, w_000_4124, w_000_4125, w_000_4126, w_000_4127, w_000_4128, w_000_4129, w_000_4130, w_000_4131, w_000_4132, w_000_4133, w_000_4134, w_000_4135, w_000_4136, w_000_4137, w_000_4138, w_000_4139, w_000_4140, w_000_4141, w_000_4142, w_000_4143, w_000_4144, w_000_4145, w_000_4146, w_000_4147, w_000_4148, w_000_4149, w_000_4150, w_000_4151, w_000_4152, w_000_4153, w_000_4154, w_000_4155, w_000_4156, w_000_4157, w_000_4158, w_000_4159, w_000_4160, w_000_4161, w_000_4162, w_000_4163, w_000_4164, w_000_4165, w_000_4166, w_000_4167, w_000_4168, w_000_4169, w_000_4170, w_000_4171, w_000_4172, w_000_4173, w_000_4174, w_000_4175, w_000_4176, w_000_4177, w_000_4178, w_000_4179, w_000_4180, w_000_4181, w_000_4182, w_000_4183, w_000_4184, w_000_4185, w_000_4186, w_000_4187, w_000_4188, w_000_4189, w_000_4190, w_000_4191, w_000_4192, w_000_4193, w_000_4194, w_000_4195, w_000_4196, w_000_4197, w_000_4198, w_000_4199, w_000_4200, w_000_4201, w_000_4202, w_000_4203, w_000_4204, w_000_4205, w_000_4206, w_000_4207, w_000_4208, w_000_4209, w_000_4210, w_000_4211, w_000_4212, w_000_4213, w_000_4214, w_000_4215, w_000_4216, w_000_4217, w_000_4218, w_000_4219, w_000_4220, w_000_4221, w_000_4222, w_000_4223, w_000_4224, w_000_4225, w_000_4226, w_000_4227, w_000_4228, w_000_4229, w_000_4230, w_000_4231, w_000_4232, w_000_4233, w_000_4234, w_000_4235, w_000_4236, w_000_4237, w_000_4238, w_000_4239, w_000_4240, w_000_4241, w_000_4242, w_000_4243, w_000_4245, w_000_4246, w_000_4247, w_000_4248, w_000_4249, w_000_4250, w_000_4251, w_000_4252, w_000_4253, w_000_4254, w_000_4255, w_000_4256, w_000_4257, w_000_4258, w_000_4259, w_000_4260, w_000_4261, w_000_4262, w_000_4263, w_000_4264, w_000_4265, w_000_4266, w_000_4267, w_000_4268, w_000_4269, w_000_4270, w_000_4271, w_000_4272, w_000_4273, w_000_4274, w_000_4275, w_000_4276, w_000_4277, w_000_4278, w_000_4279, w_000_4280, w_000_4281, w_000_4282, w_000_4283, w_000_4284, w_000_4285, w_000_4286, w_000_4287, w_000_4288, w_000_4289, w_000_4290, w_000_4291, w_000_4292, w_000_4293, w_000_4294, w_000_4295, w_000_4296, w_000_4297, w_000_4298, w_000_4299, w_000_4300, w_000_4301, w_000_4302, w_000_4303, w_000_4304, w_000_4305, w_000_4306, w_000_4307, w_000_4308, w_000_4309, w_000_4310, w_000_4311, w_000_4312, w_000_4313, w_000_4314, w_000_4315, w_000_4316, w_000_4317, w_000_4318, w_000_4319, w_000_4320, w_000_4321, w_000_4322, w_000_4323, w_000_4324, w_000_4325, w_000_4326, w_000_4327, w_000_4328, w_000_4329, w_000_4330, w_000_4331, w_000_4332, w_000_4333, w_000_4334, w_000_4335, w_000_4336, w_000_4337, w_000_4338, w_000_4339, w_000_4340, w_000_4341, w_000_4342, w_000_4343, w_000_4344, w_000_4345, w_000_4346, w_000_4347, w_000_4348, w_000_4349, w_000_4350, w_000_4351, w_000_4352, w_000_4353, w_000_4354, w_000_4355, w_000_4356, w_000_4357, w_000_4358, w_000_4359, w_000_4360, w_000_4361, w_000_4362, w_000_4363, w_000_4364, w_000_4365, w_000_4366, w_000_4367, w_000_4368, w_000_4369, w_000_4370, w_000_4371, w_000_4372, w_000_4373, w_000_4374, w_000_4375, w_000_4376, w_000_4377, w_000_4378, w_000_4379, w_000_4380, w_000_4381, w_000_4382, w_000_4383, w_000_4384, w_000_4385, w_000_4386, w_000_4387, w_000_4388, w_000_4389, w_000_4390, w_000_4391, w_000_4392, w_000_4393, w_000_4394, w_000_4395, w_000_4396, w_000_4397, w_000_4398, w_000_4399, w_000_4400, w_000_4401, w_000_4402, w_000_4403, w_000_4404, w_000_4405, w_000_4406, w_000_4407, w_000_4408, w_000_4409, w_000_4410, w_000_4411, w_000_4412, w_000_4413, w_000_4414, w_000_4415, w_000_4416, w_000_4417, w_000_4418, w_000_4419, w_000_4420, w_000_4421, w_000_4422, w_000_4423, w_000_4424, w_000_4425, w_000_4426, w_000_4427, w_000_4428, w_000_4429, w_000_4430, w_000_4431, w_000_4432, w_000_4433, w_000_4434, w_000_4435, w_000_4436, w_000_4437, w_000_4438, w_000_4439, w_000_4440, w_000_4441, w_000_4442, w_000_4443, w_000_4444, w_000_4445, w_000_4446, w_000_4447, w_000_4448, w_000_4449, w_000_4450, w_000_4451, w_000_4452, w_000_4453, w_000_4454, w_000_4455, w_000_4456, w_000_4457, w_000_4458, w_000_4459, w_000_4460, w_000_4461, w_000_4462, w_000_4463, w_000_4464, w_000_4465, w_000_4466, w_000_4467, w_000_4468, w_000_4469, w_000_4470, w_000_4471, w_000_4472, w_000_4473, w_000_4474, w_000_4475, w_000_4476, w_000_4477, w_000_4478, w_000_4479, w_000_4480, w_000_4481, w_000_4482, w_000_4483, w_000_4484, w_000_4485, w_000_4486, w_000_4487, w_000_4488, w_000_4489, w_000_4490, w_000_4491, w_000_4492, w_000_4493, w_000_4494, w_000_4495, w_000_4496, w_000_4497, w_000_4498, w_000_4499, w_000_4500, w_000_4501, w_000_4502, w_000_4503, w_000_4504, w_000_4505, w_000_4506, w_000_4507, w_000_4508, w_000_4509, w_000_4510, w_000_4511, w_000_4512, w_000_4513, w_000_4514, w_000_4515, w_000_4516, w_000_4517, w_000_4518, w_000_4519, w_000_4520, w_000_4521, w_000_4522, w_000_4523, w_000_4524, w_000_4525, w_000_4526, w_000_4527, w_000_4528, w_000_4529, w_000_4530, w_000_4531, w_000_4532, w_000_4533, w_000_4534, w_000_4535, w_000_4536, w_000_4537, w_000_4538, w_000_4539, w_000_4540, w_000_4541, w_000_4542, w_000_4543, w_000_4544, w_000_4545, w_000_4546, w_000_4547, w_000_4548, w_000_4549, w_000_4550, w_000_4551, w_000_4552, w_000_4553, w_000_4554, w_000_4555, w_000_4556, w_000_4557, w_000_4558, w_000_4559, w_000_4560, w_000_4561, w_000_4562, w_000_4563, w_000_4564, w_000_4565, w_000_4566, w_000_4567, w_000_4568, w_000_4569, w_000_4570, w_000_4571, w_000_4572, w_000_4573, w_000_4574, w_000_4575, w_000_4576, w_000_4577, w_000_4578, w_000_4579, w_000_4580, w_000_4581, w_000_4582, w_000_4583, w_000_4584, w_000_4585, w_000_4586, w_000_4588, w_000_4589, w_000_4590, w_000_4591, w_000_4592, w_000_4593, w_000_4594, w_000_4595, w_000_4596, w_000_4597, w_000_4598, w_000_4599, w_000_4600, w_000_4601, w_000_4602, w_000_4603, w_000_4604, w_000_4605, w_000_4606, w_000_4607, w_000_4608, w_000_4609, w_000_4610, w_000_4611, w_000_4612, w_000_4613, w_000_4614, w_000_4615, w_000_4616, w_000_4617, w_000_4618, w_000_4619, w_000_4620, w_000_4621, w_000_4622, w_000_4623, w_000_4624, w_000_4625, w_000_4626, w_000_4627, w_000_4628, w_000_4629, w_000_4630, w_000_4631, w_000_4632, w_000_4633, w_000_4634, w_000_4635, w_000_4636, w_000_4637, w_000_4638, w_000_4639, w_000_4640, w_000_4641, w_000_4642, w_000_4643, w_000_4644, w_000_4645, w_000_4646, w_000_4647, w_000_4648, w_000_4649, w_000_4650, w_000_4651, w_000_4652, w_000_4653, w_000_4654, w_000_4655, w_000_4656, w_000_4657, w_000_4658, w_000_4659, w_000_4660, w_000_4661, w_000_4662, w_000_4663, w_000_4664, w_000_4665, w_000_4666, w_000_4667, w_000_4668, w_000_4669, w_000_4670, w_000_4671, w_000_4672, w_000_4673, w_000_4674, w_000_4675, w_000_4676, w_000_4677, w_000_4678, w_000_4679, w_000_4680, w_000_4681, w_000_4682, w_000_4683, w_000_4684, w_000_4685, w_000_4686, w_000_4687, w_000_4688, w_000_4689, w_000_4690, w_000_4691, w_000_4692, w_000_4693, w_000_4694, w_000_4695, w_000_4696, w_000_4697, w_000_4698, w_000_4699, w_000_4700, w_000_4701, w_000_4702, w_000_4703, w_000_4704, w_000_4705, w_000_4706, w_000_4707, w_000_4708, w_000_4709, w_000_4710, w_000_4711, w_000_4712, w_000_4713, w_000_4714, w_000_4715, w_000_4716, w_000_4717, w_000_4718, w_000_4719, w_000_4720, w_000_4721, w_000_4722, w_000_4723, w_000_4724, w_000_4725, w_000_4726, w_000_4727, w_000_4728, w_000_4729, w_000_4730, w_000_4731, w_000_4732, w_000_4733, w_000_4734, w_000_4735, w_000_4736, w_000_4737, w_000_4738, w_000_4739, w_000_4740, w_000_4741, w_000_4742, w_000_4743, w_000_4744, w_000_4745, w_000_4746, w_000_4747, w_000_4748, w_000_4749, w_000_4750, w_000_4751, w_000_4752, w_000_4753, w_000_4754, w_000_4755, w_000_4756, w_000_4757, w_000_4758, w_000_4759, w_000_4760, w_000_4761, w_000_4762, w_000_4763, w_000_4764, w_000_4765, w_000_4766, w_000_4767, w_000_4768, w_000_4769, w_000_4770, w_000_4771, w_000_4772, w_000_4773, w_000_4774, w_000_4775, w_000_4776, w_000_4777, w_000_4778, w_000_4779, w_000_4780, w_000_4781, w_000_4782, w_000_4783, w_000_4784, w_000_4785, w_000_4786, w_000_4787, w_000_4788, w_000_4789, w_000_4790, w_000_4791, w_000_4792, w_000_4793, w_000_4794, w_000_4795, w_000_4796, w_000_4797, w_000_4798, w_000_4799, w_000_4800, w_000_4801, w_000_4802, w_000_4803, w_000_4804, w_000_4805, w_000_4806, w_000_4807, w_000_4808, w_000_4809, w_000_4810, w_000_4811, w_000_4812, w_000_4813, w_000_4814, w_000_4815, w_000_4816, w_000_4817, w_000_4818, w_000_4819, w_000_4820, w_000_4821, w_000_4822, w_000_4823, w_000_4824, w_000_4825, w_000_4826, w_000_4827, w_000_4828, w_000_4829, w_000_4830, w_000_4831, w_000_4832, w_000_4833, w_000_4834, w_000_4835, w_000_4836, w_000_4837, w_000_4838, w_000_4839, w_000_4840, w_000_4841, w_000_4842, w_000_4843, w_000_4844, w_000_4845, w_000_4846, w_000_4847, w_000_4848, w_000_4849, w_000_4850, w_000_4851, w_000_4852, w_000_4853, w_000_4854, w_000_4855, w_000_4856, w_000_4857, w_000_4858, w_000_4859, w_000_4860, w_000_4861, w_000_4862, w_000_4863, w_000_4864, w_000_4865, w_000_4866, w_000_4867, w_000_4868, w_000_4869, w_000_4870, w_000_4871, w_000_4872, w_000_4873, w_000_4874, w_000_4875, w_000_4876, w_000_4877, w_000_4878, w_000_4879, w_000_4880, w_000_4881, w_000_4882, w_000_4883, w_000_4884, w_000_4885, w_000_4886, w_000_4887, w_000_4888, w_000_4889, w_000_4890, w_000_4891, w_000_4892, w_000_4893, w_000_4894, w_000_4895, w_000_4896, w_000_4897, w_000_4898, w_000_4899, w_000_4900, w_000_4901, w_000_4902, w_000_4903, w_000_4904, w_000_4905, w_000_4906, w_000_4907, w_000_4908, w_000_4909, w_000_4910, w_000_4911, w_000_4912, w_000_4913, w_000_4914, w_000_4915, w_000_4916, w_000_4917, w_000_4918, w_000_4919, w_000_4920, w_000_4921, w_000_4922, w_000_4923, w_000_4924, w_000_4925, w_000_4926, w_000_4927, w_000_4928, w_000_4929, w_000_4930, w_000_4931, w_000_4932, w_000_4933, w_000_4934, w_000_4935, w_000_4936, w_000_4937, w_000_4938, w_000_4939, w_000_4940, w_000_4941, w_000_4942, w_000_4943, w_000_4944, w_000_4945, w_000_4946, w_000_4947, w_000_4948, w_000_4949, w_000_4950, w_000_4951, w_000_4952, w_000_4953, w_000_4954, w_000_4955, w_000_4956, w_000_4957, w_000_4958, w_000_4959, w_000_4960, w_000_4961, w_000_4962, w_000_4963, w_000_4964, w_000_4965, w_000_4966, w_000_4967, w_000_4968, w_000_4969, w_000_4970, w_000_4971, w_000_4972, w_000_4973, w_000_4974, w_000_4975, w_000_4976, w_000_4977, w_000_4978, w_000_4979, w_000_4980, w_000_4981, w_000_4982, w_000_4983, w_000_4984, w_000_4985, w_000_4986, w_000_4987, w_000_4988, w_000_4989, w_000_4990, w_000_4991, w_000_4992, w_000_4993, w_000_4994, w_000_4995, w_000_4996, w_000_4997, w_000_4998, w_000_4999, w_000_5000, w_000_5001, w_000_5002, w_000_5003, w_000_5004, w_000_5005, w_000_5006, w_000_5007, w_000_5008, w_000_5009, w_000_5010, w_000_5011, w_000_5012, w_000_5013, w_000_5014, w_000_5015, w_000_5016, w_000_5017, w_000_5018, w_000_5019, w_000_5020, w_000_5021, w_000_5022, w_000_5023, w_000_5024, w_000_5025, w_000_5026, w_000_5027, w_000_5028, w_000_5029, w_000_5030, w_000_5031, w_000_5032, w_000_5033, w_000_5034, w_000_5035, w_000_5036, w_000_5037, w_000_5038, w_000_5039, w_000_5040, w_000_5041, w_000_5042, w_000_5043, w_000_5044, w_000_5045, w_000_5046, w_000_5047, w_000_5048, w_000_5049, w_000_5050, w_000_5051, w_000_5052, w_000_5053, w_000_5054, w_000_5055, w_000_5056, w_000_5057, w_000_5058, w_000_5059, w_000_5060, w_000_5061, w_000_5062, w_000_5063, w_000_5064, w_000_5065, w_000_5066, w_000_5067, w_000_5068, w_000_5069, w_000_5070, w_000_5071, w_000_5072, w_000_5073, w_000_5074, w_000_5075, w_000_5076, w_000_5077, w_000_5078, w_000_5079, w_000_5080, w_000_5081, w_000_5082, w_000_5083, w_000_5084, w_000_5085, w_000_5086, w_000_5087, w_000_5088, w_000_5089, w_000_5090, w_000_5091, w_000_5092, w_000_5093, w_000_5094, w_000_5095, w_000_5096, w_000_5097, w_000_5098, w_000_5099, w_000_5100, w_000_5101, w_000_5102, w_000_5103, w_000_5104, w_000_5105, w_000_5106, w_000_5107, w_000_5108, w_000_5109, w_000_5110, w_000_5111, w_000_5112, w_000_5113, w_000_5114, w_000_5115, w_000_5116, w_000_5117, w_000_5118, w_000_5119, w_000_5120, w_000_5121, w_000_5122, w_000_5123, w_000_5124, w_000_5125, w_000_5126, w_000_5127, w_000_5128, w_000_5129, w_000_5130, w_000_5131, w_000_5132, w_000_5133, w_000_5134, w_000_5135, w_000_5136, w_000_5137, w_000_5138, w_000_5139, w_000_5140, w_000_5141, w_000_5142, w_000_5143, w_000_5144, w_000_5145, w_000_5146, w_000_5147, w_000_5148, w_000_5149, w_000_5150, w_000_5151, w_000_5152, w_000_5153, w_000_5154, w_000_5155, w_000_5156, w_000_5157, w_000_5158, w_000_5159, w_000_5160, w_000_5161, w_000_5162, w_000_5163, w_000_5164, w_000_5165, w_000_5166, w_000_5167, w_000_5168, w_000_5169, w_000_5170, w_000_5171, w_000_5172, w_000_5173, w_000_5174, w_000_5175, w_000_5176, w_000_5177, w_000_5178, w_000_5179, w_000_5180, w_000_5181, w_000_5182, w_000_5183, w_000_5184, w_000_5185, w_000_5186, w_000_5187, w_000_5188, w_000_5189, w_000_5190, w_000_5191, w_000_5192, w_000_5193, w_000_5194, w_000_5195, w_000_5196, w_000_5197, w_000_5198, w_000_5199, w_000_5200, w_000_5201, w_000_5202, w_000_5203, w_000_5204, w_000_5205, w_000_5206, w_000_5207, w_000_5208, w_000_5209, w_000_5210, w_000_5211, w_000_5212, w_000_5213, w_000_5214, w_000_5215, w_000_5216, w_000_5217, w_000_5218, w_000_5219, w_000_5220, w_000_5221, w_000_5222, w_000_5223, w_000_5224, w_000_5225, w_000_5226, w_000_5227, w_000_5228, w_000_5229, w_000_5230, w_000_5231, w_000_5232, w_000_5233, w_000_5234, w_000_5235, w_000_5236, w_000_5237, w_000_5238, w_000_5239, w_000_5240, w_000_5241, w_000_5242, w_000_5243, w_000_5244, w_000_5245, w_000_5246, w_000_5247, w_000_5248, w_000_5249, w_000_5250, w_000_5251, w_000_5252, w_000_5253, w_000_5254, w_000_5255, w_000_5256, w_000_5257, w_000_5258, w_000_5259, w_000_5260, w_000_5261, w_000_5262, w_000_5263, w_000_5264, w_000_5265, w_000_5266, w_000_5267, w_000_5268, w_000_5269, w_000_5270, w_000_5271, w_000_5272, w_000_5273, w_000_5274, w_000_5275, w_000_5276, w_000_5277, w_000_5278, w_000_5279, w_000_5280, w_000_5281, w_000_5282, w_000_5283, w_000_5284, w_000_5285, w_000_5286, w_000_5287, w_000_5288, w_000_5289, w_000_5290, w_000_5291, w_000_5292, w_000_5293, w_000_5294, w_000_5295, w_000_5296, w_000_5297, w_000_5298, w_000_5299, w_000_5300, w_000_5301, w_000_5302, w_000_5303, w_000_5304, w_000_5305, w_000_5306, w_000_5307, w_000_5308, w_000_5309, w_000_5310, w_000_5311, w_000_5312, w_000_5313, w_000_5314, w_000_5315, w_000_5316, w_000_5317, w_000_5318, w_000_5319, w_000_5320, w_000_5321, w_000_5322, w_000_5323, w_000_5324, w_000_5325, w_000_5326, w_000_5327, w_000_5328, w_000_5329, w_000_5330, w_000_5331, w_000_5332, w_000_5333, w_000_5334, w_000_5335, w_000_5336, w_000_5337, w_000_5338, w_000_5339, w_000_5340, w_000_5341, w_000_5342, w_000_5343, w_000_5344, w_000_5345, w_000_5346, w_000_5347, w_000_5348, w_000_5349, w_000_5350, w_000_5351, w_000_5352, w_000_5353, w_000_5354, w_000_5355, w_000_5356, w_000_5357, w_000_5358, w_000_5359, w_000_5360, w_000_5361, w_000_5362, w_000_5363, w_000_5364, w_000_5365, w_000_5366, w_000_5367, w_000_5368, w_000_5369, w_000_5370, w_000_5371, w_000_5372, w_000_5373, w_000_5374, w_000_5375, w_000_5376, w_000_5377, w_000_5378, w_000_5379, w_000_5380, w_000_5381, w_000_5382, w_000_5383, w_000_5384, w_000_5385, w_000_5386, w_000_5387, w_000_5388, w_000_5389, w_000_5390, w_000_5391, w_000_5392, w_000_5393, w_000_5394, w_000_5395, w_000_5396, w_000_5397, w_000_5398, w_000_5399, w_000_5400, w_000_5401, w_000_5402, w_000_5403, w_000_5404, w_000_5405, w_000_5406, w_000_5407, w_000_5408, w_000_5409, w_000_5410, w_000_5411, w_000_5412, w_000_5413, w_000_5414, w_000_5415, w_000_5416, w_000_5417, w_000_5418, w_000_5419, w_000_5420, w_000_5421, w_000_5422, w_000_5423, w_000_5424, w_000_5425, w_000_5426, w_000_5427, w_000_5428, w_000_5429, w_000_5430, w_000_5431, w_000_5432, w_000_5433, w_000_5434, w_000_5435, w_000_5436, w_000_5437, w_000_5438, w_000_5439, w_000_5440, w_000_5441, w_000_5442, w_000_5443, w_000_5444, w_000_5445, w_000_5446, w_000_5447, w_000_5448, w_000_5449, w_000_5450, w_000_5451, w_000_5452, w_000_5453, w_000_5454, w_000_5455, w_000_5456, w_000_5457, w_000_5458, w_000_5459, w_000_5460, w_000_5461, w_000_5462, w_000_5463, w_000_5464, w_000_5465, w_000_5466, w_000_5467, w_000_5468, w_000_5469, w_000_5470, w_000_5471, w_000_5472, w_000_5473, w_000_5474, w_000_5475, w_000_5476, w_000_5477, w_000_5478, w_000_5479, w_000_5480, w_000_5481, w_000_5482, w_000_5483, w_000_5484, w_000_5485, w_000_5486, w_000_5487, w_000_5488, w_000_5489, w_000_5490, w_000_5491, w_000_5492, w_000_5493, w_000_5494, w_000_5495, w_000_5496, w_000_5497, w_000_5498, w_000_5499, w_000_5500, w_000_5501, w_000_5502, w_000_5503, w_000_5504, w_000_5505, w_000_5506, w_000_5507, w_000_5508, w_000_5509, w_000_5510, w_000_5511, w_000_5512, w_000_5513, w_000_5514, w_000_5515, w_000_5516, w_000_5517, w_000_5518, w_000_5519, w_000_5520, w_000_5521, w_000_5522, w_000_5523, w_000_5524, w_000_5525, w_000_5526, w_000_5527, w_000_5528, w_000_5529, w_000_5530, w_000_5531, w_000_5532, w_000_5533, w_000_5534, w_000_5535, w_000_5536, w_000_5537, w_000_5538, w_000_5539, w_000_5540, w_000_5541, w_000_5542, w_000_5543, w_000_5544, w_000_5545, w_000_5546, w_000_5547, w_000_5548, w_000_5549, w_000_5550, w_000_5551, w_000_5552, w_000_5553, w_000_5554, w_000_5555, w_000_5556, w_000_5557, w_000_5558, w_000_5559, w_000_5560, w_000_5561, w_000_5562, w_000_5563, w_000_5564, w_000_5565, w_000_5566, w_000_5567, w_000_5568, w_000_5569, w_000_5570, w_000_5571, w_000_5572, w_000_5573, w_000_5574, w_000_5575, w_000_5576, w_000_5577, w_000_5578, w_000_5579, w_000_5580, w_000_5581, w_000_5582, w_000_5583, w_000_5584, w_000_5585, w_000_5586, w_000_5587, w_000_5588, w_000_5589, w_000_5590, w_000_5591, w_000_5592, w_000_5593, w_000_5594, w_000_5595, w_000_5596, w_000_5597, w_000_5598, w_000_5599, w_000_5600, w_000_5601, w_000_5602, w_000_5603, w_000_5604, w_000_5605, w_000_5606, w_000_5607, w_000_5608, w_000_5609, w_000_5610, w_000_5611, w_000_5612, w_000_5613, w_000_5614, w_000_5615, w_000_5616, w_000_5617, w_000_5618, w_000_5619, w_000_5620, w_000_5621, w_000_5622, w_000_5623, w_000_5624, w_000_5625, w_000_5626, w_000_5627, w_000_5628, w_000_5629, w_000_5630, w_000_5631, w_000_5632, w_000_5633, w_000_5634, w_000_5635, w_000_5636, w_000_5637, w_000_5638, w_000_5639, w_000_5640, w_000_5641, w_000_5642, w_000_5643, w_000_5644, w_000_5645, w_000_5646, w_000_5647, w_000_5648, w_000_5649, w_000_5650, w_000_5651, w_000_5652, w_000_5653, w_000_5654, w_000_5655, w_000_5656, w_000_5657, w_000_5658, w_000_5659, w_000_5660, w_000_5661, w_000_5662, w_000_5663, w_000_5664, w_000_5665, w_000_5666, w_000_5667, w_000_5668, w_000_5669, w_000_5670, w_000_5671, w_000_5672, w_000_5673, w_000_5674, w_000_5675, w_000_5676, w_000_5677, w_000_5678, w_000_5679, w_000_5680, w_000_5681, w_000_5682, w_000_5683, w_000_5684, w_000_5685, w_000_5686, w_000_5687, w_000_5688, w_000_5689, w_000_5690, w_000_5691, w_000_5692, w_000_5693, w_000_5694, w_000_5695, w_000_5696, w_000_5697, w_000_5698, w_000_5699, w_000_5700, w_000_5701, w_000_5702, w_000_5703, w_000_5704, w_000_5705, w_000_5706, w_000_5707, w_000_5708, w_000_5709, w_000_5710, w_000_5711, w_000_5712, w_000_5713, w_000_5714, w_000_5715, w_000_5716, w_000_5717, w_000_5718, w_000_5719, w_000_5720, w_000_5721, w_000_5722, w_000_5723, w_000_5724, w_000_5725, w_000_5726, w_000_5727, w_000_5728, w_000_5729, w_000_5730, w_000_5731, w_000_5732, w_000_5733, w_000_5734, w_000_5735, w_000_5736, w_000_5737, w_000_5738, w_000_5739, w_000_5740, w_000_5741, w_000_5742, w_000_5743, w_000_5744, w_000_5745, w_000_5746, w_000_5747, w_000_5748, w_000_5749, w_000_5750, w_000_5751, w_000_5752, w_000_5753, w_000_5754, w_000_5755, w_000_5756, w_000_5757, w_000_5758, w_000_5759, w_000_5760, w_000_5761, w_000_5762, w_000_5763, w_000_5764, w_000_5765, w_000_5766, w_000_5767, w_000_5768, w_000_5769, w_000_5770, w_000_5771, w_000_5772, w_000_5773, w_000_5774, w_000_5775, w_000_5776, w_000_5777, w_000_5778, w_000_5779, w_000_5780, w_000_5781, w_000_5782, w_000_5783, w_000_5784, w_000_5785, w_000_5786, w_000_5787, w_000_5788, w_000_5789, w_000_5790, w_000_5791, w_000_5792, w_000_5793, w_000_5794, w_000_5795, w_000_5796, w_000_5797, w_000_5798, w_000_5799, w_000_5800, w_000_5801, w_000_5802, w_000_5803, w_000_5804, w_000_5805, w_000_5806, w_000_5807, w_000_5808, w_000_5809, w_000_5810, w_000_5811, w_000_5812, w_000_5813, w_000_5814, w_000_5815, w_000_5816, w_000_5817, w_000_5818, w_000_5819, w_000_5820, w_000_5821, w_000_5822, w_000_5823, w_000_5824, w_000_5825, w_000_5826, w_000_5827, w_000_5828, w_000_5829, w_000_5830, w_000_5831, w_000_5832, w_000_5833, w_000_5834, w_000_5835, w_000_5836, w_000_5837, w_000_5838, w_000_5839, w_000_5840, w_000_5841, w_000_5842, w_000_5843, w_000_5844, w_000_5845, w_000_5846, w_000_5847, w_000_5848, w_000_5849, w_000_5850, w_000_5851, w_000_5852, w_000_5853, w_000_5854, w_000_5855, w_000_5856, w_000_5857, w_000_5858, w_000_5859, w_000_5860, w_000_5861, w_000_5862, w_000_5863, w_000_5864, w_000_5865, w_000_5866, w_000_5867, w_000_5868, w_000_5869, w_000_5870, w_000_5871, w_000_5872, w_000_5873, w_000_5874, w_000_5875, w_000_5876, w_000_5877, w_000_5878, w_000_5879, w_000_5880, w_000_5881, w_000_5882, w_000_5883, w_000_5884, w_000_5885, w_000_5886, w_000_5887, w_000_5888, w_000_5889, w_000_5890, w_000_5891, w_000_5892, w_000_5893, w_000_5894, w_000_5895, w_000_5896, w_000_5897, w_000_5898, w_000_5899, w_000_5900, w_000_5901, w_000_5902, w_000_5903, w_000_5904, w_000_5905, w_000_5906, w_000_5907, w_000_5908, w_000_5909, w_000_5910, w_000_5911, w_000_5912, w_000_5913, w_000_5914, w_000_5915, w_000_5916, w_000_5917, w_000_5918, w_000_5919, w_000_5920, w_000_5921, w_000_5922, w_000_5923, w_000_5924, w_000_5925, w_000_5926, w_000_5927, w_000_5928, w_000_5929, w_000_5930, w_000_5931, w_000_5932, w_000_5933, w_000_5934, w_000_5935, w_000_5936, w_000_5937, w_000_5938, w_000_5939, w_000_5940, w_000_5941, w_000_5942, w_000_5943, w_000_5944, w_000_5945, w_000_5946, w_000_5947, w_000_5948, w_000_5949, w_000_5950, w_000_5951, w_000_5952, w_000_5953, w_000_5954, w_000_5955, w_000_5956, w_000_5957, w_000_5958, w_000_5959, w_000_5960, w_000_5961, w_000_5962, w_000_5963, w_000_5964, w_000_5965, w_000_5966, w_000_5967, w_000_5968, w_000_5969, w_000_5970, w_000_5971, w_000_5972, w_000_5973, w_000_5974, w_000_5975, w_000_5976, w_000_5977, w_000_5978, w_000_5979, w_000_5980, w_000_5981, w_000_5982, w_000_5983, w_000_5984, w_000_5985, w_000_5986, w_000_5987, w_000_5988, w_000_5989, w_000_5990, w_000_5991, w_000_5992, w_000_5993, w_000_5994, w_000_5995, w_000_5996, w_000_5997, w_000_5998, w_000_5999, w_000_6000, w_000_6001, w_000_6002, w_000_6003, w_000_6004, w_000_6005, w_000_6006, w_000_6007, w_000_6008, w_000_6009, w_000_6010, w_000_6011, w_000_6012, w_000_6013, w_000_6014, w_000_6015, w_000_6016, w_000_6017, w_000_6018, w_000_6019, w_000_6020, w_000_6021, w_000_6022, w_000_6023, w_000_6024, w_000_6025, w_000_6026, w_000_6027, w_000_6028, w_000_6029, w_000_6030, w_000_6031, w_000_6032, w_000_6033, w_000_6034, w_000_6035, w_000_6036, w_000_6037, w_000_6038, w_000_6039, w_000_6040, w_000_6041, w_000_6042, w_000_6043, w_000_6044, w_000_6045, w_000_6046, w_000_6047, w_000_6048, w_000_6049, w_000_6050, w_000_6051, w_000_6052, w_000_6053, w_000_6054, w_000_6055, w_000_6056, w_000_6057, w_000_6058, w_000_6059, w_000_6060, w_000_6061, w_000_6062, w_000_6063, w_000_6064, w_000_6065, w_000_6066, w_000_6067, w_000_6068, w_000_6069, w_000_6070, w_000_6071, w_000_6072, w_000_6073, w_000_6074, w_000_6075, w_000_6076, w_000_6077, w_000_6078, w_000_6079, w_000_6080, w_000_6081, w_000_6082, w_000_6083, w_000_6084, w_000_6085, w_000_6086, w_000_6087, w_000_6088, w_000_6089, w_000_6090, w_000_6091, w_000_6092, w_000_6093, w_000_6094, w_000_6095, w_000_6096, w_000_6097, w_000_6098, w_000_6099, w_000_6100, w_000_6101, w_000_6102, w_000_6103, w_000_6104, w_000_6105, w_000_6106, w_000_6107, w_000_6108, w_000_6109, w_000_6110, w_000_6111, w_000_6112, w_000_6113, w_000_6114, w_000_6115, w_000_6116, w_000_6117, w_000_6118, w_000_6119, w_000_6120, w_000_6121, w_000_6122, w_000_6123, w_000_6124, w_000_6125, w_000_6126, w_000_6127, w_000_6128, w_000_6129, w_000_6130, w_000_6131, w_000_6132, w_000_6133, w_000_6134, w_000_6135, w_000_6136, w_000_6137, w_000_6138, w_000_6139, w_000_6140, w_000_6141, w_000_6142, w_000_6143, w_000_6144, w_000_6145, w_000_6146, w_000_6147, w_000_6148, w_000_6149, w_000_6150, w_000_6151, w_000_6152, w_000_6153, w_000_6154, w_000_6155, w_000_6156, w_000_6157, w_000_6158, w_000_6159, w_000_6160, w_000_6161, w_000_6162, w_000_6163, w_000_6164, w_000_6165, w_000_6166, w_000_6167, w_000_6168, w_000_6169, w_000_6170, w_000_6171, w_000_6172, w_000_6173, w_000_6174, w_000_6175, w_000_6176, w_000_6177, w_000_6178, w_000_6179, w_000_6180, w_000_6181, w_000_6182, w_000_6183, w_000_6184, w_000_6185, w_000_6186, w_000_6187, w_000_6188, w_000_6189, w_000_6190, w_000_6191, w_000_6192, w_000_6193, w_000_6194, w_000_6195, w_000_6196, w_000_6197, w_000_6198, w_000_6199, w_000_6200, w_000_6201, w_000_6202, w_000_6203, w_000_6204, w_000_6205, w_000_6206, w_000_6207, w_000_6208, w_000_6209, w_000_6210, w_000_6211, w_000_6212, w_000_6213, w_000_6214, w_000_6215, w_000_6216, w_000_6217, w_000_6218, w_000_6219, w_000_6220, w_000_6221, w_000_6222, w_000_6223, w_000_6224, w_000_6225, w_000_6226, w_000_6227, w_000_6228, w_000_6229, w_000_6230, w_000_6231, w_000_6232, w_000_6233, w_000_6234, w_000_6235, w_000_6236, w_000_6237, w_000_6238, w_000_6239, w_000_6240, w_000_6241, w_000_6242, w_000_6243, w_000_6244, w_000_6245, w_000_6246, w_000_6247, w_000_6248, w_000_6249, w_000_6250, w_000_6251, w_000_6252, w_000_6253, w_000_6254, w_000_6255, w_000_6256, w_000_6257, w_000_6258, w_000_6259, w_000_6260, w_000_6261, w_000_6262, w_000_6263, w_000_6264, w_000_6265, w_000_6266, w_000_6267, w_000_6268, w_000_6269, w_000_6270, w_000_6271, w_000_6272, w_000_6273, w_000_6274, w_000_6275, w_000_6276, w_000_6277, w_000_6278, w_000_6279, w_000_6280, w_000_6281, w_000_6282, w_000_6283, w_000_6284, w_000_6285, w_000_6286, w_000_6287, w_000_6288, w_000_6289, w_000_6290, w_000_6291, w_000_6293, w_000_6294, w_000_6295, w_000_6296, w_000_6297, w_000_6298, w_000_6299, w_000_6300, w_000_6301, w_000_6302, w_000_6303, w_000_6304, w_000_6305, w_000_6306, w_000_6307, w_000_6308, w_000_6309, w_000_6310, w_000_6311, w_000_6312, w_000_6313, w_000_6314, w_000_6315, w_000_6316, w_000_6317, w_000_6318, w_000_6319, w_000_6320, w_000_6321, w_000_6322, w_000_6323, w_000_6324, w_000_6325, w_000_6326, w_000_6327, w_000_6328, w_000_6329, w_000_6330, w_000_6331, w_000_6332, w_000_6333, w_000_6334, w_000_6335, w_000_6336, w_000_6337, w_000_6338, w_000_6339, w_000_6340, w_000_6341, w_000_6342, w_000_6343, w_000_6344, w_000_6345, w_000_6346, w_000_6347, w_000_6348, w_000_6349, w_000_6350, w_000_6351, w_000_6352, w_000_6353, w_000_6354, w_000_6355, w_000_6356, w_000_6357, w_000_6358, w_000_6359, w_000_6360, w_000_6361, w_000_6362, w_000_6363, w_000_6364, w_000_6365, w_000_6366, w_000_6367, w_000_6368, w_000_6369, w_000_6370, w_000_6371, w_000_6372, w_000_6373, w_000_6374, w_000_6375, w_000_6376, w_000_6377, w_000_6378, w_000_6379, w_000_6380, w_000_6381, w_000_6382, w_000_6383, w_000_6384, w_000_6385, w_000_6386, w_000_6387, w_000_6388, w_000_6389, w_000_6390, w_000_6391, w_000_6392, w_000_6393, w_000_6394, w_000_6395, w_000_6396, w_000_6397, w_000_6398, w_000_6399, w_000_6400, w_000_6401, w_000_6402, w_000_6403, w_000_6404, w_000_6405, w_000_6406, w_000_6407, w_000_6408, w_000_6409, w_000_6410, w_000_6411, w_000_6412, w_000_6413, w_000_6414, w_000_6415, w_000_6416, w_000_6417, w_000_6418, w_000_6419, w_000_6420, w_000_6421, w_000_6422, w_000_6423, w_000_6424, w_000_6425, w_000_6426, w_000_6427, w_000_6428, w_000_6429, w_000_6430, w_000_6431, w_000_6432, w_000_6433, w_000_6434, w_000_6435, w_000_6436, w_000_6437, w_000_6438, w_000_6439, w_000_6440, w_000_6441, w_000_6442, w_000_6443, w_000_6444, w_000_6445, w_000_6446, w_000_6447, w_000_6448, w_000_6449, w_000_6450, w_000_6451, w_000_6452, w_000_6453, w_000_6454, w_000_6455, w_000_6456, w_000_6457, w_000_6458, w_000_6459, w_000_6460, w_000_6461, w_000_6462, w_000_6463, w_000_6464, w_000_6465, w_000_6466, w_000_6467, w_000_6468, w_000_6469, w_000_6470, w_000_6471, w_000_6472, w_000_6473, w_000_6474, w_000_6475, w_000_6476, w_000_6477, w_000_6478, w_000_6479, w_000_6480, w_000_6481, w_000_6482, w_000_6483, w_000_6484, w_000_6485, w_000_6486, w_000_6487, w_000_6488, w_000_6489, w_000_6490, w_000_6491, w_000_6492, w_000_6493, w_000_6494, w_000_6495, w_000_6496, w_000_6497, w_000_6498, w_000_6499, w_000_6500, w_000_6501, w_000_6502, w_000_6503, w_000_6504, w_000_6505, w_000_6506, w_000_6507, w_000_6508, w_000_6509, w_000_6510, w_000_6511, w_000_6512, w_000_6513, w_000_6514, w_000_6515, w_000_6516, w_000_6517, w_000_6518, w_000_6519, w_000_6520, w_000_6521, w_000_6522, w_000_6523, w_000_6524, w_000_6525, w_000_6526, w_000_6527, w_000_6528, w_000_6529, w_000_6530, w_000_6531, w_000_6532, w_000_6533, w_000_6534, w_000_6535, w_000_6536, w_000_6537, w_000_6538, w_000_6539, w_000_6540, w_000_6541, w_000_6542, w_000_6543, w_000_6544, w_000_6545, w_000_6546, w_000_6547, w_000_6548, w_000_6549, w_000_6550, w_000_6551, w_000_6552, w_000_6553, w_000_6554, w_000_6555, w_000_6556, w_000_6557, w_000_6558, w_000_6559, w_000_6560, w_000_6561, w_000_6562, w_000_6563, w_000_6564, w_000_6565, w_000_6566, w_000_6567, w_000_6568, w_000_6569, w_000_6570, w_000_6571, w_000_6572, w_000_6573, w_000_6574, w_000_6575, w_000_6576, w_000_6577, w_000_6578, w_000_6579, w_000_6580, w_000_6581, w_000_6582, w_000_6583, w_000_6584, w_000_6585, w_000_6586, w_000_6587, w_000_6588, w_000_6589, w_000_6590, w_000_6591, w_000_6592, w_000_6593, w_000_6594, w_000_6595, w_000_6596, w_000_6597, w_000_6598, w_000_6599, w_000_6600, w_000_6601, w_000_6602, w_000_6603, w_000_6604, w_000_6605, w_000_6606, w_000_6607, w_000_6608, w_000_6609, w_000_6610, w_000_6611, w_000_6612, w_000_6613, w_000_6614, w_000_6615, w_000_6616, w_000_6617, w_000_6618, w_000_6619, w_000_6620, w_000_6621, w_000_6622, w_000_6623, w_000_6624, w_000_6625, w_000_6626, w_000_6627, w_000_6628, w_000_6629, w_000_6630, w_000_6631, w_000_6632, w_000_6633, w_000_6634, w_000_6635, w_000_6636, w_000_6637, w_000_6638, w_000_6639, w_000_6640, w_000_6641, w_000_6642, w_000_6643, w_000_6644, w_000_6645, w_000_6646, w_000_6647, w_000_6648, w_000_6649, w_000_6650, w_000_6651, w_000_6652, w_000_6653, w_000_6654, w_000_6655, w_000_6656, w_000_6657, w_000_6658, w_000_6659, w_000_6660, w_000_6661, w_000_6662, w_000_6663, w_000_6664, w_000_6665, w_000_6666, w_000_6667, w_000_6668, w_000_6669, w_000_6670, w_000_6671, w_000_6672, w_000_6673, w_000_6674, w_000_6675, w_000_6676, w_000_6677, w_000_6678, w_000_6679, w_000_6680, w_000_6681, w_000_6682, w_000_6683, w_000_6684, w_000_6685, w_000_6686, w_000_6687, w_000_6688, w_000_6689, w_000_6690, w_000_6691, w_000_6692, w_000_6693, w_000_6694, w_000_6695, w_000_6696, w_000_6697, w_000_6698, w_000_6699, w_000_6700, w_000_6701, w_000_6702, w_000_6703, w_000_6704, w_000_6705, w_000_6706, w_000_6707, w_000_6708, w_000_6709, w_000_6710, w_000_6711, w_000_6712, w_000_6714, w_000_6715, w_000_6716, w_000_6717, w_000_6718, w_000_6719, w_000_6720, w_000_6721, w_000_6722, w_000_6723, w_000_6724, w_000_6725, w_000_6726, w_000_6727, w_000_6728, w_000_6729, w_000_6730, w_000_6731, w_000_6732, w_000_6733, w_000_6734, w_000_6735, w_000_6736, w_000_6737, w_000_6738, w_000_6739, w_000_6740, w_000_6741, w_000_6742, w_000_6743, w_000_6744, w_000_6745, w_000_6746, w_000_6747, w_000_6748, w_000_6749, w_000_6750, w_000_6751, w_000_6752, w_000_6753, w_000_6754, w_000_6755, w_000_6756, w_000_6757, w_000_6758, w_000_6759, w_000_6760, w_000_6761, w_000_6762, w_000_6763, w_000_6764, w_000_6765, w_000_6766, w_000_6767, w_000_6768, w_000_6769, w_000_6770, w_000_6771, w_000_6772, w_000_6773, w_000_6774, w_000_6775, w_000_6776, w_000_6777, w_000_6778, w_000_6779, w_000_6780, w_000_6781, w_000_6782, w_000_6783, w_000_6784, w_000_6785, w_000_6786, w_000_6787, w_000_6788, w_000_6789, w_000_6790, w_000_6791, w_000_6792, w_000_6793, w_000_6794, w_000_6795, w_000_6796, w_000_6797, w_000_6798, w_000_6799, w_000_6800, w_000_6801, w_000_6802, w_000_6803, w_000_6804, w_000_6805, w_000_6806, w_000_6807, w_000_6808, w_000_6809, w_000_6810, w_000_6811, w_000_6812, w_000_6813, w_000_6814, w_000_6815, w_000_6816, w_000_6817, w_000_6818, w_000_6819, w_000_6820, w_000_6821, w_000_6822, w_000_6823, w_000_6824, w_000_6825, w_000_6826, w_000_6827, w_000_6828, w_000_6829, w_000_6830, w_000_6831, w_000_6832, w_000_6833, w_000_6834, w_000_6835, w_000_6836, w_000_6837, w_000_6838, w_000_6839, w_000_6840, w_000_6841, w_000_6842, w_000_6843, w_000_6844, w_000_6845, w_000_6846, w_000_6847, w_000_6848, w_000_6849, w_000_6850, w_000_6851, w_000_6852, w_000_6853, w_000_6854, w_000_6855, w_000_6856, w_000_6857, w_000_6858, w_000_6859, w_000_6860, w_000_6861, w_000_6862, w_000_6863, w_000_6864, w_000_6865, w_000_6866, w_000_6867, w_000_6868, w_000_6869, w_000_6870, w_000_6871, w_000_6872, w_000_6873, w_000_6874, w_000_6875, w_000_6876, w_000_6877, w_000_6878, w_000_6879, w_000_6880, w_000_6881, w_000_6882, w_000_6883, w_000_6884, w_000_6885, w_000_6886, w_000_6887, w_000_6888, w_000_6889, w_000_6890, w_000_6891, w_000_6892, w_000_6893, w_000_6894, w_000_6895, w_000_6896, w_000_6897, w_000_6898, w_000_6899, w_000_6900, w_000_6901, w_000_6902, w_000_6903, w_000_6904, w_000_6905, w_000_6906, w_000_6907, w_000_6908, w_000_6909, w_000_6910, w_000_6911, w_000_6912, w_000_6913, w_000_6914, w_000_6915, w_000_6916, w_000_6917, w_000_6918, w_000_6919, w_000_6920, w_000_6921, w_000_6922, w_000_6923, w_000_6924, w_000_6925, w_000_6926, w_000_6927, w_000_6928, w_000_6929, w_000_6930, w_000_6931, w_000_6932, w_000_6933, w_000_6934, w_000_6935, w_000_6936, w_000_6937, w_000_6938, w_000_6939, w_000_6940, w_000_6941, w_000_6942, w_000_6943, w_000_6944, w_000_6945, w_000_6946, w_000_6947, w_000_6948, w_000_6949, w_000_6950, w_000_6951, w_000_6952, w_000_6953, w_000_6954, w_000_6955, w_000_6956, w_000_6957, w_000_6958, w_000_6959, w_000_6960, w_000_6961, w_000_6962, w_000_6963, w_000_6964, w_000_6965, w_000_6966, w_000_6967, w_000_6968, w_000_6969, w_000_6970, w_000_6971, w_000_6972, w_000_6973, w_000_6974, w_000_6975, w_000_6976, w_000_6977, w_000_6978, w_000_6979, w_000_6980, w_000_6981, w_000_6982, w_000_6983, w_000_6984, w_000_6985, w_000_6986, w_000_6987, w_000_6988, w_000_6989, w_000_6990, w_000_6991, w_000_6992, w_000_6993, w_000_6994, w_000_6995, w_000_6996, w_000_6997, w_000_6998, w_000_6999, w_000_7000, w_000_7001, w_000_7002, w_000_7003, w_000_7004, w_000_7005, w_000_7006, w_000_7007, w_000_7008, w_000_7009, w_000_7010, w_000_7011, w_000_7012, w_000_7013, w_000_7014, w_000_7015, w_000_7016, w_000_7017, w_000_7018, w_000_7019, w_000_7020, w_000_7021, w_000_7022, w_000_7023, w_000_7024, w_000_7025, w_000_7026, w_000_7027, w_000_7028, w_000_7029, w_000_7030, w_000_7031, w_000_7032, w_000_7033, w_000_7034, w_000_7035, w_000_7036, w_000_7037, w_000_7038, w_000_7039, w_000_7040, w_000_7041, w_000_7042, w_000_7043, w_000_7044, w_000_7045, w_000_7046, w_000_7047, w_000_7048, w_000_7049, w_000_7050, w_000_7051, w_000_7052, w_000_7053, w_000_7054, w_000_7055, w_000_7056, w_000_7057, w_000_7058, w_000_7059, w_000_7060, w_000_7061, w_000_7062, w_000_7063, w_000_7064, w_000_7065, w_000_7066, w_000_7067, w_000_7068, w_000_7069, w_000_7070, w_000_7071, w_000_7072, w_000_7073, w_000_7074, w_000_7075, w_000_7076, w_000_7077, w_000_7078, w_000_7079, w_000_7080, w_000_7081, w_000_7082, w_000_7083, w_000_7084, w_000_7085, w_000_7086, w_000_7087, w_000_7088, w_000_7089, w_000_7090, w_000_7091, w_000_7092, w_000_7093, w_000_7094, w_000_7095, w_000_7096, w_000_7097, w_000_7098, w_000_7099, w_000_7100, w_000_7101, w_000_7102, w_000_7103, w_000_7104, w_000_7105, w_000_7106, w_000_7107, w_000_7108, w_000_7109, w_000_7110, w_000_7111, w_000_7112, w_000_7113, w_000_7114, w_000_7115, w_000_7116, w_000_7117, w_000_7118, w_000_7119, w_000_7120, w_000_7121, w_000_7122, w_000_7123, w_000_7124, w_000_7125, w_000_7126, w_000_7127, w_000_7128, w_000_7129, w_000_7130, w_000_7131, w_000_7132, w_000_7133, w_000_7134, w_000_7135, w_000_7136, w_000_7137, w_000_7138, w_000_7139, w_000_7140, w_000_7141, w_000_7142, w_000_7143, w_000_7144, w_000_7145, w_000_7146, w_000_7147, w_000_7148, w_000_7149, w_000_7150, w_000_7151, w_000_7152, w_000_7153, w_000_7154, w_000_7155, w_000_7156, w_000_7157, w_000_7158, w_000_7159, w_000_7160, w_000_7161, w_000_7162, w_000_7163, w_000_7164, w_000_7165, w_000_7166, w_000_7167, w_000_7168, w_000_7169, w_000_7170, w_000_7171, w_000_7172, w_000_7173, w_000_7174, w_000_7175, w_000_7176, w_000_7177, w_000_7178, w_000_7179, w_000_7180, w_000_7181, w_000_7182, w_000_7183, w_000_7184, w_000_7185, w_000_7186, w_000_7187, w_000_7188, w_000_7189, w_000_7190, w_000_7191, w_000_7192, w_000_7193, w_000_7194, w_000_7195, w_000_7196, w_000_7197, w_000_7198, w_000_7199, w_000_7200, w_000_7201, w_000_7202, w_000_7203, w_000_7204, w_000_7205, w_000_7206, w_000_7207, w_000_7208, w_000_7209, w_000_7210, w_000_7211, w_000_7212, w_000_7213, w_000_7214, w_000_7215, w_000_7216, w_000_7217, w_000_7218, w_000_7219, w_000_7220, w_000_7221, w_000_7222, w_000_7223, w_000_7224, w_000_7225, w_000_7226, w_000_7227, w_000_7228, w_000_7229, w_000_7230, w_000_7231, w_000_7232, w_000_7233, w_000_7234, w_000_7235, w_000_7236, w_000_7237, w_000_7238, w_000_7239, w_000_7240, w_000_7241, w_000_7242, w_000_7243, w_000_7244, w_000_7245, w_000_7246, w_000_7247, w_000_7248, w_000_7249, w_000_7250, w_000_7251, w_000_7252, w_000_7253, w_000_7254, w_000_7255, w_000_7256, w_000_7257, w_000_7258, w_000_7259, w_000_7260, w_000_7261, w_000_7262, w_000_7263, w_000_7264, w_000_7265, w_000_7266, w_000_7267, w_000_7268, w_000_7269, w_000_7270, w_000_7271, w_000_7272, w_000_7273, w_000_7274, w_000_7275, w_000_7276, w_000_7277, w_000_7278, w_000_7279, w_000_7280, w_000_7281, w_000_7282, w_000_7283, w_000_7284, w_000_7285, w_000_7286, w_000_7287, w_000_7288, w_000_7289, w_000_7290, w_000_7291, w_000_7292, w_000_7293, w_000_7294, w_000_7295, w_000_7296, w_000_7297, w_000_7298, w_000_7299, w_000_7300, w_000_7301, w_000_7302, w_000_7303, w_000_7304, w_000_7305, w_000_7306, w_000_7307, w_000_7308, w_000_7309, w_000_7310, w_000_7311, w_000_7312, w_000_7313, w_000_7314, w_000_7315, w_000_7316, w_000_7317, w_000_7318, w_000_7319, w_000_7320, w_000_7321, w_000_7322, w_000_7323, w_000_7324, w_000_7325, w_000_7326, w_000_7327, w_000_7328, w_000_7329, w_000_7330, w_000_7331, w_000_7332, w_000_7333, w_000_7334, w_000_7335, w_000_7336, w_000_7337, w_000_7338, w_000_7339, w_000_7340, w_000_7341, w_000_7342, w_000_7343, w_000_7344, w_000_7345, w_000_7346, w_000_7347, w_000_7348, w_000_7349, w_000_7350, w_000_7351, w_000_7352, w_000_7353, w_000_7354, w_000_7355, w_000_7356, w_000_7357, w_000_7358, w_000_7359, w_000_7360, w_000_7361, w_000_7362, w_000_7363, w_000_7364, w_000_7365, w_000_7366, w_000_7367, w_000_7368, w_000_7369, w_000_7370, w_000_7371, w_000_7372, w_000_7373, w_000_7374, w_000_7375, w_000_7376, w_000_7377, w_000_7378, w_000_7379, w_000_7380, w_000_7381, w_000_7382, w_000_7383, w_000_7384, w_000_7385, w_000_7386, w_000_7387, w_000_7388, w_000_7389, w_000_7390, w_000_7391, w_000_7392, w_000_7393, w_000_7394, w_000_7395, w_000_7396, w_000_7397, w_000_7398, w_000_7399, w_000_7400, w_000_7401, w_000_7402, w_000_7403, w_000_7404, w_000_7405, w_000_7406, w_000_7407, w_000_7408, w_000_7409, w_000_7410, w_000_7411, w_000_7412, w_000_7413, w_000_7414, w_000_7415, w_000_7416, w_000_7417, w_000_7418, w_000_7419, w_000_7420, w_000_7421, w_000_7422, w_000_7423, w_000_7424, w_000_7425, w_000_7426, w_000_7427, w_000_7428, w_000_7429, w_000_7430, w_000_7431, w_000_7432, w_000_7433, w_000_7434, w_000_7435, w_000_7436, w_000_7437, w_000_7438, w_000_7439, w_000_7440, w_000_7441, w_000_7442, w_000_7443, w_000_7444, w_000_7445, w_000_7446, w_000_7447, w_000_7448, w_000_7449, w_000_7450, w_000_7451, w_000_7452, w_000_7453, w_000_7454, w_000_7455, w_000_7456, w_000_7457, w_000_7458, w_000_7459, w_000_7460, w_000_7461, w_000_7462, w_000_7463, w_000_7464, w_000_7465, w_000_7466, w_000_7467, w_000_7468, w_000_7469, w_000_7470, w_000_7471, w_000_7472, w_000_7473, w_000_7474, w_000_7475, w_000_7476, w_000_7477, w_000_7478, w_000_7479, w_000_7480, w_000_7481, w_000_7482, w_000_7483, w_000_7484, w_000_7485, w_000_7486, w_000_7487, w_000_7488, w_000_7489, w_000_7490, w_000_7491, w_000_7492, w_000_7493, w_000_7494, w_000_7495, w_000_7496, w_000_7497, w_000_7498, w_000_7499, w_000_7500, w_000_7501, w_000_7502, w_000_7503, w_000_7504, w_000_7505, w_000_7506, w_000_7507, w_000_7508, w_000_7509, w_000_7510, w_000_7511, w_000_7512, w_000_7513, w_000_7514, w_000_7515, w_000_7516, w_000_7517, w_000_7518, w_000_7519, w_000_7520, w_000_7521, w_000_7522, w_000_7523, w_000_7524, w_000_7525, w_000_7526, w_000_7527, w_000_7528, w_000_7529, w_000_7530, w_000_7531, w_000_7532, w_000_7533, w_000_7534, w_000_7535, w_000_7536, w_000_7537, w_000_7538, w_000_7539, w_000_7540, w_000_7541, w_000_7542, w_000_7543, w_000_7544, w_000_7545, w_000_7546, w_000_7547, w_000_7548, w_000_7549, w_000_7550, w_000_7551, w_000_7552, w_000_7553, w_000_7554, w_000_7555, w_000_7556, w_000_7557, w_000_7558, w_000_7559, w_000_7560, w_000_7561, w_000_7562, w_000_7563, w_000_7564, w_000_7565, w_000_7566, w_000_7567, w_000_7568, w_000_7569, w_000_7570, w_000_7571, w_000_7572, w_000_7573, w_000_7574, w_000_7575, w_000_7576, w_000_7577, w_000_7578, w_000_7579, w_000_7580, w_000_7581, w_000_7582, w_000_7583, w_000_7584, w_000_7585, w_000_7586, w_000_7587, w_000_7588, w_000_7589, w_000_7590, w_000_7591, w_000_7592, w_000_7593, w_000_7594, w_000_7595, w_000_7596, w_000_7597, w_000_7598, w_000_7599, w_000_7600, w_000_7601, w_000_7602, w_000_7603, w_000_7604, w_000_7605, w_000_7606, w_000_7607, w_000_7608, w_000_7610, w_000_7611, w_000_7612, w_000_7613, w_000_7614, w_000_7615, w_000_7616, w_000_7617, w_000_7618, w_000_7619, w_000_7620, w_000_7621, w_000_7622, w_000_7623, w_000_7624, w_000_7625, w_000_7626, w_000_7627, w_000_7628, w_000_7629, w_000_7630, w_000_7631, w_000_7632, w_000_7633, w_000_7634, w_000_7635, w_000_7636, w_000_7637, w_000_7638, w_000_7639, w_000_7640, w_000_7641, w_000_7642, w_000_7643, w_000_7644, w_000_7645, w_000_7646, w_000_7647, w_000_7648, w_000_7649, w_000_7650, w_000_7651, w_000_7652, w_000_7653, w_000_7654, w_000_7655, w_000_7656, w_000_7657, w_000_7658, w_000_7659, w_000_7660, w_000_7661, w_000_7662, w_000_7663, w_000_7664, w_000_7665, w_000_7666, w_000_7667, w_000_7668, w_000_7669, w_000_7670, w_000_7671, w_000_7672, w_000_7673, w_000_7674, w_000_7675, w_000_7676, w_000_7677, w_000_7678, w_000_7679, w_000_7680, w_000_7681, w_000_7682, w_000_7683, w_000_7684, w_000_7685, w_000_7686, w_000_7687, w_000_7688, w_000_7689, w_000_7690, w_000_7692, w_000_7693, w_000_7694, w_000_7695, w_000_7696, w_000_7697, w_000_7698, w_000_7699, w_000_7700, w_000_7701, w_000_7702, w_000_7703, w_000_7704, w_000_7705, w_000_7706, w_000_7707, w_000_7708, w_000_7709, w_000_7710, w_000_7711, w_000_7712, w_000_7713, w_000_7714, w_000_7715, w_000_7716, w_000_7717, w_000_7718, w_000_7719, w_000_7720, w_000_7721, w_000_7722, w_000_7723, w_000_7724, w_000_7725, w_000_7726, w_000_7727, w_000_7728, w_000_7729, w_000_7730, w_000_7731, w_000_7732, w_000_7733, w_000_7734, w_000_7735, w_000_7736, w_000_7737, w_000_7738, w_000_7739, w_000_7740, w_000_7741, w_000_7742, w_000_7743, w_000_7744, w_000_7745, w_000_7746, w_000_7747, w_000_7748, w_000_7749, w_000_7750, w_000_7751, w_000_7752, w_000_7753, w_000_7754, w_000_7755, w_000_7756, w_000_7757, w_000_7758, w_000_7759, w_000_7760, w_000_7761, w_000_7762, w_000_7763, w_000_7764, w_000_7765, w_000_7766, w_000_7767, w_000_7768, w_000_7769, w_000_7770, w_000_7771, w_000_7772, w_000_7773, w_000_7774, w_000_7775, w_000_7776, w_000_7777, w_000_7778, w_000_7779, w_000_7780, w_000_7781, w_000_7782, w_000_7784, w_000_7785, w_000_7786, w_000_7787, w_000_7788, w_000_7789, w_000_7790, w_000_7791, w_000_7792, w_000_7793, w_000_7794, w_000_7795, w_000_7796, w_000_7797, w_000_7799, w_000_7800, w_000_7801, w_000_7802, w_000_7803, w_000_7804, w_000_7805, w_000_7806, w_000_7807, w_000_7808, w_000_7809, w_000_7810, w_000_7811, w_000_7812, w_000_7813, w_000_7814, w_000_7815, w_000_7816, w_000_7817, w_000_7818, w_000_7819, w_000_7820, w_000_7821, w_000_7822, w_000_7823, w_000_7824, w_000_7825, w_000_7826, w_000_7827, w_000_7828, w_000_7829, w_000_7830, w_000_7831, w_000_7832, w_000_7833, w_000_7834, w_000_7835, w_000_7836, w_000_7837, w_000_7838, w_000_7839, w_000_7840, w_000_7841, w_000_7842, w_000_7843, w_000_7844, w_000_7845, w_000_7846, w_000_7847, w_000_7848, w_000_7849, w_000_7850, w_000_7851, w_000_7852, w_000_7853, w_000_7854, w_000_7855, w_000_7856, w_000_7857, w_000_7858, w_000_7859, w_000_7860, w_000_7861, w_000_7862, w_000_7863, w_000_7864, w_000_7865, w_000_7866, w_000_7867, w_000_7868, w_000_7869, w_000_7870, w_000_7871, w_000_7872, w_000_7874, w_000_7875, w_000_7876, w_000_7877, w_000_7878, w_000_7879, w_000_7880, w_000_7881, w_000_7882, w_000_7883, w_000_7884, w_000_7885, w_000_7886, w_000_7887, w_000_7888, w_000_7889, w_000_7890, w_000_7891, w_000_7892, w_000_7893, w_000_7894, w_000_7895, w_000_7896, w_000_7897, w_000_7898, w_000_7899, w_000_7900, w_000_7901, w_000_7902, w_000_7903, w_000_7904, w_000_7905, w_000_7906, w_000_7907, w_000_7908, w_000_7909, w_000_7910, w_000_7911, w_000_7912, w_000_7913, w_000_7914, w_000_7915, w_000_7916, w_000_7917, w_000_7918, w_000_7919, w_000_7920, w_000_7921, w_000_7922, w_000_7923, w_000_7924, w_000_7925, w_000_7926, w_000_7927, w_000_7928, w_000_7929, w_000_7930, w_000_7931, w_000_7932, w_000_7933, w_000_7934, w_000_7935, w_000_7936, w_000_7937, w_000_7938, w_000_7939, w_000_7940, w_000_7941, w_000_7942, w_000_7943, w_000_7944, w_000_7945, w_000_7946, w_000_7947, w_000_7948, w_000_7949, w_000_7950, w_000_7951, w_000_7952, w_000_7953, w_000_7954, w_000_7955, w_000_7956, w_000_7957, w_000_7958, w_000_7959, w_000_7960, w_000_7961, w_000_7962, w_000_7963, w_000_7964, w_000_7965, w_000_7966, w_000_7967, w_000_7968, w_000_7969, w_000_7970, w_000_7971, w_000_7972, w_000_7973, w_000_7974, w_000_7975, w_000_7976, w_000_7977, w_000_7978, w_000_7979, w_000_7980, w_000_7981, w_000_7982, w_000_7983, w_000_7984, w_000_7985, w_000_7986, w_000_7987, w_000_7988, w_000_7989, w_000_7990, w_000_7991, w_000_7992, w_000_7993, w_000_7994, w_000_7995, w_000_7996, w_000_7997, w_000_7998, w_000_7999, w_000_8000, w_000_8001, w_000_8002, w_000_8003, w_000_8004, w_000_8005, w_000_8006, w_000_8007, w_000_8008, w_000_8009, w_000_8010, w_000_8011, w_000_8012, w_000_8013, w_000_8014, w_000_8015, w_000_8016, w_000_8017, w_000_8018, w_000_8019, w_000_8020, w_000_8021, w_000_8022, w_000_8023, w_000_8024, w_000_8025, w_000_8026, w_000_8027, w_000_8028, w_000_8029, w_000_8030, w_000_8031, w_000_8032, w_000_8033, w_000_8034, w_000_8035, w_000_8036, w_000_8037, w_000_8038, w_000_8039, w_000_8040, w_000_8041, w_000_8042, w_000_8043, w_000_8044, w_000_8045, w_000_8046, w_000_8047, w_000_8048, w_000_8049, w_000_8050, w_000_8051, w_000_8052, w_000_8053, w_000_8054, w_000_8055, w_000_8056, w_000_8057, w_000_8058, w_000_8059, w_000_8060, w_000_8061, w_000_8062, w_000_8063, w_000_8064, w_000_8065, w_000_8066, w_000_8067, w_000_8068, w_000_8069, w_000_8070, w_000_8071, w_000_8072, w_000_8073, w_000_8074, w_000_8075, w_000_8076, w_000_8077, w_000_8078, w_000_8079, w_000_8080, w_000_8081, w_000_8082, w_000_8083, w_000_8084, w_000_8085, w_000_8086, w_000_8087, w_000_8088, w_000_8089, w_000_8090, w_000_8091, w_000_8092, w_000_8093, w_000_8094, w_000_8095, w_000_8096, w_000_8097, w_000_8098, w_000_8099, w_000_8100, w_000_8101, w_000_8102, w_000_8103, w_000_8104, w_000_8105, w_000_8106, w_000_8107, w_000_8108, w_000_8109, w_000_8110, w_000_8111, w_000_8112, w_000_8113, w_000_8114, w_000_8115, w_000_8116, w_000_8117, w_000_8118, w_000_8119, w_000_8120, w_000_8121, w_000_8122, w_000_8123, w_000_8124, w_000_8125, w_000_8126, w_000_8127, w_000_8128, w_000_8129, w_000_8130, w_000_8131, w_000_8132, w_000_8133, w_000_8134, w_000_8135, w_000_8136, w_000_8137, w_000_8138, w_000_8139, w_000_8140, w_000_8141, w_000_8142, w_000_8143, w_000_8144, w_000_8145, w_000_8146, w_000_8147, w_000_8148, w_000_8149, w_000_8150, w_000_8151, w_000_8152, w_000_8153, w_000_8154, w_000_8155, w_000_8156, w_000_8157, w_000_8158, w_000_8159, w_000_8160, w_000_8161, w_000_8162, w_000_8163, w_000_8164, w_000_8165, w_000_8166, w_000_8167, w_000_8168, w_000_8169, w_000_8170, w_000_8171, w_000_8172, w_000_8173, w_000_8174, w_000_8175, w_000_8176, w_000_8177, w_000_8178, w_000_8179, w_000_8180, w_000_8181, w_000_8182, w_000_8183, w_000_8184, w_000_8185, w_000_8186, w_000_8187, w_000_8188, w_000_8189, w_000_8190, w_000_8191, w_000_8192, w_000_8193, w_000_8194, w_000_8195, w_000_8196, w_000_8197, w_000_8198, w_000_8199, w_000_8200, w_000_8201, w_000_8202, w_000_8203, w_000_8204, w_000_8205, w_000_8206, w_000_8207, w_000_8208, w_000_8209, w_000_8210, w_000_8211, w_000_8212, w_000_8213, w_000_8214, w_000_8215, w_000_8216, w_000_8217, w_000_8218, w_000_8219, w_000_8220, w_000_8221, w_000_8222, w_000_8223, w_000_8224, w_000_8225, w_000_8226, w_000_8227, w_000_8228, w_000_8229, w_000_8230, w_000_8231, w_000_8232, w_000_8233, w_000_8234, w_000_8235, w_000_8236, w_000_8237, w_000_8238, w_000_8239, w_000_8240, w_000_8241, w_000_8242, w_000_8243, w_000_8244, w_000_8245, w_000_8246, w_000_8247, w_000_8248, w_000_8249, w_000_8250, w_000_8251, w_000_8252, w_000_8253, w_000_8254, w_000_8255, w_000_8256, w_000_8257, w_000_8258, w_000_8259, w_000_8260, w_000_8261, w_000_8262, w_000_8263, w_000_8264, w_000_8265, w_000_8266, w_000_8267, w_000_8268, w_000_8269, w_000_8270, w_000_8271, w_000_8272, w_000_8273, w_000_8274, w_000_8275, w_000_8276, w_000_8277, w_000_8278, w_000_8279, w_000_8280, w_000_8281, w_000_8282, w_000_8283, w_000_8284, w_000_8285, w_000_8286, w_000_8287, w_000_8288, w_000_8289, w_000_8290, w_000_8291, w_000_8292, w_000_8293, w_000_8294, w_000_8295, w_000_8296, w_000_8297, w_000_8298, w_000_8299, w_000_8300, w_000_8301, w_000_8302, w_000_8303, w_000_8304, w_000_8305, w_000_8306, w_000_8307, w_000_8308, w_000_8309, w_000_8310, w_000_8311, w_000_8312, w_000_8313, w_000_8314, w_000_8315, w_000_8316, w_000_8317, w_000_8318, w_000_8319, w_000_8320, w_000_8321, w_000_8322, w_000_8323, w_000_8324, w_000_8325, w_000_8326, w_000_8327, w_000_8328, w_000_8329, w_000_8330, w_000_8331, w_000_8332, w_000_8333, w_000_8334, w_000_8335, w_000_8336, w_000_8337, w_000_8338, w_000_8339, w_000_8340, w_000_8341, w_000_8342, w_000_8343, w_000_8344, w_000_8345, w_000_8346, w_000_8347, w_000_8348, w_000_8349, w_000_8350, w_000_8351, w_000_8352, w_000_8353, w_000_8354, w_000_8355, w_000_8356, w_000_8357, w_000_8358, w_000_8359, w_000_8360, w_000_8361, w_000_8362, w_000_8363, w_000_8364, w_000_8365, w_000_8366, w_000_8367, w_000_8368, w_000_8369, w_000_8370, w_000_8371, w_000_8372, w_000_8373, w_000_8374, w_000_8375, w_000_8376, w_000_8377, w_000_8378, w_000_8379, w_000_8380, w_000_8381, w_000_8382, w_000_8383, w_000_8384, w_000_8385, w_000_8386, w_000_8387, w_000_8388, w_000_8389, w_000_8390, w_000_8391, w_000_8392, w_000_8393, w_000_8394, w_000_8395, w_000_8396, w_000_8397, w_000_8398, w_000_8399, w_000_8400, w_000_8401, w_000_8402, w_000_8403, w_000_8404, w_000_8405, w_000_8406, w_000_8407, w_000_8408, w_000_8409, w_000_8410, w_000_8411, w_000_8412, w_000_8413, w_000_8414, w_000_8415, w_000_8416, w_000_8417, w_000_8418, w_000_8419, w_000_8420, w_000_8421, w_000_8422, w_000_8423, w_000_8424, w_000_8425, w_000_8426, w_000_8427, w_000_8428, w_000_8429, w_000_8430, w_000_8431, w_000_8432, w_000_8433, w_000_8434, w_000_8435, w_000_8436, w_000_8437, w_000_8438, w_000_8439, w_000_8440, w_000_8441, w_000_8442, w_000_8443, w_000_8444, w_000_8445, w_000_8446, w_000_8447, w_000_8448, w_000_8449, w_000_8450, w_000_8451, w_000_8452, w_000_8453, w_000_8454, w_000_8455, w_000_8456, w_000_8457, w_000_8458, w_000_8459, w_000_8460, w_000_8461, w_000_8462, w_000_8463, w_000_8464, w_000_8465, w_000_8466, w_000_8467, w_000_8468, w_000_8469, w_000_8470, w_000_8471, w_000_8472, w_000_8473, w_000_8474, w_000_8475, w_000_8476, w_000_8477, w_000_8478, w_000_8479, w_000_8480, w_000_8481, w_000_8482, w_000_8483, w_000_8484, w_000_8485, w_000_8486, w_000_8487, w_000_8488, w_000_8489, w_000_8490, w_000_8491, w_000_8492, w_000_8493, w_000_8494, w_000_8495, w_000_8496, w_000_8497, w_000_8498, w_000_8499, w_000_8500, w_000_8501, w_000_8502, w_000_8503, w_000_8504, w_000_8505, w_000_8506, w_000_8507, w_000_8508, w_000_8509, w_000_8510, w_000_8511, w_000_8512, w_000_8513, w_000_8514, w_000_8515, w_000_8516, w_000_8517, w_000_8518, w_000_8519, w_000_8520, w_000_8521, w_000_8522, w_000_8523, w_000_8524, w_000_8525, w_000_8526, w_000_8527, w_000_8528, w_000_8529, w_000_8530, w_000_8531, w_000_8532, w_000_8533, w_000_8534, w_000_8535, w_000_8536, w_000_8537, w_000_8538, w_000_8539, w_000_8540, w_000_8541, w_000_8542, w_000_8543, w_000_8544, w_000_8545, w_000_8546, w_000_8547, w_000_8548, w_000_8549, w_000_8550, w_000_8551, w_000_8552, w_000_8553, w_000_8554, w_000_8555, w_000_8556, w_000_8557, w_000_8558, w_000_8559, w_000_8560, w_000_8561, w_000_8562, w_000_8563, w_000_8564, w_000_8565, w_000_8566, w_000_8567, w_000_8568, w_000_8569, w_000_8570, w_000_8571, w_000_8572, w_000_8573, w_000_8574, w_000_8575, w_000_8576, w_000_8577, w_000_8578, w_000_8579, w_000_8580, w_000_8581, w_000_8582, w_000_8583, w_000_8584, w_000_8585, w_000_8586, w_000_8587, w_000_8588, w_000_8589, w_000_8590, w_000_8591, w_000_8592, w_000_8593, w_000_8594, w_000_8595, w_000_8596, w_000_8597, w_000_8598, w_000_8599, w_000_8600, w_000_8601, w_000_8602, w_000_8603, w_000_8604, w_000_8605, w_000_8606, w_000_8607, w_000_8608, w_000_8609, w_000_8610, w_000_8611, w_000_8612, w_000_8613, w_000_8614, w_000_8615, w_000_8616, w_000_8617, w_000_8618, w_000_8619, w_000_8620, w_000_8621, w_000_8622, w_000_8623, w_000_8624, w_000_8625, w_000_8626, w_000_8627, w_000_8628, w_000_8629, w_000_8630, w_000_8631, w_000_8632, w_000_8633, w_000_8634, w_000_8635, w_000_8636, w_000_8637, w_000_8638, w_000_8639, w_000_8640, w_000_8641, w_000_8642, w_000_8643, w_000_8644, w_000_8645, w_000_8646, w_000_8647, w_000_8648, w_000_8649, w_000_8650, w_000_8651, w_000_8652, w_000_8653, w_000_8654, w_000_8655, w_000_8656, w_000_8657, w_000_8658, w_000_8659, w_000_8660, w_000_8661, w_000_8662, w_000_8663, w_000_8664, w_000_8665, w_000_8666, w_000_8667, w_000_8668, w_000_8669, w_000_8670, w_000_8671, w_000_8672, w_000_8673, w_000_8674, w_000_8675, w_000_8676, w_000_8677, w_000_8678, w_000_8679, w_000_8680, w_000_8681, w_000_8682, w_000_8683, w_000_8684, w_000_8685, w_000_8686, w_000_8687, w_000_8688, w_000_8689, w_000_8690, w_000_8691, w_000_8692, w_000_8693, w_000_8694, w_000_8695, w_000_8696, w_000_8697, w_000_8698, w_000_8699, w_000_8700, w_000_8701, w_000_8702, w_000_8703, w_000_8704, w_000_8705, w_000_8706, w_000_8707, w_000_8708, w_000_8709, w_000_8710, w_000_8711, w_000_8712, w_000_8713, w_000_8714, w_000_8715, w_000_8716, w_000_8717, w_000_8718, w_000_8719, w_000_8720, w_000_8721, w_000_8722, w_000_8723, w_000_8724, w_000_8725, w_000_8726, w_000_8728, w_000_8729, w_000_8730, w_000_8731, w_000_8732, w_000_8733, w_000_8734, w_000_8735, w_000_8736, w_000_8737, w_000_8738, w_000_8739, w_000_8740, w_000_8741, w_000_8742, w_000_8743, w_000_8744, w_000_8745, w_000_8746, w_000_8747, w_000_8748, w_000_8749, w_000_8751, w_000_8752, w_000_8753, w_000_8754, w_000_8755, w_000_8756, w_000_8757, w_000_8758, w_000_8759, w_000_8760, w_000_8761, w_000_8762, w_000_8763, w_000_8764, w_000_8765, w_000_8766, w_000_8767, w_000_8768, w_000_8769, w_000_8770, w_000_8771, w_000_8772, w_000_8773, w_000_8774, w_000_8775, w_000_8776, w_000_8777, w_000_8778, w_000_8779, w_000_8780, w_000_8781, w_000_8782, w_000_8783, w_000_8784, w_000_8785, w_000_8786, w_000_8787, w_000_8788, w_000_8789, w_000_8790, w_000_8791, w_000_8792, w_000_8793, w_000_8794, w_000_8795, w_000_8796, w_000_8797, w_000_8798, w_000_8799, w_000_8800, w_000_8801, w_000_8802, w_000_8803, w_000_8804, w_000_8805, w_000_8806, w_000_8807, w_000_8808, w_000_8809, w_000_8810, w_000_8811, w_000_8812, w_000_8813, w_000_8814, w_000_8815, w_000_8816, w_000_8817, w_000_8818, w_000_8819, w_000_8820, w_000_8821, w_000_8822, w_000_8823, w_000_8824, w_000_8825, w_000_8826, w_000_8827, w_000_8828, w_000_8829, w_000_8830, w_000_8831, w_000_8832, w_000_8833, w_000_8834, w_000_8835, w_000_8836, w_000_8837, w_000_8838, w_000_8839, w_000_8840, w_000_8841, w_000_8842, w_000_8843, w_000_8844, w_000_8845, w_000_8846, w_000_8848, w_000_8849, w_000_8850, w_000_8851, w_000_8852, w_000_8853, w_000_8854, w_000_8855, w_000_8856, w_000_8857, w_000_8858, w_000_8859, w_000_8860, w_000_8861, w_000_8862, w_000_8863, w_000_8864, w_000_8865, w_000_8866, w_000_8867, w_000_8868, w_000_8869, w_000_8870, w_000_8871, w_000_8872, w_000_8873, w_000_8874, w_000_8875, w_000_8876, w_000_8877, w_000_8878, w_000_8879, w_000_8880, w_000_8881, w_000_8882, w_000_8883, w_000_8884, w_000_8885, w_000_8886, w_000_8887, w_000_8888, w_000_8889, w_000_8891, w_000_8892, w_000_8893, w_000_8894, w_000_8895, w_000_8896, w_000_8897, w_000_8898, w_000_8899, w_000_8900, w_000_8901, w_000_8902, w_000_8903, w_000_8904, w_000_8905, w_000_8906, w_000_8907, w_000_8908, w_000_8909, w_000_8910, w_000_8911, w_000_8912, w_000_8913, w_000_8914, w_000_8916, w_000_8917, w_000_8918, w_000_8919, w_000_8920, w_000_8921, w_000_8922, w_000_8923, w_000_8924, w_000_8925, w_000_8926, w_000_8927, w_000_8928, w_000_8929, w_000_8930, w_000_8931, w_000_8932, w_000_8933, w_000_8934, w_000_8935, w_000_8936, w_000_8937, w_000_8938, w_000_8939, w_000_8940, w_000_8941, w_000_8942, w_000_8943, w_000_8944, w_000_8945, w_000_8946, w_000_8947, w_000_8948, w_000_8949, w_000_8950, w_000_8951, w_000_8952, w_000_8953, w_000_8954, w_000_8955, w_000_8956, w_000_8957, w_000_8958, w_000_8959, w_000_8960, w_000_8961, w_000_8962, w_000_8963, w_000_8964, w_000_8965, w_000_8966, w_000_8967, w_000_8968, w_000_8969, w_000_8970, w_000_8971, w_000_8972, w_000_8973, w_000_8974, w_000_8975, w_000_8976, w_000_8977, w_000_8978, w_000_8979, w_000_8980, w_000_8981, w_000_8982, w_000_8983, w_000_8984, w_000_8985, w_000_8986, w_000_8987, w_000_8988, w_000_8989, w_000_8990, w_000_8991, w_000_8992, w_000_8993, w_000_8994, w_000_8995, w_000_8996, w_000_8997, w_000_8998, w_000_8999, w_000_9000, w_000_9001, w_000_9002, w_000_9003, w_000_9004, w_000_9005, w_000_9006, w_000_9007, w_000_9008, w_000_9009, w_000_9010, w_000_9011, w_000_9012, w_000_9013, w_000_9014, w_000_9015, w_000_9016, w_000_9017, w_000_9018, w_000_9019, w_000_9020, w_000_9021, w_000_9022, w_000_9023, w_000_9024, w_000_9025, w_000_9026, w_000_9027, w_000_9028, w_000_9029, w_000_9030, w_000_9031, w_000_9032, w_000_9033, w_000_9034, w_000_9035, w_000_9036, w_000_9037, w_000_9038, w_000_9039, w_000_9040, w_000_9041, w_000_9042, w_000_9043, w_000_9044, w_000_9045, w_000_9046, w_000_9047, w_000_9048, w_000_9049, w_000_9050, w_000_9051, w_000_9052, w_000_9053, w_000_9054, w_000_9055, w_000_9056, w_000_9057, w_000_9058, w_000_9059, w_000_9060, w_000_9061, w_000_9062, w_000_9063, w_000_9064, w_000_9065, w_000_9066, w_000_9067, w_000_9068, w_000_9069, w_000_9070, w_000_9071, w_000_9072, w_000_9073, w_000_9074, w_000_9075, w_000_9076, w_000_9077, w_000_9078, w_000_9079, w_000_9080, w_000_9081, w_000_9082, w_000_9083, w_000_9084, w_000_9085, w_000_9086, w_000_9087, w_000_9088, w_000_9089, w_000_9090, w_000_9091, w_000_9092, w_000_9093, w_000_9094, w_000_9095, w_000_9096, w_000_9097, w_000_9098, w_000_9099, w_000_9100, w_000_9101, w_000_9102, w_000_9103, w_000_9104, w_000_9105, w_000_9106, w_000_9107, w_000_9108, w_000_9109, w_000_9110, w_000_9111, w_000_9112, w_000_9113, w_000_9114, w_000_9115, w_000_9116, w_000_9117, w_000_9118, w_000_9119, w_000_9120, w_000_9121, w_000_9122, w_000_9123, w_000_9124, w_000_9125, w_000_9126, w_000_9127, w_000_9128, w_000_9129, w_000_9130, w_000_9131, w_000_9132, w_000_9133, w_000_9134, w_000_9135, w_000_9136, w_000_9137, w_000_9138, w_000_9139, w_000_9140, w_000_9141, w_000_9142, w_000_9143, w_000_9144, w_000_9145, w_000_9146, w_000_9147, w_000_9148, w_000_9149, w_000_9150, w_000_9151, w_000_9152, w_000_9153, w_000_9154, w_000_9155, w_000_9156, w_000_9157, w_000_9158, w_000_9159, w_000_9160, w_000_9161, w_000_9162, w_000_9163, w_000_9164, w_000_9165, w_000_9166, w_000_9167, w_000_9168, w_000_9169, w_000_9170, w_000_9171, w_000_9172, w_000_9173, w_000_9174, w_000_9175, w_000_9176, w_000_9177, w_000_9178, w_000_9179, w_000_9180, w_000_9181, w_000_9182, w_000_9183, w_000_9184, w_000_9185, w_000_9186, w_000_9187, w_000_9188, w_000_9189, w_000_9190, w_000_9191, w_000_9192, w_000_9193, w_000_9194, w_000_9195, w_000_9196, w_000_9197, w_000_9198, w_000_9199, w_000_9200, w_000_9201, w_000_9202, w_000_9203, w_000_9204, w_000_9205, w_000_9206, w_000_9207, w_000_9208, w_000_9209, w_000_9210, w_000_9211, w_000_9212, w_000_9213, w_000_9214, w_000_9215, w_000_9216, w_000_9217, w_000_9218, w_000_9219, w_000_9220, w_000_9221, w_000_9222, w_000_9223, w_000_9224, w_000_9225, w_000_9226, w_000_9227, w_000_9228, w_000_9229, w_000_9230, w_000_9231, w_000_9232, w_000_9233, w_000_9234, w_000_9235, w_000_9236, w_000_9237, w_000_9238, w_000_9239, w_000_9240, w_000_9241, w_000_9242, w_000_9243, w_000_9244, w_000_9245, w_000_9246, w_000_9247, w_000_9248, w_000_9249, w_000_9250, w_000_9251, w_000_9252, w_000_9253, w_000_9254, w_000_9255, w_000_9256, w_000_9257, w_000_9258, w_000_9259, w_000_9260, w_000_9261, w_000_9262, w_000_9263, w_000_9264, w_000_9265, w_000_9266, w_000_9267, w_000_9268, w_000_9269, w_000_9270, w_000_9271, w_000_9272, w_000_9273, w_000_9274, w_000_9275, w_000_9276, w_000_9277, w_000_9278, w_000_9279, w_000_9280, w_000_9281, w_000_9282, w_000_9283, w_000_9284, w_000_9285, w_000_9286, w_000_9287, w_000_9288, w_000_9289, w_000_9290, w_000_9291, w_000_9292, w_000_9293, w_000_9294, w_000_9295, w_000_9296, w_000_9297, w_000_9298, w_000_9299, w_000_9300, w_000_9301, w_000_9302, w_000_9303, w_000_9304, w_000_9305, w_000_9306, w_000_9307, w_000_9308, w_000_9309, w_000_9310, w_000_9311, w_000_9312, w_000_9313, w_000_9314, w_000_9315, w_000_9316, w_000_9317, w_000_9318, w_000_9319, w_000_9320, w_000_9321, w_000_9322, w_000_9323, w_000_9324, w_000_9325, w_000_9326, w_000_9327, w_000_9328, w_000_9329, w_000_9330, w_000_9331, w_000_9332, w_000_9333, w_000_9334, w_000_9335, w_000_9336, w_000_9337, w_000_9338, w_000_9339, w_000_9340, w_000_9341, w_000_9342, w_000_9343, w_000_9344, w_000_9345, w_000_9346, w_000_9347, w_000_9348, w_000_9349, w_000_9350, w_000_9351, w_000_9352, w_000_9353, w_000_9354, w_000_9355, w_000_9356, w_000_9357, w_000_9358, w_000_9359, w_000_9360, w_000_9361, w_000_9362, w_000_9363, w_000_9364, w_000_9365, w_000_9366, w_000_9367, w_000_9368, w_000_9369, w_000_9370, w_000_9371, w_000_9372, w_000_9373, w_000_9374, w_000_9375, w_000_9376, w_000_9377, w_000_9378, w_000_9379, w_000_9380, w_000_9381, w_000_9382, w_000_9383, w_000_9384, w_000_9385, w_000_9386, w_000_9387, w_000_9388, w_000_9389, w_000_9390, w_000_9391, w_000_9392, w_000_9393, w_000_9394, w_000_9395, w_000_9396, w_000_9397, w_000_9398, w_000_9399, w_000_9400, w_000_9401, w_000_9402, w_000_9403, w_000_9404, w_000_9405, w_000_9406, w_000_9407, w_000_9408, w_000_9409, w_000_9410, w_000_9411, w_000_9412, w_000_9413, w_000_9414, w_000_9415, w_000_9416, w_000_9417, w_000_9418, w_000_9419, w_000_9420, w_000_9421, w_000_9422, w_000_9423, w_000_9424, w_000_9425, w_000_9426, w_000_9427, w_000_9428, w_000_9429, w_000_9430, w_000_9431, w_000_9432, w_000_9433, w_000_9434, w_000_9435, w_000_9436, w_000_9437, w_000_9438, w_000_9439, w_000_9440, w_000_9441, w_000_9442, w_000_9443, w_000_9444, w_000_9445, w_000_9446, w_000_9447, w_000_9448, w_000_9449, w_000_9450, w_000_9451, w_000_9452, w_000_9453, w_000_9454, w_000_9455, w_000_9456, w_000_9457, w_000_9458, w_000_9459, w_000_9460, w_000_9461, w_000_9462, w_000_9463, w_000_9464, w_000_9465, w_000_9466, w_000_9467, w_000_9468, w_000_9469, w_000_9470, w_000_9471, w_000_9472, w_000_9473, w_000_9474, w_000_9475, w_000_9476, w_000_9477, w_000_9478, w_000_9479, w_000_9480, w_000_9481, w_000_9482, w_000_9483, w_000_9484, w_000_9485, w_000_9486, w_000_9487, w_000_9488, w_000_9489, w_000_9490, w_000_9491, w_000_9492, w_000_9493, w_000_9494, w_000_9495, w_000_9496, w_000_9497, w_000_9498, w_000_9499, w_000_9500, w_000_9501, w_000_9502, w_000_9504, w_000_9505, w_000_9506, w_000_9507, w_000_9508, w_000_9509, w_000_9510, w_000_9511, w_000_9512, w_000_9513, w_000_9514, w_000_9515, w_000_9516, w_000_9517, w_000_9518, w_000_9519, w_000_9520, w_000_9521, w_000_9522, w_000_9523, w_000_9524, w_000_9525, w_000_9526, w_000_9527, w_000_9528, w_000_9529, w_000_9530, w_000_9531, w_000_9532, w_000_9533, w_000_9534, w_000_9535, w_000_9536, w_000_9537, w_000_9538, w_000_9539, w_000_9540, w_000_9541, w_000_9542, w_000_9543, w_000_9544, w_000_9545, w_000_9547, w_000_9548, w_000_9549, w_000_9550, w_000_9551, w_000_9552, w_000_9554, w_000_9555, w_000_9556, w_000_9557, w_000_9558, w_000_9559, w_000_9560, w_000_9561, w_000_9563, w_000_9564, w_000_9565, w_000_9566, w_000_9567, w_000_9569, w_000_9570, w_000_9571, w_000_9572, w_000_9573, w_000_9574, w_000_9575, w_000_9576, w_000_9577, w_000_9578, w_000_9579, w_000_9580, w_000_9581, w_000_9582, w_000_9583, w_000_9584, w_000_9585, w_000_9586, w_000_9587, w_000_9588, w_000_9589, w_000_9590, w_000_9591, w_000_9592, w_000_9593, w_000_9594, w_000_9595, w_000_9596, w_000_9597, w_000_9598, w_000_9599, w_000_9600, w_000_9601, w_000_9602, w_000_9603, w_000_9604, w_000_9605, w_000_9606, w_000_9607, w_000_9608, w_000_9609, w_000_9610, w_000_9611, w_000_9612, w_000_9613, w_000_9614, w_000_9615, w_000_9616, w_000_9617, w_000_9618, w_000_9619, w_000_9620, w_000_9621, w_000_9622, w_000_9623, w_000_9624, w_000_9625, w_000_9626, w_000_9627, w_000_9628, w_000_9629, w_000_9630, w_000_9632, w_000_9633, w_000_9634, w_000_9635, w_000_9636, w_000_9637, w_000_9639, w_000_9640, w_000_9641, w_000_9642, w_000_9643, w_000_9644, w_000_9646, w_000_9647, w_000_9648, w_000_9649, w_000_9650, w_000_9651, w_000_9652, w_000_9653, w_000_9654, w_000_9655, w_000_9656, w_000_9657, w_000_9658, w_000_9659, w_000_9660, w_000_9661, w_000_9662, w_000_9663, w_000_9664, w_000_9666, w_000_9667, w_000_9668, w_000_9669, w_000_9670, w_000_9671, w_000_9672, w_000_9673, w_000_9674, w_000_9675, w_000_9676, w_000_9677, w_000_9678, w_000_9679, w_000_9682, w_000_9683, w_000_9684, w_000_9685, w_000_9686, w_000_9687, w_000_9688, w_000_9689, w_000_9690, w_000_9691, w_000_9692, w_000_9693, w_000_9694, w_000_9695, w_000_9696, w_000_9697, w_000_9698, w_000_9699, w_000_9701, w_000_9702, w_000_9704, w_000_9706, w_000_9708, w_000_9709, w_000_9710, w_000_9711, w_000_9713, w_000_9715, w_000_9716, w_000_9717, w_000_9719, w_000_9720, w_000_9721, w_000_9723, w_000_9725, w_000_9727, w_000_9728, w_000_9729, w_000_9730, w_000_9731, w_000_9732, w_000_9733, w_000_9734, w_000_9735, w_000_9736, w_000_9737, w_000_9738, w_000_9739, w_000_9740, w_000_9741, w_000_9742, w_000_9743, w_000_9744, w_000_9745, w_000_9747, w_000_9748, w_000_9749, w_000_9750, w_000_9752, w_000_9753, w_000_9754, w_000_9755, w_000_9756, w_000_9757, w_000_9758, w_000_9759, w_000_9760, w_000_9761, w_000_9765, w_000_9766, w_000_9767, w_000_9769, w_000_9770, w_000_9771, w_000_9772, w_000_9774, w_000_9776, w_000_9777, w_000_9778, w_000_9779, w_000_9780, w_000_9781, w_000_9782, w_000_9783, w_000_9785, w_000_9786, w_000_9788, w_000_9789, w_000_9790, w_000_9791, w_000_9792, w_000_9793, w_000_9794, w_000_9795, w_000_9796, w_000_9797, w_000_9798, w_000_9799, w_000_9800, w_000_9801, w_000_9802, w_000_9803, w_000_9804, w_000_9805, w_000_9806, w_000_9807, w_000_9808, w_000_9809, w_000_9810, w_000_9811, w_000_9812, w_000_9813, w_000_9814, w_000_9815, w_000_9816, w_000_9817, w_000_9819, w_000_9820, w_000_9821, w_000_9822, w_000_9823, w_000_9824, w_000_9825, w_000_9826, w_000_9827, w_000_9828, w_000_9829, w_000_9830, w_000_9831, w_000_9832, w_000_9833, w_000_9834, w_000_9835, w_000_9837, w_000_9838, w_000_9841, w_000_9842, w_000_9843, w_000_9844, w_000_9846, w_000_9847, w_000_9848, w_000_9849, w_000_9851, w_000_9853, w_000_9854, w_000_9855, w_000_9856, w_000_9857, w_000_9858, w_000_9859, w_000_9860, w_000_9861, w_000_9862, w_000_9864, w_000_9865, w_000_9866, w_000_9867, w_000_9871, w_000_9872, w_000_9874, w_000_9875, w_000_9877, w_000_9878, w_000_9879, w_000_9880, w_000_9882, w_000_9884, w_000_9887, w_000_9889, w_000_9890, w_000_9892, w_000_9893, w_000_9894, w_000_9895, w_000_9896, w_000_9897, w_000_9898, w_000_9899, w_000_9900, w_000_9902, w_000_9904, w_000_9905, w_000_9907, w_000_9908, w_000_9910, w_000_9914, w_000_9920, w_000_9922, w_000_9925, w_000_9926, w_000_9929, w_000_9930, w_000_9934, w_000_9936, w_000_9937, w_000_9938, w_000_9941, w_000_9949, w_000_9951, w_000_9958, w_000_9970, w_000_9978, w_000_9985, w_000_9996, w_10000_000, w_10000_001, w_10000_002, w_10000_003, w_10000_004, w_10000_005, w_10000_006, w_10000_007, w_10000_008, w_10000_009, w_10000_010, w_10000_011, w_10000_012, w_10000_013, w_10000_014, w_10000_015, w_10000_016, w_10000_017, w_10000_018, w_10000_019, w_10000_020, w_10000_021, w_10000_022, w_10000_023, w_10000_024, w_10000_025, w_10000_026, w_10000_027, w_10000_028, w_10000_029, w_10000_030, w_10000_031, w_10000_032, w_10000_033, w_10000_034, w_10000_035, w_10000_036, w_10000_037, w_10000_038, w_10000_039, w_10000_040, w_10000_041, w_10000_042, w_10000_043, w_10000_044, w_10000_045, w_10000_046, w_10000_047, w_10000_048, w_10000_049, w_10000_050, w_10000_051, w_10000_052, w_10000_053, w_10000_054, w_10000_055, w_10000_056, w_10000_057, w_10000_058, w_10000_059, w_10000_060, w_10000_061, w_10000_062, w_10000_063, w_10000_064, w_10000_065, w_10000_066, w_10000_067, w_10000_068, w_10000_069, w_10000_070, w_10000_071, w_10000_072, w_10000_073, w_10000_074, w_10000_075, w_10000_076, w_10000_077, w_10000_078, w_10000_079, w_10000_080, w_10000_081, w_10000_082, w_10000_083, w_10000_084, w_10000_085, w_10000_086, w_10000_087, w_10000_088, w_10000_089, w_10000_090, w_10000_091, w_10000_092, w_10000_093, w_10000_094, w_10000_095, w_10000_096, w_10000_097, w_10000_098, w_10000_099, w_10000_100, w_10000_101, w_10000_102, w_10000_103, w_10000_104, w_10000_105, w_10000_106, w_10000_107, w_10000_108, w_10000_109, w_10000_110, w_10000_111, w_10000_112, w_10000_113, w_10000_114, w_10000_115, w_10000_116, w_10000_117, w_10000_118, w_10000_119, w_10000_120, w_10000_121, w_10000_122, w_10000_123, w_10000_124, w_10000_125, w_10000_126, w_10000_127, w_10000_128, w_10000_129, w_10000_130, w_10000_131, w_10000_132, w_10000_133, w_10000_134, w_10000_135, w_10000_136, w_10000_137, w_10000_138, w_10000_139, w_10000_140, w_10000_141, w_10000_142, w_10000_143, w_10000_144, w_10000_145, w_10000_146, w_10000_147, w_10000_148, w_10000_149, w_10000_150, w_10000_151, w_10000_152, w_10000_153, w_10000_154, w_10000_155, w_10000_156, w_10000_157, w_10000_158, w_10000_159, w_10000_160, w_10000_161, w_10000_162, w_10000_163, w_10000_164, w_10000_165, w_10000_166, w_10000_167, w_10000_168, w_10000_169, w_10000_170, w_10000_171, w_10000_172, w_10000_173, w_10000_174, w_10000_175, w_10000_176, w_10000_177, w_10000_178, w_10000_179, w_10000_180, w_10000_181, w_10000_182, w_10000_183, w_10000_184, w_10000_185, w_10000_186, w_10000_187, w_10000_188, w_10000_189, w_10000_190, w_10000_191, w_10000_192, w_10000_193, w_10000_194, w_10000_195, w_10000_196, w_10000_197, w_10000_198, w_10000_199, w_10000_200, w_10000_201, w_10000_202, w_10000_203, w_10000_204, w_10000_205, w_10000_206, w_10000_207, w_10000_208, w_10000_209, w_10000_210, w_10000_211, w_10000_212, w_10000_213, w_10000_214, w_10000_215, w_10000_216, w_10000_217, w_10000_218, w_10000_219, w_10000_220, w_10000_221, w_10000_222, w_10000_223, w_10000_224, w_10000_225, w_10000_226, w_10000_227, w_10000_228, w_10000_229, w_10000_230, w_10000_231, w_10000_232, w_10000_233, w_10000_234, w_10000_235, w_10000_236, w_10000_237, w_10000_238, w_10000_239, w_10000_240, w_10000_241, w_10000_242, w_10000_243, w_10000_244, w_10000_245, w_10000_246, w_10000_247, w_10000_248, w_10000_249, w_10000_250, w_10000_251, w_10000_252, w_10000_253, w_10000_254, w_10000_255, w_10000_256, w_10000_257, w_10000_258, w_10000_259, w_10000_260, w_10000_261, w_10000_262, w_10000_263, w_10000_264, w_10000_265, w_10000_266, w_10000_267, w_10000_268, w_10000_269, w_10000_270, w_10000_271, w_10000_272, w_10000_273, w_10000_274, w_10000_275, w_10000_276, w_10000_277, w_10000_278, w_10000_279, w_10000_280, w_10000_281, w_10000_282, w_10000_283, w_10000_284, w_10000_285, w_10000_286, w_10000_287, w_10000_288, w_10000_289, w_10000_290, w_10000_291, w_10000_292, w_10000_293, w_10000_294, w_10000_295, w_10000_296, w_10000_297, w_10000_298, w_10000_299, w_10000_300, w_10000_301, w_10000_302, w_10000_303, w_10000_304, w_10000_305, w_10000_306, w_10000_307, w_10000_308, w_10000_309, w_10000_310, w_10000_311, w_10000_312, w_10000_313, w_10000_314, w_10000_315, w_10000_316, w_10000_317, w_10000_318, w_10000_319, w_10000_320, w_10000_321, w_10000_322, w_10000_323, w_10000_324, w_10000_325, w_10000_326, w_10000_327, w_10000_328, w_10000_329, w_10000_330, w_10000_331, w_10000_332, w_10000_333, w_10000_334, w_10000_335, w_10000_336, w_10000_337, w_10000_338, w_10000_339, w_10000_340, w_10000_341, w_10000_342, w_10000_343, w_10000_344, w_10000_345, w_10000_346, w_10000_347, w_10000_348, w_10000_349, w_10000_350, w_10000_351, w_10000_352, w_10000_353, w_10000_354, w_10000_355, w_10000_356, w_10000_357, w_10000_358, w_10000_359, w_10000_360, w_10000_361, w_10000_362, w_10000_363, w_10000_364, w_10000_365, w_10000_366, w_10000_367, w_10000_368, w_10000_369, w_10000_370, w_10000_371, w_10000_372, w_10000_373, w_10000_374, w_10000_375, w_10000_376, w_10000_377, w_10000_378, w_10000_379, w_10000_380, w_10000_381, w_10000_382, w_10000_383, w_10000_384, w_10000_385, w_10000_386, w_10000_387, w_10000_388, w_10000_389, w_10000_390, w_10000_391, w_10000_392, w_10000_393, w_10000_394, w_10000_395, w_10000_396, w_10000_397, w_10000_398, w_10000_399, w_10000_400, w_10000_401, w_10000_402, w_10000_403, w_10000_404, w_10000_405, w_10000_406, w_10000_407, w_10000_408, w_10000_409, w_10000_410, w_10000_411, w_10000_412, w_10000_413, w_10000_414, w_10000_415, w_10000_416, w_10000_417, w_10000_418, w_10000_419, w_10000_420, w_10000_421, w_10000_422, w_10000_423, w_10000_424, w_10000_425, w_10000_426, w_10000_427, w_10000_428, w_10000_429, w_10000_430, w_10000_431, w_10000_432, w_10000_433, w_10000_434, w_10000_435, w_10000_436, w_10000_437, w_10000_438, w_10000_439, w_10000_440, w_10000_441, w_10000_442, w_10000_443, w_10000_444, w_10000_445, w_10000_446, w_10000_447, w_10000_448, w_10000_449, w_10000_450, w_10000_451, w_10000_452, w_10000_453, w_10000_454, w_10000_455, w_10000_456, w_10000_457, w_10000_458, w_10000_459, w_10000_460, w_10000_461, w_10000_462, w_10000_463, w_10000_464, w_10000_465, w_10000_466, w_10000_467, w_10000_468, w_10000_469, w_10000_470, w_10000_471, w_10000_472, w_10000_473, w_10000_474, w_10000_475, w_10000_476, w_10000_477, w_10000_478, w_10000_479, w_10000_480, w_10000_481, w_10000_482, w_10000_483, w_10000_484, w_10000_485, w_10000_486, w_10000_487, w_10000_488, w_10000_489, w_10000_490, w_10000_491, w_10000_492, w_10000_493, w_10000_494, w_10000_495, w_10000_496, w_10000_497, w_10000_498, w_10000_499, w_10000_500, w_10000_501, w_10000_502, w_10000_503, w_10000_504, w_10000_505, w_10000_506, w_10000_507, w_10000_508, w_10000_509, w_10000_510, w_10000_511, w_10000_512, w_10000_513, w_10000_514, w_10000_515, w_10000_516, w_10000_517, w_10000_518, w_10000_519, w_10000_520, w_10000_521, w_10000_522, w_10000_523, w_10000_524, w_10000_525, w_10000_526, w_10000_527, w_10000_528, w_10000_529, w_10000_530, w_10000_531, w_10000_532, w_10000_533, w_10000_534, w_10000_535, w_10000_536, w_10000_537, w_10000_538, w_10000_539, w_10000_540, w_10000_541, w_10000_542, w_10000_543, w_10000_544, w_10000_545, w_10000_546, w_10000_547, w_10000_548, w_10000_549, w_10000_550, w_10000_551, w_10000_552, w_10000_553, w_10000_554, w_10000_555, w_10000_556, w_10000_557, w_10000_558, w_10000_559, w_10000_560, w_10000_561, w_10000_562, w_10000_563, w_10000_564, w_10000_565, w_10000_566, w_10000_567, w_10000_568, w_10000_569, w_10000_570, w_10000_571, w_10000_572, w_10000_573, w_10000_574, w_10000_575, w_10000_576, w_10000_577, w_10000_578, w_10000_579, w_10000_580, w_10000_581, w_10000_582, w_10000_583, w_10000_584, w_10000_585, w_10000_586, w_10000_587, w_10000_588, w_10000_589, w_10000_590, w_10000_591, w_10000_592, w_10000_593, w_10000_594, w_10000_595, w_10000_596, w_10000_597, w_10000_598, w_10000_599, w_10000_600, w_10000_601, w_10000_602, w_10000_603, w_10000_604, w_10000_605, w_10000_606, w_10000_607, w_10000_608, w_10000_609, w_10000_610, w_10000_611, w_10000_612, w_10000_613, w_10000_614, w_10000_615, w_10000_616, w_10000_617, w_10000_618, w_10000_619, w_10000_620, w_10000_621, w_10000_622, w_10000_623, w_10000_624, w_10000_625, w_10000_626, w_10000_627, w_10000_628, w_10000_629, w_10000_630, w_10000_631, w_10000_632, w_10000_633, w_10000_634, w_10000_635, w_10000_636, w_10000_637, w_10000_638, w_10000_639, w_10000_640, w_10000_641, w_10000_642, w_10000_643, w_10000_644, w_10000_645, w_10000_646, w_10000_647, w_10000_648, w_10000_649, w_10000_650, w_10000_651, w_10000_652, w_10000_653, w_10000_654, w_10000_655, w_10000_656, w_10000_657, w_10000_658, w_10000_659, w_10000_660, w_10000_661, w_10000_662, w_10000_663, w_10000_664, w_10000_665, w_10000_666, w_10000_667, w_10000_668, w_10000_669, w_10000_670, w_10000_671, w_10000_672, w_10000_673, w_10000_674, w_10000_675, w_10000_676, w_10000_677, w_10000_678, w_10000_679, w_10000_680, w_10000_681, w_10000_682, w_10000_683, w_10000_684, w_10000_685, w_10000_686, w_10000_687, w_10000_688, w_10000_689, w_10000_690, w_10000_691, w_10000_692, w_10000_693, w_10000_694, w_10000_695, w_10000_696, w_10000_697, w_10000_698, w_10000_699, w_10000_700, w_10000_701, w_10000_702, w_10000_703, w_10000_704, w_10000_705, w_10000_706, w_10000_707, w_10000_708, w_10000_709, w_10000_710, w_10000_711, w_10000_712, w_10000_713, w_10000_714, w_10000_715, w_10000_716, w_10000_717, w_10000_718, w_10000_719, w_10000_720, w_10000_721, w_10000_722, w_10000_723, w_10000_724, w_10000_725, w_10000_726, w_10000_727, w_10000_728, w_10000_729, w_10000_730, w_10000_731, w_10000_732, w_10000_733, w_10000_734, w_10000_735, w_10000_736, w_10000_737, w_10000_738, w_10000_739, w_10000_740, w_10000_741, w_10000_742, w_10000_743, w_10000_744, w_10000_745, w_10000_746, w_10000_747, w_10000_748, w_10000_749, w_10000_750, w_10000_751, w_10000_752, w_10000_753, w_10000_754, w_10000_755, w_10000_756, w_10000_757, w_10000_758, w_10000_759, w_10000_760, w_10000_761, w_10000_762, w_10000_763, w_10000_764, w_10000_765, w_10000_766, w_10000_767, w_10000_768, w_10000_769, w_10000_770, w_10000_771, w_10000_772, w_10000_773, w_10000_774, w_10000_775, w_10000_776, w_10000_777, w_10000_778, w_10000_779, w_10000_780, w_10000_781, w_10000_782, w_10000_783, w_10000_784, w_10000_785, w_10000_786, w_10000_787, w_10000_788, w_10000_789, w_10000_790, w_10000_791, w_10000_792, w_10000_793, w_10000_794, w_10000_795, w_10000_796, w_10000_797, w_10000_798, w_10000_799, w_10000_800, w_10000_801, w_10000_802, w_10000_803, w_10000_804, w_10000_805, w_10000_806, w_10000_807, w_10000_808, w_10000_809, w_10000_810, w_10000_811, w_10000_812, w_10000_813, w_10000_814, w_10000_815, w_10000_816, w_10000_817, w_10000_818, w_10000_819, w_10000_820, w_10000_821, w_10000_822, w_10000_823, w_10000_824, w_10000_825, w_10000_826, w_10000_827, w_10000_828, w_10000_829, w_10000_830, w_10000_831, w_10000_832, w_10000_833, w_10000_834, w_10000_835, w_10000_836, w_10000_837, w_10000_838, w_10000_839, w_10000_840, w_10000_841, w_10000_842, w_10000_843, w_10000_844, w_10000_845, w_10000_846, w_10000_847, w_10000_848, w_10000_849, w_10000_850, w_10000_851, w_10000_852, w_10000_853, w_10000_854, w_10000_855, w_10000_856, w_10000_857, w_10000_858, w_10000_859, w_10000_860, w_10000_861, w_10000_862, w_10000_863, w_10000_864, w_10000_865, w_10000_866, w_10000_867, w_10000_868, w_10000_869, w_10000_870, w_10000_871, w_10000_872, w_10000_873, w_10000_874, w_10000_875, w_10000_876, w_10000_877, w_10000_878, w_10000_879, w_10000_880, w_10000_881, w_10000_882, w_10000_883, w_10000_884, w_10000_885, w_10000_886, w_10000_887, w_10000_888, w_10000_889, w_10000_890, w_10000_891, w_10000_892, w_10000_893, w_10000_894, w_10000_895, w_10000_896, w_10000_897, w_10000_898, w_10000_899, w_10000_900, w_10000_901, w_10000_902, w_10000_903, w_10000_904, w_10000_905, w_10000_906, w_10000_907, w_10000_908, w_10000_909, w_10000_910, w_10000_911, w_10000_912, w_10000_913, w_10000_914, w_10000_915, w_10000_916, w_10000_917, w_10000_918, w_10000_919, w_10000_920, w_10000_921, w_10000_922, w_10000_923, w_10000_924, w_10000_925, w_10000_926, w_10000_927, w_10000_928, w_10000_929, w_10000_930, w_10000_931, w_10000_932, w_10000_933, w_10000_934, w_10000_935, w_10000_936, w_10000_937, w_10000_938, w_10000_939, w_10000_940, w_10000_941, w_10000_942, w_10000_943, w_10000_944, w_10000_945, w_10000_946, w_10000_947, w_10000_948, w_10000_949, w_10000_950, w_10000_951, w_10000_952, w_10000_953, w_10000_954, w_10000_955, w_10000_956, w_10000_957, w_10000_958, w_10000_959, w_10000_960, w_10000_961, w_10000_962, w_10000_963, w_10000_964, w_10000_965, w_10000_966, w_10000_967, w_10000_968, w_10000_969, w_10000_970, w_10000_971, w_10000_972, w_10000_973, w_10000_974, w_10000_975, w_10000_976, w_10000_977, w_10000_978, w_10000_979, w_10000_980, w_10000_981, w_10000_982, w_10000_983, w_10000_984, w_10000_985, w_10000_986, w_10000_987, w_10000_988, w_10000_989, w_10000_990, w_10000_991, w_10000_992, w_10000_993, w_10000_994, w_10000_995, w_10000_996, w_10000_997, w_10000_998, w_10000_999, w_10000_1000, w_10000_1001, w_10000_1002, w_10000_1003, w_10000_1004, w_10000_1005, w_10000_1006, w_10000_1007, w_10000_1008, w_10000_1009, w_10000_1010, w_10000_1011, w_10000_1012, w_10000_1013, w_10000_1014, w_10000_1015, w_10000_1016, w_10000_1017, w_10000_1018, w_10000_1019, w_10000_1020, w_10000_1021, w_10000_1022, w_10000_1023, w_10000_1024, w_10000_1025, w_10000_1026, w_10000_1027, w_10000_1028, w_10000_1029, w_10000_1030, w_10000_1031, w_10000_1032, w_10000_1033, w_10000_1034, w_10000_1035, w_10000_1036, w_10000_1037, w_10000_1038, w_10000_1039, w_10000_1040, w_10000_1041, w_10000_1042, w_10000_1043, w_10000_1044, w_10000_1045, w_10000_1046, w_10000_1047, w_10000_1048, w_10000_1049, w_10000_1050, w_10000_1051, w_10000_1052, w_10000_1053, w_10000_1054, w_10000_1055, w_10000_1056, w_10000_1057, w_10000_1058, w_10000_1059, w_10000_1060, w_10000_1061, w_10000_1062, w_10000_1063, w_10000_1064, w_10000_1065, w_10000_1066, w_10000_1067, w_10000_1068, w_10000_1069, w_10000_1070, w_10000_1071, w_10000_1072, w_10000_1073, w_10000_1074, w_10000_1075, w_10000_1076, w_10000_1077, w_10000_1078, w_10000_1079, w_10000_1080, w_10000_1081, w_10000_1082, w_10000_1083, w_10000_1084, w_10000_1085, w_10000_1086, w_10000_1087, w_10000_1088, w_10000_1089, w_10000_1090, w_10000_1091, w_10000_1092, w_10000_1093, w_10000_1094, w_10000_1095, w_10000_1096, w_10000_1097, w_10000_1098, w_10000_1099, w_10000_1100, w_10000_1101, w_10000_1102, w_10000_1103, w_10000_1104, w_10000_1105, w_10000_1106, w_10000_1107, w_10000_1108, w_10000_1109, w_10000_1110, w_10000_1111, w_10000_1112, w_10000_1113, w_10000_1114, w_10000_1115, w_10000_1116, w_10000_1117, w_10000_1118, w_10000_1119, w_10000_1120, w_10000_1121, w_10000_1122, w_10000_1123, w_10000_1124, w_10000_1125, w_10000_1126, w_10000_1127, w_10000_1128, w_10000_1129, w_10000_1130, w_10000_1131, w_10000_1132, w_10000_1133, w_10000_1134, w_10000_1135, w_10000_1136, w_10000_1137, w_10000_1138, w_10000_1139, w_10000_1140, w_10000_1141, w_10000_1142, w_10000_1143, w_10000_1144, w_10000_1145, w_10000_1146, w_10000_1147, w_10000_1148, w_10000_1149, w_10000_1150, w_10000_1151, w_10000_1152, w_10000_1153, w_10000_1154, w_10000_1155, w_10000_1156, w_10000_1157, w_10000_1158, w_10000_1159, w_10000_1160, w_10000_1161, w_10000_1162, w_10000_1163, w_10000_1164, w_10000_1165, w_10000_1166, w_10000_1167, w_10000_1168, w_10000_1169, w_10000_1170, w_10000_1171, w_10000_1172, w_10000_1173, w_10000_1174, w_10000_1175, w_10000_1176, w_10000_1177, w_10000_1178, w_10000_1179, w_10000_1180, w_10000_1181, w_10000_1182, w_10000_1183, w_10000_1184, w_10000_1185, w_10000_1186, w_10000_1187, w_10000_1188, w_10000_1189, w_10000_1190, w_10000_1191, w_10000_1192, w_10000_1193, w_10000_1194, w_10000_1195, w_10000_1196, w_10000_1197, w_10000_1198, w_10000_1199, w_10000_1200, w_10000_1201, w_10000_1202, w_10000_1203, w_10000_1204, w_10000_1205, w_10000_1206, w_10000_1207, w_10000_1208, w_10000_1209, w_10000_1210, w_10000_1211, w_10000_1212, w_10000_1213, w_10000_1214, w_10000_1215, w_10000_1216, w_10000_1217, w_10000_1218, w_10000_1219, w_10000_1220, w_10000_1221, w_10000_1222, w_10000_1223, w_10000_1224, w_10000_1225, w_10000_1226, w_10000_1227, w_10000_1228, w_10000_1229, w_10000_1230, w_10000_1231, w_10000_1232, w_10000_1233, w_10000_1234, w_10000_1235, w_10000_1236, w_10000_1237, w_10000_1238, w_10000_1239, w_10000_1240, w_10000_1241, w_10000_1242, w_10000_1243, w_10000_1244, w_10000_1245, w_10000_1246, w_10000_1247, w_10000_1248, w_10000_1249, w_10000_1250, w_10000_1251, w_10000_1252, w_10000_1253, w_10000_1254, w_10000_1255, w_10000_1256, w_10000_1257, w_10000_1258, w_10000_1259, w_10000_1260, w_10000_1261, w_10000_1262, w_10000_1263, w_10000_1264, w_10000_1265, w_10000_1266, w_10000_1267, w_10000_1268, w_10000_1269, w_10000_1270, w_10000_1271, w_10000_1272, w_10000_1273, w_10000_1274, w_10000_1275, w_10000_1276, w_10000_1277, w_10000_1278, w_10000_1279, w_10000_1280, w_10000_1281, w_10000_1282, w_10000_1283, w_10000_1284, w_10000_1285, w_10000_1286, w_10000_1287, w_10000_1288, w_10000_1289, w_10000_1290, w_10000_1291, w_10000_1292, w_10000_1293, w_10000_1294, w_10000_1295, w_10000_1296, w_10000_1297, w_10000_1298, w_10000_1299, w_10000_1300, w_10000_1301, w_10000_1302, w_10000_1303, w_10000_1304, w_10000_1305, w_10000_1306, w_10000_1307, w_10000_1308, w_10000_1309, w_10000_1310, w_10000_1311, w_10000_1312, w_10000_1313, w_10000_1314, w_10000_1315, w_10000_1316, w_10000_1317, w_10000_1318, w_10000_1319, w_10000_1320, w_10000_1321, w_10000_1322, w_10000_1323, w_10000_1324, w_10000_1325, w_10000_1326, w_10000_1327, w_10000_1328, w_10000_1329, w_10000_1330, w_10000_1331, w_10000_1332, w_10000_1333, w_10000_1334, w_10000_1335, w_10000_1336, w_10000_1337, w_10000_1338, w_10000_1339, w_10000_1340, w_10000_1341, w_10000_1342, w_10000_1343, w_10000_1344, w_10000_1345, w_10000_1346, w_10000_1347, w_10000_1348, w_10000_1349, w_10000_1350, w_10000_1351, w_10000_1352, w_10000_1353, w_10000_1354, w_10000_1355, w_10000_1356, w_10000_1357, w_10000_1358, w_10000_1359, w_10000_1360, w_10000_1361, w_10000_1362, w_10000_1363, w_10000_1364, w_10000_1365, w_10000_1366, w_10000_1367, w_10000_1368, w_10000_1369, w_10000_1370, w_10000_1371, w_10000_1372, w_10000_1373, w_10000_1374, w_10000_1375, w_10000_1376, w_10000_1377, w_10000_1378, w_10000_1379, w_10000_1380, w_10000_1381, w_10000_1382, w_10000_1383, w_10000_1384, w_10000_1385, w_10000_1386, w_10000_1387, w_10000_1388, w_10000_1389, w_10000_1390, w_10000_1391, w_10000_1392, w_10000_1393, w_10000_1394, w_10000_1395, w_10000_1396, w_10000_1397, w_10000_1398, w_10000_1399, w_10000_1400, w_10000_1401, w_10000_1402, w_10000_1403, w_10000_1404, w_10000_1405, w_10000_1406, w_10000_1407, w_10000_1408, w_10000_1409, w_10000_1410, w_10000_1411, w_10000_1412, w_10000_1413, w_10000_1414, w_10000_1415, w_10000_1416, w_10000_1417, w_10000_1418, w_10000_1419, w_10000_1420, w_10000_1421, w_10000_1422, w_10000_1423, w_10000_1424, w_10000_1425, w_10000_1426, w_10000_1427, w_10000_1428, w_10000_1429, w_10000_1430, w_10000_1431, w_10000_1432, w_10000_1433, w_10000_1434, w_10000_1435, w_10000_1436, w_10000_1437, w_10000_1438, w_10000_1439, w_10000_1440, w_10000_1441, w_10000_1442, w_10000_1443, w_10000_1444, w_10000_1445, w_10000_1446, w_10000_1447, w_10000_1448, w_10000_1449, w_10000_1450, w_10000_1451, w_10000_1452, w_10000_1453, w_10000_1454, w_10000_1455, w_10000_1456, w_10000_1457, w_10000_1458, w_10000_1459, w_10000_1460, w_10000_1461, w_10000_1462, w_10000_1463, w_10000_1464, w_10000_1465, w_10000_1466, w_10000_1467, w_10000_1468, w_10000_1469, w_10000_1470, w_10000_1471, w_10000_1472, w_10000_1473, w_10000_1474, w_10000_1475, w_10000_1476, w_10000_1477, w_10000_1478, w_10000_1479, w_10000_1480, w_10000_1481, w_10000_1482, w_10000_1483, w_10000_1484, w_10000_1485, w_10000_1486, w_10000_1487, w_10000_1488, w_10000_1489, w_10000_1490, w_10000_1491, w_10000_1492, w_10000_1493, w_10000_1494, w_10000_1495, w_10000_1496, w_10000_1497, w_10000_1498, w_10000_1499, w_10000_1500, w_10000_1501, w_10000_1502, w_10000_1503, w_10000_1504, w_10000_1505, w_10000_1506, w_10000_1507, w_10000_1508, w_10000_1509, w_10000_1510, w_10000_1511, w_10000_1512, w_10000_1513, w_10000_1514, w_10000_1515, w_10000_1516, w_10000_1517, w_10000_1518, w_10000_1519, w_10000_1520, w_10000_1521, w_10000_1522, w_10000_1523, w_10000_1524, w_10000_1525, w_10000_1526, w_10000_1527, w_10000_1528, w_10000_1529, w_10000_1530, w_10000_1531, w_10000_1532, w_10000_1533, w_10000_1534, w_10000_1535, w_10000_1536, w_10000_1537, w_10000_1538, w_10000_1539, w_10000_1540, w_10000_1541, w_10000_1542, w_10000_1543, w_10000_1544, w_10000_1545, w_10000_1546, w_10000_1547, w_10000_1548, w_10000_1549, w_10000_1550, w_10000_1551, w_10000_1552, w_10000_1553, w_10000_1554, w_10000_1555, w_10000_1556, w_10000_1557, w_10000_1558, w_10000_1559, w_10000_1560, w_10000_1561, w_10000_1562, w_10000_1563, w_10000_1564, w_10000_1565, w_10000_1566, w_10000_1567, w_10000_1568, w_10000_1569, w_10000_1570, w_10000_1571, w_10000_1572, w_10000_1573, w_10000_1574, w_10000_1575, w_10000_1576, w_10000_1577, w_10000_1578, w_10000_1579, w_10000_1580, w_10000_1581, w_10000_1582, w_10000_1583, w_10000_1584, w_10000_1585, w_10000_1586, w_10000_1587, w_10000_1588, w_10000_1589, w_10000_1590, w_10000_1591, w_10000_1592, w_10000_1593, w_10000_1594, w_10000_1595, w_10000_1596, w_10000_1597, w_10000_1598, w_10000_1599, w_10000_1600, w_10000_1601, w_10000_1602, w_10000_1603, w_10000_1604, w_10000_1605, w_10000_1606, w_10000_1607, w_10000_1608, w_10000_1609, w_10000_1610, w_10000_1611, w_10000_1612, w_10000_1613, w_10000_1614, w_10000_1615, w_10000_1616, w_10000_1617, w_10000_1618, w_10000_1619, w_10000_1620, w_10000_1621, w_10000_1622, w_10000_1623, w_10000_1624, w_10000_1625, w_10000_1626, w_10000_1627, w_10000_1628, w_10000_1629, w_10000_1630, w_10000_1631, w_10000_1632, w_10000_1633, w_10000_1634, w_10000_1635, w_10000_1636, w_10000_1637, w_10000_1638, w_10000_1639, w_10000_1640, w_10000_1641, w_10000_1642, w_10000_1643, w_10000_1644, w_10000_1645, w_10000_1646, w_10000_1647, w_10000_1648, w_10000_1649, w_10000_1650, w_10000_1651, w_10000_1652, w_10000_1653, w_10000_1654, w_10000_1655, w_10000_1656, w_10000_1657, w_10000_1658, w_10000_1659, w_10000_1660, w_10000_1661, w_10000_1662, w_10000_1663, w_10000_1664, w_10000_1665, w_10000_1666, w_10000_1667, w_10000_1668, w_10000_1669, w_10000_1670, w_10000_1671, w_10000_1672, w_10000_1673, w_10000_1674, w_10000_1675, w_10000_1676, w_10000_1677, w_10000_1678, w_10000_1679, w_10000_1680, w_10000_1681, w_10000_1682, w_10000_1683, w_10000_1684, w_10000_1685, w_10000_1686, w_10000_1687, w_10000_1688, w_10000_1689, w_10000_1690, w_10000_1691, w_10000_1692, w_10000_1693, w_10000_1694, w_10000_1695, w_10000_1696, w_10000_1697, w_10000_1698, w_10000_1699, w_10000_1700, w_10000_1701, w_10000_1702, w_10000_1703, w_10000_1704, w_10000_1705, w_10000_1706, w_10000_1707, w_10000_1708, w_10000_1709, w_10000_1710, w_10000_1711, w_10000_1712, w_10000_1713, w_10000_1714, w_10000_1715, w_10000_1716, w_10000_1717, w_10000_1718, w_10000_1719, w_10000_1720, w_10000_1721, w_10000_1722, w_10000_1723, w_10000_1724, w_10000_1725, w_10000_1726, w_10000_1727, w_10000_1728, w_10000_1729, w_10000_1730, w_10000_1731, w_10000_1732, w_10000_1733, w_10000_1734, w_10000_1735, w_10000_1736, w_10000_1737, w_10000_1738, w_10000_1739, w_10000_1740, w_10000_1741, w_10000_1742, w_10000_1743, w_10000_1744, w_10000_1745, w_10000_1746, w_10000_1747, w_10000_1748, w_10000_1749, w_10000_1750, w_10000_1751, w_10000_1752, w_10000_1753, w_10000_1754, w_10000_1755, w_10000_1756, w_10000_1757, w_10000_1758, w_10000_1759, w_10000_1760, w_10000_1761, w_10000_1762, w_10000_1763, w_10000_1764, w_10000_1765, w_10000_1766, w_10000_1767, w_10000_1768, w_10000_1769, w_10000_1770, w_10000_1771, w_10000_1772, w_10000_1773, w_10000_1774, w_10000_1775, w_10000_1776, w_10000_1777, w_10000_1778, w_10000_1779, w_10000_1780, w_10000_1781, w_10000_1782, w_10000_1783, w_10000_1784, w_10000_1785, w_10000_1786, w_10000_1787, w_10000_1788, w_10000_1789, w_10000_1790, w_10000_1791, w_10000_1792, w_10000_1793, w_10000_1794, w_10000_1795, w_10000_1796, w_10000_1797, w_10000_1798, w_10000_1799, w_10000_1800, w_10000_1801, w_10000_1802, w_10000_1803, w_10000_1804, w_10000_1805, w_10000_1806, w_10000_1807, w_10000_1808, w_10000_1809, w_10000_1810, w_10000_1811, w_10000_1812, w_10000_1813, w_10000_1814, w_10000_1815, w_10000_1816, w_10000_1817, w_10000_1818, w_10000_1819, w_10000_1820, w_10000_1821, w_10000_1822, w_10000_1823, w_10000_1824, w_10000_1825, w_10000_1826, w_10000_1827, w_10000_1828, w_10000_1829, w_10000_1830, w_10000_1831, w_10000_1832, w_10000_1833, w_10000_1834, w_10000_1835, w_10000_1836, w_10000_1837, w_10000_1838, w_10000_1839, w_10000_1840, w_10000_1841, w_10000_1842, w_10000_1843, w_10000_1844, w_10000_1845, w_10000_1846, w_10000_1847, w_10000_1848, w_10000_1849, w_10000_1850, w_10000_1851, w_10000_1852, w_10000_1853, w_10000_1854, w_10000_1855, w_10000_1856, w_10000_1857, w_10000_1858, w_10000_1859, w_10000_1860, w_10000_1861, w_10000_1862, w_10000_1863, w_10000_1864, w_10000_1865, w_10000_1866, w_10000_1867, w_10000_1868, w_10000_1869, w_10000_1870, w_10000_1871, w_10000_1872, w_10000_1873, w_10000_1874, w_10000_1875, w_10000_1876, w_10000_1877, w_10000_1878, w_10000_1879, w_10000_1880, w_10000_1881, w_10000_1882, w_10000_1883, w_10000_1884, w_10000_1885, w_10000_1886, w_10000_1887, w_10000_1888, w_10000_1889, w_10000_1890, w_10000_1891, w_10000_1892, w_10000_1893, w_10000_1894, w_10000_1895, w_10000_1896, w_10000_1897, w_10000_1898, w_10000_1899, w_10000_1900, w_10000_1901, w_10000_1902, w_10000_1903, w_10000_1904, w_10000_1905, w_10000_1906, w_10000_1907, w_10000_1908, w_10000_1909, w_10000_1910, w_10000_1911, w_10000_1912, w_10000_1913, w_10000_1914, w_10000_1915, w_10000_1916, w_10000_1917, w_10000_1918, w_10000_1919, w_10000_1920, w_10000_1921, w_10000_1922, w_10000_1923, w_10000_1924, w_10000_1925, w_10000_1926, w_10000_1927, w_10000_1928, w_10000_1929, w_10000_1930, w_10000_1931, w_10000_1932, w_10000_1933, w_10000_1934, w_10000_1935, w_10000_1936, w_10000_1937, w_10000_1938, w_10000_1939, w_10000_1940, w_10000_1941, w_10000_1942, w_10000_1943, w_10000_1944, w_10000_1945, w_10000_1946, w_10000_1947, w_10000_1948, w_10000_1949, w_10000_1950, w_10000_1951, w_10000_1952, w_10000_1953, w_10000_1954, w_10000_1955, w_10000_1956, w_10000_1957, w_10000_1958, w_10000_1959, w_10000_1960, w_10000_1961, w_10000_1962, w_10000_1963, w_10000_1964, w_10000_1965, w_10000_1966, w_10000_1967, w_10000_1968, w_10000_1969, w_10000_1970, w_10000_1971, w_10000_1972, w_10000_1973, w_10000_1974, w_10000_1975, w_10000_1976, w_10000_1977, w_10000_1978, w_10000_1979, w_10000_1980, w_10000_1981, w_10000_1982, w_10000_1983, w_10000_1984, w_10000_1985, w_10000_1986, w_10000_1987, w_10000_1988, w_10000_1989, w_10000_1990, w_10000_1991, w_10000_1992, w_10000_1993, w_10000_1994, w_10000_1995, w_10000_1996, w_10000_1997, w_10000_1998, w_10000_1999, w_10000_2000, w_10000_2001, w_10000_2002, w_10000_2003, w_10000_2004, w_10000_2005, w_10000_2006, w_10000_2007, w_10000_2008, w_10000_2009, w_10000_2010, w_10000_2011, w_10000_2012, w_10000_2013, w_10000_2014, w_10000_2015, w_10000_2016, w_10000_2017, w_10000_2018, w_10000_2019, w_10000_2020, w_10000_2021, w_10000_2022, w_10000_2023, w_10000_2024, w_10000_2025, w_10000_2026, w_10000_2027, w_10000_2028, w_10000_2029, w_10000_2030, w_10000_2031, w_10000_2032, w_10000_2033, w_10000_2034, w_10000_2035, w_10000_2036, w_10000_2037, w_10000_2038, w_10000_2039, w_10000_2040, w_10000_2041, w_10000_2042, w_10000_2043, w_10000_2044, w_10000_2045, w_10000_2046, w_10000_2047, w_10000_2048, w_10000_2049, w_10000_2050, w_10000_2051, w_10000_2052, w_10000_2053, w_10000_2054, w_10000_2055, w_10000_2056, w_10000_2057, w_10000_2058, w_10000_2059, w_10000_2060, w_10000_2061, w_10000_2062, w_10000_2063, w_10000_2064, w_10000_2065, w_10000_2066, w_10000_2067, w_10000_2068, w_10000_2069, w_10000_2070, w_10000_2071, w_10000_2072, w_10000_2073, w_10000_2074, w_10000_2075, w_10000_2076, w_10000_2077, w_10000_2078, w_10000_2079, w_10000_2080, w_10000_2081, w_10000_2082, w_10000_2083, w_10000_2084, w_10000_2085, w_10000_2086, w_10000_2087, w_10000_2088, w_10000_2089, w_10000_2090, w_10000_2091, w_10000_2092, w_10000_2093, w_10000_2094, w_10000_2095, w_10000_2096, w_10000_2097, w_10000_2098, w_10000_2099, w_10000_2100, w_10000_2101, w_10000_2102, w_10000_2103, w_10000_2104, w_10000_2105, w_10000_2106, w_10000_2107, w_10000_2108, w_10000_2109, w_10000_2110, w_10000_2111, w_10000_2112, w_10000_2113, w_10000_2114, w_10000_2115, w_10000_2116, w_10000_2117, w_10000_2118, w_10000_2119, w_10000_2120, w_10000_2121, w_10000_2122, w_10000_2123, w_10000_2124, w_10000_2125, w_10000_2126, w_10000_2127, w_10000_2128, w_10000_2129, w_10000_2130, w_10000_2131, w_10000_2132, w_10000_2133, w_10000_2134, w_10000_2135, w_10000_2136, w_10000_2137, w_10000_2138, w_10000_2139, w_10000_2140, w_10000_2141, w_10000_2142, w_10000_2143, w_10000_2144, w_10000_2145, w_10000_2146, w_10000_2147, w_10000_2148, w_10000_2149, w_10000_2150, w_10000_2151, w_10000_2152, w_10000_2153, w_10000_2154, w_10000_2155, w_10000_2156, w_10000_2157, w_10000_2158, w_10000_2159, w_10000_2160, w_10000_2161, w_10000_2162, w_10000_2163, w_10000_2164, w_10000_2165, w_10000_2166, w_10000_2167, w_10000_2168, w_10000_2169, w_10000_2170, w_10000_2171, w_10000_2172, w_10000_2173, w_10000_2174, w_10000_2175, w_10000_2176, w_10000_2177, w_10000_2178, w_10000_2179, w_10000_2180, w_10000_2181, w_10000_2182, w_10000_2183, w_10000_2184, w_10000_2185, w_10000_2186, w_10000_2187, w_10000_2188, w_10000_2189, w_10000_2190, w_10000_2191, w_10000_2192, w_10000_2193, w_10000_2194, w_10000_2195, w_10000_2196, w_10000_2197, w_10000_2198, w_10000_2199, w_10000_2200, w_10000_2201, w_10000_2202, w_10000_2203, w_10000_2204, w_10000_2205, w_10000_2206, w_10000_2207, w_10000_2208, w_10000_2209, w_10000_2210, w_10000_2211, w_10000_2212, w_10000_2213, w_10000_2214, w_10000_2215, w_10000_2216, w_10000_2217, w_10000_2218, w_10000_2219, w_10000_2220, w_10000_2221, w_10000_2222, w_10000_2223, w_10000_2224, w_10000_2225, w_10000_2226, w_10000_2227, w_10000_2228, w_10000_2229, w_10000_2230, w_10000_2231, w_10000_2232, w_10000_2233, w_10000_2234, w_10000_2235, w_10000_2236, w_10000_2237, w_10000_2238, w_10000_2239, w_10000_2240, w_10000_2241, w_10000_2242, w_10000_2243, w_10000_2244, w_10000_2245, w_10000_2246, w_10000_2247, w_10000_2248, w_10000_2249, w_10000_2250, w_10000_2251, w_10000_2252, w_10000_2253, w_10000_2254, w_10000_2255, w_10000_2256, w_10000_2257, w_10000_2258, w_10000_2259, w_10000_2260, w_10000_2261, w_10000_2262, w_10000_2263, w_10000_2264, w_10000_2265, w_10000_2266, w_10000_2267, w_10000_2268, w_10000_2269, w_10000_2270, w_10000_2271, w_10000_2272, w_10000_2273, w_10000_2274, w_10000_2275, w_10000_2276, w_10000_2277, w_10000_2278, w_10000_2279, w_10000_2280, w_10000_2281, w_10000_2282, w_10000_2283, w_10000_2284, w_10000_2285, w_10000_2286, w_10000_2287, w_10000_2288, w_10000_2289, w_10000_2290, w_10000_2291, w_10000_2292, w_10000_2293, w_10000_2294, w_10000_2295, w_10000_2296, w_10000_2297, w_10000_2298, w_10000_2299, w_10000_2300, w_10000_2301, w_10000_2302, w_10000_2303, w_10000_2304, w_10000_2305, w_10000_2306, w_10000_2307, w_10000_2308, w_10000_2309, w_10000_2310, w_10000_2311, w_10000_2312, w_10000_2313, w_10000_2314, w_10000_2315, w_10000_2316, w_10000_2317, w_10000_2318, w_10000_2319, w_10000_2320, w_10000_2321, w_10000_2322, w_10000_2323, w_10000_2324, w_10000_2325, w_10000_2326, w_10000_2327, w_10000_2328, w_10000_2329, w_10000_2330, w_10000_2331, w_10000_2332, w_10000_2333, w_10000_2334, w_10000_2335, w_10000_2336, w_10000_2337, w_10000_2338, w_10000_2339, w_10000_2340, w_10000_2341, w_10000_2342, w_10000_2343, w_10000_2344, w_10000_2345, w_10000_2346, w_10000_2347, w_10000_2348, w_10000_2349, w_10000_2350, w_10000_2351, w_10000_2352, w_10000_2353, w_10000_2354, w_10000_2355, w_10000_2356, w_10000_2357, w_10000_2358, w_10000_2359, w_10000_2360, w_10000_2361, w_10000_2362, w_10000_2363, w_10000_2364, w_10000_2365, w_10000_2366, w_10000_2367, w_10000_2368, w_10000_2369, w_10000_2370, w_10000_2371, w_10000_2372, w_10000_2373, w_10000_2374, w_10000_2375, w_10000_2376, w_10000_2377, w_10000_2378, w_10000_2379, w_10000_2380, w_10000_2381, w_10000_2382, w_10000_2383, w_10000_2384, w_10000_2385, w_10000_2386, w_10000_2387, w_10000_2388, w_10000_2389, w_10000_2390, w_10000_2391, w_10000_2392, w_10000_2393, w_10000_2394, w_10000_2395, w_10000_2396, w_10000_2397, w_10000_2398, w_10000_2399, w_10000_2400, w_10000_2401, w_10000_2402, w_10000_2403, w_10000_2404, w_10000_2405, w_10000_2406, w_10000_2407, w_10000_2408, w_10000_2409, w_10000_2410, w_10000_2411, w_10000_2412, w_10000_2413, w_10000_2414, w_10000_2415, w_10000_2416, w_10000_2417, w_10000_2418, w_10000_2419, w_10000_2420, w_10000_2421, w_10000_2422, w_10000_2423, w_10000_2424, w_10000_2425, w_10000_2426, w_10000_2427, w_10000_2428, w_10000_2429, w_10000_2430, w_10000_2431, w_10000_2432, w_10000_2433, w_10000_2434, w_10000_2435, w_10000_2436, w_10000_2437, w_10000_2438, w_10000_2439, w_10000_2440, w_10000_2441, w_10000_2442, w_10000_2443, w_10000_2444, w_10000_2445, w_10000_2446, w_10000_2447, w_10000_2448, w_10000_2449, w_10000_2450, w_10000_2451, w_10000_2452, w_10000_2453, w_10000_2454, w_10000_2455, w_10000_2456, w_10000_2457, w_10000_2458, w_10000_2459, w_10000_2460, w_10000_2461, w_10000_2462, w_10000_2463, w_10000_2464, w_10000_2465, w_10000_2466, w_10000_2467, w_10000_2468, w_10000_2469, w_10000_2470, w_10000_2471, w_10000_2472, w_10000_2473, w_10000_2474, w_10000_2475, w_10000_2476, w_10000_2477, w_10000_2478, w_10000_2479, w_10000_2480, w_10000_2481, w_10000_2482, w_10000_2483, w_10000_2484, w_10000_2485, w_10000_2486, w_10000_2487, w_10000_2488, w_10000_2489, w_10000_2490, w_10000_2491, w_10000_2492, w_10000_2493, w_10000_2494, w_10000_2495, w_10000_2496, w_10000_2497, w_10000_2498, w_10000_2499, w_10000_2500, w_10000_2501, w_10000_2502, w_10000_2503, w_10000_2504, w_10000_2505, w_10000_2506, w_10000_2507, w_10000_2508, w_10000_2509, w_10000_2510, w_10000_2511, w_10000_2512, w_10000_2513, w_10000_2514, w_10000_2515, w_10000_2516, w_10000_2517, w_10000_2518, w_10000_2519, w_10000_2520, w_10000_2521, w_10000_2522, w_10000_2523, w_10000_2524, w_10000_2525, w_10000_2526, w_10000_2527, w_10000_2528, w_10000_2529, w_10000_2530, w_10000_2531, w_10000_2532, w_10000_2533, w_10000_2534, w_10000_2535, w_10000_2536, w_10000_2537, w_10000_2538, w_10000_2539, w_10000_2540, w_10000_2541, w_10000_2542, w_10000_2543, w_10000_2544, w_10000_2545, w_10000_2546, w_10000_2547, w_10000_2548, w_10000_2549, w_10000_2550, w_10000_2551, w_10000_2552, w_10000_2553, w_10000_2554, w_10000_2555, w_10000_2556, w_10000_2557, w_10000_2558, w_10000_2559, w_10000_2560, w_10000_2561, w_10000_2562, w_10000_2563, w_10000_2564, w_10000_2565, w_10000_2566, w_10000_2567, w_10000_2568, w_10000_2569, w_10000_2570, w_10000_2571, w_10000_2572, w_10000_2573, w_10000_2574, w_10000_2575, w_10000_2576, w_10000_2577, w_10000_2578, w_10000_2579, w_10000_2580, w_10000_2581, w_10000_2582, w_10000_2583, w_10000_2584, w_10000_2585, w_10000_2586, w_10000_2587, w_10000_2588, w_10000_2589, w_10000_2590, w_10000_2591, w_10000_2592, w_10000_2593, w_10000_2594, w_10000_2595, w_10000_2596, w_10000_2597, w_10000_2598, w_10000_2599, w_10000_2600, w_10000_2601, w_10000_2602, w_10000_2603, w_10000_2604, w_10000_2605, w_10000_2606, w_10000_2607, w_10000_2608, w_10000_2609, w_10000_2610, w_10000_2611, w_10000_2612, w_10000_2613, w_10000_2614, w_10000_2615, w_10000_2616, w_10000_2617, w_10000_2618, w_10000_2619, w_10000_2620, w_10000_2621, w_10000_2622, w_10000_2623, w_10000_2624, w_10000_2625, w_10000_2626, w_10000_2627, w_10000_2628, w_10000_2629, w_10000_2630, w_10000_2631, w_10000_2632, w_10000_2633, w_10000_2634, w_10000_2635, w_10000_2636, w_10000_2637, w_10000_2638, w_10000_2639, w_10000_2640, w_10000_2641, w_10000_2642, w_10000_2643, w_10000_2644, w_10000_2645, w_10000_2646, w_10000_2647, w_10000_2648, w_10000_2649, w_10000_2650, w_10000_2651, w_10000_2652, w_10000_2653, w_10000_2654, w_10000_2655, w_10000_2656, w_10000_2657, w_10000_2658, w_10000_2659, w_10000_2660, w_10000_2661, w_10000_2662, w_10000_2663, w_10000_2664, w_10000_2665, w_10000_2666, w_10000_2667, w_10000_2668, w_10000_2669, w_10000_2670, w_10000_2671, w_10000_2672, w_10000_2673, w_10000_2674, w_10000_2675, w_10000_2676, w_10000_2677, w_10000_2678, w_10000_2679, w_10000_2680, w_10000_2681, w_10000_2682, w_10000_2683, w_10000_2684, w_10000_2685, w_10000_2686, w_10000_2687, w_10000_2688, w_10000_2689, w_10000_2690, w_10000_2691, w_10000_2692, w_10000_2693, w_10000_2694, w_10000_2695, w_10000_2696, w_10000_2697, w_10000_2698, w_10000_2699, w_10000_2700, w_10000_2701, w_10000_2702, w_10000_2703, w_10000_2704, w_10000_2705, w_10000_2706, w_10000_2707, w_10000_2708, w_10000_2709, w_10000_2710, w_10000_2711, w_10000_2712, w_10000_2713, w_10000_2714, w_10000_2715, w_10000_2716, w_10000_2717, w_10000_2718, w_10000_2719, w_10000_2720, w_10000_2721, w_10000_2722, w_10000_2723, w_10000_2724, w_10000_2725, w_10000_2726, w_10000_2727, w_10000_2728, w_10000_2729, w_10000_2730, w_10000_2731, w_10000_2732, w_10000_2733, w_10000_2734, w_10000_2735, w_10000_2736, w_10000_2737, w_10000_2738, w_10000_2739, w_10000_2740, w_10000_2741, w_10000_2742, w_10000_2743, w_10000_2744, w_10000_2745, w_10000_2746, w_10000_2747, w_10000_2748, w_10000_2749, w_10000_2750, w_10000_2751, w_10000_2752, w_10000_2753, w_10000_2754, w_10000_2755, w_10000_2756, w_10000_2757, w_10000_2758, w_10000_2759, w_10000_2760, w_10000_2761, w_10000_2762, w_10000_2763, w_10000_2764, w_10000_2765, w_10000_2766, w_10000_2767, w_10000_2768, w_10000_2769, w_10000_2770, w_10000_2771, w_10000_2772, w_10000_2773, w_10000_2774, w_10000_2775, w_10000_2776, w_10000_2777, w_10000_2778, w_10000_2779, w_10000_2780, w_10000_2781, w_10000_2782, w_10000_2783, w_10000_2784, w_10000_2785, w_10000_2786, w_10000_2787, w_10000_2788, w_10000_2789, w_10000_2790, w_10000_2791, w_10000_2792, w_10000_2793, w_10000_2794, w_10000_2795, w_10000_2796, w_10000_2797, w_10000_2798, w_10000_2799, w_10000_2800, w_10000_2801, w_10000_2802, w_10000_2803, w_10000_2804, w_10000_2805, w_10000_2806, w_10000_2807, w_10000_2808, w_10000_2809, w_10000_2810, w_10000_2811, w_10000_2812, w_10000_2813, w_10000_2814, w_10000_2815, w_10000_2816, w_10000_2817, w_10000_2818, w_10000_2819, w_10000_2820, w_10000_2821, w_10000_2822, w_10000_2823, w_10000_2824, w_10000_2825, w_10000_2826, w_10000_2827, w_10000_2828, w_10000_2829, w_10000_2830, w_10000_2831, w_10000_2832, w_10000_2833, w_10000_2834, w_10000_2835, w_10000_2836, w_10000_2837, w_10000_2838, w_10000_2839, w_10000_2840, w_10000_2841, w_10000_2842, w_10000_2843, w_10000_2844, w_10000_2845, w_10000_2846, w_10000_2847, w_10000_2848, w_10000_2849, w_10000_2850, w_10000_2851, w_10000_2852, w_10000_2853, w_10000_2854, w_10000_2855, w_10000_2856, w_10000_2857, w_10000_2858, w_10000_2859, w_10000_2860, w_10000_2861, w_10000_2862, w_10000_2863, w_10000_2864, w_10000_2865, w_10000_2866, w_10000_2867, w_10000_2868, w_10000_2869, w_10000_2870, w_10000_2871, w_10000_2872, w_10000_2873, w_10000_2874, w_10000_2875, w_10000_2876, w_10000_2877, w_10000_2878, w_10000_2879, w_10000_2880, w_10000_2881, w_10000_2882, w_10000_2883, w_10000_2884, w_10000_2885, w_10000_2886, w_10000_2887, w_10000_2888, w_10000_2889, w_10000_2890, w_10000_2891, w_10000_2892, w_10000_2893, w_10000_2894, w_10000_2895, w_10000_2896, w_10000_2897, w_10000_2898, w_10000_2899, w_10000_2900, w_10000_2901, w_10000_2902, w_10000_2903, w_10000_2904, w_10000_2905, w_10000_2906, w_10000_2907, w_10000_2908, w_10000_2909, w_10000_2910, w_10000_2911, w_10000_2912, w_10000_2913, w_10000_2914, w_10000_2915, w_10000_2916, w_10000_2917, w_10000_2918, w_10000_2919, w_10000_2920, w_10000_2921, w_10000_2922, w_10000_2923, w_10000_2924, w_10000_2925, w_10000_2926, w_10000_2927, w_10000_2928, w_10000_2929, w_10000_2930, w_10000_2931, w_10000_2932, w_10000_2933, w_10000_2934, w_10000_2935, w_10000_2936, w_10000_2937, w_10000_2938, w_10000_2939, w_10000_2940, w_10000_2941, w_10000_2942, w_10000_2943, w_10000_2944, w_10000_2945, w_10000_2946, w_10000_2947, w_10000_2948, w_10000_2949, w_10000_2950, w_10000_2951, w_10000_2952, w_10000_2953, w_10000_2954, w_10000_2955, w_10000_2956, w_10000_2957, w_10000_2958, w_10000_2959, w_10000_2960, w_10000_2961, w_10000_2962, w_10000_2963, w_10000_2964, w_10000_2965, w_10000_2966, w_10000_2967, w_10000_2968, w_10000_2969, w_10000_2970, w_10000_2971, w_10000_2972, w_10000_2973, w_10000_2974, w_10000_2975, w_10000_2976, w_10000_2977, w_10000_2978, w_10000_2979, w_10000_2980, w_10000_2981, w_10000_2982, w_10000_2983, w_10000_2984, w_10000_2985, w_10000_2986, w_10000_2987, w_10000_2988, w_10000_2989, w_10000_2990, w_10000_2991, w_10000_2992, w_10000_2993, w_10000_2994, w_10000_2995, w_10000_2996, w_10000_2997, w_10000_2998, w_10000_2999, w_10000_3000, w_10000_3001, w_10000_3002, w_10000_3003, w_10000_3004, w_10000_3005, w_10000_3006, w_10000_3007, w_10000_3008, w_10000_3009, w_10000_3010, w_10000_3011, w_10000_3012, w_10000_3013, w_10000_3014, w_10000_3015, w_10000_3016, w_10000_3017, w_10000_3018, w_10000_3019, w_10000_3020, w_10000_3021, w_10000_3022, w_10000_3023, w_10000_3024, w_10000_3025, w_10000_3026, w_10000_3027, w_10000_3028, w_10000_3029, w_10000_3030, w_10000_3031, w_10000_3032, w_10000_3033, w_10000_3034, w_10000_3035, w_10000_3036, w_10000_3037, w_10000_3038, w_10000_3039, w_10000_3040, w_10000_3041, w_10000_3042, w_10000_3043, w_10000_3044, w_10000_3045, w_10000_3046, w_10000_3047, w_10000_3048, w_10000_3049, w_10000_3050, w_10000_3051, w_10000_3052, w_10000_3053, w_10000_3054, w_10000_3055, w_10000_3056, w_10000_3057, w_10000_3058, w_10000_3059, w_10000_3060, w_10000_3061, w_10000_3062, w_10000_3063, w_10000_3064, w_10000_3065, w_10000_3066, w_10000_3067, w_10000_3068, w_10000_3069, w_10000_3070, w_10000_3071, w_10000_3072, w_10000_3073, w_10000_3074, w_10000_3075, w_10000_3076, w_10000_3077, w_10000_3078, w_10000_3079, w_10000_3080, w_10000_3081, w_10000_3082, w_10000_3083, w_10000_3084, w_10000_3085, w_10000_3086, w_10000_3087, w_10000_3088, w_10000_3089, w_10000_3090, w_10000_3091, w_10000_3092, w_10000_3093, w_10000_3094, w_10000_3095, w_10000_3096, w_10000_3097, w_10000_3098, w_10000_3099, w_10000_3100, w_10000_3101, w_10000_3102, w_10000_3103, w_10000_3104, w_10000_3105, w_10000_3106, w_10000_3107, w_10000_3108, w_10000_3109, w_10000_3110, w_10000_3111, w_10000_3112, w_10000_3113, w_10000_3114, w_10000_3115, w_10000_3116, w_10000_3117, w_10000_3118, w_10000_3119, w_10000_3120, w_10000_3121, w_10000_3122, w_10000_3123, w_10000_3124, w_10000_3125, w_10000_3126, w_10000_3127, w_10000_3128, w_10000_3129, w_10000_3130, w_10000_3131, w_10000_3132, w_10000_3133, w_10000_3134, w_10000_3135, w_10000_3136, w_10000_3137, w_10000_3138, w_10000_3139, w_10000_3140, w_10000_3141, w_10000_3142, w_10000_3143, w_10000_3144, w_10000_3145, w_10000_3146, w_10000_3147, w_10000_3148, w_10000_3149, w_10000_3150, w_10000_3151, w_10000_3152, w_10000_3153, w_10000_3154, w_10000_3155, w_10000_3156, w_10000_3157, w_10000_3158, w_10000_3159, w_10000_3160, w_10000_3161, w_10000_3162, w_10000_3163, w_10000_3164, w_10000_3165, w_10000_3166, w_10000_3167, w_10000_3168, w_10000_3169, w_10000_3170, w_10000_3171, w_10000_3172, w_10000_3173, w_10000_3174, w_10000_3175, w_10000_3176, w_10000_3177, w_10000_3178, w_10000_3179, w_10000_3180, w_10000_3181, w_10000_3182, w_10000_3183, w_10000_3184, w_10000_3185, w_10000_3186, w_10000_3187, w_10000_3188, w_10000_3189, w_10000_3190, w_10000_3191, w_10000_3192, w_10000_3193, w_10000_3194, w_10000_3195, w_10000_3196, w_10000_3197, w_10000_3198, w_10000_3199, w_10000_3200, w_10000_3201, w_10000_3202, w_10000_3203, w_10000_3204, w_10000_3205, w_10000_3206, w_10000_3207, w_10000_3208, w_10000_3209, w_10000_3210, w_10000_3211, w_10000_3212, w_10000_3213, w_10000_3214, w_10000_3215, w_10000_3216, w_10000_3217, w_10000_3218, w_10000_3219, w_10000_3220, w_10000_3221, w_10000_3222, w_10000_3223, w_10000_3224, w_10000_3225, w_10000_3226, w_10000_3227, w_10000_3228, w_10000_3229, w_10000_3230, w_10000_3231, w_10000_3232, w_10000_3233, w_10000_3234, w_10000_3235, w_10000_3236, w_10000_3237, w_10000_3238, w_10000_3239, w_10000_3240, w_10000_3241, w_10000_3242, w_10000_3243, w_10000_3244, w_10000_3245, w_10000_3246, w_10000_3247, w_10000_3248, w_10000_3249, w_10000_3250, w_10000_3251, w_10000_3252, w_10000_3253, w_10000_3254, w_10000_3255, w_10000_3256, w_10000_3257, w_10000_3258, w_10000_3259, w_10000_3260, w_10000_3261, w_10000_3262, w_10000_3263, w_10000_3264, w_10000_3265, w_10000_3266, w_10000_3267, w_10000_3268, w_10000_3269, w_10000_3270, w_10000_3271, w_10000_3272, w_10000_3273, w_10000_3274, w_10000_3275, w_10000_3276, w_10000_3277, w_10000_3278, w_10000_3279, w_10000_3280, w_10000_3281, w_10000_3282, w_10000_3283, w_10000_3284, w_10000_3285, w_10000_3286, w_10000_3287, w_10000_3288, w_10000_3289, w_10000_3290, w_10000_3291, w_10000_3292, w_10000_3293, w_10000_3294, w_10000_3295, w_10000_3296, w_10000_3297, w_10000_3298, w_10000_3299, w_10000_3300, w_10000_3301, w_10000_3302, w_10000_3303, w_10000_3304, w_10000_3305, w_10000_3306, w_10000_3307, w_10000_3308, w_10000_3309, w_10000_3310, w_10000_3311, w_10000_3312, w_10000_3313, w_10000_3314, w_10000_3315, w_10000_3316, w_10000_3317, w_10000_3318, w_10000_3319, w_10000_3320, w_10000_3321, w_10000_3322, w_10000_3323, w_10000_3324, w_10000_3325, w_10000_3326, w_10000_3327, w_10000_3328, w_10000_3329, w_10000_3330, w_10000_3331, w_10000_3332, w_10000_3333, w_10000_3334, w_10000_3335, w_10000_3336, w_10000_3337, w_10000_3338, w_10000_3339, w_10000_3340, w_10000_3341, w_10000_3342, w_10000_3343, w_10000_3344, w_10000_3345, w_10000_3346, w_10000_3347, w_10000_3348, w_10000_3349, w_10000_3350, w_10000_3351, w_10000_3352, w_10000_3353, w_10000_3354, w_10000_3355, w_10000_3356, w_10000_3357, w_10000_3358, w_10000_3359, w_10000_3360, w_10000_3361, w_10000_3362, w_10000_3363, w_10000_3364, w_10000_3365, w_10000_3366, w_10000_3367, w_10000_3368, w_10000_3369, w_10000_3370, w_10000_3371, w_10000_3372, w_10000_3373, w_10000_3374, w_10000_3375, w_10000_3376, w_10000_3377, w_10000_3378, w_10000_3379, w_10000_3380, w_10000_3381, w_10000_3382, w_10000_3383, w_10000_3384, w_10000_3385, w_10000_3386, w_10000_3387, w_10000_3388, w_10000_3389, w_10000_3390, w_10000_3391, w_10000_3392, w_10000_3393, w_10000_3394, w_10000_3395, w_10000_3396, w_10000_3397, w_10000_3398, w_10000_3399, w_10000_3400, w_10000_3401, w_10000_3402, w_10000_3403, w_10000_3404, w_10000_3405, w_10000_3406, w_10000_3407, w_10000_3408, w_10000_3409, w_10000_3410, w_10000_3411, w_10000_3412, w_10000_3413, w_10000_3414, w_10000_3415, w_10000_3416, w_10000_3417, w_10000_3418, w_10000_3419, w_10000_3420, w_10000_3421, w_10000_3422, w_10000_3423, w_10000_3424, w_10000_3425, w_10000_3426, w_10000_3427, w_10000_3428, w_10000_3429, w_10000_3430, w_10000_3431, w_10000_3432, w_10000_3433, w_10000_3434, w_10000_3435, w_10000_3436, w_10000_3437, w_10000_3438, w_10000_3439, w_10000_3440, w_10000_3441, w_10000_3442, w_10000_3443, w_10000_3444, w_10000_3445, w_10000_3446, w_10000_3447, w_10000_3448, w_10000_3449, w_10000_3450, w_10000_3451, w_10000_3452, w_10000_3453, w_10000_3454, w_10000_3455, w_10000_3456, w_10000_3457, w_10000_3458, w_10000_3459, w_10000_3460, w_10000_3461, w_10000_3462, w_10000_3463, w_10000_3464, w_10000_3465, w_10000_3466, w_10000_3467, w_10000_3468, w_10000_3469, w_10000_3470, w_10000_3471, w_10000_3472, w_10000_3473, w_10000_3474, w_10000_3475, w_10000_3476, w_10000_3477, w_10000_3478, w_10000_3479, w_10000_3480, w_10000_3481, w_10000_3482, w_10000_3483, w_10000_3484, w_10000_3485, w_10000_3486, w_10000_3487, w_10000_3488, w_10000_3489, w_10000_3490, w_10000_3491, w_10000_3492, w_10000_3493, w_10000_3494, w_10000_3495, w_10000_3496, w_10000_3497, w_10000_3498, w_10000_3499, w_10000_3500, w_10000_3501, w_10000_3502, w_10000_3503, w_10000_3504, w_10000_3505, w_10000_3506, w_10000_3507, w_10000_3508, w_10000_3509, w_10000_3510, w_10000_3511, w_10000_3512, w_10000_3513, w_10000_3514, w_10000_3515, w_10000_3516, w_10000_3517, w_10000_3518, w_10000_3519, w_10000_3520, w_10000_3521, w_10000_3522, w_10000_3523, w_10000_3524, w_10000_3525, w_10000_3526, w_10000_3527, w_10000_3528, w_10000_3529, w_10000_3530, w_10000_3531, w_10000_3532, w_10000_3533, w_10000_3534, w_10000_3535, w_10000_3536, w_10000_3537, w_10000_3538, w_10000_3539, w_10000_3540, w_10000_3541, w_10000_3542, w_10000_3543, w_10000_3544, w_10000_3545, w_10000_3546, w_10000_3547, w_10000_3548, w_10000_3549, w_10000_3550, w_10000_3551, w_10000_3552, w_10000_3553, w_10000_3554, w_10000_3555, w_10000_3556, w_10000_3557, w_10000_3558, w_10000_3559, w_10000_3560, w_10000_3561, w_10000_3562, w_10000_3563, w_10000_3564, w_10000_3565, w_10000_3566, w_10000_3567, w_10000_3568, w_10000_3569, w_10000_3570, w_10000_3571, w_10000_3572, w_10000_3573, w_10000_3574, w_10000_3575, w_10000_3576, w_10000_3577, w_10000_3578, w_10000_3579, w_10000_3580, w_10000_3581, w_10000_3582, w_10000_3583, w_10000_3584, w_10000_3585, w_10000_3586, w_10000_3587, w_10000_3588, w_10000_3589, w_10000_3590, w_10000_3591, w_10000_3592, w_10000_3593, w_10000_3594, w_10000_3595, w_10000_3596, w_10000_3597, w_10000_3598, w_10000_3599, w_10000_3600, w_10000_3601, w_10000_3602, w_10000_3603, w_10000_3604, w_10000_3605, w_10000_3606, w_10000_3607, w_10000_3608, w_10000_3609, w_10000_3610, w_10000_3611, w_10000_3612, w_10000_3613, w_10000_3614, w_10000_3615, w_10000_3616, w_10000_3617, w_10000_3618, w_10000_3619, w_10000_3620, w_10000_3621, w_10000_3622, w_10000_3623, w_10000_3624, w_10000_3625, w_10000_3626, w_10000_3627, w_10000_3628, w_10000_3629, w_10000_3630, w_10000_3631, w_10000_3632, w_10000_3633, w_10000_3634, w_10000_3635, w_10000_3636, w_10000_3637, w_10000_3638, w_10000_3639, w_10000_3640, w_10000_3641, w_10000_3642, w_10000_3643, w_10000_3644, w_10000_3645, w_10000_3646, w_10000_3647, w_10000_3648, w_10000_3649, w_10000_3650, w_10000_3651, w_10000_3652, w_10000_3653, w_10000_3654, w_10000_3655, w_10000_3656, w_10000_3657, w_10000_3658, w_10000_3659, w_10000_3660, w_10000_3661, w_10000_3662, w_10000_3663, w_10000_3664, w_10000_3665, w_10000_3666, w_10000_3667, w_10000_3668, w_10000_3669, w_10000_3670, w_10000_3671, w_10000_3672, w_10000_3673, w_10000_3674, w_10000_3675, w_10000_3676, w_10000_3677, w_10000_3678, w_10000_3679, w_10000_3680, w_10000_3681, w_10000_3682, w_10000_3683, w_10000_3684, w_10000_3685, w_10000_3686, w_10000_3687, w_10000_3688, w_10000_3689, w_10000_3690, w_10000_3691, w_10000_3692, w_10000_3693, w_10000_3694, w_10000_3695, w_10000_3696, w_10000_3697, w_10000_3698, w_10000_3699, w_10000_3700, w_10000_3701, w_10000_3702, w_10000_3703, w_10000_3704, w_10000_3705, w_10000_3706, w_10000_3707, w_10000_3708, w_10000_3709, w_10000_3710, w_10000_3711, w_10000_3712, w_10000_3713, w_10000_3714, w_10000_3715, w_10000_3716, w_10000_3717, w_10000_3718, w_10000_3719, w_10000_3720, w_10000_3721, w_10000_3722, w_10000_3723, w_10000_3724, w_10000_3725, w_10000_3726, w_10000_3727, w_10000_3728, w_10000_3729, w_10000_3730, w_10000_3731, w_10000_3732, w_10000_3733, w_10000_3734, w_10000_3735, w_10000_3736, w_10000_3737, w_10000_3738, w_10000_3739, w_10000_3740, w_10000_3741, w_10000_3742, w_10000_3743, w_10000_3744, w_10000_3745, w_10000_3746, w_10000_3747, w_10000_3748, w_10000_3749, w_10000_3750, w_10000_3751, w_10000_3752, w_10000_3753, w_10000_3754, w_10000_3755, w_10000_3756, w_10000_3757, w_10000_3758, w_10000_3759, w_10000_3760, w_10000_3761, w_10000_3762, w_10000_3763, w_10000_3764, w_10000_3765, w_10000_3766, w_10000_3767, w_10000_3768, w_10000_3769, w_10000_3770, w_10000_3771, w_10000_3772, w_10000_3773, w_10000_3774, w_10000_3775, w_10000_3776, w_10000_3777, w_10000_3778, w_10000_3779, w_10000_3780, w_10000_3781, w_10000_3782, w_10000_3783, w_10000_3784, w_10000_3785, w_10000_3786, w_10000_3787, w_10000_3788, w_10000_3789, w_10000_3790, w_10000_3791, w_10000_3792, w_10000_3793, w_10000_3794, w_10000_3795, w_10000_3796, w_10000_3797, w_10000_3798, w_10000_3799, w_10000_3800, w_10000_3801, w_10000_3802, w_10000_3803, w_10000_3804, w_10000_3805, w_10000_3806, w_10000_3807, w_10000_3808, w_10000_3809, w_10000_3810, w_10000_3811, w_10000_3812, w_10000_3813, w_10000_3814, w_10000_3815, w_10000_3816, w_10000_3817, w_10000_3818, w_10000_3819, w_10000_3820, w_10000_3821, w_10000_3822, w_10000_3823, w_10000_3824, w_10000_3825, w_10000_3826, w_10000_3827, w_10000_3828, w_10000_3829, w_10000_3830, w_10000_3831, w_10000_3832, w_10000_3833, w_10000_3834, w_10000_3835, w_10000_3836, w_10000_3837, w_10000_3838, w_10000_3839, w_10000_3840, w_10000_3841, w_10000_3842, w_10000_3843, w_10000_3844, w_10000_3845, w_10000_3846, w_10000_3847, w_10000_3848, w_10000_3849, w_10000_3850, w_10000_3851, w_10000_3852, w_10000_3853, w_10000_3854, w_10000_3855, w_10000_3856, w_10000_3857, w_10000_3858, w_10000_3859, w_10000_3860, w_10000_3861, w_10000_3862, w_10000_3863, w_10000_3864, w_10000_3865, w_10000_3866, w_10000_3867, w_10000_3868, w_10000_3869, w_10000_3870, w_10000_3871, w_10000_3872, w_10000_3873, w_10000_3874, w_10000_3875, w_10000_3876, w_10000_3877, w_10000_3878, w_10000_3879, w_10000_3880, w_10000_3881, w_10000_3882, w_10000_3883, w_10000_3884, w_10000_3885, w_10000_3886, w_10000_3887, w_10000_3888, w_10000_3889, w_10000_3890, w_10000_3891, w_10000_3892, w_10000_3893, w_10000_3894, w_10000_3895, w_10000_3896, w_10000_3897, w_10000_3898, w_10000_3899, w_10000_3900, w_10000_3901, w_10000_3902, w_10000_3903, w_10000_3904, w_10000_3905, w_10000_3906, w_10000_3907, w_10000_3908, w_10000_3909, w_10000_3910, w_10000_3911, w_10000_3912, w_10000_3913, w_10000_3914, w_10000_3915, w_10000_3916, w_10000_3917, w_10000_3918, w_10000_3919, w_10000_3920, w_10000_3921, w_10000_3922, w_10000_3923, w_10000_3924, w_10000_3925, w_10000_3926, w_10000_3927, w_10000_3928, w_10000_3929, w_10000_3930, w_10000_3931, w_10000_3932, w_10000_3933, w_10000_3934, w_10000_3935, w_10000_3936, w_10000_3937, w_10000_3938, w_10000_3939, w_10000_3940, w_10000_3941, w_10000_3942, w_10000_3943, w_10000_3944, w_10000_3945, w_10000_3946, w_10000_3947, w_10000_3948, w_10000_3949, w_10000_3950, w_10000_3951, w_10000_3952, w_10000_3953, w_10000_3954, w_10000_3955, w_10000_3956, w_10000_3957, w_10000_3958, w_10000_3959, w_10000_3960, w_10000_3961, w_10000_3962, w_10000_3963, w_10000_3964, w_10000_3965, w_10000_3966, w_10000_3967, w_10000_3968, w_10000_3969, w_10000_3970, w_10000_3971, w_10000_3972, w_10000_3973, w_10000_3974, w_10000_3975, w_10000_3976, w_10000_3977, w_10000_3978, w_10000_3979, w_10000_3980, w_10000_3981, w_10000_3982, w_10000_3983, w_10000_3984, w_10000_3985, w_10000_3986, w_10000_3987, w_10000_3988, w_10000_3989, w_10000_3990, w_10000_3991, w_10000_3992, w_10000_3993, w_10000_3994, w_10000_3995, w_10000_3996, w_10000_3997, w_10000_3998, w_10000_3999, w_10000_4000, w_10000_4001, w_10000_4002, w_10000_4003, w_10000_4004, w_10000_4005, w_10000_4006, w_10000_4007, w_10000_4008, w_10000_4009, w_10000_4010, w_10000_4011, w_10000_4012, w_10000_4013, w_10000_4014, w_10000_4015, w_10000_4016, w_10000_4017, w_10000_4018, w_10000_4019, w_10000_4020, w_10000_4021, w_10000_4022, w_10000_4023, w_10000_4024, w_10000_4025, w_10000_4026, w_10000_4027, w_10000_4028, w_10000_4029, w_10000_4030, w_10000_4031, w_10000_4032, w_10000_4033, w_10000_4034, w_10000_4035, w_10000_4036, w_10000_4037, w_10000_4038, w_10000_4039, w_10000_4040, w_10000_4041, w_10000_4042, w_10000_4043, w_10000_4044, w_10000_4045, w_10000_4046, w_10000_4047, w_10000_4048, w_10000_4049, w_10000_4050, w_10000_4051, w_10000_4052, w_10000_4053, w_10000_4054, w_10000_4055, w_10000_4056, w_10000_4057, w_10000_4058, w_10000_4059, w_10000_4060, w_10000_4061, w_10000_4062, w_10000_4063, w_10000_4064, w_10000_4065, w_10000_4066, w_10000_4067, w_10000_4068, w_10000_4069, w_10000_4070, w_10000_4071, w_10000_4072, w_10000_4073, w_10000_4074, w_10000_4075, w_10000_4076, w_10000_4077, w_10000_4078, w_10000_4079, w_10000_4080, w_10000_4081, w_10000_4082, w_10000_4083, w_10000_4084, w_10000_4085, w_10000_4086, w_10000_4087, w_10000_4088, w_10000_4089, w_10000_4090, w_10000_4091, w_10000_4092, w_10000_4093, w_10000_4094, w_10000_4095, w_10000_4096, w_10000_4097, w_10000_4098, w_10000_4099, w_10000_4100, w_10000_4101, w_10000_4102, w_10000_4103, w_10000_4104, w_10000_4105, w_10000_4106, w_10000_4107, w_10000_4108, w_10000_4109, w_10000_4110, w_10000_4111, w_10000_4112, w_10000_4113, w_10000_4114, w_10000_4115, w_10000_4116, w_10000_4117, w_10000_4118, w_10000_4119, w_10000_4120, w_10000_4121, w_10000_4122, w_10000_4123, w_10000_4124, w_10000_4125, w_10000_4126, w_10000_4127, w_10000_4128, w_10000_4129, w_10000_4130, w_10000_4131, w_10000_4132, w_10000_4133, w_10000_4134, w_10000_4135, w_10000_4136, w_10000_4137, w_10000_4138, w_10000_4139, w_10000_4140, w_10000_4141, w_10000_4142, w_10000_4143, w_10000_4144, w_10000_4145, w_10000_4146, w_10000_4147, w_10000_4148, w_10000_4149, w_10000_4150, w_10000_4151, w_10000_4152, w_10000_4153, w_10000_4154, w_10000_4155, w_10000_4156, w_10000_4157, w_10000_4158, w_10000_4159, w_10000_4160, w_10000_4161, w_10000_4162, w_10000_4163, w_10000_4164, w_10000_4165, w_10000_4166, w_10000_4167, w_10000_4168, w_10000_4169, w_10000_4170, w_10000_4171, w_10000_4172, w_10000_4173, w_10000_4174, w_10000_4175, w_10000_4176, w_10000_4177, w_10000_4178, w_10000_4179, w_10000_4180, w_10000_4181, w_10000_4182, w_10000_4183, w_10000_4184, w_10000_4185, w_10000_4186, w_10000_4187, w_10000_4188, w_10000_4189, w_10000_4190, w_10000_4191, w_10000_4192, w_10000_4193, w_10000_4194, w_10000_4195, w_10000_4196, w_10000_4197, w_10000_4198, w_10000_4199, w_10000_4200, w_10000_4201, w_10000_4202, w_10000_4203, w_10000_4204, w_10000_4205, w_10000_4206, w_10000_4207, w_10000_4208, w_10000_4209, w_10000_4210, w_10000_4211, w_10000_4212, w_10000_4213, w_10000_4214, w_10000_4215, w_10000_4216, w_10000_4217, w_10000_4218, w_10000_4219, w_10000_4220, w_10000_4221, w_10000_4222, w_10000_4223, w_10000_4224, w_10000_4225, w_10000_4226, w_10000_4227, w_10000_4228, w_10000_4229, w_10000_4230, w_10000_4231, w_10000_4232, w_10000_4233, w_10000_4234, w_10000_4235, w_10000_4236, w_10000_4237, w_10000_4238, w_10000_4239, w_10000_4240, w_10000_4241, w_10000_4242, w_10000_4243, w_10000_4244, w_10000_4245, w_10000_4246, w_10000_4247, w_10000_4248, w_10000_4249, w_10000_4250, w_10000_4251, w_10000_4252, w_10000_4253, w_10000_4254, w_10000_4255, w_10000_4256, w_10000_4257, w_10000_4258, w_10000_4259, w_10000_4260, w_10000_4261, w_10000_4262, w_10000_4263, w_10000_4264, w_10000_4265, w_10000_4266, w_10000_4267, w_10000_4268, w_10000_4269, w_10000_4270, w_10000_4271, w_10000_4272, w_10000_4273, w_10000_4274, w_10000_4275, w_10000_4276, w_10000_4277, w_10000_4278, w_10000_4279, w_10000_4280, w_10000_4281, w_10000_4282, w_10000_4283, w_10000_4284, w_10000_4285, w_10000_4286, w_10000_4287, w_10000_4288, w_10000_4289, w_10000_4290, w_10000_4291, w_10000_4292, w_10000_4293, w_10000_4294, w_10000_4295, w_10000_4296, w_10000_4297, w_10000_4298, w_10000_4299, w_10000_4300, w_10000_4301, w_10000_4302, w_10000_4303, w_10000_4304, w_10000_4305, w_10000_4306, w_10000_4307, w_10000_4308, w_10000_4309, w_10000_4310, w_10000_4311, w_10000_4312, w_10000_4313, w_10000_4314, w_10000_4315, w_10000_4316, w_10000_4317, w_10000_4318, w_10000_4319, w_10000_4320, w_10000_4321, w_10000_4322, w_10000_4323, w_10000_4324, w_10000_4325, w_10000_4326, w_10000_4327, w_10000_4328, w_10000_4329, w_10000_4330, w_10000_4331, w_10000_4332, w_10000_4333, w_10000_4334, w_10000_4335, w_10000_4336, w_10000_4337, w_10000_4338, w_10000_4339, w_10000_4340, w_10000_4341, w_10000_4342, w_10000_4343, w_10000_4344, w_10000_4345, w_10000_4346, w_10000_4347, w_10000_4348, w_10000_4349, w_10000_4350, w_10000_4351, w_10000_4352, w_10000_4353, w_10000_4354, w_10000_4355, w_10000_4356, w_10000_4357, w_10000_4358, w_10000_4359, w_10000_4360, w_10000_4361, w_10000_4362, w_10000_4363, w_10000_4364, w_10000_4365, w_10000_4366, w_10000_4367, w_10000_4368, w_10000_4369, w_10000_4370, w_10000_4371, w_10000_4372, w_10000_4373, w_10000_4374, w_10000_4375, w_10000_4376, w_10000_4377, w_10000_4378, w_10000_4379, w_10000_4380, w_10000_4381, w_10000_4382, w_10000_4383, w_10000_4384, w_10000_4385, w_10000_4386, w_10000_4387, w_10000_4388, w_10000_4389, w_10000_4390, w_10000_4391, w_10000_4392, w_10000_4393, w_10000_4394, w_10000_4395, w_10000_4396, w_10000_4397, w_10000_4398, w_10000_4399, w_10000_4400, w_10000_4401, w_10000_4402, w_10000_4403, w_10000_4404, w_10000_4405, w_10000_4406, w_10000_4407, w_10000_4408, w_10000_4409, w_10000_4410, w_10000_4411, w_10000_4412, w_10000_4413, w_10000_4414, w_10000_4415, w_10000_4416, w_10000_4417, w_10000_4418, w_10000_4419, w_10000_4420, w_10000_4421, w_10000_4422, w_10000_4423, w_10000_4424, w_10000_4425, w_10000_4426, w_10000_4427, w_10000_4428, w_10000_4429, w_10000_4430, w_10000_4431, w_10000_4432, w_10000_4433, w_10000_4434, w_10000_4435, w_10000_4436, w_10000_4437, w_10000_4438, w_10000_4439, w_10000_4440, w_10000_4441, w_10000_4442, w_10000_4443, w_10000_4444, w_10000_4445, w_10000_4446, w_10000_4447, w_10000_4448, w_10000_4449, w_10000_4450, w_10000_4451, w_10000_4452, w_10000_4453, w_10000_4454, w_10000_4455, w_10000_4456, w_10000_4457, w_10000_4458, w_10000_4459, w_10000_4460, w_10000_4461, w_10000_4462, w_10000_4463, w_10000_4464, w_10000_4465, w_10000_4466, w_10000_4467, w_10000_4468, w_10000_4469, w_10000_4470, w_10000_4471, w_10000_4472, w_10000_4473, w_10000_4474, w_10000_4475, w_10000_4476, w_10000_4477, w_10000_4478, w_10000_4479, w_10000_4480, w_10000_4481, w_10000_4482, w_10000_4483, w_10000_4484, w_10000_4485, w_10000_4486, w_10000_4487, w_10000_4488, w_10000_4489, w_10000_4490, w_10000_4491, w_10000_4492, w_10000_4493, w_10000_4494, w_10000_4495, w_10000_4496, w_10000_4497, w_10000_4498, w_10000_4499, w_10000_4500, w_10000_4501, w_10000_4502, w_10000_4503, w_10000_4504, w_10000_4505, w_10000_4506, w_10000_4507, w_10000_4508, w_10000_4509, w_10000_4510, w_10000_4511, w_10000_4512, w_10000_4513, w_10000_4514, w_10000_4515, w_10000_4516, w_10000_4517, w_10000_4518, w_10000_4519, w_10000_4520, w_10000_4521, w_10000_4522, w_10000_4523, w_10000_4524, w_10000_4525, w_10000_4526, w_10000_4527, w_10000_4528, w_10000_4529, w_10000_4530, w_10000_4531, w_10000_4532, w_10000_4533, w_10000_4534, w_10000_4535, w_10000_4536, w_10000_4537, w_10000_4538, w_10000_4539, w_10000_4540, w_10000_4541, w_10000_4542, w_10000_4543, w_10000_4544, w_10000_4545, w_10000_4546, w_10000_4547, w_10000_4548, w_10000_4549, w_10000_4550, w_10000_4551, w_10000_4552, w_10000_4553, w_10000_4554, w_10000_4555, w_10000_4556, w_10000_4557, w_10000_4558, w_10000_4559, w_10000_4560, w_10000_4561, w_10000_4562, w_10000_4563, w_10000_4564, w_10000_4565, w_10000_4566, w_10000_4567, w_10000_4568, w_10000_4569, w_10000_4570, w_10000_4571, w_10000_4572, w_10000_4573, w_10000_4574, w_10000_4575, w_10000_4576, w_10000_4577, w_10000_4578, w_10000_4579, w_10000_4580, w_10000_4581, w_10000_4582, w_10000_4583, w_10000_4584, w_10000_4585, w_10000_4586, w_10000_4587, w_10000_4588, w_10000_4589, w_10000_4590, w_10000_4591, w_10000_4592, w_10000_4593, w_10000_4594, w_10000_4595, w_10000_4596, w_10000_4597, w_10000_4598, w_10000_4599, w_10000_4600, w_10000_4601, w_10000_4602, w_10000_4603, w_10000_4604, w_10000_4605, w_10000_4606, w_10000_4607, w_10000_4608, w_10000_4609, w_10000_4610, w_10000_4611, w_10000_4612, w_10000_4613, w_10000_4614, w_10000_4615, w_10000_4616, w_10000_4617, w_10000_4618, w_10000_4619, w_10000_4620, w_10000_4621, w_10000_4622, w_10000_4623, w_10000_4624, w_10000_4625, w_10000_4626, w_10000_4627, w_10000_4628, w_10000_4629, w_10000_4630, w_10000_4631, w_10000_4632, w_10000_4633, w_10000_4634, w_10000_4635, w_10000_4636, w_10000_4637, w_10000_4638, w_10000_4639, w_10000_4640, w_10000_4641, w_10000_4642, w_10000_4643, w_10000_4644, w_10000_4645, w_10000_4646, w_10000_4647, w_10000_4648, w_10000_4649, w_10000_4650, w_10000_4651, w_10000_4652, w_10000_4653, w_10000_4654, w_10000_4655, w_10000_4656, w_10000_4657, w_10000_4658, w_10000_4659, w_10000_4660, w_10000_4661, w_10000_4662, w_10000_4663, w_10000_4664, w_10000_4665, w_10000_4666, w_10000_4667, w_10000_4668, w_10000_4669, w_10000_4670, w_10000_4671, w_10000_4672, w_10000_4673, w_10000_4674, w_10000_4675, w_10000_4676, w_10000_4677, w_10000_4678, w_10000_4679, w_10000_4680, w_10000_4681, w_10000_4682, w_10000_4683, w_10000_4684, w_10000_4685, w_10000_4686, w_10000_4687, w_10000_4688, w_10000_4689, w_10000_4690, w_10000_4691, w_10000_4692, w_10000_4693, w_10000_4694, w_10000_4695, w_10000_4696, w_10000_4697, w_10000_4698, w_10000_4699, w_10000_4700, w_10000_4701, w_10000_4702, w_10000_4703, w_10000_4704, w_10000_4705, w_10000_4706, w_10000_4707, w_10000_4708, w_10000_4709, w_10000_4710, w_10000_4711, w_10000_4712, w_10000_4713, w_10000_4714, w_10000_4715, w_10000_4716, w_10000_4717, w_10000_4718, w_10000_4719, w_10000_4720, w_10000_4721, w_10000_4722, w_10000_4723, w_10000_4724, w_10000_4725, w_10000_4726, w_10000_4727, w_10000_4728, w_10000_4729, w_10000_4730, w_10000_4731, w_10000_4732, w_10000_4733, w_10000_4734, w_10000_4735, w_10000_4736, w_10000_4737, w_10000_4738, w_10000_4739, w_10000_4740, w_10000_4741, w_10000_4742, w_10000_4743, w_10000_4744, w_10000_4745, w_10000_4746, w_10000_4747, w_10000_4748, w_10000_4749, w_10000_4750, w_10000_4751, w_10000_4752, w_10000_4753, w_10000_4754, w_10000_4755, w_10000_4756, w_10000_4757, w_10000_4758, w_10000_4759, w_10000_4760, w_10000_4761, w_10000_4762, w_10000_4763, w_10000_4764, w_10000_4765, w_10000_4766, w_10000_4767, w_10000_4768, w_10000_4769, w_10000_4770, w_10000_4771, w_10000_4772, w_10000_4773, w_10000_4774, w_10000_4775, w_10000_4776, w_10000_4777, w_10000_4778, w_10000_4779, w_10000_4780, w_10000_4781, w_10000_4782, w_10000_4783, w_10000_4784, w_10000_4785, w_10000_4786, w_10000_4787, w_10000_4788, w_10000_4789, w_10000_4790, w_10000_4791, w_10000_4792, w_10000_4793, w_10000_4794, w_10000_4795, w_10000_4796, w_10000_4797, w_10000_4798, w_10000_4799, w_10000_4800, w_10000_4801, w_10000_4802, w_10000_4803, w_10000_4804, w_10000_4805, w_10000_4806, w_10000_4807, w_10000_4808, w_10000_4809, w_10000_4810, w_10000_4811, w_10000_4812, w_10000_4813, w_10000_4814, w_10000_4815, w_10000_4816, w_10000_4817, w_10000_4818, w_10000_4819, w_10000_4820, w_10000_4821, w_10000_4822, w_10000_4823, w_10000_4824, w_10000_4825, w_10000_4826, w_10000_4827, w_10000_4828, w_10000_4829, w_10000_4830, w_10000_4831, w_10000_4832, w_10000_4833, w_10000_4834, w_10000_4835, w_10000_4836, w_10000_4837, w_10000_4838, w_10000_4839, w_10000_4840, w_10000_4841, w_10000_4842, w_10000_4843, w_10000_4844, w_10000_4845, w_10000_4846, w_10000_4847, w_10000_4848, w_10000_4849, w_10000_4850, w_10000_4851, w_10000_4852, w_10000_4853, w_10000_4854, w_10000_4855, w_10000_4856, w_10000_4857, w_10000_4858, w_10000_4859, w_10000_4860, w_10000_4861, w_10000_4862, w_10000_4863, w_10000_4864, w_10000_4865, w_10000_4866, w_10000_4867, w_10000_4868, w_10000_4869, w_10000_4870, w_10000_4871, w_10000_4872, w_10000_4873, w_10000_4874, w_10000_4875, w_10000_4876, w_10000_4877, w_10000_4878, w_10000_4879, w_10000_4880, w_10000_4881, w_10000_4882, w_10000_4883, w_10000_4884, w_10000_4885, w_10000_4886, w_10000_4887, w_10000_4888, w_10000_4889, w_10000_4890, w_10000_4891, w_10000_4892, w_10000_4893, w_10000_4894, w_10000_4895, w_10000_4896, w_10000_4897, w_10000_4898, w_10000_4899, w_10000_4900, w_10000_4901, w_10000_4902, w_10000_4903, w_10000_4904, w_10000_4905, w_10000_4906, w_10000_4907, w_10000_4908, w_10000_4909, w_10000_4910, w_10000_4911, w_10000_4912, w_10000_4913, w_10000_4914, w_10000_4915, w_10000_4916, w_10000_4917, w_10000_4918, w_10000_4919, w_10000_4920, w_10000_4921, w_10000_4922, w_10000_4923, w_10000_4924, w_10000_4925, w_10000_4926, w_10000_4927, w_10000_4928, w_10000_4929, w_10000_4930, w_10000_4931, w_10000_4932, w_10000_4933, w_10000_4934, w_10000_4935, w_10000_4936, w_10000_4937, w_10000_4938, w_10000_4939, w_10000_4940, w_10000_4941, w_10000_4942, w_10000_4943, w_10000_4944, w_10000_4945, w_10000_4946, w_10000_4947, w_10000_4948, w_10000_4949, w_10000_4950, w_10000_4951, w_10000_4952, w_10000_4953, w_10000_4954, w_10000_4955, w_10000_4956, w_10000_4957, w_10000_4958, w_10000_4959, w_10000_4960, w_10000_4961, w_10000_4962, w_10000_4963, w_10000_4964, w_10000_4965, w_10000_4966, w_10000_4967, w_10000_4968, w_10000_4969, w_10000_4970, w_10000_4971, w_10000_4972, w_10000_4973, w_10000_4974, w_10000_4975, w_10000_4976, w_10000_4977, w_10000_4978, w_10000_4979, w_10000_4980, w_10000_4981, w_10000_4982, w_10000_4983, w_10000_4984, w_10000_4985, w_10000_4986, w_10000_4987, w_10000_4988, w_10000_4989, w_10000_4990, w_10000_4991, w_10000_4992, w_10000_4993, w_10000_4994, w_10000_4995, w_10000_4996, w_10000_4997, w_10000_4998, w_10000_4999, w_10000_5000, w_10000_5001, w_10000_5002, w_10000_5003, w_10000_5004, w_10000_5005, w_10000_5006, w_10000_5007, w_10000_5008, w_10000_5009, w_10000_5010, w_10000_5011, w_10000_5012, w_10000_5013, w_10000_5014, w_10000_5015, w_10000_5016, w_10000_5017, w_10000_5018, w_10000_5019, w_10000_5020, w_10000_5021, w_10000_5022, w_10000_5023, w_10000_5024, w_10000_5025, w_10000_5026, w_10000_5027, w_10000_5028, w_10000_5029, w_10000_5030, w_10000_5031, w_10000_5032, w_10000_5033, w_10000_5034, w_10000_5035, w_10000_5036, w_10000_5037, w_10000_5038, w_10000_5039, w_10000_5040, w_10000_5041, w_10000_5042, w_10000_5043, w_10000_5044, w_10000_5045, w_10000_5046, w_10000_5047, w_10000_5048, w_10000_5049, w_10000_5050, w_10000_5051, w_10000_5052, w_10000_5053, w_10000_5054, w_10000_5055, w_10000_5056, w_10000_5057, w_10000_5058, w_10000_5059, w_10000_5060, w_10000_5061, w_10000_5062, w_10000_5063, w_10000_5064, w_10000_5065, w_10000_5066, w_10000_5067, w_10000_5068, w_10000_5069, w_10000_5070, w_10000_5071, w_10000_5072, w_10000_5073, w_10000_5074, w_10000_5075, w_10000_5076, w_10000_5077, w_10000_5078, w_10000_5079, w_10000_5080, w_10000_5081, w_10000_5082, w_10000_5083, w_10000_5084, w_10000_5085, w_10000_5086, w_10000_5087, w_10000_5088, w_10000_5089, w_10000_5090, w_10000_5091, w_10000_5092, w_10000_5093, w_10000_5094, w_10000_5095, w_10000_5096, w_10000_5097, w_10000_5098, w_10000_5099, w_10000_5100, w_10000_5101, w_10000_5102, w_10000_5103, w_10000_5104, w_10000_5105, w_10000_5106, w_10000_5107, w_10000_5108, w_10000_5109, w_10000_5110, w_10000_5111, w_10000_5112, w_10000_5113, w_10000_5114, w_10000_5115, w_10000_5116, w_10000_5117, w_10000_5118, w_10000_5119, w_10000_5120, w_10000_5121, w_10000_5122, w_10000_5123, w_10000_5124, w_10000_5125, w_10000_5126, w_10000_5127, w_10000_5128, w_10000_5129, w_10000_5130, w_10000_5131, w_10000_5132, w_10000_5133, w_10000_5134, w_10000_5135, w_10000_5136, w_10000_5137, w_10000_5138, w_10000_5139, w_10000_5140, w_10000_5141, w_10000_5142, w_10000_5143, w_10000_5144, w_10000_5145, w_10000_5146, w_10000_5147, w_10000_5148, w_10000_5149, w_10000_5150, w_10000_5151, w_10000_5152, w_10000_5153, w_10000_5154, w_10000_5155, w_10000_5156, w_10000_5157, w_10000_5158, w_10000_5159, w_10000_5160, w_10000_5161, w_10000_5162, w_10000_5163, w_10000_5164, w_10000_5165, w_10000_5166, w_10000_5167, w_10000_5168, w_10000_5169, w_10000_5170, w_10000_5171, w_10000_5172, w_10000_5173, w_10000_5174, w_10000_5175, w_10000_5176, w_10000_5177, w_10000_5178, w_10000_5179, w_10000_5180, w_10000_5181, w_10000_5182, w_10000_5183, w_10000_5184, w_10000_5185, w_10000_5186, w_10000_5187, w_10000_5188, w_10000_5189, w_10000_5190, w_10000_5191, w_10000_5192, w_10000_5193, w_10000_5194, w_10000_5195, w_10000_5196, w_10000_5197, w_10000_5198, w_10000_5199, w_10000_5200, w_10000_5201, w_10000_5202, w_10000_5203, w_10000_5204, w_10000_5205, w_10000_5206, w_10000_5207, w_10000_5208, w_10000_5209, w_10000_5210, w_10000_5211, w_10000_5212, w_10000_5213, w_10000_5214, w_10000_5215, w_10000_5216, w_10000_5217, w_10000_5218, w_10000_5219, w_10000_5220, w_10000_5221, w_10000_5222, w_10000_5223, w_10000_5224, w_10000_5225, w_10000_5226, w_10000_5227, w_10000_5228, w_10000_5229, w_10000_5230, w_10000_5231, w_10000_5232, w_10000_5233, w_10000_5234, w_10000_5235, w_10000_5236, w_10000_5237, w_10000_5238, w_10000_5239, w_10000_5240, w_10000_5241, w_10000_5242, w_10000_5243, w_10000_5244, w_10000_5245, w_10000_5246, w_10000_5247, w_10000_5248, w_10000_5249, w_10000_5250, w_10000_5251, w_10000_5252, w_10000_5253, w_10000_5254, w_10000_5255, w_10000_5256, w_10000_5257, w_10000_5258, w_10000_5259, w_10000_5260, w_10000_5261, w_10000_5262, w_10000_5263, w_10000_5264, w_10000_5265, w_10000_5266, w_10000_5267, w_10000_5268, w_10000_5269, w_10000_5270, w_10000_5271, w_10000_5272, w_10000_5273, w_10000_5274, w_10000_5275, w_10000_5276, w_10000_5277, w_10000_5278, w_10000_5279, w_10000_5280, w_10000_5281, w_10000_5282, w_10000_5283, w_10000_5284, w_10000_5285, w_10000_5286, w_10000_5287, w_10000_5288, w_10000_5289, w_10000_5290, w_10000_5291, w_10000_5292, w_10000_5293, w_10000_5294, w_10000_5295, w_10000_5296, w_10000_5297, w_10000_5298, w_10000_5299, w_10000_5300, w_10000_5301, w_10000_5302, w_10000_5303, w_10000_5304, w_10000_5305, w_10000_5306, w_10000_5307, w_10000_5308, w_10000_5309, w_10000_5310, w_10000_5311, w_10000_5312, w_10000_5313, w_10000_5314, w_10000_5315, w_10000_5316, w_10000_5317, w_10000_5318, w_10000_5319, w_10000_5320, w_10000_5321, w_10000_5322, w_10000_5323, w_10000_5324, w_10000_5325, w_10000_5326, w_10000_5327, w_10000_5328, w_10000_5329, w_10000_5330, w_10000_5331, w_10000_5332, w_10000_5333, w_10000_5334, w_10000_5335, w_10000_5336, w_10000_5337, w_10000_5338, w_10000_5339, w_10000_5340, w_10000_5341, w_10000_5342, w_10000_5343, w_10000_5344, w_10000_5345, w_10000_5346, w_10000_5347, w_10000_5348, w_10000_5349, w_10000_5350, w_10000_5351, w_10000_5352, w_10000_5353, w_10000_5354, w_10000_5355, w_10000_5356, w_10000_5357, w_10000_5358, w_10000_5359, w_10000_5360, w_10000_5361, w_10000_5362, w_10000_5363, w_10000_5364, w_10000_5365, w_10000_5366, w_10000_5367, w_10000_5368, w_10000_5369, w_10000_5370, w_10000_5371, w_10000_5372, w_10000_5373, w_10000_5374, w_10000_5375, w_10000_5376, w_10000_5377, w_10000_5378, w_10000_5379, w_10000_5380, w_10000_5381, w_10000_5382, w_10000_5383, w_10000_5384, w_10000_5385, w_10000_5386, w_10000_5387, w_10000_5388, w_10000_5389, w_10000_5390, w_10000_5391, w_10000_5392, w_10000_5393, w_10000_5394, w_10000_5395, w_10000_5396, w_10000_5397, w_10000_5398, w_10000_5399, w_10000_5400, w_10000_5401, w_10000_5402, w_10000_5403, w_10000_5404, w_10000_5405, w_10000_5406, w_10000_5407, w_10000_5408, w_10000_5409, w_10000_5410, w_10000_5411, w_10000_5412, w_10000_5413, w_10000_5414, w_10000_5415, w_10000_5416, w_10000_5417, w_10000_5418, w_10000_5419, w_10000_5420, w_10000_5421, w_10000_5422, w_10000_5423, w_10000_5424, w_10000_5425, w_10000_5426, w_10000_5427, w_10000_5428, w_10000_5429, w_10000_5430, w_10000_5431, w_10000_5432, w_10000_5433, w_10000_5434, w_10000_5435, w_10000_5436, w_10000_5437, w_10000_5438, w_10000_5439, w_10000_5440, w_10000_5441, w_10000_5442, w_10000_5443, w_10000_5444, w_10000_5445, w_10000_5446, w_10000_5447, w_10000_5448, w_10000_5449, w_10000_5450, w_10000_5451, w_10000_5452, w_10000_5453, w_10000_5454, w_10000_5455, w_10000_5456, w_10000_5457, w_10000_5458, w_10000_5459, w_10000_5460, w_10000_5461, w_10000_5462, w_10000_5463, w_10000_5464, w_10000_5465, w_10000_5466, w_10000_5467, w_10000_5468, w_10000_5469, w_10000_5470, w_10000_5471, w_10000_5472, w_10000_5473, w_10000_5474, w_10000_5475, w_10000_5476, w_10000_5477, w_10000_5478, w_10000_5479, w_10000_5480, w_10000_5481, w_10000_5482, w_10000_5483, w_10000_5484, w_10000_5485, w_10000_5486, w_10000_5487, w_10000_5488, w_10000_5489, w_10000_5490, w_10000_5491, w_10000_5492, w_10000_5493, w_10000_5494, w_10000_5495, w_10000_5496, w_10000_5497, w_10000_5498, w_10000_5499, w_10000_5500, w_10000_5501, w_10000_5502, w_10000_5503, w_10000_5504, w_10000_5505, w_10000_5506, w_10000_5507, w_10000_5508, w_10000_5509, w_10000_5510, w_10000_5511, w_10000_5512, w_10000_5513, w_10000_5514, w_10000_5515, w_10000_5516, w_10000_5517, w_10000_5518, w_10000_5519, w_10000_5520, w_10000_5521, w_10000_5522, w_10000_5523, w_10000_5524, w_10000_5525, w_10000_5526, w_10000_5527, w_10000_5528, w_10000_5529, w_10000_5530, w_10000_5531, w_10000_5532, w_10000_5533, w_10000_5534, w_10000_5535, w_10000_5536, w_10000_5537, w_10000_5538, w_10000_5539, w_10000_5540, w_10000_5541, w_10000_5542, w_10000_5543, w_10000_5544, w_10000_5545, w_10000_5546, w_10000_5547, w_10000_5548, w_10000_5549, w_10000_5550, w_10000_5551, w_10000_5552, w_10000_5553, w_10000_5554, w_10000_5555, w_10000_5556, w_10000_5557, w_10000_5558, w_10000_5559, w_10000_5560, w_10000_5561, w_10000_5562, w_10000_5563, w_10000_5564, w_10000_5565, w_10000_5566, w_10000_5567, w_10000_5568, w_10000_5569, w_10000_5570, w_10000_5571, w_10000_5572, w_10000_5573, w_10000_5574, w_10000_5575, w_10000_5576, w_10000_5577, w_10000_5578, w_10000_5579, w_10000_5580, w_10000_5581, w_10000_5582, w_10000_5583, w_10000_5584, w_10000_5585, w_10000_5586, w_10000_5587, w_10000_5588, w_10000_5589, w_10000_5590, w_10000_5591, w_10000_5592, w_10000_5593, w_10000_5594, w_10000_5595, w_10000_5596, w_10000_5597, w_10000_5598, w_10000_5599, w_10000_5600, w_10000_5601, w_10000_5602, w_10000_5603, w_10000_5604, w_10000_5605, w_10000_5606, w_10000_5607, w_10000_5608, w_10000_5609, w_10000_5610, w_10000_5611, w_10000_5612, w_10000_5613, w_10000_5614, w_10000_5615, w_10000_5616, w_10000_5617, w_10000_5618, w_10000_5619, w_10000_5620, w_10000_5621, w_10000_5622, w_10000_5623, w_10000_5624, w_10000_5625, w_10000_5626, w_10000_5627, w_10000_5628, w_10000_5629, w_10000_5630, w_10000_5631, w_10000_5632, w_10000_5633, w_10000_5634, w_10000_5635, w_10000_5636, w_10000_5637, w_10000_5638, w_10000_5639, w_10000_5640, w_10000_5641, w_10000_5642, w_10000_5643, w_10000_5644, w_10000_5645, w_10000_5646, w_10000_5647, w_10000_5648, w_10000_5649, w_10000_5650, w_10000_5651, w_10000_5652, w_10000_5653, w_10000_5654, w_10000_5655, w_10000_5656, w_10000_5657, w_10000_5658, w_10000_5659, w_10000_5660, w_10000_5661, w_10000_5662, w_10000_5663, w_10000_5664, w_10000_5665, w_10000_5666, w_10000_5667, w_10000_5668, w_10000_5669, w_10000_5670, w_10000_5671, w_10000_5672, w_10000_5673, w_10000_5674, w_10000_5675, w_10000_5676, w_10000_5677, w_10000_5678, w_10000_5679, w_10000_5680, w_10000_5681, w_10000_5682, w_10000_5683, w_10000_5684, w_10000_5685, w_10000_5686, w_10000_5687, w_10000_5688, w_10000_5689, w_10000_5690, w_10000_5691, w_10000_5692, w_10000_5693, w_10000_5694, w_10000_5695, w_10000_5696, w_10000_5697, w_10000_5698, w_10000_5699, w_10000_5700, w_10000_5701, w_10000_5702, w_10000_5703, w_10000_5704, w_10000_5705, w_10000_5706, w_10000_5707, w_10000_5708, w_10000_5709, w_10000_5710, w_10000_5711, w_10000_5712, w_10000_5713, w_10000_5714, w_10000_5715, w_10000_5716, w_10000_5717, w_10000_5718, w_10000_5719, w_10000_5720, w_10000_5721, w_10000_5722, w_10000_5723, w_10000_5724, w_10000_5725, w_10000_5726, w_10000_5727, w_10000_5728, w_10000_5729, w_10000_5730, w_10000_5731, w_10000_5732, w_10000_5733, w_10000_5734, w_10000_5735, w_10000_5736, w_10000_5737, w_10000_5738, w_10000_5739, w_10000_5740, w_10000_5741, w_10000_5742, w_10000_5743, w_10000_5744, w_10000_5745, w_10000_5746, w_10000_5747, w_10000_5748, w_10000_5749, w_10000_5750, w_10000_5751, w_10000_5752, w_10000_5753, w_10000_5754, w_10000_5755, w_10000_5756, w_10000_5757, w_10000_5758, w_10000_5759, w_10000_5760, w_10000_5761, w_10000_5762, w_10000_5763, w_10000_5764, w_10000_5765, w_10000_5766, w_10000_5767, w_10000_5768, w_10000_5769, w_10000_5770, w_10000_5771, w_10000_5772, w_10000_5773, w_10000_5774, w_10000_5775, w_10000_5776, w_10000_5777, w_10000_5778, w_10000_5779, w_10000_5780, w_10000_5781, w_10000_5782, w_10000_5783, w_10000_5784, w_10000_5785, w_10000_5786, w_10000_5787, w_10000_5788, w_10000_5789, w_10000_5790, w_10000_5791, w_10000_5792, w_10000_5793, w_10000_5794, w_10000_5795, w_10000_5796, w_10000_5797, w_10000_5798, w_10000_5799, w_10000_5800, w_10000_5801, w_10000_5802, w_10000_5803, w_10000_5804, w_10000_5805, w_10000_5806, w_10000_5807, w_10000_5808, w_10000_5809, w_10000_5810, w_10000_5811, w_10000_5812, w_10000_5813, w_10000_5814, w_10000_5815, w_10000_5816, w_10000_5817, w_10000_5818, w_10000_5819, w_10000_5820, w_10000_5821, w_10000_5822, w_10000_5823, w_10000_5824, w_10000_5825, w_10000_5826, w_10000_5827, w_10000_5828, w_10000_5829, w_10000_5830, w_10000_5831, w_10000_5832, w_10000_5833, w_10000_5834, w_10000_5835, w_10000_5836, w_10000_5837, w_10000_5838, w_10000_5839, w_10000_5840, w_10000_5841, w_10000_5842, w_10000_5843, w_10000_5844, w_10000_5845, w_10000_5846, w_10000_5847, w_10000_5848, w_10000_5849, w_10000_5850, w_10000_5851, w_10000_5852, w_10000_5853, w_10000_5854, w_10000_5855, w_10000_5856, w_10000_5857, w_10000_5858, w_10000_5859, w_10000_5860, w_10000_5861, w_10000_5862, w_10000_5863, w_10000_5864, w_10000_5865, w_10000_5866, w_10000_5867, w_10000_5868, w_10000_5869, w_10000_5870, w_10000_5871, w_10000_5872, w_10000_5873, w_10000_5874, w_10000_5875, w_10000_5876, w_10000_5877, w_10000_5878, w_10000_5879, w_10000_5880, w_10000_5881, w_10000_5882, w_10000_5883, w_10000_5884, w_10000_5885, w_10000_5886, w_10000_5887, w_10000_5888, w_10000_5889, w_10000_5890, w_10000_5891, w_10000_5892, w_10000_5893, w_10000_5894, w_10000_5895, w_10000_5896, w_10000_5897, w_10000_5898, w_10000_5899, w_10000_5900, w_10000_5901, w_10000_5902, w_10000_5903, w_10000_5904, w_10000_5905, w_10000_5906, w_10000_5907, w_10000_5908, w_10000_5909, w_10000_5910, w_10000_5911, w_10000_5912, w_10000_5913, w_10000_5914, w_10000_5915, w_10000_5916, w_10000_5917, w_10000_5918, w_10000_5919, w_10000_5920, w_10000_5921, w_10000_5922, w_10000_5923, w_10000_5924, w_10000_5925, w_10000_5926, w_10000_5927, w_10000_5928, w_10000_5929, w_10000_5930, w_10000_5931, w_10000_5932, w_10000_5933, w_10000_5934, w_10000_5935, w_10000_5936, w_10000_5937, w_10000_5938, w_10000_5939, w_10000_5940, w_10000_5941, w_10000_5942, w_10000_5943, w_10000_5944, w_10000_5945, w_10000_5946, w_10000_5947, w_10000_5948, w_10000_5949, w_10000_5950, w_10000_5951, w_10000_5952, w_10000_5953, w_10000_5954, w_10000_5955, w_10000_5956, w_10000_5957, w_10000_5958, w_10000_5959, w_10000_5960, w_10000_5961, w_10000_5962, w_10000_5963, w_10000_5964, w_10000_5965, w_10000_5966, w_10000_5967, w_10000_5968, w_10000_5969, w_10000_5970, w_10000_5971, w_10000_5972, w_10000_5973, w_10000_5974, w_10000_5975, w_10000_5976, w_10000_5977, w_10000_5978, w_10000_5979, w_10000_5980, w_10000_5981, w_10000_5982, w_10000_5983, w_10000_5984, w_10000_5985, w_10000_5986, w_10000_5987, w_10000_5988, w_10000_5989, w_10000_5990, w_10000_5991, w_10000_5992, w_10000_5993, w_10000_5994, w_10000_5995, w_10000_5996, w_10000_5997, w_10000_5998, w_10000_5999, w_10000_6000, w_10000_6001, w_10000_6002, w_10000_6003, w_10000_6004, w_10000_6005, w_10000_6006, w_10000_6007, w_10000_6008, w_10000_6009, w_10000_6010, w_10000_6011, w_10000_6012, w_10000_6013, w_10000_6014, w_10000_6015, w_10000_6016, w_10000_6017, w_10000_6018, w_10000_6019, w_10000_6020, w_10000_6021, w_10000_6022, w_10000_6023, w_10000_6024, w_10000_6025, w_10000_6026, w_10000_6027, w_10000_6028, w_10000_6029, w_10000_6030, w_10000_6031, w_10000_6032, w_10000_6033, w_10000_6034, w_10000_6035, w_10000_6036, w_10000_6037, w_10000_6038, w_10000_6039, w_10000_6040, w_10000_6041, w_10000_6042, w_10000_6043, w_10000_6044, w_10000_6045, w_10000_6046, w_10000_6047, w_10000_6048, w_10000_6049, w_10000_6050, w_10000_6051, w_10000_6052, w_10000_6053, w_10000_6054, w_10000_6055, w_10000_6056, w_10000_6057, w_10000_6058, w_10000_6059, w_10000_6060, w_10000_6061, w_10000_6062, w_10000_6063, w_10000_6064, w_10000_6065, w_10000_6066, w_10000_6067, w_10000_6068, w_10000_6069, w_10000_6070, w_10000_6071, w_10000_6072, w_10000_6073, w_10000_6074, w_10000_6075, w_10000_6076, w_10000_6077, w_10000_6078, w_10000_6079, w_10000_6080, w_10000_6081, w_10000_6082, w_10000_6083, w_10000_6084, w_10000_6085, w_10000_6086, w_10000_6087, w_10000_6088, w_10000_6089, w_10000_6090, w_10000_6091, w_10000_6092, w_10000_6093, w_10000_6094, w_10000_6095, w_10000_6096, w_10000_6097, w_10000_6098, w_10000_6099, w_10000_6100, w_10000_6101, w_10000_6102, w_10000_6103, w_10000_6104, w_10000_6105, w_10000_6106, w_10000_6107, w_10000_6108, w_10000_6109, w_10000_6110, w_10000_6111, w_10000_6112, w_10000_6113, w_10000_6114, w_10000_6115, w_10000_6116, w_10000_6117, w_10000_6118, w_10000_6119, w_10000_6120, w_10000_6121, w_10000_6122, w_10000_6123, w_10000_6124, w_10000_6125, w_10000_6126, w_10000_6127, w_10000_6128, w_10000_6129, w_10000_6130, w_10000_6131, w_10000_6132, w_10000_6133, w_10000_6134, w_10000_6135, w_10000_6136, w_10000_6137, w_10000_6138, w_10000_6139, w_10000_6140, w_10000_6141, w_10000_6142, w_10000_6143, w_10000_6144, w_10000_6145, w_10000_6146, w_10000_6147, w_10000_6148, w_10000_6149, w_10000_6150, w_10000_6151, w_10000_6152, w_10000_6153, w_10000_6154, w_10000_6155, w_10000_6156, w_10000_6157, w_10000_6158, w_10000_6159, w_10000_6160, w_10000_6161, w_10000_6162, w_10000_6163, w_10000_6164, w_10000_6165, w_10000_6166, w_10000_6167, w_10000_6168, w_10000_6169, w_10000_6170, w_10000_6171, w_10000_6172, w_10000_6173, w_10000_6174, w_10000_6175, w_10000_6176, w_10000_6177, w_10000_6178, w_10000_6179, w_10000_6180, w_10000_6181, w_10000_6182, w_10000_6183, w_10000_6184, w_10000_6185, w_10000_6186, w_10000_6187, w_10000_6188, w_10000_6189, w_10000_6190, w_10000_6191, w_10000_6192, w_10000_6193, w_10000_6194, w_10000_6195, w_10000_6196, w_10000_6197, w_10000_6198, w_10000_6199, w_10000_6200, w_10000_6201, w_10000_6202, w_10000_6203, w_10000_6204, w_10000_6205, w_10000_6206, w_10000_6207, w_10000_6208, w_10000_6209, w_10000_6210, w_10000_6211, w_10000_6212, w_10000_6213, w_10000_6214, w_10000_6215, w_10000_6216, w_10000_6217, w_10000_6218, w_10000_6219, w_10000_6220, w_10000_6221, w_10000_6222, w_10000_6223, w_10000_6224, w_10000_6225, w_10000_6226, w_10000_6227, w_10000_6228, w_10000_6229, w_10000_6230, w_10000_6231, w_10000_6232, w_10000_6233, w_10000_6234, w_10000_6235, w_10000_6236, w_10000_6237, w_10000_6238, w_10000_6239, w_10000_6240, w_10000_6241, w_10000_6242, w_10000_6243, w_10000_6244, w_10000_6245, w_10000_6246, w_10000_6247, w_10000_6248, w_10000_6249, w_10000_6250, w_10000_6251, w_10000_6252, w_10000_6253, w_10000_6254, w_10000_6255, w_10000_6256, w_10000_6257, w_10000_6258, w_10000_6259, w_10000_6260, w_10000_6261, w_10000_6262, w_10000_6263, w_10000_6264, w_10000_6265, w_10000_6266, w_10000_6267, w_10000_6268, w_10000_6269, w_10000_6270, w_10000_6271, w_10000_6272, w_10000_6273, w_10000_6274, w_10000_6275, w_10000_6276, w_10000_6277, w_10000_6278, w_10000_6279, w_10000_6280, w_10000_6281, w_10000_6282, w_10000_6283, w_10000_6284, w_10000_6285, w_10000_6286, w_10000_6287, w_10000_6288, w_10000_6289, w_10000_6290, w_10000_6291, w_10000_6292, w_10000_6293, w_10000_6294, w_10000_6295, w_10000_6296, w_10000_6297, w_10000_6298, w_10000_6299, w_10000_6300, w_10000_6301, w_10000_6302, w_10000_6303, w_10000_6304, w_10000_6305, w_10000_6306, w_10000_6307, w_10000_6308, w_10000_6309, w_10000_6310, w_10000_6311, w_10000_6312, w_10000_6313, w_10000_6314, w_10000_6315, w_10000_6316, w_10000_6317, w_10000_6318, w_10000_6319, w_10000_6320, w_10000_6321, w_10000_6322, w_10000_6323, w_10000_6324, w_10000_6325, w_10000_6326, w_10000_6327, w_10000_6328, w_10000_6329, w_10000_6330, w_10000_6331, w_10000_6332, w_10000_6333, w_10000_6334, w_10000_6335, w_10000_6336, w_10000_6337, w_10000_6338, w_10000_6339, w_10000_6340, w_10000_6341, w_10000_6342, w_10000_6343, w_10000_6344, w_10000_6345, w_10000_6346, w_10000_6347, w_10000_6348, w_10000_6349, w_10000_6350, w_10000_6351, w_10000_6352, w_10000_6353, w_10000_6354, w_10000_6355, w_10000_6356, w_10000_6357, w_10000_6358, w_10000_6359, w_10000_6360, w_10000_6361, w_10000_6362, w_10000_6363, w_10000_6364, w_10000_6365, w_10000_6366, w_10000_6367, w_10000_6368, w_10000_6369, w_10000_6370, w_10000_6371, w_10000_6372, w_10000_6373, w_10000_6374, w_10000_6375, w_10000_6376, w_10000_6377, w_10000_6378, w_10000_6379, w_10000_6380, w_10000_6381, w_10000_6382, w_10000_6383, w_10000_6384, w_10000_6385, w_10000_6386, w_10000_6387, w_10000_6388, w_10000_6389, w_10000_6390, w_10000_6391, w_10000_6392, w_10000_6393, w_10000_6394, w_10000_6395, w_10000_6396, w_10000_6397, w_10000_6398, w_10000_6399, w_10000_6400, w_10000_6401, w_10000_6402, w_10000_6403, w_10000_6404, w_10000_6405, w_10000_6406, w_10000_6407, w_10000_6408, w_10000_6409, w_10000_6410, w_10000_6411, w_10000_6412, w_10000_6413, w_10000_6414, w_10000_6415, w_10000_6416, w_10000_6417, w_10000_6418, w_10000_6419, w_10000_6420, w_10000_6421, w_10000_6422, w_10000_6423, w_10000_6424, w_10000_6425, w_10000_6426, w_10000_6427, w_10000_6428, w_10000_6429, w_10000_6430, w_10000_6431, w_10000_6432, w_10000_6433, w_10000_6434, w_10000_6435, w_10000_6436, w_10000_6437, w_10000_6438, w_10000_6439, w_10000_6440, w_10000_6441, w_10000_6442, w_10000_6443, w_10000_6444, w_10000_6445, w_10000_6446, w_10000_6447, w_10000_6448, w_10000_6449, w_10000_6450, w_10000_6451, w_10000_6452, w_10000_6453, w_10000_6454, w_10000_6455, w_10000_6456, w_10000_6457, w_10000_6458, w_10000_6459, w_10000_6460, w_10000_6461, w_10000_6462, w_10000_6463, w_10000_6464, w_10000_6465, w_10000_6466, w_10000_6467, w_10000_6468, w_10000_6469, w_10000_6470, w_10000_6471, w_10000_6472, w_10000_6473, w_10000_6474, w_10000_6475, w_10000_6476, w_10000_6477, w_10000_6478, w_10000_6479, w_10000_6480, w_10000_6481, w_10000_6482, w_10000_6483, w_10000_6484, w_10000_6485, w_10000_6486, w_10000_6487, w_10000_6488, w_10000_6489, w_10000_6490, w_10000_6491, w_10000_6492, w_10000_6493, w_10000_6494, w_10000_6495, w_10000_6496, w_10000_6497, w_10000_6498, w_10000_6499, w_10000_6500, w_10000_6501, w_10000_6502, w_10000_6503, w_10000_6504, w_10000_6505, w_10000_6506, w_10000_6507, w_10000_6508, w_10000_6509, w_10000_6510, w_10000_6511, w_10000_6512, w_10000_6513, w_10000_6514, w_10000_6515, w_10000_6516, w_10000_6517, w_10000_6518, w_10000_6519, w_10000_6520, w_10000_6521, w_10000_6522, w_10000_6523, w_10000_6524, w_10000_6525, w_10000_6526, w_10000_6527, w_10000_6528, w_10000_6529, w_10000_6530, w_10000_6531, w_10000_6532, w_10000_6533, w_10000_6534, w_10000_6535, w_10000_6536, w_10000_6537, w_10000_6538, w_10000_6539, w_10000_6540, w_10000_6541, w_10000_6542, w_10000_6543, w_10000_6544, w_10000_6545, w_10000_6546, w_10000_6547, w_10000_6548, w_10000_6549, w_10000_6550, w_10000_6551, w_10000_6552, w_10000_6553, w_10000_6554, w_10000_6555, w_10000_6556, w_10000_6557, w_10000_6558, w_10000_6559, w_10000_6560, w_10000_6561, w_10000_6562, w_10000_6563, w_10000_6564, w_10000_6565, w_10000_6566, w_10000_6567, w_10000_6568, w_10000_6569, w_10000_6570, w_10000_6571, w_10000_6572, w_10000_6573, w_10000_6574, w_10000_6575, w_10000_6576, w_10000_6577, w_10000_6578, w_10000_6579, w_10000_6580, w_10000_6581, w_10000_6582, w_10000_6583, w_10000_6584, w_10000_6585, w_10000_6586, w_10000_6587, w_10000_6588, w_10000_6589, w_10000_6590, w_10000_6591, w_10000_6592, w_10000_6593, w_10000_6594, w_10000_6595, w_10000_6596, w_10000_6597, w_10000_6598, w_10000_6599, w_10000_6600, w_10000_6601, w_10000_6602, w_10000_6603, w_10000_6604, w_10000_6605, w_10000_6606, w_10000_6607, w_10000_6608, w_10000_6609, w_10000_6610, w_10000_6611, w_10000_6612, w_10000_6613, w_10000_6614, w_10000_6615, w_10000_6616, w_10000_6617, w_10000_6618, w_10000_6619, w_10000_6620, w_10000_6621, w_10000_6622, w_10000_6623, w_10000_6624, w_10000_6625, w_10000_6626, w_10000_6627, w_10000_6628, w_10000_6629, w_10000_6630, w_10000_6631, w_10000_6632, w_10000_6633, w_10000_6634, w_10000_6635, w_10000_6636, w_10000_6637, w_10000_6638, w_10000_6639, w_10000_6640, w_10000_6641, w_10000_6642, w_10000_6643, w_10000_6644, w_10000_6645, w_10000_6646, w_10000_6647, w_10000_6648, w_10000_6649, w_10000_6650, w_10000_6651, w_10000_6652, w_10000_6653, w_10000_6654, w_10000_6655, w_10000_6656, w_10000_6657, w_10000_6658, w_10000_6659, w_10000_6660, w_10000_6661, w_10000_6662, w_10000_6663, w_10000_6664, w_10000_6665, w_10000_6666, w_10000_6667, w_10000_6668, w_10000_6669, w_10000_6670, w_10000_6671, w_10000_6672, w_10000_6673, w_10000_6674, w_10000_6675, w_10000_6676, w_10000_6677, w_10000_6678, w_10000_6679, w_10000_6680, w_10000_6681, w_10000_6682, w_10000_6683, w_10000_6684, w_10000_6685, w_10000_6686, w_10000_6687, w_10000_6688, w_10000_6689, w_10000_6690, w_10000_6691, w_10000_6692, w_10000_6693, w_10000_6694, w_10000_6695, w_10000_6696, w_10000_6697, w_10000_6698, w_10000_6699, w_10000_6700, w_10000_6701, w_10000_6702, w_10000_6703, w_10000_6704, w_10000_6705, w_10000_6706, w_10000_6707, w_10000_6708, w_10000_6709, w_10000_6710, w_10000_6711, w_10000_6712, w_10000_6713, w_10000_6714, w_10000_6715, w_10000_6716, w_10000_6717, w_10000_6718, w_10000_6719, w_10000_6720, w_10000_6721, w_10000_6722, w_10000_6723, w_10000_6724, w_10000_6725, w_10000_6726, w_10000_6727, w_10000_6728, w_10000_6729, w_10000_6730, w_10000_6731, w_10000_6732, w_10000_6733, w_10000_6734, w_10000_6735, w_10000_6736, w_10000_6737, w_10000_6738, w_10000_6739, w_10000_6740, w_10000_6741, w_10000_6742, w_10000_6743, w_10000_6744, w_10000_6745, w_10000_6746, w_10000_6747, w_10000_6748, w_10000_6749, w_10000_6750, w_10000_6751, w_10000_6752, w_10000_6753, w_10000_6754, w_10000_6755, w_10000_6756, w_10000_6757, w_10000_6758, w_10000_6759, w_10000_6760, w_10000_6761, w_10000_6762, w_10000_6763, w_10000_6764, w_10000_6765, w_10000_6766, w_10000_6767, w_10000_6768, w_10000_6769, w_10000_6770, w_10000_6771, w_10000_6772, w_10000_6773, w_10000_6774, w_10000_6775, w_10000_6776, w_10000_6777, w_10000_6778, w_10000_6779, w_10000_6780, w_10000_6781, w_10000_6782, w_10000_6783, w_10000_6784, w_10000_6785, w_10000_6786, w_10000_6787, w_10000_6788, w_10000_6789, w_10000_6790, w_10000_6791, w_10000_6792, w_10000_6793, w_10000_6794, w_10000_6795, w_10000_6796, w_10000_6797, w_10000_6798, w_10000_6799, w_10000_6800, w_10000_6801, w_10000_6802, w_10000_6803, w_10000_6804, w_10000_6805, w_10000_6806, w_10000_6807, w_10000_6808, w_10000_6809, w_10000_6810, w_10000_6811, w_10000_6812, w_10000_6813, w_10000_6814, w_10000_6815, w_10000_6816, w_10000_6817, w_10000_6818, w_10000_6819, w_10000_6820, w_10000_6821, w_10000_6822, w_10000_6823, w_10000_6824, w_10000_6825, w_10000_6826, w_10000_6827, w_10000_6828, w_10000_6829, w_10000_6830, w_10000_6831, w_10000_6832, w_10000_6833, w_10000_6834, w_10000_6835, w_10000_6836, w_10000_6837, w_10000_6838, w_10000_6839, w_10000_6840, w_10000_6841, w_10000_6842, w_10000_6843, w_10000_6844, w_10000_6845, w_10000_6846, w_10000_6847, w_10000_6848, w_10000_6849, w_10000_6850, w_10000_6851, w_10000_6852, w_10000_6853, w_10000_6854, w_10000_6855, w_10000_6856, w_10000_6857, w_10000_6858, w_10000_6859, w_10000_6860, w_10000_6861, w_10000_6862, w_10000_6863, w_10000_6864, w_10000_6865, w_10000_6866, w_10000_6867, w_10000_6868, w_10000_6869, w_10000_6870, w_10000_6871, w_10000_6872, w_10000_6873, w_10000_6874, w_10000_6875, w_10000_6876, w_10000_6877, w_10000_6878, w_10000_6879, w_10000_6880, w_10000_6881, w_10000_6882, w_10000_6883, w_10000_6884, w_10000_6885, w_10000_6886, w_10000_6887, w_10000_6888, w_10000_6889, w_10000_6890, w_10000_6891, w_10000_6892, w_10000_6893, w_10000_6894, w_10000_6895, w_10000_6896, w_10000_6897, w_10000_6898, w_10000_6899, w_10000_6900, w_10000_6901, w_10000_6902, w_10000_6903, w_10000_6904, w_10000_6905, w_10000_6906, w_10000_6907, w_10000_6908, w_10000_6909, w_10000_6910, w_10000_6911, w_10000_6912, w_10000_6913, w_10000_6914, w_10000_6915, w_10000_6916, w_10000_6917, w_10000_6918, w_10000_6919, w_10000_6920, w_10000_6921, w_10000_6922, w_10000_6923, w_10000_6924, w_10000_6925, w_10000_6926, w_10000_6927, w_10000_6928, w_10000_6929, w_10000_6930, w_10000_6931, w_10000_6932, w_10000_6933, w_10000_6934, w_10000_6935, w_10000_6936, w_10000_6937, w_10000_6938, w_10000_6939, w_10000_6940, w_10000_6941, w_10000_6942, w_10000_6943, w_10000_6944, w_10000_6945, w_10000_6946, w_10000_6947, w_10000_6948, w_10000_6949, w_10000_6950, w_10000_6951, w_10000_6952, w_10000_6953, w_10000_6954, w_10000_6955, w_10000_6956, w_10000_6957, w_10000_6958, w_10000_6959, w_10000_6960, w_10000_6961, w_10000_6962, w_10000_6963, w_10000_6964, w_10000_6965, w_10000_6966, w_10000_6967, w_10000_6968, w_10000_6969, w_10000_6970, w_10000_6971, w_10000_6972, w_10000_6973, w_10000_6974, w_10000_6975, w_10000_6976, w_10000_6977, w_10000_6978, w_10000_6979, w_10000_6980, w_10000_6981, w_10000_6982, w_10000_6983, w_10000_6984, w_10000_6985, w_10000_6986, w_10000_6987, w_10000_6988, w_10000_6989, w_10000_6990, w_10000_6991, w_10000_6992, w_10000_6993, w_10000_6994, w_10000_6995, w_10000_6996, w_10000_6997, w_10000_6998, w_10000_6999, w_10000_7000, w_10000_7001, w_10000_7002, w_10000_7003, w_10000_7004, w_10000_7005, w_10000_7006, w_10000_7007, w_10000_7008, w_10000_7009, w_10000_7010, w_10000_7011, w_10000_7012, w_10000_7013, w_10000_7014, w_10000_7015, w_10000_7016, w_10000_7017, w_10000_7018, w_10000_7019, w_10000_7020, w_10000_7021, w_10000_7022, w_10000_7023, w_10000_7024, w_10000_7025, w_10000_7026, w_10000_7027, w_10000_7028, w_10000_7029, w_10000_7030, w_10000_7031, w_10000_7032, w_10000_7033, w_10000_7034, w_10000_7035, w_10000_7036, w_10000_7037, w_10000_7038, w_10000_7039, w_10000_7040, w_10000_7041, w_10000_7042, w_10000_7043, w_10000_7044, w_10000_7045, w_10000_7046, w_10000_7047, w_10000_7048, w_10000_7049, w_10000_7050, w_10000_7051, w_10000_7052, w_10000_7053, w_10000_7054, w_10000_7055, w_10000_7056, w_10000_7057, w_10000_7058, w_10000_7059, w_10000_7060, w_10000_7061, w_10000_7062, w_10000_7063, w_10000_7064, w_10000_7065, w_10000_7066, w_10000_7067, w_10000_7068, w_10000_7069, w_10000_7070, w_10000_7071, w_10000_7072, w_10000_7073, w_10000_7074, w_10000_7075, w_10000_7076, w_10000_7077, w_10000_7078, w_10000_7079, w_10000_7080, w_10000_7081, w_10000_7082, w_10000_7083, w_10000_7084, w_10000_7085, w_10000_7086, w_10000_7087, w_10000_7088, w_10000_7089, w_10000_7090, w_10000_7091, w_10000_7092, w_10000_7093, w_10000_7094, w_10000_7095, w_10000_7096, w_10000_7097, w_10000_7098, w_10000_7099, w_10000_7100, w_10000_7101, w_10000_7102, w_10000_7103, w_10000_7104, w_10000_7105, w_10000_7106, w_10000_7107, w_10000_7108, w_10000_7109, w_10000_7110, w_10000_7111, w_10000_7112, w_10000_7113, w_10000_7114, w_10000_7115, w_10000_7116, w_10000_7117, w_10000_7118, w_10000_7119, w_10000_7120, w_10000_7121, w_10000_7122, w_10000_7123, w_10000_7124, w_10000_7125, w_10000_7126, w_10000_7127, w_10000_7128, w_10000_7129, w_10000_7130, w_10000_7131, w_10000_7132, w_10000_7133, w_10000_7134, w_10000_7135, w_10000_7136, w_10000_7137, w_10000_7138, w_10000_7139, w_10000_7140, w_10000_7141, w_10000_7142, w_10000_7143, w_10000_7144, w_10000_7145, w_10000_7146, w_10000_7147, w_10000_7148, w_10000_7149, w_10000_7150, w_10000_7151, w_10000_7152, w_10000_7153, w_10000_7154, w_10000_7155, w_10000_7156, w_10000_7157, w_10000_7158, w_10000_7159, w_10000_7160, w_10000_7161, w_10000_7162, w_10000_7163, w_10000_7164, w_10000_7165, w_10000_7166, w_10000_7167, w_10000_7168, w_10000_7169, w_10000_7170, w_10000_7171, w_10000_7172, w_10000_7173, w_10000_7174, w_10000_7175, w_10000_7176, w_10000_7177, w_10000_7178, w_10000_7179, w_10000_7180, w_10000_7181, w_10000_7182, w_10000_7183, w_10000_7184, w_10000_7185, w_10000_7186, w_10000_7187, w_10000_7188, w_10000_7189, w_10000_7190, w_10000_7191, w_10000_7192, w_10000_7193, w_10000_7194, w_10000_7195, w_10000_7196, w_10000_7197, w_10000_7198, w_10000_7199, w_10000_7200, w_10000_7201, w_10000_7202, w_10000_7203, w_10000_7204, w_10000_7205, w_10000_7206, w_10000_7207, w_10000_7208, w_10000_7209, w_10000_7210, w_10000_7211, w_10000_7212, w_10000_7213, w_10000_7214, w_10000_7215, w_10000_7216, w_10000_7217, w_10000_7218, w_10000_7219, w_10000_7220, w_10000_7221, w_10000_7222, w_10000_7223, w_10000_7224, w_10000_7225, w_10000_7226, w_10000_7227, w_10000_7228, w_10000_7229, w_10000_7230, w_10000_7231, w_10000_7232, w_10000_7233, w_10000_7234, w_10000_7235, w_10000_7236, w_10000_7237, w_10000_7238, w_10000_7239, w_10000_7240, w_10000_7241, w_10000_7242, w_10000_7243, w_10000_7244, w_10000_7245, w_10000_7246, w_10000_7247, w_10000_7248, w_10000_7249, w_10000_7250, w_10000_7251, w_10000_7252, w_10000_7253, w_10000_7254, w_10000_7255, w_10000_7256, w_10000_7257, w_10000_7258, w_10000_7259, w_10000_7260, w_10000_7261, w_10000_7262, w_10000_7263, w_10000_7264, w_10000_7265, w_10000_7266, w_10000_7267, w_10000_7268, w_10000_7269, w_10000_7270, w_10000_7271, w_10000_7272, w_10000_7273, w_10000_7274, w_10000_7275, w_10000_7276, w_10000_7277, w_10000_7278, w_10000_7279, w_10000_7280, w_10000_7281, w_10000_7282, w_10000_7283, w_10000_7284, w_10000_7285, w_10000_7286, w_10000_7287, w_10000_7288 );
  inout w_000_000, w_000_001, w_000_002, w_000_003, w_000_004, w_000_005, w_000_006, w_000_007, w_000_008, w_000_009, w_000_010, w_000_011, w_000_012, w_000_013, w_000_014, w_000_015, w_000_016, w_000_017, w_000_018, w_000_019, w_000_020, w_000_021, w_000_022, w_000_023, w_000_024, w_000_025, w_000_026, w_000_027, w_000_028, w_000_029, w_000_030, w_000_031, w_000_032, w_000_033, w_000_034, w_000_035, w_000_036, w_000_037, w_000_038, w_000_039, w_000_040, w_000_041, w_000_042, w_000_043, w_000_044, w_000_045, w_000_046, w_000_047, w_000_048, w_000_049, w_000_050, w_000_051, w_000_052, w_000_053, w_000_054, w_000_055, w_000_056, w_000_057, w_000_058, w_000_059, w_000_060, w_000_061, w_000_062, w_000_063, w_000_064, w_000_065, w_000_066, w_000_067, w_000_068, w_000_069, w_000_070, w_000_071, w_000_072, w_000_073, w_000_074, w_000_075, w_000_076, w_000_077, w_000_078, w_000_079, w_000_080, w_000_081, w_000_082, w_000_083, w_000_084, w_000_085, w_000_086, w_000_087, w_000_088, w_000_089, w_000_090, w_000_091, w_000_092, w_000_093, w_000_094, w_000_095, w_000_096, w_000_097, w_000_098, w_000_099, w_000_100, w_000_101, w_000_102, w_000_103, w_000_104, w_000_105, w_000_106, w_000_107, w_000_108, w_000_109, w_000_110, w_000_111, w_000_112, w_000_113, w_000_114, w_000_115, w_000_116, w_000_117, w_000_118, w_000_119, w_000_120, w_000_121, w_000_122, w_000_123, w_000_124, w_000_125, w_000_126, w_000_127, w_000_128, w_000_129, w_000_130, w_000_131, w_000_132, w_000_133, w_000_134, w_000_135, w_000_136, w_000_137, w_000_138, w_000_139, w_000_140, w_000_141, w_000_142, w_000_143, w_000_144, w_000_145, w_000_146, w_000_147, w_000_148, w_000_149, w_000_150, w_000_151, w_000_152, w_000_153, w_000_154, w_000_155, w_000_156, w_000_157, w_000_158, w_000_159, w_000_160, w_000_161, w_000_162, w_000_163, w_000_164, w_000_165, w_000_166, w_000_167, w_000_168, w_000_169, w_000_170, w_000_171, w_000_172, w_000_173, w_000_174, w_000_175, w_000_176, w_000_177, w_000_178, w_000_179, w_000_180, w_000_181, w_000_182, w_000_183, w_000_184, w_000_185, w_000_186, w_000_187, w_000_188, w_000_189, w_000_190, w_000_191, w_000_192, w_000_193, w_000_194, w_000_195, w_000_196, w_000_197, w_000_198, w_000_199, w_000_200, w_000_201, w_000_202, w_000_203, w_000_204, w_000_205, w_000_206, w_000_207, w_000_208, w_000_209, w_000_210, w_000_211, w_000_212, w_000_213, w_000_214, w_000_215, w_000_216, w_000_217, w_000_218, w_000_219, w_000_220, w_000_221, w_000_222, w_000_223, w_000_224, w_000_225, w_000_226, w_000_227, w_000_228, w_000_229, w_000_230, w_000_231, w_000_232, w_000_233, w_000_234, w_000_235, w_000_236, w_000_237, w_000_238, w_000_239, w_000_240, w_000_241, w_000_242, w_000_243, w_000_244, w_000_245, w_000_246, w_000_247, w_000_248, w_000_249, w_000_250, w_000_251, w_000_252, w_000_253, w_000_254, w_000_255, w_000_256, w_000_257, w_000_258, w_000_259, w_000_260, w_000_261, w_000_262, w_000_263, w_000_264, w_000_265, w_000_266, w_000_267, w_000_268, w_000_269, w_000_270, w_000_271, w_000_272, w_000_273, w_000_274, w_000_275, w_000_276, w_000_277, w_000_278, w_000_279, w_000_280, w_000_281, w_000_282, w_000_283, w_000_284, w_000_285, w_000_286, w_000_287, w_000_288, w_000_289, w_000_290, w_000_291, w_000_292, w_000_293, w_000_294, w_000_295, w_000_296, w_000_297, w_000_298, w_000_299, w_000_300, w_000_301, w_000_302, w_000_303, w_000_304, w_000_305, w_000_306, w_000_307, w_000_308, w_000_309, w_000_310, w_000_311, w_000_312, w_000_313, w_000_314, w_000_315, w_000_316, w_000_317, w_000_318, w_000_319, w_000_320, w_000_321, w_000_322, w_000_323, w_000_324, w_000_325, w_000_326, w_000_327, w_000_328, w_000_329, w_000_330, w_000_331, w_000_332, w_000_333, w_000_334, w_000_335, w_000_336, w_000_337, w_000_338, w_000_339, w_000_340, w_000_341, w_000_342, w_000_343, w_000_344, w_000_345, w_000_346, w_000_347, w_000_348, w_000_349, w_000_350, w_000_351, w_000_352, w_000_353, w_000_354, w_000_355, w_000_356, w_000_357, w_000_358, w_000_359, w_000_360, w_000_361, w_000_362, w_000_363, w_000_364, w_000_365, w_000_366, w_000_367, w_000_368, w_000_369, w_000_370, w_000_371, w_000_372, w_000_373, w_000_374, w_000_375, w_000_376, w_000_377, w_000_378, w_000_379, w_000_380, w_000_381, w_000_382, w_000_383, w_000_384, w_000_385, w_000_386, w_000_387, w_000_388, w_000_389, w_000_390, w_000_391, w_000_392, w_000_393, w_000_394, w_000_395, w_000_396, w_000_397, w_000_398, w_000_399, w_000_400, w_000_401, w_000_402, w_000_403, w_000_404, w_000_405, w_000_406, w_000_407, w_000_408, w_000_409, w_000_410, w_000_411, w_000_412, w_000_413, w_000_414, w_000_415, w_000_416, w_000_417, w_000_418, w_000_419, w_000_420, w_000_421, w_000_422, w_000_423, w_000_424, w_000_425, w_000_426, w_000_427, w_000_428, w_000_429, w_000_430, w_000_431, w_000_432, w_000_433, w_000_434, w_000_435, w_000_436, w_000_437, w_000_438, w_000_439, w_000_440, w_000_441, w_000_442, w_000_443, w_000_444, w_000_445, w_000_446, w_000_447, w_000_448, w_000_449, w_000_450, w_000_451, w_000_452, w_000_453, w_000_454, w_000_455, w_000_456, w_000_457, w_000_458, w_000_459, w_000_460, w_000_461, w_000_462, w_000_463, w_000_464, w_000_465, w_000_466, w_000_467, w_000_468, w_000_469, w_000_470, w_000_471, w_000_472, w_000_473, w_000_474, w_000_475, w_000_476, w_000_477, w_000_478, w_000_479, w_000_480, w_000_481, w_000_482, w_000_483, w_000_484, w_000_485, w_000_486, w_000_487, w_000_488, w_000_489, w_000_490, w_000_491, w_000_492, w_000_493, w_000_494, w_000_495, w_000_496, w_000_497, w_000_498, w_000_499, w_000_500, w_000_501, w_000_502, w_000_503, w_000_504, w_000_505, w_000_506, w_000_507, w_000_508, w_000_509, w_000_510, w_000_511, w_000_512, w_000_513, w_000_514, w_000_515, w_000_516, w_000_517, w_000_518, w_000_519, w_000_520, w_000_521, w_000_522, w_000_523, w_000_524, w_000_525, w_000_526, w_000_527, w_000_528, w_000_529, w_000_530, w_000_531, w_000_532, w_000_533, w_000_534, w_000_535, w_000_536, w_000_537, w_000_538, w_000_539, w_000_540, w_000_541, w_000_542, w_000_543, w_000_544, w_000_545, w_000_546, w_000_547, w_000_548, w_000_549, w_000_550, w_000_551, w_000_552, w_000_553, w_000_554, w_000_555, w_000_556, w_000_557, w_000_558, w_000_559, w_000_560, w_000_561, w_000_562, w_000_563, w_000_564, w_000_565, w_000_566, w_000_567, w_000_568, w_000_569, w_000_570, w_000_571, w_000_572, w_000_573, w_000_574, w_000_575, w_000_576, w_000_577, w_000_578, w_000_579, w_000_580, w_000_581, w_000_582, w_000_583, w_000_584, w_000_585, w_000_586, w_000_587, w_000_588, w_000_589, w_000_590, w_000_591, w_000_592, w_000_593, w_000_594, w_000_595, w_000_596, w_000_597, w_000_598, w_000_599, w_000_600, w_000_601, w_000_602, w_000_603, w_000_604, w_000_605, w_000_606, w_000_607, w_000_608, w_000_609, w_000_610, w_000_611, w_000_612, w_000_613, w_000_614, w_000_615, w_000_616, w_000_617, w_000_618, w_000_619, w_000_620, w_000_621, w_000_622, w_000_623, w_000_624, w_000_625, w_000_626, w_000_627, w_000_628, w_000_629, w_000_630, w_000_631, w_000_632, w_000_633, w_000_634, w_000_635, w_000_636, w_000_637, w_000_638, w_000_639, w_000_640, w_000_641, w_000_642, w_000_643, w_000_644, w_000_645, w_000_646, w_000_647, w_000_648, w_000_649, w_000_650, w_000_651, w_000_652, w_000_653, w_000_654, w_000_655, w_000_656, w_000_657, w_000_658, w_000_659, w_000_660, w_000_661, w_000_662, w_000_663, w_000_664, w_000_665, w_000_666, w_000_667, w_000_668, w_000_669, w_000_670, w_000_671, w_000_672, w_000_673, w_000_674, w_000_675, w_000_676, w_000_677, w_000_678, w_000_679, w_000_680, w_000_681, w_000_682, w_000_683, w_000_684, w_000_685, w_000_686, w_000_687, w_000_688, w_000_689, w_000_690, w_000_691, w_000_692, w_000_693, w_000_694, w_000_695, w_000_696, w_000_697, w_000_698, w_000_699, w_000_700, w_000_701, w_000_702, w_000_703, w_000_704, w_000_705, w_000_706, w_000_707, w_000_708, w_000_709, w_000_710, w_000_711, w_000_712, w_000_713, w_000_714, w_000_715, w_000_716, w_000_717, w_000_718, w_000_719, w_000_720, w_000_721, w_000_722, w_000_723, w_000_724, w_000_725, w_000_726, w_000_727, w_000_728, w_000_729, w_000_730, w_000_731, w_000_732, w_000_733, w_000_734, w_000_735, w_000_736, w_000_737, w_000_738, w_000_739, w_000_740, w_000_741, w_000_742, w_000_743, w_000_744, w_000_745, w_000_746, w_000_747, w_000_748, w_000_749, w_000_750, w_000_751, w_000_752, w_000_753, w_000_754, w_000_755, w_000_756, w_000_757, w_000_758, w_000_759, w_000_760, w_000_761, w_000_762, w_000_763, w_000_764, w_000_765, w_000_766, w_000_767, w_000_768, w_000_769, w_000_770, w_000_771, w_000_772, w_000_773, w_000_774, w_000_775, w_000_776, w_000_777, w_000_778, w_000_779, w_000_780, w_000_781, w_000_782, w_000_783, w_000_784, w_000_785, w_000_786, w_000_787, w_000_788, w_000_789, w_000_790, w_000_791, w_000_792, w_000_793, w_000_794, w_000_795, w_000_796, w_000_797, w_000_798, w_000_799, w_000_800, w_000_801, w_000_802, w_000_803, w_000_804, w_000_805, w_000_806, w_000_807, w_000_808, w_000_809, w_000_810, w_000_811, w_000_812, w_000_813, w_000_814, w_000_815, w_000_816, w_000_817, w_000_818, w_000_819, w_000_820, w_000_821, w_000_822, w_000_823, w_000_824, w_000_825, w_000_826, w_000_827, w_000_828, w_000_829, w_000_830, w_000_831, w_000_832, w_000_833, w_000_834, w_000_835, w_000_836, w_000_837, w_000_838, w_000_839, w_000_840, w_000_841, w_000_842, w_000_843, w_000_844, w_000_845, w_000_846, w_000_847, w_000_848, w_000_849, w_000_850, w_000_851, w_000_852, w_000_853, w_000_854, w_000_855, w_000_856, w_000_857, w_000_858, w_000_859, w_000_860, w_000_861, w_000_862, w_000_863, w_000_864, w_000_865, w_000_866, w_000_867, w_000_868, w_000_869, w_000_870, w_000_871, w_000_872, w_000_873, w_000_874, w_000_875, w_000_876, w_000_877, w_000_878, w_000_879, w_000_880, w_000_881, w_000_882, w_000_883, w_000_884, w_000_885, w_000_886, w_000_887, w_000_888, w_000_889, w_000_890, w_000_891, w_000_892, w_000_893, w_000_894, w_000_895, w_000_896, w_000_897, w_000_898, w_000_899, w_000_900, w_000_901, w_000_902, w_000_903, w_000_904, w_000_905, w_000_906, w_000_907, w_000_908, w_000_909, w_000_910, w_000_911, w_000_912, w_000_913, w_000_914, w_000_915, w_000_916, w_000_917, w_000_918, w_000_919, w_000_920, w_000_921, w_000_922, w_000_923, w_000_924, w_000_925, w_000_926, w_000_927, w_000_928, w_000_929, w_000_930, w_000_931, w_000_932, w_000_933, w_000_934, w_000_935, w_000_936, w_000_937, w_000_938, w_000_939, w_000_940, w_000_941, w_000_942, w_000_943, w_000_944, w_000_945, w_000_946, w_000_947, w_000_948, w_000_949, w_000_950, w_000_951, w_000_952, w_000_953, w_000_954, w_000_955, w_000_956, w_000_957, w_000_958, w_000_959, w_000_960, w_000_961, w_000_962, w_000_963, w_000_964, w_000_965, w_000_966, w_000_967, w_000_968, w_000_969, w_000_970, w_000_971, w_000_972, w_000_973, w_000_974, w_000_975, w_000_976, w_000_977, w_000_978, w_000_979, w_000_980, w_000_981, w_000_982, w_000_983, w_000_984, w_000_985, w_000_986, w_000_987, w_000_988, w_000_989, w_000_990, w_000_991, w_000_992, w_000_993, w_000_994, w_000_995, w_000_996, w_000_997, w_000_998, w_000_999, w_000_1000, w_000_1001, w_000_1002, w_000_1003, w_000_1004, w_000_1005, w_000_1006, w_000_1007, w_000_1008, w_000_1009, w_000_1010, w_000_1011, w_000_1012, w_000_1013, w_000_1014, w_000_1015, w_000_1016, w_000_1017, w_000_1018, w_000_1019, w_000_1020, w_000_1021, w_000_1022, w_000_1023, w_000_1024, w_000_1025, w_000_1026, w_000_1027, w_000_1028, w_000_1029, w_000_1030, w_000_1031, w_000_1032, w_000_1033, w_000_1034, w_000_1035, w_000_1036, w_000_1037, w_000_1038, w_000_1039, w_000_1040, w_000_1041, w_000_1042, w_000_1043, w_000_1044, w_000_1045, w_000_1046, w_000_1047, w_000_1048, w_000_1049, w_000_1050, w_000_1051, w_000_1052, w_000_1053, w_000_1054, w_000_1055, w_000_1056, w_000_1057, w_000_1058, w_000_1059, w_000_1060, w_000_1061, w_000_1062, w_000_1063, w_000_1064, w_000_1065, w_000_1066, w_000_1067, w_000_1068, w_000_1069, w_000_1070, w_000_1071, w_000_1072, w_000_1073, w_000_1074, w_000_1075, w_000_1076, w_000_1077, w_000_1078, w_000_1079, w_000_1080, w_000_1081, w_000_1082, w_000_1083, w_000_1084, w_000_1085, w_000_1086, w_000_1087, w_000_1088, w_000_1089, w_000_1090, w_000_1091, w_000_1092, w_000_1093, w_000_1094, w_000_1095, w_000_1096, w_000_1097, w_000_1098, w_000_1099, w_000_1100, w_000_1101, w_000_1102, w_000_1103, w_000_1104, w_000_1105, w_000_1106, w_000_1107, w_000_1108, w_000_1109, w_000_1110, w_000_1111, w_000_1112, w_000_1113, w_000_1114, w_000_1115, w_000_1116, w_000_1117, w_000_1118, w_000_1119, w_000_1120, w_000_1121, w_000_1122, w_000_1123, w_000_1124, w_000_1125, w_000_1126, w_000_1127, w_000_1128, w_000_1129, w_000_1130, w_000_1131, w_000_1132, w_000_1133, w_000_1134, w_000_1135, w_000_1136, w_000_1137, w_000_1138, w_000_1139, w_000_1140, w_000_1141, w_000_1142, w_000_1143, w_000_1144, w_000_1145, w_000_1146, w_000_1147, w_000_1148, w_000_1149, w_000_1150, w_000_1151, w_000_1152, w_000_1153, w_000_1154, w_000_1155, w_000_1156, w_000_1157, w_000_1158, w_000_1159, w_000_1160, w_000_1161, w_000_1162, w_000_1163, w_000_1164, w_000_1165, w_000_1166, w_000_1167, w_000_1168, w_000_1169, w_000_1170, w_000_1171, w_000_1172, w_000_1173, w_000_1174, w_000_1175, w_000_1176, w_000_1177, w_000_1178, w_000_1179, w_000_1180, w_000_1181, w_000_1182, w_000_1183, w_000_1184, w_000_1185, w_000_1186, w_000_1187, w_000_1188, w_000_1189, w_000_1190, w_000_1191, w_000_1192, w_000_1193, w_000_1194, w_000_1195, w_000_1196, w_000_1197, w_000_1198, w_000_1199, w_000_1200, w_000_1201, w_000_1202, w_000_1203, w_000_1204, w_000_1205, w_000_1206, w_000_1207, w_000_1208, w_000_1209, w_000_1210, w_000_1211, w_000_1212, w_000_1213, w_000_1214, w_000_1215, w_000_1216, w_000_1217, w_000_1218, w_000_1219, w_000_1220, w_000_1221, w_000_1222, w_000_1223, w_000_1224, w_000_1225, w_000_1226, w_000_1227, w_000_1228, w_000_1229, w_000_1230, w_000_1231, w_000_1232, w_000_1233, w_000_1234, w_000_1235, w_000_1236, w_000_1237, w_000_1238, w_000_1239, w_000_1240, w_000_1241, w_000_1242, w_000_1243, w_000_1244, w_000_1245, w_000_1246, w_000_1247, w_000_1248, w_000_1249, w_000_1250, w_000_1251, w_000_1252, w_000_1253, w_000_1254, w_000_1255, w_000_1256, w_000_1257, w_000_1258, w_000_1259, w_000_1260, w_000_1261, w_000_1262, w_000_1263, w_000_1264, w_000_1265, w_000_1266, w_000_1267, w_000_1268, w_000_1269, w_000_1270, w_000_1271, w_000_1272, w_000_1273, w_000_1274, w_000_1275, w_000_1276, w_000_1277, w_000_1278, w_000_1279, w_000_1280, w_000_1281, w_000_1282, w_000_1283, w_000_1284, w_000_1285, w_000_1286, w_000_1287, w_000_1288, w_000_1289, w_000_1290, w_000_1291, w_000_1292, w_000_1293, w_000_1294, w_000_1295, w_000_1296, w_000_1297, w_000_1298, w_000_1299, w_000_1300, w_000_1301, w_000_1302, w_000_1303, w_000_1304, w_000_1305, w_000_1306, w_000_1307, w_000_1308, w_000_1309, w_000_1310, w_000_1311, w_000_1312, w_000_1313, w_000_1314, w_000_1315, w_000_1316, w_000_1317, w_000_1318, w_000_1319, w_000_1320, w_000_1321, w_000_1322, w_000_1323, w_000_1324, w_000_1325, w_000_1326, w_000_1327, w_000_1328, w_000_1329, w_000_1330, w_000_1331, w_000_1332, w_000_1333, w_000_1334, w_000_1335, w_000_1336, w_000_1337, w_000_1338, w_000_1339, w_000_1340, w_000_1341, w_000_1342, w_000_1343, w_000_1344, w_000_1345, w_000_1346, w_000_1347, w_000_1348, w_000_1349, w_000_1350, w_000_1351, w_000_1352, w_000_1353, w_000_1354, w_000_1355, w_000_1356, w_000_1357, w_000_1358, w_000_1359, w_000_1360, w_000_1361, w_000_1362, w_000_1363, w_000_1364, w_000_1365, w_000_1366, w_000_1367, w_000_1368, w_000_1369, w_000_1370, w_000_1371, w_000_1372, w_000_1373, w_000_1374, w_000_1375, w_000_1376, w_000_1377, w_000_1378, w_000_1379, w_000_1380, w_000_1381, w_000_1382, w_000_1383, w_000_1384, w_000_1385, w_000_1386, w_000_1387, w_000_1388, w_000_1389, w_000_1390, w_000_1391, w_000_1392, w_000_1393, w_000_1394, w_000_1395, w_000_1396, w_000_1397, w_000_1398, w_000_1399, w_000_1400, w_000_1401, w_000_1402, w_000_1403, w_000_1404, w_000_1405, w_000_1406, w_000_1407, w_000_1408, w_000_1409, w_000_1410, w_000_1411, w_000_1412, w_000_1413, w_000_1414, w_000_1415, w_000_1416, w_000_1417, w_000_1418, w_000_1419, w_000_1420, w_000_1421, w_000_1422, w_000_1423, w_000_1424, w_000_1425, w_000_1426, w_000_1427, w_000_1428, w_000_1429, w_000_1430, w_000_1431, w_000_1432, w_000_1433, w_000_1434, w_000_1435, w_000_1436, w_000_1437, w_000_1438, w_000_1439, w_000_1440, w_000_1441, w_000_1442, w_000_1443, w_000_1444, w_000_1445, w_000_1446, w_000_1447, w_000_1448, w_000_1449, w_000_1450, w_000_1451, w_000_1452, w_000_1453, w_000_1454, w_000_1455, w_000_1456, w_000_1457, w_000_1458, w_000_1459, w_000_1460, w_000_1461, w_000_1462, w_000_1463, w_000_1464, w_000_1465, w_000_1466, w_000_1467, w_000_1468, w_000_1469, w_000_1470, w_000_1471, w_000_1472, w_000_1473, w_000_1474, w_000_1475, w_000_1476, w_000_1477, w_000_1478, w_000_1479, w_000_1480, w_000_1481, w_000_1482, w_000_1483, w_000_1484, w_000_1485, w_000_1486, w_000_1487, w_000_1488, w_000_1489, w_000_1490, w_000_1491, w_000_1492, w_000_1493, w_000_1494, w_000_1495, w_000_1496, w_000_1497, w_000_1498, w_000_1499, w_000_1500, w_000_1501, w_000_1502, w_000_1503, w_000_1504, w_000_1505, w_000_1506, w_000_1507, w_000_1508, w_000_1509, w_000_1510, w_000_1511, w_000_1512, w_000_1513, w_000_1514, w_000_1515, w_000_1516, w_000_1517, w_000_1518, w_000_1519, w_000_1520, w_000_1521, w_000_1522, w_000_1523, w_000_1524, w_000_1525, w_000_1526, w_000_1527, w_000_1528, w_000_1529, w_000_1530, w_000_1531, w_000_1532, w_000_1533, w_000_1534, w_000_1535, w_000_1536, w_000_1537, w_000_1538, w_000_1539, w_000_1540, w_000_1541, w_000_1542, w_000_1543, w_000_1544, w_000_1545, w_000_1546, w_000_1547, w_000_1548, w_000_1549, w_000_1550, w_000_1551, w_000_1552, w_000_1553, w_000_1554, w_000_1555, w_000_1556, w_000_1557, w_000_1558, w_000_1559, w_000_1560, w_000_1561, w_000_1562, w_000_1563, w_000_1564, w_000_1565, w_000_1566, w_000_1567, w_000_1568, w_000_1569, w_000_1570, w_000_1571, w_000_1572, w_000_1573, w_000_1574, w_000_1575, w_000_1576, w_000_1577, w_000_1578, w_000_1579, w_000_1580, w_000_1581, w_000_1582, w_000_1583, w_000_1584, w_000_1585, w_000_1586, w_000_1587, w_000_1588, w_000_1589, w_000_1590, w_000_1591, w_000_1592, w_000_1593, w_000_1594, w_000_1595, w_000_1596, w_000_1597, w_000_1598, w_000_1599, w_000_1600, w_000_1601, w_000_1602, w_000_1603, w_000_1604, w_000_1605, w_000_1606, w_000_1607, w_000_1608, w_000_1609, w_000_1610, w_000_1611, w_000_1612, w_000_1613, w_000_1614, w_000_1615, w_000_1616, w_000_1617, w_000_1618, w_000_1619, w_000_1620, w_000_1621, w_000_1622, w_000_1623, w_000_1624, w_000_1625, w_000_1626, w_000_1627, w_000_1628, w_000_1629, w_000_1630, w_000_1631, w_000_1632, w_000_1633, w_000_1634, w_000_1635, w_000_1636, w_000_1637, w_000_1638, w_000_1639, w_000_1640, w_000_1641, w_000_1642, w_000_1643, w_000_1644, w_000_1645, w_000_1646, w_000_1647, w_000_1648, w_000_1649, w_000_1650, w_000_1651, w_000_1652, w_000_1653, w_000_1654, w_000_1655, w_000_1656, w_000_1657, w_000_1658, w_000_1659, w_000_1660, w_000_1661, w_000_1662, w_000_1663, w_000_1664, w_000_1665, w_000_1666, w_000_1667, w_000_1668, w_000_1669, w_000_1670, w_000_1671, w_000_1672, w_000_1673, w_000_1674, w_000_1675, w_000_1676, w_000_1677, w_000_1678, w_000_1679, w_000_1680, w_000_1681, w_000_1682, w_000_1683, w_000_1684, w_000_1685, w_000_1686, w_000_1687, w_000_1688, w_000_1689, w_000_1690, w_000_1691, w_000_1692, w_000_1693, w_000_1694, w_000_1695, w_000_1696, w_000_1697, w_000_1698, w_000_1699, w_000_1700, w_000_1701, w_000_1702, w_000_1703, w_000_1704, w_000_1705, w_000_1706, w_000_1707, w_000_1708, w_000_1709, w_000_1710, w_000_1711, w_000_1712, w_000_1713, w_000_1714, w_000_1715, w_000_1716, w_000_1717, w_000_1718, w_000_1719, w_000_1720, w_000_1721, w_000_1722, w_000_1723, w_000_1724, w_000_1725, w_000_1726, w_000_1727, w_000_1728, w_000_1729, w_000_1730, w_000_1731, w_000_1732, w_000_1733, w_000_1734, w_000_1735, w_000_1736, w_000_1737, w_000_1738, w_000_1739, w_000_1740, w_000_1741, w_000_1742, w_000_1743, w_000_1744, w_000_1745, w_000_1746, w_000_1747, w_000_1748, w_000_1749, w_000_1750, w_000_1751, w_000_1752, w_000_1753, w_000_1754, w_000_1755, w_000_1756, w_000_1757, w_000_1758, w_000_1759, w_000_1760, w_000_1761, w_000_1762, w_000_1763, w_000_1764, w_000_1765, w_000_1766, w_000_1767, w_000_1768, w_000_1769, w_000_1770, w_000_1771, w_000_1772, w_000_1773, w_000_1774, w_000_1775, w_000_1776, w_000_1777, w_000_1778, w_000_1779, w_000_1780, w_000_1781, w_000_1782, w_000_1783, w_000_1784, w_000_1785, w_000_1786, w_000_1787, w_000_1788, w_000_1789, w_000_1790, w_000_1791, w_000_1792, w_000_1793, w_000_1794, w_000_1795, w_000_1796, w_000_1797, w_000_1798, w_000_1799, w_000_1800, w_000_1801, w_000_1802, w_000_1803, w_000_1804, w_000_1805, w_000_1806, w_000_1807, w_000_1808, w_000_1809, w_000_1810, w_000_1811, w_000_1812, w_000_1813, w_000_1814, w_000_1815, w_000_1816, w_000_1817, w_000_1818, w_000_1819, w_000_1820, w_000_1821, w_000_1822, w_000_1823, w_000_1824, w_000_1825, w_000_1826, w_000_1827, w_000_1828, w_000_1829, w_000_1830, w_000_1831, w_000_1832, w_000_1833, w_000_1834, w_000_1835, w_000_1836, w_000_1837, w_000_1838, w_000_1839, w_000_1840, w_000_1841, w_000_1842, w_000_1843, w_000_1844, w_000_1845, w_000_1846, w_000_1847, w_000_1848, w_000_1849, w_000_1850, w_000_1851, w_000_1852, w_000_1853, w_000_1854, w_000_1855, w_000_1856, w_000_1857, w_000_1858, w_000_1859, w_000_1860, w_000_1861, w_000_1862, w_000_1863, w_000_1864, w_000_1865, w_000_1866, w_000_1867, w_000_1868, w_000_1869, w_000_1870, w_000_1871, w_000_1872, w_000_1873, w_000_1874, w_000_1875, w_000_1876, w_000_1877, w_000_1878, w_000_1879, w_000_1880, w_000_1881, w_000_1882, w_000_1883, w_000_1884, w_000_1885, w_000_1886, w_000_1887, w_000_1888, w_000_1889, w_000_1890, w_000_1891, w_000_1892, w_000_1893, w_000_1894, w_000_1895, w_000_1896, w_000_1897, w_000_1898, w_000_1899, w_000_1900, w_000_1901, w_000_1902, w_000_1903, w_000_1904, w_000_1905, w_000_1906, w_000_1907, w_000_1908, w_000_1909, w_000_1910, w_000_1911, w_000_1912, w_000_1913, w_000_1914, w_000_1915, w_000_1916, w_000_1917, w_000_1918, w_000_1919, w_000_1920, w_000_1921, w_000_1922, w_000_1923, w_000_1924, w_000_1925, w_000_1926, w_000_1927, w_000_1928, w_000_1929, w_000_1930, w_000_1931, w_000_1932, w_000_1933, w_000_1934, w_000_1935, w_000_1936, w_000_1937, w_000_1938, w_000_1939, w_000_1940, w_000_1941, w_000_1942, w_000_1943, w_000_1944, w_000_1945, w_000_1946, w_000_1947, w_000_1948, w_000_1949, w_000_1950, w_000_1951, w_000_1952, w_000_1953, w_000_1954, w_000_1955, w_000_1956, w_000_1957, w_000_1958, w_000_1959, w_000_1960, w_000_1961, w_000_1962, w_000_1963, w_000_1964, w_000_1965, w_000_1966, w_000_1967, w_000_1968, w_000_1969, w_000_1970, w_000_1971, w_000_1972, w_000_1973, w_000_1974, w_000_1975, w_000_1976, w_000_1977, w_000_1978, w_000_1979, w_000_1980, w_000_1981, w_000_1982, w_000_1983, w_000_1984, w_000_1985, w_000_1986, w_000_1987, w_000_1988, w_000_1989, w_000_1990, w_000_1991, w_000_1992, w_000_1993, w_000_1994, w_000_1995, w_000_1996, w_000_1997, w_000_1998, w_000_1999, w_000_2000, w_000_2001, w_000_2002, w_000_2003, w_000_2004, w_000_2005, w_000_2006, w_000_2007, w_000_2008, w_000_2009, w_000_2010, w_000_2011, w_000_2012, w_000_2013, w_000_2014, w_000_2015, w_000_2016, w_000_2017, w_000_2018, w_000_2019, w_000_2020, w_000_2021, w_000_2022, w_000_2023, w_000_2024, w_000_2025, w_000_2026, w_000_2027, w_000_2028, w_000_2029, w_000_2030, w_000_2031, w_000_2032, w_000_2033, w_000_2034, w_000_2035, w_000_2036, w_000_2037, w_000_2038, w_000_2039, w_000_2040, w_000_2041, w_000_2042, w_000_2043, w_000_2044, w_000_2045, w_000_2046, w_000_2047, w_000_2048, w_000_2049, w_000_2050, w_000_2051, w_000_2052, w_000_2053, w_000_2054, w_000_2055, w_000_2056, w_000_2057, w_000_2058, w_000_2059, w_000_2060, w_000_2061, w_000_2062, w_000_2063, w_000_2064, w_000_2065, w_000_2066, w_000_2067, w_000_2068, w_000_2069, w_000_2070, w_000_2071, w_000_2072, w_000_2073, w_000_2074, w_000_2075, w_000_2076, w_000_2077, w_000_2078, w_000_2079, w_000_2080, w_000_2081, w_000_2082, w_000_2083, w_000_2084, w_000_2085, w_000_2086, w_000_2087, w_000_2088, w_000_2089, w_000_2090, w_000_2091, w_000_2092, w_000_2093, w_000_2094, w_000_2095, w_000_2096, w_000_2097, w_000_2098, w_000_2099, w_000_2100, w_000_2101, w_000_2102, w_000_2103, w_000_2104, w_000_2105, w_000_2106, w_000_2107, w_000_2108, w_000_2109, w_000_2110, w_000_2111, w_000_2112, w_000_2113, w_000_2114, w_000_2115, w_000_2116, w_000_2117, w_000_2118, w_000_2119, w_000_2120, w_000_2121, w_000_2122, w_000_2123, w_000_2124, w_000_2125, w_000_2126, w_000_2127, w_000_2128, w_000_2129, w_000_2130, w_000_2131, w_000_2132, w_000_2133, w_000_2134, w_000_2135, w_000_2136, w_000_2137, w_000_2138, w_000_2139, w_000_2140, w_000_2141, w_000_2142, w_000_2143, w_000_2144, w_000_2145, w_000_2146, w_000_2147, w_000_2148, w_000_2149, w_000_2150, w_000_2151, w_000_2152, w_000_2153, w_000_2154, w_000_2155, w_000_2156, w_000_2157, w_000_2158, w_000_2160, w_000_2161, w_000_2162, w_000_2163, w_000_2164, w_000_2165, w_000_2166, w_000_2167, w_000_2168, w_000_2169, w_000_2170, w_000_2171, w_000_2172, w_000_2173, w_000_2174, w_000_2175, w_000_2176, w_000_2177, w_000_2178, w_000_2179, w_000_2180, w_000_2181, w_000_2182, w_000_2183, w_000_2184, w_000_2185, w_000_2186, w_000_2187, w_000_2188, w_000_2189, w_000_2190, w_000_2191, w_000_2192, w_000_2193, w_000_2194, w_000_2195, w_000_2196, w_000_2197, w_000_2198, w_000_2199, w_000_2200, w_000_2201, w_000_2202, w_000_2203, w_000_2204, w_000_2205, w_000_2206, w_000_2207, w_000_2208, w_000_2209, w_000_2210, w_000_2211, w_000_2212, w_000_2213, w_000_2214, w_000_2215, w_000_2216, w_000_2217, w_000_2218, w_000_2219, w_000_2220, w_000_2221, w_000_2222, w_000_2223, w_000_2224, w_000_2225, w_000_2226, w_000_2227, w_000_2228, w_000_2229, w_000_2230, w_000_2231, w_000_2232, w_000_2233, w_000_2234, w_000_2235, w_000_2236, w_000_2237, w_000_2238, w_000_2239, w_000_2240, w_000_2241, w_000_2242, w_000_2243, w_000_2244, w_000_2245, w_000_2246, w_000_2247, w_000_2248, w_000_2249, w_000_2250, w_000_2251, w_000_2252, w_000_2253, w_000_2254, w_000_2255, w_000_2256, w_000_2257, w_000_2258, w_000_2259, w_000_2260, w_000_2261, w_000_2262, w_000_2263, w_000_2264, w_000_2265, w_000_2266, w_000_2267, w_000_2268, w_000_2269, w_000_2270, w_000_2271, w_000_2272, w_000_2273, w_000_2274, w_000_2275, w_000_2276, w_000_2277, w_000_2278, w_000_2279, w_000_2280, w_000_2281, w_000_2282, w_000_2283, w_000_2284, w_000_2285, w_000_2286, w_000_2287, w_000_2288, w_000_2289, w_000_2290, w_000_2291, w_000_2292, w_000_2293, w_000_2294, w_000_2295, w_000_2296, w_000_2297, w_000_2298, w_000_2299, w_000_2300, w_000_2301, w_000_2302, w_000_2303, w_000_2304, w_000_2305, w_000_2306, w_000_2307, w_000_2308, w_000_2309, w_000_2310, w_000_2311, w_000_2312, w_000_2313, w_000_2314, w_000_2315, w_000_2316, w_000_2317, w_000_2318, w_000_2319, w_000_2320, w_000_2321, w_000_2322, w_000_2323, w_000_2324, w_000_2325, w_000_2326, w_000_2327, w_000_2328, w_000_2329, w_000_2330, w_000_2331, w_000_2332, w_000_2333, w_000_2334, w_000_2335, w_000_2336, w_000_2337, w_000_2338, w_000_2339, w_000_2340, w_000_2341, w_000_2342, w_000_2343, w_000_2344, w_000_2345, w_000_2346, w_000_2347, w_000_2348, w_000_2349, w_000_2350, w_000_2351, w_000_2352, w_000_2353, w_000_2354, w_000_2355, w_000_2356, w_000_2357, w_000_2358, w_000_2359, w_000_2360, w_000_2361, w_000_2362, w_000_2363, w_000_2364, w_000_2365, w_000_2366, w_000_2367, w_000_2368, w_000_2369, w_000_2370, w_000_2371, w_000_2372, w_000_2373, w_000_2374, w_000_2375, w_000_2376, w_000_2377, w_000_2378, w_000_2379, w_000_2380, w_000_2381, w_000_2382, w_000_2383, w_000_2384, w_000_2385, w_000_2386, w_000_2387, w_000_2388, w_000_2389, w_000_2390, w_000_2391, w_000_2392, w_000_2393, w_000_2394, w_000_2395, w_000_2396, w_000_2397, w_000_2398, w_000_2399, w_000_2400, w_000_2401, w_000_2402, w_000_2403, w_000_2404, w_000_2405, w_000_2406, w_000_2407, w_000_2408, w_000_2410, w_000_2411, w_000_2412, w_000_2413, w_000_2414, w_000_2415, w_000_2416, w_000_2417, w_000_2418, w_000_2419, w_000_2420, w_000_2421, w_000_2422, w_000_2423, w_000_2424, w_000_2425, w_000_2426, w_000_2427, w_000_2428, w_000_2429, w_000_2430, w_000_2431, w_000_2432, w_000_2433, w_000_2434, w_000_2435, w_000_2436, w_000_2437, w_000_2438, w_000_2439, w_000_2440, w_000_2441, w_000_2442, w_000_2443, w_000_2444, w_000_2445, w_000_2446, w_000_2447, w_000_2448, w_000_2449, w_000_2450, w_000_2451, w_000_2452, w_000_2453, w_000_2454, w_000_2455, w_000_2456, w_000_2457, w_000_2458, w_000_2459, w_000_2460, w_000_2461, w_000_2462, w_000_2463, w_000_2464, w_000_2465, w_000_2466, w_000_2467, w_000_2468, w_000_2469, w_000_2470, w_000_2471, w_000_2472, w_000_2473, w_000_2474, w_000_2475, w_000_2476, w_000_2477, w_000_2478, w_000_2479, w_000_2480, w_000_2481, w_000_2482, w_000_2483, w_000_2484, w_000_2485, w_000_2486, w_000_2487, w_000_2488, w_000_2489, w_000_2490, w_000_2491, w_000_2492, w_000_2493, w_000_2494, w_000_2495, w_000_2496, w_000_2497, w_000_2498, w_000_2499, w_000_2500, w_000_2501, w_000_2502, w_000_2503, w_000_2504, w_000_2505, w_000_2506, w_000_2507, w_000_2508, w_000_2509, w_000_2510, w_000_2511, w_000_2512, w_000_2513, w_000_2514, w_000_2515, w_000_2516, w_000_2517, w_000_2518, w_000_2519, w_000_2520, w_000_2521, w_000_2522, w_000_2523, w_000_2524, w_000_2525, w_000_2526, w_000_2527, w_000_2528, w_000_2529, w_000_2530, w_000_2531, w_000_2532, w_000_2533, w_000_2534, w_000_2535, w_000_2536, w_000_2537, w_000_2538, w_000_2539, w_000_2540, w_000_2541, w_000_2542, w_000_2543, w_000_2544, w_000_2545, w_000_2546, w_000_2547, w_000_2548, w_000_2549, w_000_2550, w_000_2551, w_000_2552, w_000_2553, w_000_2554, w_000_2555, w_000_2556, w_000_2557, w_000_2558, w_000_2559, w_000_2560, w_000_2561, w_000_2562, w_000_2563, w_000_2564, w_000_2565, w_000_2566, w_000_2567, w_000_2568, w_000_2569, w_000_2570, w_000_2571, w_000_2572, w_000_2573, w_000_2574, w_000_2575, w_000_2576, w_000_2577, w_000_2578, w_000_2579, w_000_2580, w_000_2581, w_000_2582, w_000_2583, w_000_2584, w_000_2585, w_000_2586, w_000_2587, w_000_2588, w_000_2589, w_000_2590, w_000_2591, w_000_2592, w_000_2593, w_000_2594, w_000_2595, w_000_2596, w_000_2597, w_000_2598, w_000_2599, w_000_2600, w_000_2601, w_000_2602, w_000_2603, w_000_2604, w_000_2605, w_000_2606, w_000_2607, w_000_2608, w_000_2609, w_000_2610, w_000_2611, w_000_2612, w_000_2613, w_000_2614, w_000_2615, w_000_2616, w_000_2617, w_000_2618, w_000_2619, w_000_2620, w_000_2621, w_000_2622, w_000_2623, w_000_2624, w_000_2625, w_000_2626, w_000_2627, w_000_2628, w_000_2629, w_000_2630, w_000_2631, w_000_2632, w_000_2633, w_000_2634, w_000_2635, w_000_2636, w_000_2637, w_000_2638, w_000_2639, w_000_2640, w_000_2641, w_000_2642, w_000_2643, w_000_2644, w_000_2645, w_000_2646, w_000_2647, w_000_2648, w_000_2649, w_000_2650, w_000_2651, w_000_2652, w_000_2653, w_000_2654, w_000_2655, w_000_2656, w_000_2657, w_000_2658, w_000_2659, w_000_2660, w_000_2661, w_000_2662, w_000_2663, w_000_2664, w_000_2665, w_000_2666, w_000_2667, w_000_2668, w_000_2669, w_000_2670, w_000_2671, w_000_2672, w_000_2673, w_000_2674, w_000_2675, w_000_2676, w_000_2677, w_000_2678, w_000_2679, w_000_2680, w_000_2681, w_000_2682, w_000_2683, w_000_2684, w_000_2685, w_000_2686, w_000_2687, w_000_2688, w_000_2689, w_000_2690, w_000_2691, w_000_2692, w_000_2693, w_000_2694, w_000_2695, w_000_2696, w_000_2697, w_000_2698, w_000_2699, w_000_2700, w_000_2701, w_000_2702, w_000_2703, w_000_2704, w_000_2705, w_000_2706, w_000_2707, w_000_2708, w_000_2709, w_000_2710, w_000_2711, w_000_2712, w_000_2713, w_000_2714, w_000_2715, w_000_2716, w_000_2717, w_000_2718, w_000_2719, w_000_2720, w_000_2721, w_000_2722, w_000_2723, w_000_2724, w_000_2725, w_000_2726, w_000_2727, w_000_2728, w_000_2729, w_000_2730, w_000_2731, w_000_2732, w_000_2733, w_000_2734, w_000_2735, w_000_2736, w_000_2737, w_000_2738, w_000_2739, w_000_2740, w_000_2741, w_000_2742, w_000_2743, w_000_2744, w_000_2745, w_000_2746, w_000_2747, w_000_2748, w_000_2749, w_000_2750, w_000_2751, w_000_2752, w_000_2753, w_000_2754, w_000_2755, w_000_2756, w_000_2757, w_000_2758, w_000_2759, w_000_2760, w_000_2761, w_000_2762, w_000_2763, w_000_2764, w_000_2765, w_000_2766, w_000_2767, w_000_2768, w_000_2769, w_000_2770, w_000_2771, w_000_2772, w_000_2773, w_000_2774, w_000_2775, w_000_2776, w_000_2777, w_000_2778, w_000_2779, w_000_2780, w_000_2781, w_000_2782, w_000_2783, w_000_2784, w_000_2785, w_000_2786, w_000_2787, w_000_2788, w_000_2789, w_000_2790, w_000_2791, w_000_2792, w_000_2793, w_000_2794, w_000_2795, w_000_2796, w_000_2797, w_000_2798, w_000_2799, w_000_2800, w_000_2801, w_000_2802, w_000_2803, w_000_2804, w_000_2805, w_000_2806, w_000_2807, w_000_2808, w_000_2809, w_000_2810, w_000_2811, w_000_2812, w_000_2813, w_000_2814, w_000_2815, w_000_2816, w_000_2817, w_000_2818, w_000_2819, w_000_2820, w_000_2821, w_000_2822, w_000_2823, w_000_2824, w_000_2825, w_000_2826, w_000_2827, w_000_2828, w_000_2829, w_000_2830, w_000_2831, w_000_2832, w_000_2834, w_000_2835, w_000_2836, w_000_2837, w_000_2838, w_000_2839, w_000_2840, w_000_2841, w_000_2842, w_000_2843, w_000_2844, w_000_2845, w_000_2846, w_000_2847, w_000_2848, w_000_2849, w_000_2850, w_000_2851, w_000_2852, w_000_2853, w_000_2854, w_000_2855, w_000_2856, w_000_2857, w_000_2858, w_000_2859, w_000_2860, w_000_2861, w_000_2862, w_000_2863, w_000_2864, w_000_2865, w_000_2866, w_000_2867, w_000_2868, w_000_2869, w_000_2870, w_000_2871, w_000_2872, w_000_2873, w_000_2874, w_000_2875, w_000_2876, w_000_2877, w_000_2878, w_000_2879, w_000_2880, w_000_2881, w_000_2882, w_000_2883, w_000_2884, w_000_2885, w_000_2886, w_000_2887, w_000_2888, w_000_2889, w_000_2890, w_000_2891, w_000_2892, w_000_2893, w_000_2894, w_000_2895, w_000_2896, w_000_2897, w_000_2898, w_000_2899, w_000_2900, w_000_2901, w_000_2902, w_000_2903, w_000_2904, w_000_2905, w_000_2906, w_000_2907, w_000_2908, w_000_2909, w_000_2910, w_000_2911, w_000_2912, w_000_2913, w_000_2914, w_000_2915, w_000_2916, w_000_2917, w_000_2918, w_000_2919, w_000_2920, w_000_2921, w_000_2922, w_000_2923, w_000_2924, w_000_2925, w_000_2926, w_000_2927, w_000_2928, w_000_2929, w_000_2930, w_000_2931, w_000_2932, w_000_2933, w_000_2934, w_000_2935, w_000_2936, w_000_2937, w_000_2938, w_000_2939, w_000_2940, w_000_2941, w_000_2942, w_000_2943, w_000_2944, w_000_2945, w_000_2946, w_000_2947, w_000_2948, w_000_2949, w_000_2950, w_000_2951, w_000_2952, w_000_2953, w_000_2954, w_000_2955, w_000_2956, w_000_2957, w_000_2958, w_000_2959, w_000_2960, w_000_2961, w_000_2962, w_000_2963, w_000_2964, w_000_2965, w_000_2966, w_000_2967, w_000_2968, w_000_2969, w_000_2970, w_000_2971, w_000_2972, w_000_2973, w_000_2974, w_000_2975, w_000_2976, w_000_2977, w_000_2978, w_000_2979, w_000_2980, w_000_2981, w_000_2982, w_000_2983, w_000_2984, w_000_2985, w_000_2986, w_000_2987, w_000_2988, w_000_2989, w_000_2990, w_000_2991, w_000_2992, w_000_2993, w_000_2994, w_000_2995, w_000_2996, w_000_2997, w_000_2998, w_000_2999, w_000_3000, w_000_3001, w_000_3002, w_000_3003, w_000_3004, w_000_3005, w_000_3006, w_000_3007, w_000_3008, w_000_3009, w_000_3010, w_000_3011, w_000_3012, w_000_3013, w_000_3014, w_000_3015, w_000_3016, w_000_3017, w_000_3018, w_000_3019, w_000_3020, w_000_3021, w_000_3022, w_000_3023, w_000_3024, w_000_3025, w_000_3026, w_000_3027, w_000_3028, w_000_3029, w_000_3030, w_000_3031, w_000_3032, w_000_3033, w_000_3034, w_000_3035, w_000_3036, w_000_3037, w_000_3038, w_000_3039, w_000_3040, w_000_3041, w_000_3042, w_000_3043, w_000_3044, w_000_3045, w_000_3046, w_000_3047, w_000_3048, w_000_3049, w_000_3050, w_000_3051, w_000_3052, w_000_3053, w_000_3054, w_000_3055, w_000_3056, w_000_3057, w_000_3058, w_000_3059, w_000_3060, w_000_3061, w_000_3062, w_000_3063, w_000_3064, w_000_3065, w_000_3066, w_000_3067, w_000_3068, w_000_3069, w_000_3070, w_000_3071, w_000_3072, w_000_3073, w_000_3074, w_000_3075, w_000_3076, w_000_3077, w_000_3078, w_000_3079, w_000_3080, w_000_3081, w_000_3082, w_000_3083, w_000_3084, w_000_3085, w_000_3086, w_000_3087, w_000_3088, w_000_3089, w_000_3090, w_000_3091, w_000_3092, w_000_3093, w_000_3094, w_000_3095, w_000_3096, w_000_3097, w_000_3098, w_000_3099, w_000_3100, w_000_3101, w_000_3102, w_000_3103, w_000_3104, w_000_3105, w_000_3106, w_000_3107, w_000_3108, w_000_3109, w_000_3110, w_000_3111, w_000_3112, w_000_3113, w_000_3114, w_000_3115, w_000_3116, w_000_3117, w_000_3118, w_000_3119, w_000_3120, w_000_3121, w_000_3122, w_000_3123, w_000_3124, w_000_3125, w_000_3126, w_000_3127, w_000_3128, w_000_3129, w_000_3130, w_000_3131, w_000_3132, w_000_3133, w_000_3134, w_000_3135, w_000_3136, w_000_3137, w_000_3138, w_000_3139, w_000_3140, w_000_3141, w_000_3142, w_000_3143, w_000_3144, w_000_3145, w_000_3146, w_000_3147, w_000_3148, w_000_3149, w_000_3150, w_000_3151, w_000_3152, w_000_3153, w_000_3154, w_000_3155, w_000_3156, w_000_3157, w_000_3158, w_000_3159, w_000_3160, w_000_3161, w_000_3162, w_000_3163, w_000_3164, w_000_3165, w_000_3166, w_000_3167, w_000_3168, w_000_3169, w_000_3170, w_000_3171, w_000_3172, w_000_3173, w_000_3174, w_000_3175, w_000_3176, w_000_3177, w_000_3178, w_000_3179, w_000_3180, w_000_3181, w_000_3182, w_000_3183, w_000_3184, w_000_3185, w_000_3186, w_000_3187, w_000_3188, w_000_3189, w_000_3190, w_000_3191, w_000_3192, w_000_3193, w_000_3194, w_000_3195, w_000_3196, w_000_3197, w_000_3198, w_000_3199, w_000_3200, w_000_3201, w_000_3202, w_000_3203, w_000_3204, w_000_3205, w_000_3206, w_000_3207, w_000_3208, w_000_3209, w_000_3210, w_000_3211, w_000_3212, w_000_3213, w_000_3214, w_000_3215, w_000_3216, w_000_3217, w_000_3218, w_000_3219, w_000_3220, w_000_3221, w_000_3222, w_000_3223, w_000_3224, w_000_3225, w_000_3226, w_000_3227, w_000_3228, w_000_3229, w_000_3230, w_000_3231, w_000_3232, w_000_3233, w_000_3234, w_000_3235, w_000_3236, w_000_3237, w_000_3238, w_000_3239, w_000_3240, w_000_3241, w_000_3242, w_000_3243, w_000_3244, w_000_3245, w_000_3246, w_000_3247, w_000_3248, w_000_3249, w_000_3250, w_000_3251, w_000_3252, w_000_3253, w_000_3254, w_000_3255, w_000_3256, w_000_3257, w_000_3258, w_000_3259, w_000_3260, w_000_3261, w_000_3262, w_000_3263, w_000_3264, w_000_3265, w_000_3266, w_000_3267, w_000_3268, w_000_3269, w_000_3270, w_000_3271, w_000_3272, w_000_3273, w_000_3274, w_000_3275, w_000_3276, w_000_3277, w_000_3278, w_000_3279, w_000_3280, w_000_3281, w_000_3282, w_000_3283, w_000_3284, w_000_3285, w_000_3286, w_000_3287, w_000_3288, w_000_3289, w_000_3290, w_000_3291, w_000_3292, w_000_3293, w_000_3294, w_000_3295, w_000_3296, w_000_3297, w_000_3298, w_000_3299, w_000_3300, w_000_3301, w_000_3302, w_000_3303, w_000_3304, w_000_3305, w_000_3306, w_000_3307, w_000_3308, w_000_3309, w_000_3310, w_000_3311, w_000_3312, w_000_3313, w_000_3314, w_000_3315, w_000_3316, w_000_3317, w_000_3318, w_000_3319, w_000_3320, w_000_3321, w_000_3322, w_000_3323, w_000_3324, w_000_3325, w_000_3326, w_000_3327, w_000_3328, w_000_3329, w_000_3330, w_000_3331, w_000_3332, w_000_3333, w_000_3334, w_000_3335, w_000_3336, w_000_3337, w_000_3338, w_000_3339, w_000_3340, w_000_3341, w_000_3342, w_000_3343, w_000_3344, w_000_3345, w_000_3346, w_000_3347, w_000_3348, w_000_3349, w_000_3350, w_000_3351, w_000_3352, w_000_3353, w_000_3354, w_000_3355, w_000_3356, w_000_3357, w_000_3358, w_000_3359, w_000_3360, w_000_3361, w_000_3362, w_000_3363, w_000_3364, w_000_3365, w_000_3366, w_000_3367, w_000_3368, w_000_3369, w_000_3370, w_000_3371, w_000_3372, w_000_3373, w_000_3374, w_000_3375, w_000_3376, w_000_3377, w_000_3378, w_000_3379, w_000_3380, w_000_3381, w_000_3382, w_000_3383, w_000_3384, w_000_3385, w_000_3386, w_000_3387, w_000_3388, w_000_3389, w_000_3390, w_000_3391, w_000_3392, w_000_3393, w_000_3394, w_000_3395, w_000_3396, w_000_3397, w_000_3398, w_000_3399, w_000_3400, w_000_3401, w_000_3402, w_000_3403, w_000_3404, w_000_3405, w_000_3406, w_000_3407, w_000_3408, w_000_3409, w_000_3410, w_000_3411, w_000_3412, w_000_3413, w_000_3414, w_000_3415, w_000_3416, w_000_3417, w_000_3418, w_000_3419, w_000_3420, w_000_3421, w_000_3422, w_000_3423, w_000_3424, w_000_3425, w_000_3426, w_000_3427, w_000_3428, w_000_3429, w_000_3430, w_000_3431, w_000_3432, w_000_3433, w_000_3434, w_000_3435, w_000_3436, w_000_3437, w_000_3438, w_000_3439, w_000_3440, w_000_3441, w_000_3442, w_000_3443, w_000_3444, w_000_3445, w_000_3446, w_000_3447, w_000_3448, w_000_3449, w_000_3450, w_000_3451, w_000_3452, w_000_3453, w_000_3454, w_000_3455, w_000_3456, w_000_3457, w_000_3458, w_000_3459, w_000_3460, w_000_3461, w_000_3462, w_000_3463, w_000_3464, w_000_3465, w_000_3466, w_000_3467, w_000_3468, w_000_3469, w_000_3470, w_000_3471, w_000_3472, w_000_3473, w_000_3474, w_000_3475, w_000_3476, w_000_3477, w_000_3478, w_000_3479, w_000_3480, w_000_3481, w_000_3482, w_000_3483, w_000_3484, w_000_3485, w_000_3486, w_000_3487, w_000_3488, w_000_3489, w_000_3490, w_000_3491, w_000_3492, w_000_3493, w_000_3494, w_000_3495, w_000_3496, w_000_3497, w_000_3498, w_000_3499, w_000_3500, w_000_3501, w_000_3502, w_000_3503, w_000_3504, w_000_3505, w_000_3506, w_000_3507, w_000_3508, w_000_3509, w_000_3510, w_000_3511, w_000_3512, w_000_3513, w_000_3514, w_000_3515, w_000_3516, w_000_3517, w_000_3518, w_000_3519, w_000_3520, w_000_3521, w_000_3522, w_000_3523, w_000_3524, w_000_3525, w_000_3526, w_000_3527, w_000_3528, w_000_3529, w_000_3530, w_000_3531, w_000_3532, w_000_3533, w_000_3534, w_000_3535, w_000_3536, w_000_3537, w_000_3538, w_000_3539, w_000_3540, w_000_3541, w_000_3542, w_000_3543, w_000_3544, w_000_3545, w_000_3546, w_000_3547, w_000_3548, w_000_3549, w_000_3550, w_000_3551, w_000_3552, w_000_3553, w_000_3554, w_000_3555, w_000_3556, w_000_3557, w_000_3558, w_000_3559, w_000_3560, w_000_3561, w_000_3562, w_000_3563, w_000_3564, w_000_3565, w_000_3566, w_000_3567, w_000_3568, w_000_3569, w_000_3570, w_000_3571, w_000_3572, w_000_3573, w_000_3574, w_000_3575, w_000_3576, w_000_3577, w_000_3578, w_000_3579, w_000_3580, w_000_3581, w_000_3582, w_000_3583, w_000_3584, w_000_3585, w_000_3586, w_000_3587, w_000_3588, w_000_3589, w_000_3590, w_000_3591, w_000_3592, w_000_3593, w_000_3594, w_000_3595, w_000_3596, w_000_3597, w_000_3598, w_000_3599, w_000_3600, w_000_3601, w_000_3602, w_000_3603, w_000_3604, w_000_3605, w_000_3606, w_000_3607, w_000_3608, w_000_3609, w_000_3610, w_000_3611, w_000_3612, w_000_3613, w_000_3614, w_000_3615, w_000_3616, w_000_3617, w_000_3618, w_000_3619, w_000_3620, w_000_3621, w_000_3622, w_000_3623, w_000_3624, w_000_3625, w_000_3626, w_000_3627, w_000_3628, w_000_3629, w_000_3630, w_000_3631, w_000_3632, w_000_3633, w_000_3634, w_000_3635, w_000_3636, w_000_3637, w_000_3638, w_000_3639, w_000_3640, w_000_3641, w_000_3642, w_000_3643, w_000_3644, w_000_3645, w_000_3646, w_000_3647, w_000_3648, w_000_3649, w_000_3650, w_000_3651, w_000_3652, w_000_3653, w_000_3654, w_000_3655, w_000_3656, w_000_3657, w_000_3658, w_000_3659, w_000_3660, w_000_3661, w_000_3662, w_000_3663, w_000_3664, w_000_3665, w_000_3666, w_000_3667, w_000_3668, w_000_3669, w_000_3670, w_000_3671, w_000_3672, w_000_3673, w_000_3674, w_000_3675, w_000_3676, w_000_3677, w_000_3678, w_000_3679, w_000_3680, w_000_3681, w_000_3682, w_000_3683, w_000_3684, w_000_3685, w_000_3686, w_000_3687, w_000_3688, w_000_3689, w_000_3690, w_000_3691, w_000_3692, w_000_3693, w_000_3694, w_000_3695, w_000_3696, w_000_3697, w_000_3698, w_000_3699, w_000_3700, w_000_3701, w_000_3702, w_000_3703, w_000_3704, w_000_3705, w_000_3706, w_000_3707, w_000_3708, w_000_3709, w_000_3710, w_000_3711, w_000_3712, w_000_3713, w_000_3714, w_000_3715, w_000_3716, w_000_3717, w_000_3718, w_000_3719, w_000_3720, w_000_3721, w_000_3722, w_000_3723, w_000_3724, w_000_3725, w_000_3726, w_000_3727, w_000_3728, w_000_3729, w_000_3730, w_000_3731, w_000_3732, w_000_3733, w_000_3734, w_000_3735, w_000_3736, w_000_3737, w_000_3738, w_000_3739, w_000_3740, w_000_3741, w_000_3742, w_000_3743, w_000_3744, w_000_3745, w_000_3746, w_000_3747, w_000_3748, w_000_3749, w_000_3750, w_000_3751, w_000_3752, w_000_3753, w_000_3754, w_000_3755, w_000_3756, w_000_3757, w_000_3758, w_000_3759, w_000_3760, w_000_3761, w_000_3762, w_000_3763, w_000_3764, w_000_3765, w_000_3766, w_000_3767, w_000_3768, w_000_3769, w_000_3770, w_000_3771, w_000_3772, w_000_3773, w_000_3774, w_000_3775, w_000_3776, w_000_3777, w_000_3778, w_000_3779, w_000_3780, w_000_3781, w_000_3782, w_000_3783, w_000_3784, w_000_3785, w_000_3786, w_000_3787, w_000_3788, w_000_3789, w_000_3790, w_000_3791, w_000_3792, w_000_3793, w_000_3794, w_000_3795, w_000_3796, w_000_3797, w_000_3798, w_000_3799, w_000_3800, w_000_3801, w_000_3802, w_000_3803, w_000_3804, w_000_3805, w_000_3806, w_000_3807, w_000_3808, w_000_3809, w_000_3810, w_000_3811, w_000_3812, w_000_3813, w_000_3814, w_000_3815, w_000_3816, w_000_3817, w_000_3818, w_000_3819, w_000_3820, w_000_3821, w_000_3822, w_000_3823, w_000_3824, w_000_3825, w_000_3826, w_000_3827, w_000_3828, w_000_3829, w_000_3830, w_000_3831, w_000_3832, w_000_3833, w_000_3834, w_000_3835, w_000_3836, w_000_3837, w_000_3838, w_000_3839, w_000_3840, w_000_3841, w_000_3842, w_000_3843, w_000_3844, w_000_3845, w_000_3846, w_000_3847, w_000_3848, w_000_3849, w_000_3850, w_000_3851, w_000_3852, w_000_3853, w_000_3854, w_000_3855, w_000_3856, w_000_3857, w_000_3858, w_000_3859, w_000_3860, w_000_3861, w_000_3862, w_000_3863, w_000_3864, w_000_3865, w_000_3866, w_000_3867, w_000_3868, w_000_3869, w_000_3870, w_000_3871, w_000_3872, w_000_3873, w_000_3874, w_000_3875, w_000_3876, w_000_3877, w_000_3878, w_000_3879, w_000_3880, w_000_3881, w_000_3882, w_000_3883, w_000_3884, w_000_3885, w_000_3886, w_000_3887, w_000_3888, w_000_3889, w_000_3890, w_000_3891, w_000_3892, w_000_3893, w_000_3894, w_000_3895, w_000_3896, w_000_3897, w_000_3898, w_000_3899, w_000_3900, w_000_3901, w_000_3902, w_000_3903, w_000_3904, w_000_3905, w_000_3906, w_000_3907, w_000_3908, w_000_3909, w_000_3910, w_000_3911, w_000_3912, w_000_3913, w_000_3914, w_000_3915, w_000_3916, w_000_3917, w_000_3918, w_000_3919, w_000_3920, w_000_3921, w_000_3922, w_000_3923, w_000_3924, w_000_3925, w_000_3926, w_000_3927, w_000_3928, w_000_3929, w_000_3930, w_000_3931, w_000_3932, w_000_3933, w_000_3934, w_000_3935, w_000_3936, w_000_3937, w_000_3938, w_000_3939, w_000_3940, w_000_3941, w_000_3942, w_000_3943, w_000_3944, w_000_3945, w_000_3946, w_000_3947, w_000_3948, w_000_3949, w_000_3950, w_000_3951, w_000_3952, w_000_3953, w_000_3954, w_000_3955, w_000_3956, w_000_3957, w_000_3958, w_000_3959, w_000_3960, w_000_3961, w_000_3962, w_000_3963, w_000_3964, w_000_3965, w_000_3966, w_000_3967, w_000_3968, w_000_3969, w_000_3970, w_000_3971, w_000_3972, w_000_3973, w_000_3974, w_000_3975, w_000_3976, w_000_3977, w_000_3978, w_000_3979, w_000_3980, w_000_3981, w_000_3982, w_000_3983, w_000_3984, w_000_3985, w_000_3986, w_000_3987, w_000_3988, w_000_3989, w_000_3990, w_000_3991, w_000_3992, w_000_3993, w_000_3994, w_000_3995, w_000_3996, w_000_3997, w_000_3998, w_000_3999, w_000_4000, w_000_4001, w_000_4002, w_000_4003, w_000_4004, w_000_4005, w_000_4006, w_000_4007, w_000_4008, w_000_4009, w_000_4010, w_000_4011, w_000_4012, w_000_4013, w_000_4014, w_000_4015, w_000_4016, w_000_4017, w_000_4018, w_000_4019, w_000_4020, w_000_4022, w_000_4023, w_000_4024, w_000_4025, w_000_4026, w_000_4027, w_000_4028, w_000_4029, w_000_4030, w_000_4031, w_000_4032, w_000_4033, w_000_4034, w_000_4035, w_000_4036, w_000_4037, w_000_4038, w_000_4039, w_000_4040, w_000_4041, w_000_4042, w_000_4043, w_000_4044, w_000_4045, w_000_4046, w_000_4047, w_000_4048, w_000_4049, w_000_4050, w_000_4051, w_000_4052, w_000_4053, w_000_4054, w_000_4055, w_000_4056, w_000_4057, w_000_4058, w_000_4059, w_000_4060, w_000_4061, w_000_4062, w_000_4063, w_000_4064, w_000_4065, w_000_4066, w_000_4067, w_000_4068, w_000_4069, w_000_4070, w_000_4071, w_000_4072, w_000_4073, w_000_4074, w_000_4075, w_000_4076, w_000_4077, w_000_4078, w_000_4079, w_000_4080, w_000_4081, w_000_4082, w_000_4083, w_000_4084, w_000_4085, w_000_4086, w_000_4087, w_000_4088, w_000_4089, w_000_4090, w_000_4091, w_000_4092, w_000_4093, w_000_4094, w_000_4095, w_000_4096, w_000_4097, w_000_4098, w_000_4099, w_000_4100, w_000_4101, w_000_4102, w_000_4103, w_000_4104, w_000_4105, w_000_4106, w_000_4107, w_000_4108, w_000_4109, w_000_4110, w_000_4111, w_000_4112, w_000_4113, w_000_4114, w_000_4115, w_000_4116, w_000_4117, w_000_4118, w_000_4119, w_000_4120, w_000_4121, w_000_4122, w_000_4123, w_000_4124, w_000_4125, w_000_4126, w_000_4127, w_000_4128, w_000_4129, w_000_4130, w_000_4131, w_000_4132, w_000_4133, w_000_4134, w_000_4135, w_000_4136, w_000_4137, w_000_4138, w_000_4139, w_000_4140, w_000_4141, w_000_4142, w_000_4143, w_000_4144, w_000_4145, w_000_4146, w_000_4147, w_000_4148, w_000_4149, w_000_4150, w_000_4151, w_000_4152, w_000_4153, w_000_4154, w_000_4155, w_000_4156, w_000_4157, w_000_4158, w_000_4159, w_000_4160, w_000_4161, w_000_4162, w_000_4163, w_000_4164, w_000_4165, w_000_4166, w_000_4167, w_000_4168, w_000_4169, w_000_4170, w_000_4171, w_000_4172, w_000_4173, w_000_4174, w_000_4175, w_000_4176, w_000_4177, w_000_4178, w_000_4179, w_000_4180, w_000_4181, w_000_4182, w_000_4183, w_000_4184, w_000_4185, w_000_4186, w_000_4187, w_000_4188, w_000_4189, w_000_4190, w_000_4191, w_000_4192, w_000_4193, w_000_4194, w_000_4195, w_000_4196, w_000_4197, w_000_4198, w_000_4199, w_000_4200, w_000_4201, w_000_4202, w_000_4203, w_000_4204, w_000_4205, w_000_4206, w_000_4207, w_000_4208, w_000_4209, w_000_4210, w_000_4211, w_000_4212, w_000_4213, w_000_4214, w_000_4215, w_000_4216, w_000_4217, w_000_4218, w_000_4219, w_000_4220, w_000_4221, w_000_4222, w_000_4223, w_000_4224, w_000_4225, w_000_4226, w_000_4227, w_000_4228, w_000_4229, w_000_4230, w_000_4231, w_000_4232, w_000_4233, w_000_4234, w_000_4235, w_000_4236, w_000_4237, w_000_4238, w_000_4239, w_000_4240, w_000_4241, w_000_4242, w_000_4243, w_000_4245, w_000_4246, w_000_4247, w_000_4248, w_000_4249, w_000_4250, w_000_4251, w_000_4252, w_000_4253, w_000_4254, w_000_4255, w_000_4256, w_000_4257, w_000_4258, w_000_4259, w_000_4260, w_000_4261, w_000_4262, w_000_4263, w_000_4264, w_000_4265, w_000_4266, w_000_4267, w_000_4268, w_000_4269, w_000_4270, w_000_4271, w_000_4272, w_000_4273, w_000_4274, w_000_4275, w_000_4276, w_000_4277, w_000_4278, w_000_4279, w_000_4280, w_000_4281, w_000_4282, w_000_4283, w_000_4284, w_000_4285, w_000_4286, w_000_4287, w_000_4288, w_000_4289, w_000_4290, w_000_4291, w_000_4292, w_000_4293, w_000_4294, w_000_4295, w_000_4296, w_000_4297, w_000_4298, w_000_4299, w_000_4300, w_000_4301, w_000_4302, w_000_4303, w_000_4304, w_000_4305, w_000_4306, w_000_4307, w_000_4308, w_000_4309, w_000_4310, w_000_4311, w_000_4312, w_000_4313, w_000_4314, w_000_4315, w_000_4316, w_000_4317, w_000_4318, w_000_4319, w_000_4320, w_000_4321, w_000_4322, w_000_4323, w_000_4324, w_000_4325, w_000_4326, w_000_4327, w_000_4328, w_000_4329, w_000_4330, w_000_4331, w_000_4332, w_000_4333, w_000_4334, w_000_4335, w_000_4336, w_000_4337, w_000_4338, w_000_4339, w_000_4340, w_000_4341, w_000_4342, w_000_4343, w_000_4344, w_000_4345, w_000_4346, w_000_4347, w_000_4348, w_000_4349, w_000_4350, w_000_4351, w_000_4352, w_000_4353, w_000_4354, w_000_4355, w_000_4356, w_000_4357, w_000_4358, w_000_4359, w_000_4360, w_000_4361, w_000_4362, w_000_4363, w_000_4364, w_000_4365, w_000_4366, w_000_4367, w_000_4368, w_000_4369, w_000_4370, w_000_4371, w_000_4372, w_000_4373, w_000_4374, w_000_4375, w_000_4376, w_000_4377, w_000_4378, w_000_4379, w_000_4380, w_000_4381, w_000_4382, w_000_4383, w_000_4384, w_000_4385, w_000_4386, w_000_4387, w_000_4388, w_000_4389, w_000_4390, w_000_4391, w_000_4392, w_000_4393, w_000_4394, w_000_4395, w_000_4396, w_000_4397, w_000_4398, w_000_4399, w_000_4400, w_000_4401, w_000_4402, w_000_4403, w_000_4404, w_000_4405, w_000_4406, w_000_4407, w_000_4408, w_000_4409, w_000_4410, w_000_4411, w_000_4412, w_000_4413, w_000_4414, w_000_4415, w_000_4416, w_000_4417, w_000_4418, w_000_4419, w_000_4420, w_000_4421, w_000_4422, w_000_4423, w_000_4424, w_000_4425, w_000_4426, w_000_4427, w_000_4428, w_000_4429, w_000_4430, w_000_4431, w_000_4432, w_000_4433, w_000_4434, w_000_4435, w_000_4436, w_000_4437, w_000_4438, w_000_4439, w_000_4440, w_000_4441, w_000_4442, w_000_4443, w_000_4444, w_000_4445, w_000_4446, w_000_4447, w_000_4448, w_000_4449, w_000_4450, w_000_4451, w_000_4452, w_000_4453, w_000_4454, w_000_4455, w_000_4456, w_000_4457, w_000_4458, w_000_4459, w_000_4460, w_000_4461, w_000_4462, w_000_4463, w_000_4464, w_000_4465, w_000_4466, w_000_4467, w_000_4468, w_000_4469, w_000_4470, w_000_4471, w_000_4472, w_000_4473, w_000_4474, w_000_4475, w_000_4476, w_000_4477, w_000_4478, w_000_4479, w_000_4480, w_000_4481, w_000_4482, w_000_4483, w_000_4484, w_000_4485, w_000_4486, w_000_4487, w_000_4488, w_000_4489, w_000_4490, w_000_4491, w_000_4492, w_000_4493, w_000_4494, w_000_4495, w_000_4496, w_000_4497, w_000_4498, w_000_4499, w_000_4500, w_000_4501, w_000_4502, w_000_4503, w_000_4504, w_000_4505, w_000_4506, w_000_4507, w_000_4508, w_000_4509, w_000_4510, w_000_4511, w_000_4512, w_000_4513, w_000_4514, w_000_4515, w_000_4516, w_000_4517, w_000_4518, w_000_4519, w_000_4520, w_000_4521, w_000_4522, w_000_4523, w_000_4524, w_000_4525, w_000_4526, w_000_4527, w_000_4528, w_000_4529, w_000_4530, w_000_4531, w_000_4532, w_000_4533, w_000_4534, w_000_4535, w_000_4536, w_000_4537, w_000_4538, w_000_4539, w_000_4540, w_000_4541, w_000_4542, w_000_4543, w_000_4544, w_000_4545, w_000_4546, w_000_4547, w_000_4548, w_000_4549, w_000_4550, w_000_4551, w_000_4552, w_000_4553, w_000_4554, w_000_4555, w_000_4556, w_000_4557, w_000_4558, w_000_4559, w_000_4560, w_000_4561, w_000_4562, w_000_4563, w_000_4564, w_000_4565, w_000_4566, w_000_4567, w_000_4568, w_000_4569, w_000_4570, w_000_4571, w_000_4572, w_000_4573, w_000_4574, w_000_4575, w_000_4576, w_000_4577, w_000_4578, w_000_4579, w_000_4580, w_000_4581, w_000_4582, w_000_4583, w_000_4584, w_000_4585, w_000_4586, w_000_4588, w_000_4589, w_000_4590, w_000_4591, w_000_4592, w_000_4593, w_000_4594, w_000_4595, w_000_4596, w_000_4597, w_000_4598, w_000_4599, w_000_4600, w_000_4601, w_000_4602, w_000_4603, w_000_4604, w_000_4605, w_000_4606, w_000_4607, w_000_4608, w_000_4609, w_000_4610, w_000_4611, w_000_4612, w_000_4613, w_000_4614, w_000_4615, w_000_4616, w_000_4617, w_000_4618, w_000_4619, w_000_4620, w_000_4621, w_000_4622, w_000_4623, w_000_4624, w_000_4625, w_000_4626, w_000_4627, w_000_4628, w_000_4629, w_000_4630, w_000_4631, w_000_4632, w_000_4633, w_000_4634, w_000_4635, w_000_4636, w_000_4637, w_000_4638, w_000_4639, w_000_4640, w_000_4641, w_000_4642, w_000_4643, w_000_4644, w_000_4645, w_000_4646, w_000_4647, w_000_4648, w_000_4649, w_000_4650, w_000_4651, w_000_4652, w_000_4653, w_000_4654, w_000_4655, w_000_4656, w_000_4657, w_000_4658, w_000_4659, w_000_4660, w_000_4661, w_000_4662, w_000_4663, w_000_4664, w_000_4665, w_000_4666, w_000_4667, w_000_4668, w_000_4669, w_000_4670, w_000_4671, w_000_4672, w_000_4673, w_000_4674, w_000_4675, w_000_4676, w_000_4677, w_000_4678, w_000_4679, w_000_4680, w_000_4681, w_000_4682, w_000_4683, w_000_4684, w_000_4685, w_000_4686, w_000_4687, w_000_4688, w_000_4689, w_000_4690, w_000_4691, w_000_4692, w_000_4693, w_000_4694, w_000_4695, w_000_4696, w_000_4697, w_000_4698, w_000_4699, w_000_4700, w_000_4701, w_000_4702, w_000_4703, w_000_4704, w_000_4705, w_000_4706, w_000_4707, w_000_4708, w_000_4709, w_000_4710, w_000_4711, w_000_4712, w_000_4713, w_000_4714, w_000_4715, w_000_4716, w_000_4717, w_000_4718, w_000_4719, w_000_4720, w_000_4721, w_000_4722, w_000_4723, w_000_4724, w_000_4725, w_000_4726, w_000_4727, w_000_4728, w_000_4729, w_000_4730, w_000_4731, w_000_4732, w_000_4733, w_000_4734, w_000_4735, w_000_4736, w_000_4737, w_000_4738, w_000_4739, w_000_4740, w_000_4741, w_000_4742, w_000_4743, w_000_4744, w_000_4745, w_000_4746, w_000_4747, w_000_4748, w_000_4749, w_000_4750, w_000_4751, w_000_4752, w_000_4753, w_000_4754, w_000_4755, w_000_4756, w_000_4757, w_000_4758, w_000_4759, w_000_4760, w_000_4761, w_000_4762, w_000_4763, w_000_4764, w_000_4765, w_000_4766, w_000_4767, w_000_4768, w_000_4769, w_000_4770, w_000_4771, w_000_4772, w_000_4773, w_000_4774, w_000_4775, w_000_4776, w_000_4777, w_000_4778, w_000_4779, w_000_4780, w_000_4781, w_000_4782, w_000_4783, w_000_4784, w_000_4785, w_000_4786, w_000_4787, w_000_4788, w_000_4789, w_000_4790, w_000_4791, w_000_4792, w_000_4793, w_000_4794, w_000_4795, w_000_4796, w_000_4797, w_000_4798, w_000_4799, w_000_4800, w_000_4801, w_000_4802, w_000_4803, w_000_4804, w_000_4805, w_000_4806, w_000_4807, w_000_4808, w_000_4809, w_000_4810, w_000_4811, w_000_4812, w_000_4813, w_000_4814, w_000_4815, w_000_4816, w_000_4817, w_000_4818, w_000_4819, w_000_4820, w_000_4821, w_000_4822, w_000_4823, w_000_4824, w_000_4825, w_000_4826, w_000_4827, w_000_4828, w_000_4829, w_000_4830, w_000_4831, w_000_4832, w_000_4833, w_000_4834, w_000_4835, w_000_4836, w_000_4837, w_000_4838, w_000_4839, w_000_4840, w_000_4841, w_000_4842, w_000_4843, w_000_4844, w_000_4845, w_000_4846, w_000_4847, w_000_4848, w_000_4849, w_000_4850, w_000_4851, w_000_4852, w_000_4853, w_000_4854, w_000_4855, w_000_4856, w_000_4857, w_000_4858, w_000_4859, w_000_4860, w_000_4861, w_000_4862, w_000_4863, w_000_4864, w_000_4865, w_000_4866, w_000_4867, w_000_4868, w_000_4869, w_000_4870, w_000_4871, w_000_4872, w_000_4873, w_000_4874, w_000_4875, w_000_4876, w_000_4877, w_000_4878, w_000_4879, w_000_4880, w_000_4881, w_000_4882, w_000_4883, w_000_4884, w_000_4885, w_000_4886, w_000_4887, w_000_4888, w_000_4889, w_000_4890, w_000_4891, w_000_4892, w_000_4893, w_000_4894, w_000_4895, w_000_4896, w_000_4897, w_000_4898, w_000_4899, w_000_4900, w_000_4901, w_000_4902, w_000_4903, w_000_4904, w_000_4905, w_000_4906, w_000_4907, w_000_4908, w_000_4909, w_000_4910, w_000_4911, w_000_4912, w_000_4913, w_000_4914, w_000_4915, w_000_4916, w_000_4917, w_000_4918, w_000_4919, w_000_4920, w_000_4921, w_000_4922, w_000_4923, w_000_4924, w_000_4925, w_000_4926, w_000_4927, w_000_4928, w_000_4929, w_000_4930, w_000_4931, w_000_4932, w_000_4933, w_000_4934, w_000_4935, w_000_4936, w_000_4937, w_000_4938, w_000_4939, w_000_4940, w_000_4941, w_000_4942, w_000_4943, w_000_4944, w_000_4945, w_000_4946, w_000_4947, w_000_4948, w_000_4949, w_000_4950, w_000_4951, w_000_4952, w_000_4953, w_000_4954, w_000_4955, w_000_4956, w_000_4957, w_000_4958, w_000_4959, w_000_4960, w_000_4961, w_000_4962, w_000_4963, w_000_4964, w_000_4965, w_000_4966, w_000_4967, w_000_4968, w_000_4969, w_000_4970, w_000_4971, w_000_4972, w_000_4973, w_000_4974, w_000_4975, w_000_4976, w_000_4977, w_000_4978, w_000_4979, w_000_4980, w_000_4981, w_000_4982, w_000_4983, w_000_4984, w_000_4985, w_000_4986, w_000_4987, w_000_4988, w_000_4989, w_000_4990, w_000_4991, w_000_4992, w_000_4993, w_000_4994, w_000_4995, w_000_4996, w_000_4997, w_000_4998, w_000_4999, w_000_5000, w_000_5001, w_000_5002, w_000_5003, w_000_5004, w_000_5005, w_000_5006, w_000_5007, w_000_5008, w_000_5009, w_000_5010, w_000_5011, w_000_5012, w_000_5013, w_000_5014, w_000_5015, w_000_5016, w_000_5017, w_000_5018, w_000_5019, w_000_5020, w_000_5021, w_000_5022, w_000_5023, w_000_5024, w_000_5025, w_000_5026, w_000_5027, w_000_5028, w_000_5029, w_000_5030, w_000_5031, w_000_5032, w_000_5033, w_000_5034, w_000_5035, w_000_5036, w_000_5037, w_000_5038, w_000_5039, w_000_5040, w_000_5041, w_000_5042, w_000_5043, w_000_5044, w_000_5045, w_000_5046, w_000_5047, w_000_5048, w_000_5049, w_000_5050, w_000_5051, w_000_5052, w_000_5053, w_000_5054, w_000_5055, w_000_5056, w_000_5057, w_000_5058, w_000_5059, w_000_5060, w_000_5061, w_000_5062, w_000_5063, w_000_5064, w_000_5065, w_000_5066, w_000_5067, w_000_5068, w_000_5069, w_000_5070, w_000_5071, w_000_5072, w_000_5073, w_000_5074, w_000_5075, w_000_5076, w_000_5077, w_000_5078, w_000_5079, w_000_5080, w_000_5081, w_000_5082, w_000_5083, w_000_5084, w_000_5085, w_000_5086, w_000_5087, w_000_5088, w_000_5089, w_000_5090, w_000_5091, w_000_5092, w_000_5093, w_000_5094, w_000_5095, w_000_5096, w_000_5097, w_000_5098, w_000_5099, w_000_5100, w_000_5101, w_000_5102, w_000_5103, w_000_5104, w_000_5105, w_000_5106, w_000_5107, w_000_5108, w_000_5109, w_000_5110, w_000_5111, w_000_5112, w_000_5113, w_000_5114, w_000_5115, w_000_5116, w_000_5117, w_000_5118, w_000_5119, w_000_5120, w_000_5121, w_000_5122, w_000_5123, w_000_5124, w_000_5125, w_000_5126, w_000_5127, w_000_5128, w_000_5129, w_000_5130, w_000_5131, w_000_5132, w_000_5133, w_000_5134, w_000_5135, w_000_5136, w_000_5137, w_000_5138, w_000_5139, w_000_5140, w_000_5141, w_000_5142, w_000_5143, w_000_5144, w_000_5145, w_000_5146, w_000_5147, w_000_5148, w_000_5149, w_000_5150, w_000_5151, w_000_5152, w_000_5153, w_000_5154, w_000_5155, w_000_5156, w_000_5157, w_000_5158, w_000_5159, w_000_5160, w_000_5161, w_000_5162, w_000_5163, w_000_5164, w_000_5165, w_000_5166, w_000_5167, w_000_5168, w_000_5169, w_000_5170, w_000_5171, w_000_5172, w_000_5173, w_000_5174, w_000_5175, w_000_5176, w_000_5177, w_000_5178, w_000_5179, w_000_5180, w_000_5181, w_000_5182, w_000_5183, w_000_5184, w_000_5185, w_000_5186, w_000_5187, w_000_5188, w_000_5189, w_000_5190, w_000_5191, w_000_5192, w_000_5193, w_000_5194, w_000_5195, w_000_5196, w_000_5197, w_000_5198, w_000_5199, w_000_5200, w_000_5201, w_000_5202, w_000_5203, w_000_5204, w_000_5205, w_000_5206, w_000_5207, w_000_5208, w_000_5209, w_000_5210, w_000_5211, w_000_5212, w_000_5213, w_000_5214, w_000_5215, w_000_5216, w_000_5217, w_000_5218, w_000_5219, w_000_5220, w_000_5221, w_000_5222, w_000_5223, w_000_5224, w_000_5225, w_000_5226, w_000_5227, w_000_5228, w_000_5229, w_000_5230, w_000_5231, w_000_5232, w_000_5233, w_000_5234, w_000_5235, w_000_5236, w_000_5237, w_000_5238, w_000_5239, w_000_5240, w_000_5241, w_000_5242, w_000_5243, w_000_5244, w_000_5245, w_000_5246, w_000_5247, w_000_5248, w_000_5249, w_000_5250, w_000_5251, w_000_5252, w_000_5253, w_000_5254, w_000_5255, w_000_5256, w_000_5257, w_000_5258, w_000_5259, w_000_5260, w_000_5261, w_000_5262, w_000_5263, w_000_5264, w_000_5265, w_000_5266, w_000_5267, w_000_5268, w_000_5269, w_000_5270, w_000_5271, w_000_5272, w_000_5273, w_000_5274, w_000_5275, w_000_5276, w_000_5277, w_000_5278, w_000_5279, w_000_5280, w_000_5281, w_000_5282, w_000_5283, w_000_5284, w_000_5285, w_000_5286, w_000_5287, w_000_5288, w_000_5289, w_000_5290, w_000_5291, w_000_5292, w_000_5293, w_000_5294, w_000_5295, w_000_5296, w_000_5297, w_000_5298, w_000_5299, w_000_5300, w_000_5301, w_000_5302, w_000_5303, w_000_5304, w_000_5305, w_000_5306, w_000_5307, w_000_5308, w_000_5309, w_000_5310, w_000_5311, w_000_5312, w_000_5313, w_000_5314, w_000_5315, w_000_5316, w_000_5317, w_000_5318, w_000_5319, w_000_5320, w_000_5321, w_000_5322, w_000_5323, w_000_5324, w_000_5325, w_000_5326, w_000_5327, w_000_5328, w_000_5329, w_000_5330, w_000_5331, w_000_5332, w_000_5333, w_000_5334, w_000_5335, w_000_5336, w_000_5337, w_000_5338, w_000_5339, w_000_5340, w_000_5341, w_000_5342, w_000_5343, w_000_5344, w_000_5345, w_000_5346, w_000_5347, w_000_5348, w_000_5349, w_000_5350, w_000_5351, w_000_5352, w_000_5353, w_000_5354, w_000_5355, w_000_5356, w_000_5357, w_000_5358, w_000_5359, w_000_5360, w_000_5361, w_000_5362, w_000_5363, w_000_5364, w_000_5365, w_000_5366, w_000_5367, w_000_5368, w_000_5369, w_000_5370, w_000_5371, w_000_5372, w_000_5373, w_000_5374, w_000_5375, w_000_5376, w_000_5377, w_000_5378, w_000_5379, w_000_5380, w_000_5381, w_000_5382, w_000_5383, w_000_5384, w_000_5385, w_000_5386, w_000_5387, w_000_5388, w_000_5389, w_000_5390, w_000_5391, w_000_5392, w_000_5393, w_000_5394, w_000_5395, w_000_5396, w_000_5397, w_000_5398, w_000_5399, w_000_5400, w_000_5401, w_000_5402, w_000_5403, w_000_5404, w_000_5405, w_000_5406, w_000_5407, w_000_5408, w_000_5409, w_000_5410, w_000_5411, w_000_5412, w_000_5413, w_000_5414, w_000_5415, w_000_5416, w_000_5417, w_000_5418, w_000_5419, w_000_5420, w_000_5421, w_000_5422, w_000_5423, w_000_5424, w_000_5425, w_000_5426, w_000_5427, w_000_5428, w_000_5429, w_000_5430, w_000_5431, w_000_5432, w_000_5433, w_000_5434, w_000_5435, w_000_5436, w_000_5437, w_000_5438, w_000_5439, w_000_5440, w_000_5441, w_000_5442, w_000_5443, w_000_5444, w_000_5445, w_000_5446, w_000_5447, w_000_5448, w_000_5449, w_000_5450, w_000_5451, w_000_5452, w_000_5453, w_000_5454, w_000_5455, w_000_5456, w_000_5457, w_000_5458, w_000_5459, w_000_5460, w_000_5461, w_000_5462, w_000_5463, w_000_5464, w_000_5465, w_000_5466, w_000_5467, w_000_5468, w_000_5469, w_000_5470, w_000_5471, w_000_5472, w_000_5473, w_000_5474, w_000_5475, w_000_5476, w_000_5477, w_000_5478, w_000_5479, w_000_5480, w_000_5481, w_000_5482, w_000_5483, w_000_5484, w_000_5485, w_000_5486, w_000_5487, w_000_5488, w_000_5489, w_000_5490, w_000_5491, w_000_5492, w_000_5493, w_000_5494, w_000_5495, w_000_5496, w_000_5497, w_000_5498, w_000_5499, w_000_5500, w_000_5501, w_000_5502, w_000_5503, w_000_5504, w_000_5505, w_000_5506, w_000_5507, w_000_5508, w_000_5509, w_000_5510, w_000_5511, w_000_5512, w_000_5513, w_000_5514, w_000_5515, w_000_5516, w_000_5517, w_000_5518, w_000_5519, w_000_5520, w_000_5521, w_000_5522, w_000_5523, w_000_5524, w_000_5525, w_000_5526, w_000_5527, w_000_5528, w_000_5529, w_000_5530, w_000_5531, w_000_5532, w_000_5533, w_000_5534, w_000_5535, w_000_5536, w_000_5537, w_000_5538, w_000_5539, w_000_5540, w_000_5541, w_000_5542, w_000_5543, w_000_5544, w_000_5545, w_000_5546, w_000_5547, w_000_5548, w_000_5549, w_000_5550, w_000_5551, w_000_5552, w_000_5553, w_000_5554, w_000_5555, w_000_5556, w_000_5557, w_000_5558, w_000_5559, w_000_5560, w_000_5561, w_000_5562, w_000_5563, w_000_5564, w_000_5565, w_000_5566, w_000_5567, w_000_5568, w_000_5569, w_000_5570, w_000_5571, w_000_5572, w_000_5573, w_000_5574, w_000_5575, w_000_5576, w_000_5577, w_000_5578, w_000_5579, w_000_5580, w_000_5581, w_000_5582, w_000_5583, w_000_5584, w_000_5585, w_000_5586, w_000_5587, w_000_5588, w_000_5589, w_000_5590, w_000_5591, w_000_5592, w_000_5593, w_000_5594, w_000_5595, w_000_5596, w_000_5597, w_000_5598, w_000_5599, w_000_5600, w_000_5601, w_000_5602, w_000_5603, w_000_5604, w_000_5605, w_000_5606, w_000_5607, w_000_5608, w_000_5609, w_000_5610, w_000_5611, w_000_5612, w_000_5613, w_000_5614, w_000_5615, w_000_5616, w_000_5617, w_000_5618, w_000_5619, w_000_5620, w_000_5621, w_000_5622, w_000_5623, w_000_5624, w_000_5625, w_000_5626, w_000_5627, w_000_5628, w_000_5629, w_000_5630, w_000_5631, w_000_5632, w_000_5633, w_000_5634, w_000_5635, w_000_5636, w_000_5637, w_000_5638, w_000_5639, w_000_5640, w_000_5641, w_000_5642, w_000_5643, w_000_5644, w_000_5645, w_000_5646, w_000_5647, w_000_5648, w_000_5649, w_000_5650, w_000_5651, w_000_5652, w_000_5653, w_000_5654, w_000_5655, w_000_5656, w_000_5657, w_000_5658, w_000_5659, w_000_5660, w_000_5661, w_000_5662, w_000_5663, w_000_5664, w_000_5665, w_000_5666, w_000_5667, w_000_5668, w_000_5669, w_000_5670, w_000_5671, w_000_5672, w_000_5673, w_000_5674, w_000_5675, w_000_5676, w_000_5677, w_000_5678, w_000_5679, w_000_5680, w_000_5681, w_000_5682, w_000_5683, w_000_5684, w_000_5685, w_000_5686, w_000_5687, w_000_5688, w_000_5689, w_000_5690, w_000_5691, w_000_5692, w_000_5693, w_000_5694, w_000_5695, w_000_5696, w_000_5697, w_000_5698, w_000_5699, w_000_5700, w_000_5701, w_000_5702, w_000_5703, w_000_5704, w_000_5705, w_000_5706, w_000_5707, w_000_5708, w_000_5709, w_000_5710, w_000_5711, w_000_5712, w_000_5713, w_000_5714, w_000_5715, w_000_5716, w_000_5717, w_000_5718, w_000_5719, w_000_5720, w_000_5721, w_000_5722, w_000_5723, w_000_5724, w_000_5725, w_000_5726, w_000_5727, w_000_5728, w_000_5729, w_000_5730, w_000_5731, w_000_5732, w_000_5733, w_000_5734, w_000_5735, w_000_5736, w_000_5737, w_000_5738, w_000_5739, w_000_5740, w_000_5741, w_000_5742, w_000_5743, w_000_5744, w_000_5745, w_000_5746, w_000_5747, w_000_5748, w_000_5749, w_000_5750, w_000_5751, w_000_5752, w_000_5753, w_000_5754, w_000_5755, w_000_5756, w_000_5757, w_000_5758, w_000_5759, w_000_5760, w_000_5761, w_000_5762, w_000_5763, w_000_5764, w_000_5765, w_000_5766, w_000_5767, w_000_5768, w_000_5769, w_000_5770, w_000_5771, w_000_5772, w_000_5773, w_000_5774, w_000_5775, w_000_5776, w_000_5777, w_000_5778, w_000_5779, w_000_5780, w_000_5781, w_000_5782, w_000_5783, w_000_5784, w_000_5785, w_000_5786, w_000_5787, w_000_5788, w_000_5789, w_000_5790, w_000_5791, w_000_5792, w_000_5793, w_000_5794, w_000_5795, w_000_5796, w_000_5797, w_000_5798, w_000_5799, w_000_5800, w_000_5801, w_000_5802, w_000_5803, w_000_5804, w_000_5805, w_000_5806, w_000_5807, w_000_5808, w_000_5809, w_000_5810, w_000_5811, w_000_5812, w_000_5813, w_000_5814, w_000_5815, w_000_5816, w_000_5817, w_000_5818, w_000_5819, w_000_5820, w_000_5821, w_000_5822, w_000_5823, w_000_5824, w_000_5825, w_000_5826, w_000_5827, w_000_5828, w_000_5829, w_000_5830, w_000_5831, w_000_5832, w_000_5833, w_000_5834, w_000_5835, w_000_5836, w_000_5837, w_000_5838, w_000_5839, w_000_5840, w_000_5841, w_000_5842, w_000_5843, w_000_5844, w_000_5845, w_000_5846, w_000_5847, w_000_5848, w_000_5849, w_000_5850, w_000_5851, w_000_5852, w_000_5853, w_000_5854, w_000_5855, w_000_5856, w_000_5857, w_000_5858, w_000_5859, w_000_5860, w_000_5861, w_000_5862, w_000_5863, w_000_5864, w_000_5865, w_000_5866, w_000_5867, w_000_5868, w_000_5869, w_000_5870, w_000_5871, w_000_5872, w_000_5873, w_000_5874, w_000_5875, w_000_5876, w_000_5877, w_000_5878, w_000_5879, w_000_5880, w_000_5881, w_000_5882, w_000_5883, w_000_5884, w_000_5885, w_000_5886, w_000_5887, w_000_5888, w_000_5889, w_000_5890, w_000_5891, w_000_5892, w_000_5893, w_000_5894, w_000_5895, w_000_5896, w_000_5897, w_000_5898, w_000_5899, w_000_5900, w_000_5901, w_000_5902, w_000_5903, w_000_5904, w_000_5905, w_000_5906, w_000_5907, w_000_5908, w_000_5909, w_000_5910, w_000_5911, w_000_5912, w_000_5913, w_000_5914, w_000_5915, w_000_5916, w_000_5917, w_000_5918, w_000_5919, w_000_5920, w_000_5921, w_000_5922, w_000_5923, w_000_5924, w_000_5925, w_000_5926, w_000_5927, w_000_5928, w_000_5929, w_000_5930, w_000_5931, w_000_5932, w_000_5933, w_000_5934, w_000_5935, w_000_5936, w_000_5937, w_000_5938, w_000_5939, w_000_5940, w_000_5941, w_000_5942, w_000_5943, w_000_5944, w_000_5945, w_000_5946, w_000_5947, w_000_5948, w_000_5949, w_000_5950, w_000_5951, w_000_5952, w_000_5953, w_000_5954, w_000_5955, w_000_5956, w_000_5957, w_000_5958, w_000_5959, w_000_5960, w_000_5961, w_000_5962, w_000_5963, w_000_5964, w_000_5965, w_000_5966, w_000_5967, w_000_5968, w_000_5969, w_000_5970, w_000_5971, w_000_5972, w_000_5973, w_000_5974, w_000_5975, w_000_5976, w_000_5977, w_000_5978, w_000_5979, w_000_5980, w_000_5981, w_000_5982, w_000_5983, w_000_5984, w_000_5985, w_000_5986, w_000_5987, w_000_5988, w_000_5989, w_000_5990, w_000_5991, w_000_5992, w_000_5993, w_000_5994, w_000_5995, w_000_5996, w_000_5997, w_000_5998, w_000_5999, w_000_6000, w_000_6001, w_000_6002, w_000_6003, w_000_6004, w_000_6005, w_000_6006, w_000_6007, w_000_6008, w_000_6009, w_000_6010, w_000_6011, w_000_6012, w_000_6013, w_000_6014, w_000_6015, w_000_6016, w_000_6017, w_000_6018, w_000_6019, w_000_6020, w_000_6021, w_000_6022, w_000_6023, w_000_6024, w_000_6025, w_000_6026, w_000_6027, w_000_6028, w_000_6029, w_000_6030, w_000_6031, w_000_6032, w_000_6033, w_000_6034, w_000_6035, w_000_6036, w_000_6037, w_000_6038, w_000_6039, w_000_6040, w_000_6041, w_000_6042, w_000_6043, w_000_6044, w_000_6045, w_000_6046, w_000_6047, w_000_6048, w_000_6049, w_000_6050, w_000_6051, w_000_6052, w_000_6053, w_000_6054, w_000_6055, w_000_6056, w_000_6057, w_000_6058, w_000_6059, w_000_6060, w_000_6061, w_000_6062, w_000_6063, w_000_6064, w_000_6065, w_000_6066, w_000_6067, w_000_6068, w_000_6069, w_000_6070, w_000_6071, w_000_6072, w_000_6073, w_000_6074, w_000_6075, w_000_6076, w_000_6077, w_000_6078, w_000_6079, w_000_6080, w_000_6081, w_000_6082, w_000_6083, w_000_6084, w_000_6085, w_000_6086, w_000_6087, w_000_6088, w_000_6089, w_000_6090, w_000_6091, w_000_6092, w_000_6093, w_000_6094, w_000_6095, w_000_6096, w_000_6097, w_000_6098, w_000_6099, w_000_6100, w_000_6101, w_000_6102, w_000_6103, w_000_6104, w_000_6105, w_000_6106, w_000_6107, w_000_6108, w_000_6109, w_000_6110, w_000_6111, w_000_6112, w_000_6113, w_000_6114, w_000_6115, w_000_6116, w_000_6117, w_000_6118, w_000_6119, w_000_6120, w_000_6121, w_000_6122, w_000_6123, w_000_6124, w_000_6125, w_000_6126, w_000_6127, w_000_6128, w_000_6129, w_000_6130, w_000_6131, w_000_6132, w_000_6133, w_000_6134, w_000_6135, w_000_6136, w_000_6137, w_000_6138, w_000_6139, w_000_6140, w_000_6141, w_000_6142, w_000_6143, w_000_6144, w_000_6145, w_000_6146, w_000_6147, w_000_6148, w_000_6149, w_000_6150, w_000_6151, w_000_6152, w_000_6153, w_000_6154, w_000_6155, w_000_6156, w_000_6157, w_000_6158, w_000_6159, w_000_6160, w_000_6161, w_000_6162, w_000_6163, w_000_6164, w_000_6165, w_000_6166, w_000_6167, w_000_6168, w_000_6169, w_000_6170, w_000_6171, w_000_6172, w_000_6173, w_000_6174, w_000_6175, w_000_6176, w_000_6177, w_000_6178, w_000_6179, w_000_6180, w_000_6181, w_000_6182, w_000_6183, w_000_6184, w_000_6185, w_000_6186, w_000_6187, w_000_6188, w_000_6189, w_000_6190, w_000_6191, w_000_6192, w_000_6193, w_000_6194, w_000_6195, w_000_6196, w_000_6197, w_000_6198, w_000_6199, w_000_6200, w_000_6201, w_000_6202, w_000_6203, w_000_6204, w_000_6205, w_000_6206, w_000_6207, w_000_6208, w_000_6209, w_000_6210, w_000_6211, w_000_6212, w_000_6213, w_000_6214, w_000_6215, w_000_6216, w_000_6217, w_000_6218, w_000_6219, w_000_6220, w_000_6221, w_000_6222, w_000_6223, w_000_6224, w_000_6225, w_000_6226, w_000_6227, w_000_6228, w_000_6229, w_000_6230, w_000_6231, w_000_6232, w_000_6233, w_000_6234, w_000_6235, w_000_6236, w_000_6237, w_000_6238, w_000_6239, w_000_6240, w_000_6241, w_000_6242, w_000_6243, w_000_6244, w_000_6245, w_000_6246, w_000_6247, w_000_6248, w_000_6249, w_000_6250, w_000_6251, w_000_6252, w_000_6253, w_000_6254, w_000_6255, w_000_6256, w_000_6257, w_000_6258, w_000_6259, w_000_6260, w_000_6261, w_000_6262, w_000_6263, w_000_6264, w_000_6265, w_000_6266, w_000_6267, w_000_6268, w_000_6269, w_000_6270, w_000_6271, w_000_6272, w_000_6273, w_000_6274, w_000_6275, w_000_6276, w_000_6277, w_000_6278, w_000_6279, w_000_6280, w_000_6281, w_000_6282, w_000_6283, w_000_6284, w_000_6285, w_000_6286, w_000_6287, w_000_6288, w_000_6289, w_000_6290, w_000_6291, w_000_6293, w_000_6294, w_000_6295, w_000_6296, w_000_6297, w_000_6298, w_000_6299, w_000_6300, w_000_6301, w_000_6302, w_000_6303, w_000_6304, w_000_6305, w_000_6306, w_000_6307, w_000_6308, w_000_6309, w_000_6310, w_000_6311, w_000_6312, w_000_6313, w_000_6314, w_000_6315, w_000_6316, w_000_6317, w_000_6318, w_000_6319, w_000_6320, w_000_6321, w_000_6322, w_000_6323, w_000_6324, w_000_6325, w_000_6326, w_000_6327, w_000_6328, w_000_6329, w_000_6330, w_000_6331, w_000_6332, w_000_6333, w_000_6334, w_000_6335, w_000_6336, w_000_6337, w_000_6338, w_000_6339, w_000_6340, w_000_6341, w_000_6342, w_000_6343, w_000_6344, w_000_6345, w_000_6346, w_000_6347, w_000_6348, w_000_6349, w_000_6350, w_000_6351, w_000_6352, w_000_6353, w_000_6354, w_000_6355, w_000_6356, w_000_6357, w_000_6358, w_000_6359, w_000_6360, w_000_6361, w_000_6362, w_000_6363, w_000_6364, w_000_6365, w_000_6366, w_000_6367, w_000_6368, w_000_6369, w_000_6370, w_000_6371, w_000_6372, w_000_6373, w_000_6374, w_000_6375, w_000_6376, w_000_6377, w_000_6378, w_000_6379, w_000_6380, w_000_6381, w_000_6382, w_000_6383, w_000_6384, w_000_6385, w_000_6386, w_000_6387, w_000_6388, w_000_6389, w_000_6390, w_000_6391, w_000_6392, w_000_6393, w_000_6394, w_000_6395, w_000_6396, w_000_6397, w_000_6398, w_000_6399, w_000_6400, w_000_6401, w_000_6402, w_000_6403, w_000_6404, w_000_6405, w_000_6406, w_000_6407, w_000_6408, w_000_6409, w_000_6410, w_000_6411, w_000_6412, w_000_6413, w_000_6414, w_000_6415, w_000_6416, w_000_6417, w_000_6418, w_000_6419, w_000_6420, w_000_6421, w_000_6422, w_000_6423, w_000_6424, w_000_6425, w_000_6426, w_000_6427, w_000_6428, w_000_6429, w_000_6430, w_000_6431, w_000_6432, w_000_6433, w_000_6434, w_000_6435, w_000_6436, w_000_6437, w_000_6438, w_000_6439, w_000_6440, w_000_6441, w_000_6442, w_000_6443, w_000_6444, w_000_6445, w_000_6446, w_000_6447, w_000_6448, w_000_6449, w_000_6450, w_000_6451, w_000_6452, w_000_6453, w_000_6454, w_000_6455, w_000_6456, w_000_6457, w_000_6458, w_000_6459, w_000_6460, w_000_6461, w_000_6462, w_000_6463, w_000_6464, w_000_6465, w_000_6466, w_000_6467, w_000_6468, w_000_6469, w_000_6470, w_000_6471, w_000_6472, w_000_6473, w_000_6474, w_000_6475, w_000_6476, w_000_6477, w_000_6478, w_000_6479, w_000_6480, w_000_6481, w_000_6482, w_000_6483, w_000_6484, w_000_6485, w_000_6486, w_000_6487, w_000_6488, w_000_6489, w_000_6490, w_000_6491, w_000_6492, w_000_6493, w_000_6494, w_000_6495, w_000_6496, w_000_6497, w_000_6498, w_000_6499, w_000_6500, w_000_6501, w_000_6502, w_000_6503, w_000_6504, w_000_6505, w_000_6506, w_000_6507, w_000_6508, w_000_6509, w_000_6510, w_000_6511, w_000_6512, w_000_6513, w_000_6514, w_000_6515, w_000_6516, w_000_6517, w_000_6518, w_000_6519, w_000_6520, w_000_6521, w_000_6522, w_000_6523, w_000_6524, w_000_6525, w_000_6526, w_000_6527, w_000_6528, w_000_6529, w_000_6530, w_000_6531, w_000_6532, w_000_6533, w_000_6534, w_000_6535, w_000_6536, w_000_6537, w_000_6538, w_000_6539, w_000_6540, w_000_6541, w_000_6542, w_000_6543, w_000_6544, w_000_6545, w_000_6546, w_000_6547, w_000_6548, w_000_6549, w_000_6550, w_000_6551, w_000_6552, w_000_6553, w_000_6554, w_000_6555, w_000_6556, w_000_6557, w_000_6558, w_000_6559, w_000_6560, w_000_6561, w_000_6562, w_000_6563, w_000_6564, w_000_6565, w_000_6566, w_000_6567, w_000_6568, w_000_6569, w_000_6570, w_000_6571, w_000_6572, w_000_6573, w_000_6574, w_000_6575, w_000_6576, w_000_6577, w_000_6578, w_000_6579, w_000_6580, w_000_6581, w_000_6582, w_000_6583, w_000_6584, w_000_6585, w_000_6586, w_000_6587, w_000_6588, w_000_6589, w_000_6590, w_000_6591, w_000_6592, w_000_6593, w_000_6594, w_000_6595, w_000_6596, w_000_6597, w_000_6598, w_000_6599, w_000_6600, w_000_6601, w_000_6602, w_000_6603, w_000_6604, w_000_6605, w_000_6606, w_000_6607, w_000_6608, w_000_6609, w_000_6610, w_000_6611, w_000_6612, w_000_6613, w_000_6614, w_000_6615, w_000_6616, w_000_6617, w_000_6618, w_000_6619, w_000_6620, w_000_6621, w_000_6622, w_000_6623, w_000_6624, w_000_6625, w_000_6626, w_000_6627, w_000_6628, w_000_6629, w_000_6630, w_000_6631, w_000_6632, w_000_6633, w_000_6634, w_000_6635, w_000_6636, w_000_6637, w_000_6638, w_000_6639, w_000_6640, w_000_6641, w_000_6642, w_000_6643, w_000_6644, w_000_6645, w_000_6646, w_000_6647, w_000_6648, w_000_6649, w_000_6650, w_000_6651, w_000_6652, w_000_6653, w_000_6654, w_000_6655, w_000_6656, w_000_6657, w_000_6658, w_000_6659, w_000_6660, w_000_6661, w_000_6662, w_000_6663, w_000_6664, w_000_6665, w_000_6666, w_000_6667, w_000_6668, w_000_6669, w_000_6670, w_000_6671, w_000_6672, w_000_6673, w_000_6674, w_000_6675, w_000_6676, w_000_6677, w_000_6678, w_000_6679, w_000_6680, w_000_6681, w_000_6682, w_000_6683, w_000_6684, w_000_6685, w_000_6686, w_000_6687, w_000_6688, w_000_6689, w_000_6690, w_000_6691, w_000_6692, w_000_6693, w_000_6694, w_000_6695, w_000_6696, w_000_6697, w_000_6698, w_000_6699, w_000_6700, w_000_6701, w_000_6702, w_000_6703, w_000_6704, w_000_6705, w_000_6706, w_000_6707, w_000_6708, w_000_6709, w_000_6710, w_000_6711, w_000_6712, w_000_6714, w_000_6715, w_000_6716, w_000_6717, w_000_6718, w_000_6719, w_000_6720, w_000_6721, w_000_6722, w_000_6723, w_000_6724, w_000_6725, w_000_6726, w_000_6727, w_000_6728, w_000_6729, w_000_6730, w_000_6731, w_000_6732, w_000_6733, w_000_6734, w_000_6735, w_000_6736, w_000_6737, w_000_6738, w_000_6739, w_000_6740, w_000_6741, w_000_6742, w_000_6743, w_000_6744, w_000_6745, w_000_6746, w_000_6747, w_000_6748, w_000_6749, w_000_6750, w_000_6751, w_000_6752, w_000_6753, w_000_6754, w_000_6755, w_000_6756, w_000_6757, w_000_6758, w_000_6759, w_000_6760, w_000_6761, w_000_6762, w_000_6763, w_000_6764, w_000_6765, w_000_6766, w_000_6767, w_000_6768, w_000_6769, w_000_6770, w_000_6771, w_000_6772, w_000_6773, w_000_6774, w_000_6775, w_000_6776, w_000_6777, w_000_6778, w_000_6779, w_000_6780, w_000_6781, w_000_6782, w_000_6783, w_000_6784, w_000_6785, w_000_6786, w_000_6787, w_000_6788, w_000_6789, w_000_6790, w_000_6791, w_000_6792, w_000_6793, w_000_6794, w_000_6795, w_000_6796, w_000_6797, w_000_6798, w_000_6799, w_000_6800, w_000_6801, w_000_6802, w_000_6803, w_000_6804, w_000_6805, w_000_6806, w_000_6807, w_000_6808, w_000_6809, w_000_6810, w_000_6811, w_000_6812, w_000_6813, w_000_6814, w_000_6815, w_000_6816, w_000_6817, w_000_6818, w_000_6819, w_000_6820, w_000_6821, w_000_6822, w_000_6823, w_000_6824, w_000_6825, w_000_6826, w_000_6827, w_000_6828, w_000_6829, w_000_6830, w_000_6831, w_000_6832, w_000_6833, w_000_6834, w_000_6835, w_000_6836, w_000_6837, w_000_6838, w_000_6839, w_000_6840, w_000_6841, w_000_6842, w_000_6843, w_000_6844, w_000_6845, w_000_6846, w_000_6847, w_000_6848, w_000_6849, w_000_6850, w_000_6851, w_000_6852, w_000_6853, w_000_6854, w_000_6855, w_000_6856, w_000_6857, w_000_6858, w_000_6859, w_000_6860, w_000_6861, w_000_6862, w_000_6863, w_000_6864, w_000_6865, w_000_6866, w_000_6867, w_000_6868, w_000_6869, w_000_6870, w_000_6871, w_000_6872, w_000_6873, w_000_6874, w_000_6875, w_000_6876, w_000_6877, w_000_6878, w_000_6879, w_000_6880, w_000_6881, w_000_6882, w_000_6883, w_000_6884, w_000_6885, w_000_6886, w_000_6887, w_000_6888, w_000_6889, w_000_6890, w_000_6891, w_000_6892, w_000_6893, w_000_6894, w_000_6895, w_000_6896, w_000_6897, w_000_6898, w_000_6899, w_000_6900, w_000_6901, w_000_6902, w_000_6903, w_000_6904, w_000_6905, w_000_6906, w_000_6907, w_000_6908, w_000_6909, w_000_6910, w_000_6911, w_000_6912, w_000_6913, w_000_6914, w_000_6915, w_000_6916, w_000_6917, w_000_6918, w_000_6919, w_000_6920, w_000_6921, w_000_6922, w_000_6923, w_000_6924, w_000_6925, w_000_6926, w_000_6927, w_000_6928, w_000_6929, w_000_6930, w_000_6931, w_000_6932, w_000_6933, w_000_6934, w_000_6935, w_000_6936, w_000_6937, w_000_6938, w_000_6939, w_000_6940, w_000_6941, w_000_6942, w_000_6943, w_000_6944, w_000_6945, w_000_6946, w_000_6947, w_000_6948, w_000_6949, w_000_6950, w_000_6951, w_000_6952, w_000_6953, w_000_6954, w_000_6955, w_000_6956, w_000_6957, w_000_6958, w_000_6959, w_000_6960, w_000_6961, w_000_6962, w_000_6963, w_000_6964, w_000_6965, w_000_6966, w_000_6967, w_000_6968, w_000_6969, w_000_6970, w_000_6971, w_000_6972, w_000_6973, w_000_6974, w_000_6975, w_000_6976, w_000_6977, w_000_6978, w_000_6979, w_000_6980, w_000_6981, w_000_6982, w_000_6983, w_000_6984, w_000_6985, w_000_6986, w_000_6987, w_000_6988, w_000_6989, w_000_6990, w_000_6991, w_000_6992, w_000_6993, w_000_6994, w_000_6995, w_000_6996, w_000_6997, w_000_6998, w_000_6999, w_000_7000, w_000_7001, w_000_7002, w_000_7003, w_000_7004, w_000_7005, w_000_7006, w_000_7007, w_000_7008, w_000_7009, w_000_7010, w_000_7011, w_000_7012, w_000_7013, w_000_7014, w_000_7015, w_000_7016, w_000_7017, w_000_7018, w_000_7019, w_000_7020, w_000_7021, w_000_7022, w_000_7023, w_000_7024, w_000_7025, w_000_7026, w_000_7027, w_000_7028, w_000_7029, w_000_7030, w_000_7031, w_000_7032, w_000_7033, w_000_7034, w_000_7035, w_000_7036, w_000_7037, w_000_7038, w_000_7039, w_000_7040, w_000_7041, w_000_7042, w_000_7043, w_000_7044, w_000_7045, w_000_7046, w_000_7047, w_000_7048, w_000_7049, w_000_7050, w_000_7051, w_000_7052, w_000_7053, w_000_7054, w_000_7055, w_000_7056, w_000_7057, w_000_7058, w_000_7059, w_000_7060, w_000_7061, w_000_7062, w_000_7063, w_000_7064, w_000_7065, w_000_7066, w_000_7067, w_000_7068, w_000_7069, w_000_7070, w_000_7071, w_000_7072, w_000_7073, w_000_7074, w_000_7075, w_000_7076, w_000_7077, w_000_7078, w_000_7079, w_000_7080, w_000_7081, w_000_7082, w_000_7083, w_000_7084, w_000_7085, w_000_7086, w_000_7087, w_000_7088, w_000_7089, w_000_7090, w_000_7091, w_000_7092, w_000_7093, w_000_7094, w_000_7095, w_000_7096, w_000_7097, w_000_7098, w_000_7099, w_000_7100, w_000_7101, w_000_7102, w_000_7103, w_000_7104, w_000_7105, w_000_7106, w_000_7107, w_000_7108, w_000_7109, w_000_7110, w_000_7111, w_000_7112, w_000_7113, w_000_7114, w_000_7115, w_000_7116, w_000_7117, w_000_7118, w_000_7119, w_000_7120, w_000_7121, w_000_7122, w_000_7123, w_000_7124, w_000_7125, w_000_7126, w_000_7127, w_000_7128, w_000_7129, w_000_7130, w_000_7131, w_000_7132, w_000_7133, w_000_7134, w_000_7135, w_000_7136, w_000_7137, w_000_7138, w_000_7139, w_000_7140, w_000_7141, w_000_7142, w_000_7143, w_000_7144, w_000_7145, w_000_7146, w_000_7147, w_000_7148, w_000_7149, w_000_7150, w_000_7151, w_000_7152, w_000_7153, w_000_7154, w_000_7155, w_000_7156, w_000_7157, w_000_7158, w_000_7159, w_000_7160, w_000_7161, w_000_7162, w_000_7163, w_000_7164, w_000_7165, w_000_7166, w_000_7167, w_000_7168, w_000_7169, w_000_7170, w_000_7171, w_000_7172, w_000_7173, w_000_7174, w_000_7175, w_000_7176, w_000_7177, w_000_7178, w_000_7179, w_000_7180, w_000_7181, w_000_7182, w_000_7183, w_000_7184, w_000_7185, w_000_7186, w_000_7187, w_000_7188, w_000_7189, w_000_7190, w_000_7191, w_000_7192, w_000_7193, w_000_7194, w_000_7195, w_000_7196, w_000_7197, w_000_7198, w_000_7199, w_000_7200, w_000_7201, w_000_7202, w_000_7203, w_000_7204, w_000_7205, w_000_7206, w_000_7207, w_000_7208, w_000_7209, w_000_7210, w_000_7211, w_000_7212, w_000_7213, w_000_7214, w_000_7215, w_000_7216, w_000_7217, w_000_7218, w_000_7219, w_000_7220, w_000_7221, w_000_7222, w_000_7223, w_000_7224, w_000_7225, w_000_7226, w_000_7227, w_000_7228, w_000_7229, w_000_7230, w_000_7231, w_000_7232, w_000_7233, w_000_7234, w_000_7235, w_000_7236, w_000_7237, w_000_7238, w_000_7239, w_000_7240, w_000_7241, w_000_7242, w_000_7243, w_000_7244, w_000_7245, w_000_7246, w_000_7247, w_000_7248, w_000_7249, w_000_7250, w_000_7251, w_000_7252, w_000_7253, w_000_7254, w_000_7255, w_000_7256, w_000_7257, w_000_7258, w_000_7259, w_000_7260, w_000_7261, w_000_7262, w_000_7263, w_000_7264, w_000_7265, w_000_7266, w_000_7267, w_000_7268, w_000_7269, w_000_7270, w_000_7271, w_000_7272, w_000_7273, w_000_7274, w_000_7275, w_000_7276, w_000_7277, w_000_7278, w_000_7279, w_000_7280, w_000_7281, w_000_7282, w_000_7283, w_000_7284, w_000_7285, w_000_7286, w_000_7287, w_000_7288, w_000_7289, w_000_7290, w_000_7291, w_000_7292, w_000_7293, w_000_7294, w_000_7295, w_000_7296, w_000_7297, w_000_7298, w_000_7299, w_000_7300, w_000_7301, w_000_7302, w_000_7303, w_000_7304, w_000_7305, w_000_7306, w_000_7307, w_000_7308, w_000_7309, w_000_7310, w_000_7311, w_000_7312, w_000_7313, w_000_7314, w_000_7315, w_000_7316, w_000_7317, w_000_7318, w_000_7319, w_000_7320, w_000_7321, w_000_7322, w_000_7323, w_000_7324, w_000_7325, w_000_7326, w_000_7327, w_000_7328, w_000_7329, w_000_7330, w_000_7331, w_000_7332, w_000_7333, w_000_7334, w_000_7335, w_000_7336, w_000_7337, w_000_7338, w_000_7339, w_000_7340, w_000_7341, w_000_7342, w_000_7343, w_000_7344, w_000_7345, w_000_7346, w_000_7347, w_000_7348, w_000_7349, w_000_7350, w_000_7351, w_000_7352, w_000_7353, w_000_7354, w_000_7355, w_000_7356, w_000_7357, w_000_7358, w_000_7359, w_000_7360, w_000_7361, w_000_7362, w_000_7363, w_000_7364, w_000_7365, w_000_7366, w_000_7367, w_000_7368, w_000_7369, w_000_7370, w_000_7371, w_000_7372, w_000_7373, w_000_7374, w_000_7375, w_000_7376, w_000_7377, w_000_7378, w_000_7379, w_000_7380, w_000_7381, w_000_7382, w_000_7383, w_000_7384, w_000_7385, w_000_7386, w_000_7387, w_000_7388, w_000_7389, w_000_7390, w_000_7391, w_000_7392, w_000_7393, w_000_7394, w_000_7395, w_000_7396, w_000_7397, w_000_7398, w_000_7399, w_000_7400, w_000_7401, w_000_7402, w_000_7403, w_000_7404, w_000_7405, w_000_7406, w_000_7407, w_000_7408, w_000_7409, w_000_7410, w_000_7411, w_000_7412, w_000_7413, w_000_7414, w_000_7415, w_000_7416, w_000_7417, w_000_7418, w_000_7419, w_000_7420, w_000_7421, w_000_7422, w_000_7423, w_000_7424, w_000_7425, w_000_7426, w_000_7427, w_000_7428, w_000_7429, w_000_7430, w_000_7431, w_000_7432, w_000_7433, w_000_7434, w_000_7435, w_000_7436, w_000_7437, w_000_7438, w_000_7439, w_000_7440, w_000_7441, w_000_7442, w_000_7443, w_000_7444, w_000_7445, w_000_7446, w_000_7447, w_000_7448, w_000_7449, w_000_7450, w_000_7451, w_000_7452, w_000_7453, w_000_7454, w_000_7455, w_000_7456, w_000_7457, w_000_7458, w_000_7459, w_000_7460, w_000_7461, w_000_7462, w_000_7463, w_000_7464, w_000_7465, w_000_7466, w_000_7467, w_000_7468, w_000_7469, w_000_7470, w_000_7471, w_000_7472, w_000_7473, w_000_7474, w_000_7475, w_000_7476, w_000_7477, w_000_7478, w_000_7479, w_000_7480, w_000_7481, w_000_7482, w_000_7483, w_000_7484, w_000_7485, w_000_7486, w_000_7487, w_000_7488, w_000_7489, w_000_7490, w_000_7491, w_000_7492, w_000_7493, w_000_7494, w_000_7495, w_000_7496, w_000_7497, w_000_7498, w_000_7499, w_000_7500, w_000_7501, w_000_7502, w_000_7503, w_000_7504, w_000_7505, w_000_7506, w_000_7507, w_000_7508, w_000_7509, w_000_7510, w_000_7511, w_000_7512, w_000_7513, w_000_7514, w_000_7515, w_000_7516, w_000_7517, w_000_7518, w_000_7519, w_000_7520, w_000_7521, w_000_7522, w_000_7523, w_000_7524, w_000_7525, w_000_7526, w_000_7527, w_000_7528, w_000_7529, w_000_7530, w_000_7531, w_000_7532, w_000_7533, w_000_7534, w_000_7535, w_000_7536, w_000_7537, w_000_7538, w_000_7539, w_000_7540, w_000_7541, w_000_7542, w_000_7543, w_000_7544, w_000_7545, w_000_7546, w_000_7547, w_000_7548, w_000_7549, w_000_7550, w_000_7551, w_000_7552, w_000_7553, w_000_7554, w_000_7555, w_000_7556, w_000_7557, w_000_7558, w_000_7559, w_000_7560, w_000_7561, w_000_7562, w_000_7563, w_000_7564, w_000_7565, w_000_7566, w_000_7567, w_000_7568, w_000_7569, w_000_7570, w_000_7571, w_000_7572, w_000_7573, w_000_7574, w_000_7575, w_000_7576, w_000_7577, w_000_7578, w_000_7579, w_000_7580, w_000_7581, w_000_7582, w_000_7583, w_000_7584, w_000_7585, w_000_7586, w_000_7587, w_000_7588, w_000_7589, w_000_7590, w_000_7591, w_000_7592, w_000_7593, w_000_7594, w_000_7595, w_000_7596, w_000_7597, w_000_7598, w_000_7599, w_000_7600, w_000_7601, w_000_7602, w_000_7603, w_000_7604, w_000_7605, w_000_7606, w_000_7607, w_000_7608, w_000_7610, w_000_7611, w_000_7612, w_000_7613, w_000_7614, w_000_7615, w_000_7616, w_000_7617, w_000_7618, w_000_7619, w_000_7620, w_000_7621, w_000_7622, w_000_7623, w_000_7624, w_000_7625, w_000_7626, w_000_7627, w_000_7628, w_000_7629, w_000_7630, w_000_7631, w_000_7632, w_000_7633, w_000_7634, w_000_7635, w_000_7636, w_000_7637, w_000_7638, w_000_7639, w_000_7640, w_000_7641, w_000_7642, w_000_7643, w_000_7644, w_000_7645, w_000_7646, w_000_7647, w_000_7648, w_000_7649, w_000_7650, w_000_7651, w_000_7652, w_000_7653, w_000_7654, w_000_7655, w_000_7656, w_000_7657, w_000_7658, w_000_7659, w_000_7660, w_000_7661, w_000_7662, w_000_7663, w_000_7664, w_000_7665, w_000_7666, w_000_7667, w_000_7668, w_000_7669, w_000_7670, w_000_7671, w_000_7672, w_000_7673, w_000_7674, w_000_7675, w_000_7676, w_000_7677, w_000_7678, w_000_7679, w_000_7680, w_000_7681, w_000_7682, w_000_7683, w_000_7684, w_000_7685, w_000_7686, w_000_7687, w_000_7688, w_000_7689, w_000_7690, w_000_7692, w_000_7693, w_000_7694, w_000_7695, w_000_7696, w_000_7697, w_000_7698, w_000_7699, w_000_7700, w_000_7701, w_000_7702, w_000_7703, w_000_7704, w_000_7705, w_000_7706, w_000_7707, w_000_7708, w_000_7709, w_000_7710, w_000_7711, w_000_7712, w_000_7713, w_000_7714, w_000_7715, w_000_7716, w_000_7717, w_000_7718, w_000_7719, w_000_7720, w_000_7721, w_000_7722, w_000_7723, w_000_7724, w_000_7725, w_000_7726, w_000_7727, w_000_7728, w_000_7729, w_000_7730, w_000_7731, w_000_7732, w_000_7733, w_000_7734, w_000_7735, w_000_7736, w_000_7737, w_000_7738, w_000_7739, w_000_7740, w_000_7741, w_000_7742, w_000_7743, w_000_7744, w_000_7745, w_000_7746, w_000_7747, w_000_7748, w_000_7749, w_000_7750, w_000_7751, w_000_7752, w_000_7753, w_000_7754, w_000_7755, w_000_7756, w_000_7757, w_000_7758, w_000_7759, w_000_7760, w_000_7761, w_000_7762, w_000_7763, w_000_7764, w_000_7765, w_000_7766, w_000_7767, w_000_7768, w_000_7769, w_000_7770, w_000_7771, w_000_7772, w_000_7773, w_000_7774, w_000_7775, w_000_7776, w_000_7777, w_000_7778, w_000_7779, w_000_7780, w_000_7781, w_000_7782, w_000_7784, w_000_7785, w_000_7786, w_000_7787, w_000_7788, w_000_7789, w_000_7790, w_000_7791, w_000_7792, w_000_7793, w_000_7794, w_000_7795, w_000_7796, w_000_7797, w_000_7799, w_000_7800, w_000_7801, w_000_7802, w_000_7803, w_000_7804, w_000_7805, w_000_7806, w_000_7807, w_000_7808, w_000_7809, w_000_7810, w_000_7811, w_000_7812, w_000_7813, w_000_7814, w_000_7815, w_000_7816, w_000_7817, w_000_7818, w_000_7819, w_000_7820, w_000_7821, w_000_7822, w_000_7823, w_000_7824, w_000_7825, w_000_7826, w_000_7827, w_000_7828, w_000_7829, w_000_7830, w_000_7831, w_000_7832, w_000_7833, w_000_7834, w_000_7835, w_000_7836, w_000_7837, w_000_7838, w_000_7839, w_000_7840, w_000_7841, w_000_7842, w_000_7843, w_000_7844, w_000_7845, w_000_7846, w_000_7847, w_000_7848, w_000_7849, w_000_7850, w_000_7851, w_000_7852, w_000_7853, w_000_7854, w_000_7855, w_000_7856, w_000_7857, w_000_7858, w_000_7859, w_000_7860, w_000_7861, w_000_7862, w_000_7863, w_000_7864, w_000_7865, w_000_7866, w_000_7867, w_000_7868, w_000_7869, w_000_7870, w_000_7871, w_000_7872, w_000_7874, w_000_7875, w_000_7876, w_000_7877, w_000_7878, w_000_7879, w_000_7880, w_000_7881, w_000_7882, w_000_7883, w_000_7884, w_000_7885, w_000_7886, w_000_7887, w_000_7888, w_000_7889, w_000_7890, w_000_7891, w_000_7892, w_000_7893, w_000_7894, w_000_7895, w_000_7896, w_000_7897, w_000_7898, w_000_7899, w_000_7900, w_000_7901, w_000_7902, w_000_7903, w_000_7904, w_000_7905, w_000_7906, w_000_7907, w_000_7908, w_000_7909, w_000_7910, w_000_7911, w_000_7912, w_000_7913, w_000_7914, w_000_7915, w_000_7916, w_000_7917, w_000_7918, w_000_7919, w_000_7920, w_000_7921, w_000_7922, w_000_7923, w_000_7924, w_000_7925, w_000_7926, w_000_7927, w_000_7928, w_000_7929, w_000_7930, w_000_7931, w_000_7932, w_000_7933, w_000_7934, w_000_7935, w_000_7936, w_000_7937, w_000_7938, w_000_7939, w_000_7940, w_000_7941, w_000_7942, w_000_7943, w_000_7944, w_000_7945, w_000_7946, w_000_7947, w_000_7948, w_000_7949, w_000_7950, w_000_7951, w_000_7952, w_000_7953, w_000_7954, w_000_7955, w_000_7956, w_000_7957, w_000_7958, w_000_7959, w_000_7960, w_000_7961, w_000_7962, w_000_7963, w_000_7964, w_000_7965, w_000_7966, w_000_7967, w_000_7968, w_000_7969, w_000_7970, w_000_7971, w_000_7972, w_000_7973, w_000_7974, w_000_7975, w_000_7976, w_000_7977, w_000_7978, w_000_7979, w_000_7980, w_000_7981, w_000_7982, w_000_7983, w_000_7984, w_000_7985, w_000_7986, w_000_7987, w_000_7988, w_000_7989, w_000_7990, w_000_7991, w_000_7992, w_000_7993, w_000_7994, w_000_7995, w_000_7996, w_000_7997, w_000_7998, w_000_7999, w_000_8000, w_000_8001, w_000_8002, w_000_8003, w_000_8004, w_000_8005, w_000_8006, w_000_8007, w_000_8008, w_000_8009, w_000_8010, w_000_8011, w_000_8012, w_000_8013, w_000_8014, w_000_8015, w_000_8016, w_000_8017, w_000_8018, w_000_8019, w_000_8020, w_000_8021, w_000_8022, w_000_8023, w_000_8024, w_000_8025, w_000_8026, w_000_8027, w_000_8028, w_000_8029, w_000_8030, w_000_8031, w_000_8032, w_000_8033, w_000_8034, w_000_8035, w_000_8036, w_000_8037, w_000_8038, w_000_8039, w_000_8040, w_000_8041, w_000_8042, w_000_8043, w_000_8044, w_000_8045, w_000_8046, w_000_8047, w_000_8048, w_000_8049, w_000_8050, w_000_8051, w_000_8052, w_000_8053, w_000_8054, w_000_8055, w_000_8056, w_000_8057, w_000_8058, w_000_8059, w_000_8060, w_000_8061, w_000_8062, w_000_8063, w_000_8064, w_000_8065, w_000_8066, w_000_8067, w_000_8068, w_000_8069, w_000_8070, w_000_8071, w_000_8072, w_000_8073, w_000_8074, w_000_8075, w_000_8076, w_000_8077, w_000_8078, w_000_8079, w_000_8080, w_000_8081, w_000_8082, w_000_8083, w_000_8084, w_000_8085, w_000_8086, w_000_8087, w_000_8088, w_000_8089, w_000_8090, w_000_8091, w_000_8092, w_000_8093, w_000_8094, w_000_8095, w_000_8096, w_000_8097, w_000_8098, w_000_8099, w_000_8100, w_000_8101, w_000_8102, w_000_8103, w_000_8104, w_000_8105, w_000_8106, w_000_8107, w_000_8108, w_000_8109, w_000_8110, w_000_8111, w_000_8112, w_000_8113, w_000_8114, w_000_8115, w_000_8116, w_000_8117, w_000_8118, w_000_8119, w_000_8120, w_000_8121, w_000_8122, w_000_8123, w_000_8124, w_000_8125, w_000_8126, w_000_8127, w_000_8128, w_000_8129, w_000_8130, w_000_8131, w_000_8132, w_000_8133, w_000_8134, w_000_8135, w_000_8136, w_000_8137, w_000_8138, w_000_8139, w_000_8140, w_000_8141, w_000_8142, w_000_8143, w_000_8144, w_000_8145, w_000_8146, w_000_8147, w_000_8148, w_000_8149, w_000_8150, w_000_8151, w_000_8152, w_000_8153, w_000_8154, w_000_8155, w_000_8156, w_000_8157, w_000_8158, w_000_8159, w_000_8160, w_000_8161, w_000_8162, w_000_8163, w_000_8164, w_000_8165, w_000_8166, w_000_8167, w_000_8168, w_000_8169, w_000_8170, w_000_8171, w_000_8172, w_000_8173, w_000_8174, w_000_8175, w_000_8176, w_000_8177, w_000_8178, w_000_8179, w_000_8180, w_000_8181, w_000_8182, w_000_8183, w_000_8184, w_000_8185, w_000_8186, w_000_8187, w_000_8188, w_000_8189, w_000_8190, w_000_8191, w_000_8192, w_000_8193, w_000_8194, w_000_8195, w_000_8196, w_000_8197, w_000_8198, w_000_8199, w_000_8200, w_000_8201, w_000_8202, w_000_8203, w_000_8204, w_000_8205, w_000_8206, w_000_8207, w_000_8208, w_000_8209, w_000_8210, w_000_8211, w_000_8212, w_000_8213, w_000_8214, w_000_8215, w_000_8216, w_000_8217, w_000_8218, w_000_8219, w_000_8220, w_000_8221, w_000_8222, w_000_8223, w_000_8224, w_000_8225, w_000_8226, w_000_8227, w_000_8228, w_000_8229, w_000_8230, w_000_8231, w_000_8232, w_000_8233, w_000_8234, w_000_8235, w_000_8236, w_000_8237, w_000_8238, w_000_8239, w_000_8240, w_000_8241, w_000_8242, w_000_8243, w_000_8244, w_000_8245, w_000_8246, w_000_8247, w_000_8248, w_000_8249, w_000_8250, w_000_8251, w_000_8252, w_000_8253, w_000_8254, w_000_8255, w_000_8256, w_000_8257, w_000_8258, w_000_8259, w_000_8260, w_000_8261, w_000_8262, w_000_8263, w_000_8264, w_000_8265, w_000_8266, w_000_8267, w_000_8268, w_000_8269, w_000_8270, w_000_8271, w_000_8272, w_000_8273, w_000_8274, w_000_8275, w_000_8276, w_000_8277, w_000_8278, w_000_8279, w_000_8280, w_000_8281, w_000_8282, w_000_8283, w_000_8284, w_000_8285, w_000_8286, w_000_8287, w_000_8288, w_000_8289, w_000_8290, w_000_8291, w_000_8292, w_000_8293, w_000_8294, w_000_8295, w_000_8296, w_000_8297, w_000_8298, w_000_8299, w_000_8300, w_000_8301, w_000_8302, w_000_8303, w_000_8304, w_000_8305, w_000_8306, w_000_8307, w_000_8308, w_000_8309, w_000_8310, w_000_8311, w_000_8312, w_000_8313, w_000_8314, w_000_8315, w_000_8316, w_000_8317, w_000_8318, w_000_8319, w_000_8320, w_000_8321, w_000_8322, w_000_8323, w_000_8324, w_000_8325, w_000_8326, w_000_8327, w_000_8328, w_000_8329, w_000_8330, w_000_8331, w_000_8332, w_000_8333, w_000_8334, w_000_8335, w_000_8336, w_000_8337, w_000_8338, w_000_8339, w_000_8340, w_000_8341, w_000_8342, w_000_8343, w_000_8344, w_000_8345, w_000_8346, w_000_8347, w_000_8348, w_000_8349, w_000_8350, w_000_8351, w_000_8352, w_000_8353, w_000_8354, w_000_8355, w_000_8356, w_000_8357, w_000_8358, w_000_8359, w_000_8360, w_000_8361, w_000_8362, w_000_8363, w_000_8364, w_000_8365, w_000_8366, w_000_8367, w_000_8368, w_000_8369, w_000_8370, w_000_8371, w_000_8372, w_000_8373, w_000_8374, w_000_8375, w_000_8376, w_000_8377, w_000_8378, w_000_8379, w_000_8380, w_000_8381, w_000_8382, w_000_8383, w_000_8384, w_000_8385, w_000_8386, w_000_8387, w_000_8388, w_000_8389, w_000_8390, w_000_8391, w_000_8392, w_000_8393, w_000_8394, w_000_8395, w_000_8396, w_000_8397, w_000_8398, w_000_8399, w_000_8400, w_000_8401, w_000_8402, w_000_8403, w_000_8404, w_000_8405, w_000_8406, w_000_8407, w_000_8408, w_000_8409, w_000_8410, w_000_8411, w_000_8412, w_000_8413, w_000_8414, w_000_8415, w_000_8416, w_000_8417, w_000_8418, w_000_8419, w_000_8420, w_000_8421, w_000_8422, w_000_8423, w_000_8424, w_000_8425, w_000_8426, w_000_8427, w_000_8428, w_000_8429, w_000_8430, w_000_8431, w_000_8432, w_000_8433, w_000_8434, w_000_8435, w_000_8436, w_000_8437, w_000_8438, w_000_8439, w_000_8440, w_000_8441, w_000_8442, w_000_8443, w_000_8444, w_000_8445, w_000_8446, w_000_8447, w_000_8448, w_000_8449, w_000_8450, w_000_8451, w_000_8452, w_000_8453, w_000_8454, w_000_8455, w_000_8456, w_000_8457, w_000_8458, w_000_8459, w_000_8460, w_000_8461, w_000_8462, w_000_8463, w_000_8464, w_000_8465, w_000_8466, w_000_8467, w_000_8468, w_000_8469, w_000_8470, w_000_8471, w_000_8472, w_000_8473, w_000_8474, w_000_8475, w_000_8476, w_000_8477, w_000_8478, w_000_8479, w_000_8480, w_000_8481, w_000_8482, w_000_8483, w_000_8484, w_000_8485, w_000_8486, w_000_8487, w_000_8488, w_000_8489, w_000_8490, w_000_8491, w_000_8492, w_000_8493, w_000_8494, w_000_8495, w_000_8496, w_000_8497, w_000_8498, w_000_8499, w_000_8500, w_000_8501, w_000_8502, w_000_8503, w_000_8504, w_000_8505, w_000_8506, w_000_8507, w_000_8508, w_000_8509, w_000_8510, w_000_8511, w_000_8512, w_000_8513, w_000_8514, w_000_8515, w_000_8516, w_000_8517, w_000_8518, w_000_8519, w_000_8520, w_000_8521, w_000_8522, w_000_8523, w_000_8524, w_000_8525, w_000_8526, w_000_8527, w_000_8528, w_000_8529, w_000_8530, w_000_8531, w_000_8532, w_000_8533, w_000_8534, w_000_8535, w_000_8536, w_000_8537, w_000_8538, w_000_8539, w_000_8540, w_000_8541, w_000_8542, w_000_8543, w_000_8544, w_000_8545, w_000_8546, w_000_8547, w_000_8548, w_000_8549, w_000_8550, w_000_8551, w_000_8552, w_000_8553, w_000_8554, w_000_8555, w_000_8556, w_000_8557, w_000_8558, w_000_8559, w_000_8560, w_000_8561, w_000_8562, w_000_8563, w_000_8564, w_000_8565, w_000_8566, w_000_8567, w_000_8568, w_000_8569, w_000_8570, w_000_8571, w_000_8572, w_000_8573, w_000_8574, w_000_8575, w_000_8576, w_000_8577, w_000_8578, w_000_8579, w_000_8580, w_000_8581, w_000_8582, w_000_8583, w_000_8584, w_000_8585, w_000_8586, w_000_8587, w_000_8588, w_000_8589, w_000_8590, w_000_8591, w_000_8592, w_000_8593, w_000_8594, w_000_8595, w_000_8596, w_000_8597, w_000_8598, w_000_8599, w_000_8600, w_000_8601, w_000_8602, w_000_8603, w_000_8604, w_000_8605, w_000_8606, w_000_8607, w_000_8608, w_000_8609, w_000_8610, w_000_8611, w_000_8612, w_000_8613, w_000_8614, w_000_8615, w_000_8616, w_000_8617, w_000_8618, w_000_8619, w_000_8620, w_000_8621, w_000_8622, w_000_8623, w_000_8624, w_000_8625, w_000_8626, w_000_8627, w_000_8628, w_000_8629, w_000_8630, w_000_8631, w_000_8632, w_000_8633, w_000_8634, w_000_8635, w_000_8636, w_000_8637, w_000_8638, w_000_8639, w_000_8640, w_000_8641, w_000_8642, w_000_8643, w_000_8644, w_000_8645, w_000_8646, w_000_8647, w_000_8648, w_000_8649, w_000_8650, w_000_8651, w_000_8652, w_000_8653, w_000_8654, w_000_8655, w_000_8656, w_000_8657, w_000_8658, w_000_8659, w_000_8660, w_000_8661, w_000_8662, w_000_8663, w_000_8664, w_000_8665, w_000_8666, w_000_8667, w_000_8668, w_000_8669, w_000_8670, w_000_8671, w_000_8672, w_000_8673, w_000_8674, w_000_8675, w_000_8676, w_000_8677, w_000_8678, w_000_8679, w_000_8680, w_000_8681, w_000_8682, w_000_8683, w_000_8684, w_000_8685, w_000_8686, w_000_8687, w_000_8688, w_000_8689, w_000_8690, w_000_8691, w_000_8692, w_000_8693, w_000_8694, w_000_8695, w_000_8696, w_000_8697, w_000_8698, w_000_8699, w_000_8700, w_000_8701, w_000_8702, w_000_8703, w_000_8704, w_000_8705, w_000_8706, w_000_8707, w_000_8708, w_000_8709, w_000_8710, w_000_8711, w_000_8712, w_000_8713, w_000_8714, w_000_8715, w_000_8716, w_000_8717, w_000_8718, w_000_8719, w_000_8720, w_000_8721, w_000_8722, w_000_8723, w_000_8724, w_000_8725, w_000_8726, w_000_8728, w_000_8729, w_000_8730, w_000_8731, w_000_8732, w_000_8733, w_000_8734, w_000_8735, w_000_8736, w_000_8737, w_000_8738, w_000_8739, w_000_8740, w_000_8741, w_000_8742, w_000_8743, w_000_8744, w_000_8745, w_000_8746, w_000_8747, w_000_8748, w_000_8749, w_000_8751, w_000_8752, w_000_8753, w_000_8754, w_000_8755, w_000_8756, w_000_8757, w_000_8758, w_000_8759, w_000_8760, w_000_8761, w_000_8762, w_000_8763, w_000_8764, w_000_8765, w_000_8766, w_000_8767, w_000_8768, w_000_8769, w_000_8770, w_000_8771, w_000_8772, w_000_8773, w_000_8774, w_000_8775, w_000_8776, w_000_8777, w_000_8778, w_000_8779, w_000_8780, w_000_8781, w_000_8782, w_000_8783, w_000_8784, w_000_8785, w_000_8786, w_000_8787, w_000_8788, w_000_8789, w_000_8790, w_000_8791, w_000_8792, w_000_8793, w_000_8794, w_000_8795, w_000_8796, w_000_8797, w_000_8798, w_000_8799, w_000_8800, w_000_8801, w_000_8802, w_000_8803, w_000_8804, w_000_8805, w_000_8806, w_000_8807, w_000_8808, w_000_8809, w_000_8810, w_000_8811, w_000_8812, w_000_8813, w_000_8814, w_000_8815, w_000_8816, w_000_8817, w_000_8818, w_000_8819, w_000_8820, w_000_8821, w_000_8822, w_000_8823, w_000_8824, w_000_8825, w_000_8826, w_000_8827, w_000_8828, w_000_8829, w_000_8830, w_000_8831, w_000_8832, w_000_8833, w_000_8834, w_000_8835, w_000_8836, w_000_8837, w_000_8838, w_000_8839, w_000_8840, w_000_8841, w_000_8842, w_000_8843, w_000_8844, w_000_8845, w_000_8846, w_000_8848, w_000_8849, w_000_8850, w_000_8851, w_000_8852, w_000_8853, w_000_8854, w_000_8855, w_000_8856, w_000_8857, w_000_8858, w_000_8859, w_000_8860, w_000_8861, w_000_8862, w_000_8863, w_000_8864, w_000_8865, w_000_8866, w_000_8867, w_000_8868, w_000_8869, w_000_8870, w_000_8871, w_000_8872, w_000_8873, w_000_8874, w_000_8875, w_000_8876, w_000_8877, w_000_8878, w_000_8879, w_000_8880, w_000_8881, w_000_8882, w_000_8883, w_000_8884, w_000_8885, w_000_8886, w_000_8887, w_000_8888, w_000_8889, w_000_8891, w_000_8892, w_000_8893, w_000_8894, w_000_8895, w_000_8896, w_000_8897, w_000_8898, w_000_8899, w_000_8900, w_000_8901, w_000_8902, w_000_8903, w_000_8904, w_000_8905, w_000_8906, w_000_8907, w_000_8908, w_000_8909, w_000_8910, w_000_8911, w_000_8912, w_000_8913, w_000_8914, w_000_8916, w_000_8917, w_000_8918, w_000_8919, w_000_8920, w_000_8921, w_000_8922, w_000_8923, w_000_8924, w_000_8925, w_000_8926, w_000_8927, w_000_8928, w_000_8929, w_000_8930, w_000_8931, w_000_8932, w_000_8933, w_000_8934, w_000_8935, w_000_8936, w_000_8937, w_000_8938, w_000_8939, w_000_8940, w_000_8941, w_000_8942, w_000_8943, w_000_8944, w_000_8945, w_000_8946, w_000_8947, w_000_8948, w_000_8949, w_000_8950, w_000_8951, w_000_8952, w_000_8953, w_000_8954, w_000_8955, w_000_8956, w_000_8957, w_000_8958, w_000_8959, w_000_8960, w_000_8961, w_000_8962, w_000_8963, w_000_8964, w_000_8965, w_000_8966, w_000_8967, w_000_8968, w_000_8969, w_000_8970, w_000_8971, w_000_8972, w_000_8973, w_000_8974, w_000_8975, w_000_8976, w_000_8977, w_000_8978, w_000_8979, w_000_8980, w_000_8981, w_000_8982, w_000_8983, w_000_8984, w_000_8985, w_000_8986, w_000_8987, w_000_8988, w_000_8989, w_000_8990, w_000_8991, w_000_8992, w_000_8993, w_000_8994, w_000_8995, w_000_8996, w_000_8997, w_000_8998, w_000_8999, w_000_9000, w_000_9001, w_000_9002, w_000_9003, w_000_9004, w_000_9005, w_000_9006, w_000_9007, w_000_9008, w_000_9009, w_000_9010, w_000_9011, w_000_9012, w_000_9013, w_000_9014, w_000_9015, w_000_9016, w_000_9017, w_000_9018, w_000_9019, w_000_9020, w_000_9021, w_000_9022, w_000_9023, w_000_9024, w_000_9025, w_000_9026, w_000_9027, w_000_9028, w_000_9029, w_000_9030, w_000_9031, w_000_9032, w_000_9033, w_000_9034, w_000_9035, w_000_9036, w_000_9037, w_000_9038, w_000_9039, w_000_9040, w_000_9041, w_000_9042, w_000_9043, w_000_9044, w_000_9045, w_000_9046, w_000_9047, w_000_9048, w_000_9049, w_000_9050, w_000_9051, w_000_9052, w_000_9053, w_000_9054, w_000_9055, w_000_9056, w_000_9057, w_000_9058, w_000_9059, w_000_9060, w_000_9061, w_000_9062, w_000_9063, w_000_9064, w_000_9065, w_000_9066, w_000_9067, w_000_9068, w_000_9069, w_000_9070, w_000_9071, w_000_9072, w_000_9073, w_000_9074, w_000_9075, w_000_9076, w_000_9077, w_000_9078, w_000_9079, w_000_9080, w_000_9081, w_000_9082, w_000_9083, w_000_9084, w_000_9085, w_000_9086, w_000_9087, w_000_9088, w_000_9089, w_000_9090, w_000_9091, w_000_9092, w_000_9093, w_000_9094, w_000_9095, w_000_9096, w_000_9097, w_000_9098, w_000_9099, w_000_9100, w_000_9101, w_000_9102, w_000_9103, w_000_9104, w_000_9105, w_000_9106, w_000_9107, w_000_9108, w_000_9109, w_000_9110, w_000_9111, w_000_9112, w_000_9113, w_000_9114, w_000_9115, w_000_9116, w_000_9117, w_000_9118, w_000_9119, w_000_9120, w_000_9121, w_000_9122, w_000_9123, w_000_9124, w_000_9125, w_000_9126, w_000_9127, w_000_9128, w_000_9129, w_000_9130, w_000_9131, w_000_9132, w_000_9133, w_000_9134, w_000_9135, w_000_9136, w_000_9137, w_000_9138, w_000_9139, w_000_9140, w_000_9141, w_000_9142, w_000_9143, w_000_9144, w_000_9145, w_000_9146, w_000_9147, w_000_9148, w_000_9149, w_000_9150, w_000_9151, w_000_9152, w_000_9153, w_000_9154, w_000_9155, w_000_9156, w_000_9157, w_000_9158, w_000_9159, w_000_9160, w_000_9161, w_000_9162, w_000_9163, w_000_9164, w_000_9165, w_000_9166, w_000_9167, w_000_9168, w_000_9169, w_000_9170, w_000_9171, w_000_9172, w_000_9173, w_000_9174, w_000_9175, w_000_9176, w_000_9177, w_000_9178, w_000_9179, w_000_9180, w_000_9181, w_000_9182, w_000_9183, w_000_9184, w_000_9185, w_000_9186, w_000_9187, w_000_9188, w_000_9189, w_000_9190, w_000_9191, w_000_9192, w_000_9193, w_000_9194, w_000_9195, w_000_9196, w_000_9197, w_000_9198, w_000_9199, w_000_9200, w_000_9201, w_000_9202, w_000_9203, w_000_9204, w_000_9205, w_000_9206, w_000_9207, w_000_9208, w_000_9209, w_000_9210, w_000_9211, w_000_9212, w_000_9213, w_000_9214, w_000_9215, w_000_9216, w_000_9217, w_000_9218, w_000_9219, w_000_9220, w_000_9221, w_000_9222, w_000_9223, w_000_9224, w_000_9225, w_000_9226, w_000_9227, w_000_9228, w_000_9229, w_000_9230, w_000_9231, w_000_9232, w_000_9233, w_000_9234, w_000_9235, w_000_9236, w_000_9237, w_000_9238, w_000_9239, w_000_9240, w_000_9241, w_000_9242, w_000_9243, w_000_9244, w_000_9245, w_000_9246, w_000_9247, w_000_9248, w_000_9249, w_000_9250, w_000_9251, w_000_9252, w_000_9253, w_000_9254, w_000_9255, w_000_9256, w_000_9257, w_000_9258, w_000_9259, w_000_9260, w_000_9261, w_000_9262, w_000_9263, w_000_9264, w_000_9265, w_000_9266, w_000_9267, w_000_9268, w_000_9269, w_000_9270, w_000_9271, w_000_9272, w_000_9273, w_000_9274, w_000_9275, w_000_9276, w_000_9277, w_000_9278, w_000_9279, w_000_9280, w_000_9281, w_000_9282, w_000_9283, w_000_9284, w_000_9285, w_000_9286, w_000_9287, w_000_9288, w_000_9289, w_000_9290, w_000_9291, w_000_9292, w_000_9293, w_000_9294, w_000_9295, w_000_9296, w_000_9297, w_000_9298, w_000_9299, w_000_9300, w_000_9301, w_000_9302, w_000_9303, w_000_9304, w_000_9305, w_000_9306, w_000_9307, w_000_9308, w_000_9309, w_000_9310, w_000_9311, w_000_9312, w_000_9313, w_000_9314, w_000_9315, w_000_9316, w_000_9317, w_000_9318, w_000_9319, w_000_9320, w_000_9321, w_000_9322, w_000_9323, w_000_9324, w_000_9325, w_000_9326, w_000_9327, w_000_9328, w_000_9329, w_000_9330, w_000_9331, w_000_9332, w_000_9333, w_000_9334, w_000_9335, w_000_9336, w_000_9337, w_000_9338, w_000_9339, w_000_9340, w_000_9341, w_000_9342, w_000_9343, w_000_9344, w_000_9345, w_000_9346, w_000_9347, w_000_9348, w_000_9349, w_000_9350, w_000_9351, w_000_9352, w_000_9353, w_000_9354, w_000_9355, w_000_9356, w_000_9357, w_000_9358, w_000_9359, w_000_9360, w_000_9361, w_000_9362, w_000_9363, w_000_9364, w_000_9365, w_000_9366, w_000_9367, w_000_9368, w_000_9369, w_000_9370, w_000_9371, w_000_9372, w_000_9373, w_000_9374, w_000_9375, w_000_9376, w_000_9377, w_000_9378, w_000_9379, w_000_9380, w_000_9381, w_000_9382, w_000_9383, w_000_9384, w_000_9385, w_000_9386, w_000_9387, w_000_9388, w_000_9389, w_000_9390, w_000_9391, w_000_9392, w_000_9393, w_000_9394, w_000_9395, w_000_9396, w_000_9397, w_000_9398, w_000_9399, w_000_9400, w_000_9401, w_000_9402, w_000_9403, w_000_9404, w_000_9405, w_000_9406, w_000_9407, w_000_9408, w_000_9409, w_000_9410, w_000_9411, w_000_9412, w_000_9413, w_000_9414, w_000_9415, w_000_9416, w_000_9417, w_000_9418, w_000_9419, w_000_9420, w_000_9421, w_000_9422, w_000_9423, w_000_9424, w_000_9425, w_000_9426, w_000_9427, w_000_9428, w_000_9429, w_000_9430, w_000_9431, w_000_9432, w_000_9433, w_000_9434, w_000_9435, w_000_9436, w_000_9437, w_000_9438, w_000_9439, w_000_9440, w_000_9441, w_000_9442, w_000_9443, w_000_9444, w_000_9445, w_000_9446, w_000_9447, w_000_9448, w_000_9449, w_000_9450, w_000_9451, w_000_9452, w_000_9453, w_000_9454, w_000_9455, w_000_9456, w_000_9457, w_000_9458, w_000_9459, w_000_9460, w_000_9461, w_000_9462, w_000_9463, w_000_9464, w_000_9465, w_000_9466, w_000_9467, w_000_9468, w_000_9469, w_000_9470, w_000_9471, w_000_9472, w_000_9473, w_000_9474, w_000_9475, w_000_9476, w_000_9477, w_000_9478, w_000_9479, w_000_9480, w_000_9481, w_000_9482, w_000_9483, w_000_9484, w_000_9485, w_000_9486, w_000_9487, w_000_9488, w_000_9489, w_000_9490, w_000_9491, w_000_9492, w_000_9493, w_000_9494, w_000_9495, w_000_9496, w_000_9497, w_000_9498, w_000_9499, w_000_9500, w_000_9501, w_000_9502, w_000_9504, w_000_9505, w_000_9506, w_000_9507, w_000_9508, w_000_9509, w_000_9510, w_000_9511, w_000_9512, w_000_9513, w_000_9514, w_000_9515, w_000_9516, w_000_9517, w_000_9518, w_000_9519, w_000_9520, w_000_9521, w_000_9522, w_000_9523, w_000_9524, w_000_9525, w_000_9526, w_000_9527, w_000_9528, w_000_9529, w_000_9530, w_000_9531, w_000_9532, w_000_9533, w_000_9534, w_000_9535, w_000_9536, w_000_9537, w_000_9538, w_000_9539, w_000_9540, w_000_9541, w_000_9542, w_000_9543, w_000_9544, w_000_9545, w_000_9547, w_000_9548, w_000_9549, w_000_9550, w_000_9551, w_000_9552, w_000_9554, w_000_9555, w_000_9556, w_000_9557, w_000_9558, w_000_9559, w_000_9560, w_000_9561, w_000_9563, w_000_9564, w_000_9565, w_000_9566, w_000_9567, w_000_9569, w_000_9570, w_000_9571, w_000_9572, w_000_9573, w_000_9574, w_000_9575, w_000_9576, w_000_9577, w_000_9578, w_000_9579, w_000_9580, w_000_9581, w_000_9582, w_000_9583, w_000_9584, w_000_9585, w_000_9586, w_000_9587, w_000_9588, w_000_9589, w_000_9590, w_000_9591, w_000_9592, w_000_9593, w_000_9594, w_000_9595, w_000_9596, w_000_9597, w_000_9598, w_000_9599, w_000_9600, w_000_9601, w_000_9602, w_000_9603, w_000_9604, w_000_9605, w_000_9606, w_000_9607, w_000_9608, w_000_9609, w_000_9610, w_000_9611, w_000_9612, w_000_9613, w_000_9614, w_000_9615, w_000_9616, w_000_9617, w_000_9618, w_000_9619, w_000_9620, w_000_9621, w_000_9622, w_000_9623, w_000_9624, w_000_9625, w_000_9626, w_000_9627, w_000_9628, w_000_9629, w_000_9630, w_000_9632, w_000_9633, w_000_9634, w_000_9635, w_000_9636, w_000_9637, w_000_9639, w_000_9640, w_000_9641, w_000_9642, w_000_9643, w_000_9644, w_000_9646, w_000_9647, w_000_9648, w_000_9649, w_000_9650, w_000_9651, w_000_9652, w_000_9653, w_000_9654, w_000_9655, w_000_9656, w_000_9657, w_000_9658, w_000_9659, w_000_9660, w_000_9661, w_000_9662, w_000_9663, w_000_9664, w_000_9666, w_000_9667, w_000_9668, w_000_9669, w_000_9670, w_000_9671, w_000_9672, w_000_9673, w_000_9674, w_000_9675, w_000_9676, w_000_9677, w_000_9678, w_000_9679, w_000_9682, w_000_9683, w_000_9684, w_000_9685, w_000_9686, w_000_9687, w_000_9688, w_000_9689, w_000_9690, w_000_9691, w_000_9692, w_000_9693, w_000_9694, w_000_9695, w_000_9696, w_000_9697, w_000_9698, w_000_9699, w_000_9701, w_000_9702, w_000_9704, w_000_9706, w_000_9708, w_000_9709, w_000_9710, w_000_9711, w_000_9713, w_000_9715, w_000_9716, w_000_9717, w_000_9719, w_000_9720, w_000_9721, w_000_9723, w_000_9725, w_000_9727, w_000_9728, w_000_9729, w_000_9730, w_000_9731, w_000_9732, w_000_9733, w_000_9734, w_000_9735, w_000_9736, w_000_9737, w_000_9738, w_000_9739, w_000_9740, w_000_9741, w_000_9742, w_000_9743, w_000_9744, w_000_9745, w_000_9747, w_000_9748, w_000_9749, w_000_9750, w_000_9752, w_000_9753, w_000_9754, w_000_9755, w_000_9756, w_000_9757, w_000_9758, w_000_9759, w_000_9760, w_000_9761, w_000_9765, w_000_9766, w_000_9767, w_000_9769, w_000_9770, w_000_9771, w_000_9772, w_000_9774, w_000_9776, w_000_9777, w_000_9778, w_000_9779, w_000_9780, w_000_9781, w_000_9782, w_000_9783, w_000_9785, w_000_9786, w_000_9788, w_000_9789, w_000_9790, w_000_9791, w_000_9792, w_000_9793, w_000_9794, w_000_9795, w_000_9796, w_000_9797, w_000_9798, w_000_9799, w_000_9800, w_000_9801, w_000_9802, w_000_9803, w_000_9804, w_000_9805, w_000_9806, w_000_9807, w_000_9808, w_000_9809, w_000_9810, w_000_9811, w_000_9812, w_000_9813, w_000_9814, w_000_9815, w_000_9816, w_000_9817, w_000_9819, w_000_9820, w_000_9821, w_000_9822, w_000_9823, w_000_9824, w_000_9825, w_000_9826, w_000_9827, w_000_9828, w_000_9829, w_000_9830, w_000_9831, w_000_9832, w_000_9833, w_000_9834, w_000_9835, w_000_9837, w_000_9838, w_000_9841, w_000_9842, w_000_9843, w_000_9844, w_000_9846, w_000_9847, w_000_9848, w_000_9849, w_000_9851, w_000_9853, w_000_9854, w_000_9855, w_000_9856, w_000_9857, w_000_9858, w_000_9859, w_000_9860, w_000_9861, w_000_9862, w_000_9864, w_000_9865, w_000_9866, w_000_9867, w_000_9871, w_000_9872, w_000_9874, w_000_9875, w_000_9877, w_000_9878, w_000_9879, w_000_9880, w_000_9882, w_000_9884, w_000_9887, w_000_9889, w_000_9890, w_000_9892, w_000_9893, w_000_9894, w_000_9895, w_000_9896, w_000_9897, w_000_9898, w_000_9899, w_000_9900, w_000_9902, w_000_9904, w_000_9905, w_000_9907, w_000_9908, w_000_9910, w_000_9914, w_000_9920, w_000_9922, w_000_9925, w_000_9926, w_000_9929, w_000_9930, w_000_9934, w_000_9936, w_000_9937, w_000_9938, w_000_9941, w_000_9949, w_000_9951, w_000_9958, w_000_9970, w_000_9978, w_000_9985, w_000_9996;
  output w_10000_000, w_10000_001, w_10000_002, w_10000_003, w_10000_004, w_10000_005, w_10000_006, w_10000_007, w_10000_008, w_10000_009, w_10000_010, w_10000_011, w_10000_012, w_10000_013, w_10000_014, w_10000_015, w_10000_016, w_10000_017, w_10000_018, w_10000_019, w_10000_020, w_10000_021, w_10000_022, w_10000_023, w_10000_024, w_10000_025, w_10000_026, w_10000_027, w_10000_028, w_10000_029, w_10000_030, w_10000_031, w_10000_032, w_10000_033, w_10000_034, w_10000_035, w_10000_036, w_10000_037, w_10000_038, w_10000_039, w_10000_040, w_10000_041, w_10000_042, w_10000_043, w_10000_044, w_10000_045, w_10000_046, w_10000_047, w_10000_048, w_10000_049, w_10000_050, w_10000_051, w_10000_052, w_10000_053, w_10000_054, w_10000_055, w_10000_056, w_10000_057, w_10000_058, w_10000_059, w_10000_060, w_10000_061, w_10000_062, w_10000_063, w_10000_064, w_10000_065, w_10000_066, w_10000_067, w_10000_068, w_10000_069, w_10000_070, w_10000_071, w_10000_072, w_10000_073, w_10000_074, w_10000_075, w_10000_076, w_10000_077, w_10000_078, w_10000_079, w_10000_080, w_10000_081, w_10000_082, w_10000_083, w_10000_084, w_10000_085, w_10000_086, w_10000_087, w_10000_088, w_10000_089, w_10000_090, w_10000_091, w_10000_092, w_10000_093, w_10000_094, w_10000_095, w_10000_096, w_10000_097, w_10000_098, w_10000_099, w_10000_100, w_10000_101, w_10000_102, w_10000_103, w_10000_104, w_10000_105, w_10000_106, w_10000_107, w_10000_108, w_10000_109, w_10000_110, w_10000_111, w_10000_112, w_10000_113, w_10000_114, w_10000_115, w_10000_116, w_10000_117, w_10000_118, w_10000_119, w_10000_120, w_10000_121, w_10000_122, w_10000_123, w_10000_124, w_10000_125, w_10000_126, w_10000_127, w_10000_128, w_10000_129, w_10000_130, w_10000_131, w_10000_132, w_10000_133, w_10000_134, w_10000_135, w_10000_136, w_10000_137, w_10000_138, w_10000_139, w_10000_140, w_10000_141, w_10000_142, w_10000_143, w_10000_144, w_10000_145, w_10000_146, w_10000_147, w_10000_148, w_10000_149, w_10000_150, w_10000_151, w_10000_152, w_10000_153, w_10000_154, w_10000_155, w_10000_156, w_10000_157, w_10000_158, w_10000_159, w_10000_160, w_10000_161, w_10000_162, w_10000_163, w_10000_164, w_10000_165, w_10000_166, w_10000_167, w_10000_168, w_10000_169, w_10000_170, w_10000_171, w_10000_172, w_10000_173, w_10000_174, w_10000_175, w_10000_176, w_10000_177, w_10000_178, w_10000_179, w_10000_180, w_10000_181, w_10000_182, w_10000_183, w_10000_184, w_10000_185, w_10000_186, w_10000_187, w_10000_188, w_10000_189, w_10000_190, w_10000_191, w_10000_192, w_10000_193, w_10000_194, w_10000_195, w_10000_196, w_10000_197, w_10000_198, w_10000_199, w_10000_200, w_10000_201, w_10000_202, w_10000_203, w_10000_204, w_10000_205, w_10000_206, w_10000_207, w_10000_208, w_10000_209, w_10000_210, w_10000_211, w_10000_212, w_10000_213, w_10000_214, w_10000_215, w_10000_216, w_10000_217, w_10000_218, w_10000_219, w_10000_220, w_10000_221, w_10000_222, w_10000_223, w_10000_224, w_10000_225, w_10000_226, w_10000_227, w_10000_228, w_10000_229, w_10000_230, w_10000_231, w_10000_232, w_10000_233, w_10000_234, w_10000_235, w_10000_236, w_10000_237, w_10000_238, w_10000_239, w_10000_240, w_10000_241, w_10000_242, w_10000_243, w_10000_244, w_10000_245, w_10000_246, w_10000_247, w_10000_248, w_10000_249, w_10000_250, w_10000_251, w_10000_252, w_10000_253, w_10000_254, w_10000_255, w_10000_256, w_10000_257, w_10000_258, w_10000_259, w_10000_260, w_10000_261, w_10000_262, w_10000_263, w_10000_264, w_10000_265, w_10000_266, w_10000_267, w_10000_268, w_10000_269, w_10000_270, w_10000_271, w_10000_272, w_10000_273, w_10000_274, w_10000_275, w_10000_276, w_10000_277, w_10000_278, w_10000_279, w_10000_280, w_10000_281, w_10000_282, w_10000_283, w_10000_284, w_10000_285, w_10000_286, w_10000_287, w_10000_288, w_10000_289, w_10000_290, w_10000_291, w_10000_292, w_10000_293, w_10000_294, w_10000_295, w_10000_296, w_10000_297, w_10000_298, w_10000_299, w_10000_300, w_10000_301, w_10000_302, w_10000_303, w_10000_304, w_10000_305, w_10000_306, w_10000_307, w_10000_308, w_10000_309, w_10000_310, w_10000_311, w_10000_312, w_10000_313, w_10000_314, w_10000_315, w_10000_316, w_10000_317, w_10000_318, w_10000_319, w_10000_320, w_10000_321, w_10000_322, w_10000_323, w_10000_324, w_10000_325, w_10000_326, w_10000_327, w_10000_328, w_10000_329, w_10000_330, w_10000_331, w_10000_332, w_10000_333, w_10000_334, w_10000_335, w_10000_336, w_10000_337, w_10000_338, w_10000_339, w_10000_340, w_10000_341, w_10000_342, w_10000_343, w_10000_344, w_10000_345, w_10000_346, w_10000_347, w_10000_348, w_10000_349, w_10000_350, w_10000_351, w_10000_352, w_10000_353, w_10000_354, w_10000_355, w_10000_356, w_10000_357, w_10000_358, w_10000_359, w_10000_360, w_10000_361, w_10000_362, w_10000_363, w_10000_364, w_10000_365, w_10000_366, w_10000_367, w_10000_368, w_10000_369, w_10000_370, w_10000_371, w_10000_372, w_10000_373, w_10000_374, w_10000_375, w_10000_376, w_10000_377, w_10000_378, w_10000_379, w_10000_380, w_10000_381, w_10000_382, w_10000_383, w_10000_384, w_10000_385, w_10000_386, w_10000_387, w_10000_388, w_10000_389, w_10000_390, w_10000_391, w_10000_392, w_10000_393, w_10000_394, w_10000_395, w_10000_396, w_10000_397, w_10000_398, w_10000_399, w_10000_400, w_10000_401, w_10000_402, w_10000_403, w_10000_404, w_10000_405, w_10000_406, w_10000_407, w_10000_408, w_10000_409, w_10000_410, w_10000_411, w_10000_412, w_10000_413, w_10000_414, w_10000_415, w_10000_416, w_10000_417, w_10000_418, w_10000_419, w_10000_420, w_10000_421, w_10000_422, w_10000_423, w_10000_424, w_10000_425, w_10000_426, w_10000_427, w_10000_428, w_10000_429, w_10000_430, w_10000_431, w_10000_432, w_10000_433, w_10000_434, w_10000_435, w_10000_436, w_10000_437, w_10000_438, w_10000_439, w_10000_440, w_10000_441, w_10000_442, w_10000_443, w_10000_444, w_10000_445, w_10000_446, w_10000_447, w_10000_448, w_10000_449, w_10000_450, w_10000_451, w_10000_452, w_10000_453, w_10000_454, w_10000_455, w_10000_456, w_10000_457, w_10000_458, w_10000_459, w_10000_460, w_10000_461, w_10000_462, w_10000_463, w_10000_464, w_10000_465, w_10000_466, w_10000_467, w_10000_468, w_10000_469, w_10000_470, w_10000_471, w_10000_472, w_10000_473, w_10000_474, w_10000_475, w_10000_476, w_10000_477, w_10000_478, w_10000_479, w_10000_480, w_10000_481, w_10000_482, w_10000_483, w_10000_484, w_10000_485, w_10000_486, w_10000_487, w_10000_488, w_10000_489, w_10000_490, w_10000_491, w_10000_492, w_10000_493, w_10000_494, w_10000_495, w_10000_496, w_10000_497, w_10000_498, w_10000_499, w_10000_500, w_10000_501, w_10000_502, w_10000_503, w_10000_504, w_10000_505, w_10000_506, w_10000_507, w_10000_508, w_10000_509, w_10000_510, w_10000_511, w_10000_512, w_10000_513, w_10000_514, w_10000_515, w_10000_516, w_10000_517, w_10000_518, w_10000_519, w_10000_520, w_10000_521, w_10000_522, w_10000_523, w_10000_524, w_10000_525, w_10000_526, w_10000_527, w_10000_528, w_10000_529, w_10000_530, w_10000_531, w_10000_532, w_10000_533, w_10000_534, w_10000_535, w_10000_536, w_10000_537, w_10000_538, w_10000_539, w_10000_540, w_10000_541, w_10000_542, w_10000_543, w_10000_544, w_10000_545, w_10000_546, w_10000_547, w_10000_548, w_10000_549, w_10000_550, w_10000_551, w_10000_552, w_10000_553, w_10000_554, w_10000_555, w_10000_556, w_10000_557, w_10000_558, w_10000_559, w_10000_560, w_10000_561, w_10000_562, w_10000_563, w_10000_564, w_10000_565, w_10000_566, w_10000_567, w_10000_568, w_10000_569, w_10000_570, w_10000_571, w_10000_572, w_10000_573, w_10000_574, w_10000_575, w_10000_576, w_10000_577, w_10000_578, w_10000_579, w_10000_580, w_10000_581, w_10000_582, w_10000_583, w_10000_584, w_10000_585, w_10000_586, w_10000_587, w_10000_588, w_10000_589, w_10000_590, w_10000_591, w_10000_592, w_10000_593, w_10000_594, w_10000_595, w_10000_596, w_10000_597, w_10000_598, w_10000_599, w_10000_600, w_10000_601, w_10000_602, w_10000_603, w_10000_604, w_10000_605, w_10000_606, w_10000_607, w_10000_608, w_10000_609, w_10000_610, w_10000_611, w_10000_612, w_10000_613, w_10000_614, w_10000_615, w_10000_616, w_10000_617, w_10000_618, w_10000_619, w_10000_620, w_10000_621, w_10000_622, w_10000_623, w_10000_624, w_10000_625, w_10000_626, w_10000_627, w_10000_628, w_10000_629, w_10000_630, w_10000_631, w_10000_632, w_10000_633, w_10000_634, w_10000_635, w_10000_636, w_10000_637, w_10000_638, w_10000_639, w_10000_640, w_10000_641, w_10000_642, w_10000_643, w_10000_644, w_10000_645, w_10000_646, w_10000_647, w_10000_648, w_10000_649, w_10000_650, w_10000_651, w_10000_652, w_10000_653, w_10000_654, w_10000_655, w_10000_656, w_10000_657, w_10000_658, w_10000_659, w_10000_660, w_10000_661, w_10000_662, w_10000_663, w_10000_664, w_10000_665, w_10000_666, w_10000_667, w_10000_668, w_10000_669, w_10000_670, w_10000_671, w_10000_672, w_10000_673, w_10000_674, w_10000_675, w_10000_676, w_10000_677, w_10000_678, w_10000_679, w_10000_680, w_10000_681, w_10000_682, w_10000_683, w_10000_684, w_10000_685, w_10000_686, w_10000_687, w_10000_688, w_10000_689, w_10000_690, w_10000_691, w_10000_692, w_10000_693, w_10000_694, w_10000_695, w_10000_696, w_10000_697, w_10000_698, w_10000_699, w_10000_700, w_10000_701, w_10000_702, w_10000_703, w_10000_704, w_10000_705, w_10000_706, w_10000_707, w_10000_708, w_10000_709, w_10000_710, w_10000_711, w_10000_712, w_10000_713, w_10000_714, w_10000_715, w_10000_716, w_10000_717, w_10000_718, w_10000_719, w_10000_720, w_10000_721, w_10000_722, w_10000_723, w_10000_724, w_10000_725, w_10000_726, w_10000_727, w_10000_728, w_10000_729, w_10000_730, w_10000_731, w_10000_732, w_10000_733, w_10000_734, w_10000_735, w_10000_736, w_10000_737, w_10000_738, w_10000_739, w_10000_740, w_10000_741, w_10000_742, w_10000_743, w_10000_744, w_10000_745, w_10000_746, w_10000_747, w_10000_748, w_10000_749, w_10000_750, w_10000_751, w_10000_752, w_10000_753, w_10000_754, w_10000_755, w_10000_756, w_10000_757, w_10000_758, w_10000_759, w_10000_760, w_10000_761, w_10000_762, w_10000_763, w_10000_764, w_10000_765, w_10000_766, w_10000_767, w_10000_768, w_10000_769, w_10000_770, w_10000_771, w_10000_772, w_10000_773, w_10000_774, w_10000_775, w_10000_776, w_10000_777, w_10000_778, w_10000_779, w_10000_780, w_10000_781, w_10000_782, w_10000_783, w_10000_784, w_10000_785, w_10000_786, w_10000_787, w_10000_788, w_10000_789, w_10000_790, w_10000_791, w_10000_792, w_10000_793, w_10000_794, w_10000_795, w_10000_796, w_10000_797, w_10000_798, w_10000_799, w_10000_800, w_10000_801, w_10000_802, w_10000_803, w_10000_804, w_10000_805, w_10000_806, w_10000_807, w_10000_808, w_10000_809, w_10000_810, w_10000_811, w_10000_812, w_10000_813, w_10000_814, w_10000_815, w_10000_816, w_10000_817, w_10000_818, w_10000_819, w_10000_820, w_10000_821, w_10000_822, w_10000_823, w_10000_824, w_10000_825, w_10000_826, w_10000_827, w_10000_828, w_10000_829, w_10000_830, w_10000_831, w_10000_832, w_10000_833, w_10000_834, w_10000_835, w_10000_836, w_10000_837, w_10000_838, w_10000_839, w_10000_840, w_10000_841, w_10000_842, w_10000_843, w_10000_844, w_10000_845, w_10000_846, w_10000_847, w_10000_848, w_10000_849, w_10000_850, w_10000_851, w_10000_852, w_10000_853, w_10000_854, w_10000_855, w_10000_856, w_10000_857, w_10000_858, w_10000_859, w_10000_860, w_10000_861, w_10000_862, w_10000_863, w_10000_864, w_10000_865, w_10000_866, w_10000_867, w_10000_868, w_10000_869, w_10000_870, w_10000_871, w_10000_872, w_10000_873, w_10000_874, w_10000_875, w_10000_876, w_10000_877, w_10000_878, w_10000_879, w_10000_880, w_10000_881, w_10000_882, w_10000_883, w_10000_884, w_10000_885, w_10000_886, w_10000_887, w_10000_888, w_10000_889, w_10000_890, w_10000_891, w_10000_892, w_10000_893, w_10000_894, w_10000_895, w_10000_896, w_10000_897, w_10000_898, w_10000_899, w_10000_900, w_10000_901, w_10000_902, w_10000_903, w_10000_904, w_10000_905, w_10000_906, w_10000_907, w_10000_908, w_10000_909, w_10000_910, w_10000_911, w_10000_912, w_10000_913, w_10000_914, w_10000_915, w_10000_916, w_10000_917, w_10000_918, w_10000_919, w_10000_920, w_10000_921, w_10000_922, w_10000_923, w_10000_924, w_10000_925, w_10000_926, w_10000_927, w_10000_928, w_10000_929, w_10000_930, w_10000_931, w_10000_932, w_10000_933, w_10000_934, w_10000_935, w_10000_936, w_10000_937, w_10000_938, w_10000_939, w_10000_940, w_10000_941, w_10000_942, w_10000_943, w_10000_944, w_10000_945, w_10000_946, w_10000_947, w_10000_948, w_10000_949, w_10000_950, w_10000_951, w_10000_952, w_10000_953, w_10000_954, w_10000_955, w_10000_956, w_10000_957, w_10000_958, w_10000_959, w_10000_960, w_10000_961, w_10000_962, w_10000_963, w_10000_964, w_10000_965, w_10000_966, w_10000_967, w_10000_968, w_10000_969, w_10000_970, w_10000_971, w_10000_972, w_10000_973, w_10000_974, w_10000_975, w_10000_976, w_10000_977, w_10000_978, w_10000_979, w_10000_980, w_10000_981, w_10000_982, w_10000_983, w_10000_984, w_10000_985, w_10000_986, w_10000_987, w_10000_988, w_10000_989, w_10000_990, w_10000_991, w_10000_992, w_10000_993, w_10000_994, w_10000_995, w_10000_996, w_10000_997, w_10000_998, w_10000_999, w_10000_1000, w_10000_1001, w_10000_1002, w_10000_1003, w_10000_1004, w_10000_1005, w_10000_1006, w_10000_1007, w_10000_1008, w_10000_1009, w_10000_1010, w_10000_1011, w_10000_1012, w_10000_1013, w_10000_1014, w_10000_1015, w_10000_1016, w_10000_1017, w_10000_1018, w_10000_1019, w_10000_1020, w_10000_1021, w_10000_1022, w_10000_1023, w_10000_1024, w_10000_1025, w_10000_1026, w_10000_1027, w_10000_1028, w_10000_1029, w_10000_1030, w_10000_1031, w_10000_1032, w_10000_1033, w_10000_1034, w_10000_1035, w_10000_1036, w_10000_1037, w_10000_1038, w_10000_1039, w_10000_1040, w_10000_1041, w_10000_1042, w_10000_1043, w_10000_1044, w_10000_1045, w_10000_1046, w_10000_1047, w_10000_1048, w_10000_1049, w_10000_1050, w_10000_1051, w_10000_1052, w_10000_1053, w_10000_1054, w_10000_1055, w_10000_1056, w_10000_1057, w_10000_1058, w_10000_1059, w_10000_1060, w_10000_1061, w_10000_1062, w_10000_1063, w_10000_1064, w_10000_1065, w_10000_1066, w_10000_1067, w_10000_1068, w_10000_1069, w_10000_1070, w_10000_1071, w_10000_1072, w_10000_1073, w_10000_1074, w_10000_1075, w_10000_1076, w_10000_1077, w_10000_1078, w_10000_1079, w_10000_1080, w_10000_1081, w_10000_1082, w_10000_1083, w_10000_1084, w_10000_1085, w_10000_1086, w_10000_1087, w_10000_1088, w_10000_1089, w_10000_1090, w_10000_1091, w_10000_1092, w_10000_1093, w_10000_1094, w_10000_1095, w_10000_1096, w_10000_1097, w_10000_1098, w_10000_1099, w_10000_1100, w_10000_1101, w_10000_1102, w_10000_1103, w_10000_1104, w_10000_1105, w_10000_1106, w_10000_1107, w_10000_1108, w_10000_1109, w_10000_1110, w_10000_1111, w_10000_1112, w_10000_1113, w_10000_1114, w_10000_1115, w_10000_1116, w_10000_1117, w_10000_1118, w_10000_1119, w_10000_1120, w_10000_1121, w_10000_1122, w_10000_1123, w_10000_1124, w_10000_1125, w_10000_1126, w_10000_1127, w_10000_1128, w_10000_1129, w_10000_1130, w_10000_1131, w_10000_1132, w_10000_1133, w_10000_1134, w_10000_1135, w_10000_1136, w_10000_1137, w_10000_1138, w_10000_1139, w_10000_1140, w_10000_1141, w_10000_1142, w_10000_1143, w_10000_1144, w_10000_1145, w_10000_1146, w_10000_1147, w_10000_1148, w_10000_1149, w_10000_1150, w_10000_1151, w_10000_1152, w_10000_1153, w_10000_1154, w_10000_1155, w_10000_1156, w_10000_1157, w_10000_1158, w_10000_1159, w_10000_1160, w_10000_1161, w_10000_1162, w_10000_1163, w_10000_1164, w_10000_1165, w_10000_1166, w_10000_1167, w_10000_1168, w_10000_1169, w_10000_1170, w_10000_1171, w_10000_1172, w_10000_1173, w_10000_1174, w_10000_1175, w_10000_1176, w_10000_1177, w_10000_1178, w_10000_1179, w_10000_1180, w_10000_1181, w_10000_1182, w_10000_1183, w_10000_1184, w_10000_1185, w_10000_1186, w_10000_1187, w_10000_1188, w_10000_1189, w_10000_1190, w_10000_1191, w_10000_1192, w_10000_1193, w_10000_1194, w_10000_1195, w_10000_1196, w_10000_1197, w_10000_1198, w_10000_1199, w_10000_1200, w_10000_1201, w_10000_1202, w_10000_1203, w_10000_1204, w_10000_1205, w_10000_1206, w_10000_1207, w_10000_1208, w_10000_1209, w_10000_1210, w_10000_1211, w_10000_1212, w_10000_1213, w_10000_1214, w_10000_1215, w_10000_1216, w_10000_1217, w_10000_1218, w_10000_1219, w_10000_1220, w_10000_1221, w_10000_1222, w_10000_1223, w_10000_1224, w_10000_1225, w_10000_1226, w_10000_1227, w_10000_1228, w_10000_1229, w_10000_1230, w_10000_1231, w_10000_1232, w_10000_1233, w_10000_1234, w_10000_1235, w_10000_1236, w_10000_1237, w_10000_1238, w_10000_1239, w_10000_1240, w_10000_1241, w_10000_1242, w_10000_1243, w_10000_1244, w_10000_1245, w_10000_1246, w_10000_1247, w_10000_1248, w_10000_1249, w_10000_1250, w_10000_1251, w_10000_1252, w_10000_1253, w_10000_1254, w_10000_1255, w_10000_1256, w_10000_1257, w_10000_1258, w_10000_1259, w_10000_1260, w_10000_1261, w_10000_1262, w_10000_1263, w_10000_1264, w_10000_1265, w_10000_1266, w_10000_1267, w_10000_1268, w_10000_1269, w_10000_1270, w_10000_1271, w_10000_1272, w_10000_1273, w_10000_1274, w_10000_1275, w_10000_1276, w_10000_1277, w_10000_1278, w_10000_1279, w_10000_1280, w_10000_1281, w_10000_1282, w_10000_1283, w_10000_1284, w_10000_1285, w_10000_1286, w_10000_1287, w_10000_1288, w_10000_1289, w_10000_1290, w_10000_1291, w_10000_1292, w_10000_1293, w_10000_1294, w_10000_1295, w_10000_1296, w_10000_1297, w_10000_1298, w_10000_1299, w_10000_1300, w_10000_1301, w_10000_1302, w_10000_1303, w_10000_1304, w_10000_1305, w_10000_1306, w_10000_1307, w_10000_1308, w_10000_1309, w_10000_1310, w_10000_1311, w_10000_1312, w_10000_1313, w_10000_1314, w_10000_1315, w_10000_1316, w_10000_1317, w_10000_1318, w_10000_1319, w_10000_1320, w_10000_1321, w_10000_1322, w_10000_1323, w_10000_1324, w_10000_1325, w_10000_1326, w_10000_1327, w_10000_1328, w_10000_1329, w_10000_1330, w_10000_1331, w_10000_1332, w_10000_1333, w_10000_1334, w_10000_1335, w_10000_1336, w_10000_1337, w_10000_1338, w_10000_1339, w_10000_1340, w_10000_1341, w_10000_1342, w_10000_1343, w_10000_1344, w_10000_1345, w_10000_1346, w_10000_1347, w_10000_1348, w_10000_1349, w_10000_1350, w_10000_1351, w_10000_1352, w_10000_1353, w_10000_1354, w_10000_1355, w_10000_1356, w_10000_1357, w_10000_1358, w_10000_1359, w_10000_1360, w_10000_1361, w_10000_1362, w_10000_1363, w_10000_1364, w_10000_1365, w_10000_1366, w_10000_1367, w_10000_1368, w_10000_1369, w_10000_1370, w_10000_1371, w_10000_1372, w_10000_1373, w_10000_1374, w_10000_1375, w_10000_1376, w_10000_1377, w_10000_1378, w_10000_1379, w_10000_1380, w_10000_1381, w_10000_1382, w_10000_1383, w_10000_1384, w_10000_1385, w_10000_1386, w_10000_1387, w_10000_1388, w_10000_1389, w_10000_1390, w_10000_1391, w_10000_1392, w_10000_1393, w_10000_1394, w_10000_1395, w_10000_1396, w_10000_1397, w_10000_1398, w_10000_1399, w_10000_1400, w_10000_1401, w_10000_1402, w_10000_1403, w_10000_1404, w_10000_1405, w_10000_1406, w_10000_1407, w_10000_1408, w_10000_1409, w_10000_1410, w_10000_1411, w_10000_1412, w_10000_1413, w_10000_1414, w_10000_1415, w_10000_1416, w_10000_1417, w_10000_1418, w_10000_1419, w_10000_1420, w_10000_1421, w_10000_1422, w_10000_1423, w_10000_1424, w_10000_1425, w_10000_1426, w_10000_1427, w_10000_1428, w_10000_1429, w_10000_1430, w_10000_1431, w_10000_1432, w_10000_1433, w_10000_1434, w_10000_1435, w_10000_1436, w_10000_1437, w_10000_1438, w_10000_1439, w_10000_1440, w_10000_1441, w_10000_1442, w_10000_1443, w_10000_1444, w_10000_1445, w_10000_1446, w_10000_1447, w_10000_1448, w_10000_1449, w_10000_1450, w_10000_1451, w_10000_1452, w_10000_1453, w_10000_1454, w_10000_1455, w_10000_1456, w_10000_1457, w_10000_1458, w_10000_1459, w_10000_1460, w_10000_1461, w_10000_1462, w_10000_1463, w_10000_1464, w_10000_1465, w_10000_1466, w_10000_1467, w_10000_1468, w_10000_1469, w_10000_1470, w_10000_1471, w_10000_1472, w_10000_1473, w_10000_1474, w_10000_1475, w_10000_1476, w_10000_1477, w_10000_1478, w_10000_1479, w_10000_1480, w_10000_1481, w_10000_1482, w_10000_1483, w_10000_1484, w_10000_1485, w_10000_1486, w_10000_1487, w_10000_1488, w_10000_1489, w_10000_1490, w_10000_1491, w_10000_1492, w_10000_1493, w_10000_1494, w_10000_1495, w_10000_1496, w_10000_1497, w_10000_1498, w_10000_1499, w_10000_1500, w_10000_1501, w_10000_1502, w_10000_1503, w_10000_1504, w_10000_1505, w_10000_1506, w_10000_1507, w_10000_1508, w_10000_1509, w_10000_1510, w_10000_1511, w_10000_1512, w_10000_1513, w_10000_1514, w_10000_1515, w_10000_1516, w_10000_1517, w_10000_1518, w_10000_1519, w_10000_1520, w_10000_1521, w_10000_1522, w_10000_1523, w_10000_1524, w_10000_1525, w_10000_1526, w_10000_1527, w_10000_1528, w_10000_1529, w_10000_1530, w_10000_1531, w_10000_1532, w_10000_1533, w_10000_1534, w_10000_1535, w_10000_1536, w_10000_1537, w_10000_1538, w_10000_1539, w_10000_1540, w_10000_1541, w_10000_1542, w_10000_1543, w_10000_1544, w_10000_1545, w_10000_1546, w_10000_1547, w_10000_1548, w_10000_1549, w_10000_1550, w_10000_1551, w_10000_1552, w_10000_1553, w_10000_1554, w_10000_1555, w_10000_1556, w_10000_1557, w_10000_1558, w_10000_1559, w_10000_1560, w_10000_1561, w_10000_1562, w_10000_1563, w_10000_1564, w_10000_1565, w_10000_1566, w_10000_1567, w_10000_1568, w_10000_1569, w_10000_1570, w_10000_1571, w_10000_1572, w_10000_1573, w_10000_1574, w_10000_1575, w_10000_1576, w_10000_1577, w_10000_1578, w_10000_1579, w_10000_1580, w_10000_1581, w_10000_1582, w_10000_1583, w_10000_1584, w_10000_1585, w_10000_1586, w_10000_1587, w_10000_1588, w_10000_1589, w_10000_1590, w_10000_1591, w_10000_1592, w_10000_1593, w_10000_1594, w_10000_1595, w_10000_1596, w_10000_1597, w_10000_1598, w_10000_1599, w_10000_1600, w_10000_1601, w_10000_1602, w_10000_1603, w_10000_1604, w_10000_1605, w_10000_1606, w_10000_1607, w_10000_1608, w_10000_1609, w_10000_1610, w_10000_1611, w_10000_1612, w_10000_1613, w_10000_1614, w_10000_1615, w_10000_1616, w_10000_1617, w_10000_1618, w_10000_1619, w_10000_1620, w_10000_1621, w_10000_1622, w_10000_1623, w_10000_1624, w_10000_1625, w_10000_1626, w_10000_1627, w_10000_1628, w_10000_1629, w_10000_1630, w_10000_1631, w_10000_1632, w_10000_1633, w_10000_1634, w_10000_1635, w_10000_1636, w_10000_1637, w_10000_1638, w_10000_1639, w_10000_1640, w_10000_1641, w_10000_1642, w_10000_1643, w_10000_1644, w_10000_1645, w_10000_1646, w_10000_1647, w_10000_1648, w_10000_1649, w_10000_1650, w_10000_1651, w_10000_1652, w_10000_1653, w_10000_1654, w_10000_1655, w_10000_1656, w_10000_1657, w_10000_1658, w_10000_1659, w_10000_1660, w_10000_1661, w_10000_1662, w_10000_1663, w_10000_1664, w_10000_1665, w_10000_1666, w_10000_1667, w_10000_1668, w_10000_1669, w_10000_1670, w_10000_1671, w_10000_1672, w_10000_1673, w_10000_1674, w_10000_1675, w_10000_1676, w_10000_1677, w_10000_1678, w_10000_1679, w_10000_1680, w_10000_1681, w_10000_1682, w_10000_1683, w_10000_1684, w_10000_1685, w_10000_1686, w_10000_1687, w_10000_1688, w_10000_1689, w_10000_1690, w_10000_1691, w_10000_1692, w_10000_1693, w_10000_1694, w_10000_1695, w_10000_1696, w_10000_1697, w_10000_1698, w_10000_1699, w_10000_1700, w_10000_1701, w_10000_1702, w_10000_1703, w_10000_1704, w_10000_1705, w_10000_1706, w_10000_1707, w_10000_1708, w_10000_1709, w_10000_1710, w_10000_1711, w_10000_1712, w_10000_1713, w_10000_1714, w_10000_1715, w_10000_1716, w_10000_1717, w_10000_1718, w_10000_1719, w_10000_1720, w_10000_1721, w_10000_1722, w_10000_1723, w_10000_1724, w_10000_1725, w_10000_1726, w_10000_1727, w_10000_1728, w_10000_1729, w_10000_1730, w_10000_1731, w_10000_1732, w_10000_1733, w_10000_1734, w_10000_1735, w_10000_1736, w_10000_1737, w_10000_1738, w_10000_1739, w_10000_1740, w_10000_1741, w_10000_1742, w_10000_1743, w_10000_1744, w_10000_1745, w_10000_1746, w_10000_1747, w_10000_1748, w_10000_1749, w_10000_1750, w_10000_1751, w_10000_1752, w_10000_1753, w_10000_1754, w_10000_1755, w_10000_1756, w_10000_1757, w_10000_1758, w_10000_1759, w_10000_1760, w_10000_1761, w_10000_1762, w_10000_1763, w_10000_1764, w_10000_1765, w_10000_1766, w_10000_1767, w_10000_1768, w_10000_1769, w_10000_1770, w_10000_1771, w_10000_1772, w_10000_1773, w_10000_1774, w_10000_1775, w_10000_1776, w_10000_1777, w_10000_1778, w_10000_1779, w_10000_1780, w_10000_1781, w_10000_1782, w_10000_1783, w_10000_1784, w_10000_1785, w_10000_1786, w_10000_1787, w_10000_1788, w_10000_1789, w_10000_1790, w_10000_1791, w_10000_1792, w_10000_1793, w_10000_1794, w_10000_1795, w_10000_1796, w_10000_1797, w_10000_1798, w_10000_1799, w_10000_1800, w_10000_1801, w_10000_1802, w_10000_1803, w_10000_1804, w_10000_1805, w_10000_1806, w_10000_1807, w_10000_1808, w_10000_1809, w_10000_1810, w_10000_1811, w_10000_1812, w_10000_1813, w_10000_1814, w_10000_1815, w_10000_1816, w_10000_1817, w_10000_1818, w_10000_1819, w_10000_1820, w_10000_1821, w_10000_1822, w_10000_1823, w_10000_1824, w_10000_1825, w_10000_1826, w_10000_1827, w_10000_1828, w_10000_1829, w_10000_1830, w_10000_1831, w_10000_1832, w_10000_1833, w_10000_1834, w_10000_1835, w_10000_1836, w_10000_1837, w_10000_1838, w_10000_1839, w_10000_1840, w_10000_1841, w_10000_1842, w_10000_1843, w_10000_1844, w_10000_1845, w_10000_1846, w_10000_1847, w_10000_1848, w_10000_1849, w_10000_1850, w_10000_1851, w_10000_1852, w_10000_1853, w_10000_1854, w_10000_1855, w_10000_1856, w_10000_1857, w_10000_1858, w_10000_1859, w_10000_1860, w_10000_1861, w_10000_1862, w_10000_1863, w_10000_1864, w_10000_1865, w_10000_1866, w_10000_1867, w_10000_1868, w_10000_1869, w_10000_1870, w_10000_1871, w_10000_1872, w_10000_1873, w_10000_1874, w_10000_1875, w_10000_1876, w_10000_1877, w_10000_1878, w_10000_1879, w_10000_1880, w_10000_1881, w_10000_1882, w_10000_1883, w_10000_1884, w_10000_1885, w_10000_1886, w_10000_1887, w_10000_1888, w_10000_1889, w_10000_1890, w_10000_1891, w_10000_1892, w_10000_1893, w_10000_1894, w_10000_1895, w_10000_1896, w_10000_1897, w_10000_1898, w_10000_1899, w_10000_1900, w_10000_1901, w_10000_1902, w_10000_1903, w_10000_1904, w_10000_1905, w_10000_1906, w_10000_1907, w_10000_1908, w_10000_1909, w_10000_1910, w_10000_1911, w_10000_1912, w_10000_1913, w_10000_1914, w_10000_1915, w_10000_1916, w_10000_1917, w_10000_1918, w_10000_1919, w_10000_1920, w_10000_1921, w_10000_1922, w_10000_1923, w_10000_1924, w_10000_1925, w_10000_1926, w_10000_1927, w_10000_1928, w_10000_1929, w_10000_1930, w_10000_1931, w_10000_1932, w_10000_1933, w_10000_1934, w_10000_1935, w_10000_1936, w_10000_1937, w_10000_1938, w_10000_1939, w_10000_1940, w_10000_1941, w_10000_1942, w_10000_1943, w_10000_1944, w_10000_1945, w_10000_1946, w_10000_1947, w_10000_1948, w_10000_1949, w_10000_1950, w_10000_1951, w_10000_1952, w_10000_1953, w_10000_1954, w_10000_1955, w_10000_1956, w_10000_1957, w_10000_1958, w_10000_1959, w_10000_1960, w_10000_1961, w_10000_1962, w_10000_1963, w_10000_1964, w_10000_1965, w_10000_1966, w_10000_1967, w_10000_1968, w_10000_1969, w_10000_1970, w_10000_1971, w_10000_1972, w_10000_1973, w_10000_1974, w_10000_1975, w_10000_1976, w_10000_1977, w_10000_1978, w_10000_1979, w_10000_1980, w_10000_1981, w_10000_1982, w_10000_1983, w_10000_1984, w_10000_1985, w_10000_1986, w_10000_1987, w_10000_1988, w_10000_1989, w_10000_1990, w_10000_1991, w_10000_1992, w_10000_1993, w_10000_1994, w_10000_1995, w_10000_1996, w_10000_1997, w_10000_1998, w_10000_1999, w_10000_2000, w_10000_2001, w_10000_2002, w_10000_2003, w_10000_2004, w_10000_2005, w_10000_2006, w_10000_2007, w_10000_2008, w_10000_2009, w_10000_2010, w_10000_2011, w_10000_2012, w_10000_2013, w_10000_2014, w_10000_2015, w_10000_2016, w_10000_2017, w_10000_2018, w_10000_2019, w_10000_2020, w_10000_2021, w_10000_2022, w_10000_2023, w_10000_2024, w_10000_2025, w_10000_2026, w_10000_2027, w_10000_2028, w_10000_2029, w_10000_2030, w_10000_2031, w_10000_2032, w_10000_2033, w_10000_2034, w_10000_2035, w_10000_2036, w_10000_2037, w_10000_2038, w_10000_2039, w_10000_2040, w_10000_2041, w_10000_2042, w_10000_2043, w_10000_2044, w_10000_2045, w_10000_2046, w_10000_2047, w_10000_2048, w_10000_2049, w_10000_2050, w_10000_2051, w_10000_2052, w_10000_2053, w_10000_2054, w_10000_2055, w_10000_2056, w_10000_2057, w_10000_2058, w_10000_2059, w_10000_2060, w_10000_2061, w_10000_2062, w_10000_2063, w_10000_2064, w_10000_2065, w_10000_2066, w_10000_2067, w_10000_2068, w_10000_2069, w_10000_2070, w_10000_2071, w_10000_2072, w_10000_2073, w_10000_2074, w_10000_2075, w_10000_2076, w_10000_2077, w_10000_2078, w_10000_2079, w_10000_2080, w_10000_2081, w_10000_2082, w_10000_2083, w_10000_2084, w_10000_2085, w_10000_2086, w_10000_2087, w_10000_2088, w_10000_2089, w_10000_2090, w_10000_2091, w_10000_2092, w_10000_2093, w_10000_2094, w_10000_2095, w_10000_2096, w_10000_2097, w_10000_2098, w_10000_2099, w_10000_2100, w_10000_2101, w_10000_2102, w_10000_2103, w_10000_2104, w_10000_2105, w_10000_2106, w_10000_2107, w_10000_2108, w_10000_2109, w_10000_2110, w_10000_2111, w_10000_2112, w_10000_2113, w_10000_2114, w_10000_2115, w_10000_2116, w_10000_2117, w_10000_2118, w_10000_2119, w_10000_2120, w_10000_2121, w_10000_2122, w_10000_2123, w_10000_2124, w_10000_2125, w_10000_2126, w_10000_2127, w_10000_2128, w_10000_2129, w_10000_2130, w_10000_2131, w_10000_2132, w_10000_2133, w_10000_2134, w_10000_2135, w_10000_2136, w_10000_2137, w_10000_2138, w_10000_2139, w_10000_2140, w_10000_2141, w_10000_2142, w_10000_2143, w_10000_2144, w_10000_2145, w_10000_2146, w_10000_2147, w_10000_2148, w_10000_2149, w_10000_2150, w_10000_2151, w_10000_2152, w_10000_2153, w_10000_2154, w_10000_2155, w_10000_2156, w_10000_2157, w_10000_2158, w_10000_2159, w_10000_2160, w_10000_2161, w_10000_2162, w_10000_2163, w_10000_2164, w_10000_2165, w_10000_2166, w_10000_2167, w_10000_2168, w_10000_2169, w_10000_2170, w_10000_2171, w_10000_2172, w_10000_2173, w_10000_2174, w_10000_2175, w_10000_2176, w_10000_2177, w_10000_2178, w_10000_2179, w_10000_2180, w_10000_2181, w_10000_2182, w_10000_2183, w_10000_2184, w_10000_2185, w_10000_2186, w_10000_2187, w_10000_2188, w_10000_2189, w_10000_2190, w_10000_2191, w_10000_2192, w_10000_2193, w_10000_2194, w_10000_2195, w_10000_2196, w_10000_2197, w_10000_2198, w_10000_2199, w_10000_2200, w_10000_2201, w_10000_2202, w_10000_2203, w_10000_2204, w_10000_2205, w_10000_2206, w_10000_2207, w_10000_2208, w_10000_2209, w_10000_2210, w_10000_2211, w_10000_2212, w_10000_2213, w_10000_2214, w_10000_2215, w_10000_2216, w_10000_2217, w_10000_2218, w_10000_2219, w_10000_2220, w_10000_2221, w_10000_2222, w_10000_2223, w_10000_2224, w_10000_2225, w_10000_2226, w_10000_2227, w_10000_2228, w_10000_2229, w_10000_2230, w_10000_2231, w_10000_2232, w_10000_2233, w_10000_2234, w_10000_2235, w_10000_2236, w_10000_2237, w_10000_2238, w_10000_2239, w_10000_2240, w_10000_2241, w_10000_2242, w_10000_2243, w_10000_2244, w_10000_2245, w_10000_2246, w_10000_2247, w_10000_2248, w_10000_2249, w_10000_2250, w_10000_2251, w_10000_2252, w_10000_2253, w_10000_2254, w_10000_2255, w_10000_2256, w_10000_2257, w_10000_2258, w_10000_2259, w_10000_2260, w_10000_2261, w_10000_2262, w_10000_2263, w_10000_2264, w_10000_2265, w_10000_2266, w_10000_2267, w_10000_2268, w_10000_2269, w_10000_2270, w_10000_2271, w_10000_2272, w_10000_2273, w_10000_2274, w_10000_2275, w_10000_2276, w_10000_2277, w_10000_2278, w_10000_2279, w_10000_2280, w_10000_2281, w_10000_2282, w_10000_2283, w_10000_2284, w_10000_2285, w_10000_2286, w_10000_2287, w_10000_2288, w_10000_2289, w_10000_2290, w_10000_2291, w_10000_2292, w_10000_2293, w_10000_2294, w_10000_2295, w_10000_2296, w_10000_2297, w_10000_2298, w_10000_2299, w_10000_2300, w_10000_2301, w_10000_2302, w_10000_2303, w_10000_2304, w_10000_2305, w_10000_2306, w_10000_2307, w_10000_2308, w_10000_2309, w_10000_2310, w_10000_2311, w_10000_2312, w_10000_2313, w_10000_2314, w_10000_2315, w_10000_2316, w_10000_2317, w_10000_2318, w_10000_2319, w_10000_2320, w_10000_2321, w_10000_2322, w_10000_2323, w_10000_2324, w_10000_2325, w_10000_2326, w_10000_2327, w_10000_2328, w_10000_2329, w_10000_2330, w_10000_2331, w_10000_2332, w_10000_2333, w_10000_2334, w_10000_2335, w_10000_2336, w_10000_2337, w_10000_2338, w_10000_2339, w_10000_2340, w_10000_2341, w_10000_2342, w_10000_2343, w_10000_2344, w_10000_2345, w_10000_2346, w_10000_2347, w_10000_2348, w_10000_2349, w_10000_2350, w_10000_2351, w_10000_2352, w_10000_2353, w_10000_2354, w_10000_2355, w_10000_2356, w_10000_2357, w_10000_2358, w_10000_2359, w_10000_2360, w_10000_2361, w_10000_2362, w_10000_2363, w_10000_2364, w_10000_2365, w_10000_2366, w_10000_2367, w_10000_2368, w_10000_2369, w_10000_2370, w_10000_2371, w_10000_2372, w_10000_2373, w_10000_2374, w_10000_2375, w_10000_2376, w_10000_2377, w_10000_2378, w_10000_2379, w_10000_2380, w_10000_2381, w_10000_2382, w_10000_2383, w_10000_2384, w_10000_2385, w_10000_2386, w_10000_2387, w_10000_2388, w_10000_2389, w_10000_2390, w_10000_2391, w_10000_2392, w_10000_2393, w_10000_2394, w_10000_2395, w_10000_2396, w_10000_2397, w_10000_2398, w_10000_2399, w_10000_2400, w_10000_2401, w_10000_2402, w_10000_2403, w_10000_2404, w_10000_2405, w_10000_2406, w_10000_2407, w_10000_2408, w_10000_2409, w_10000_2410, w_10000_2411, w_10000_2412, w_10000_2413, w_10000_2414, w_10000_2415, w_10000_2416, w_10000_2417, w_10000_2418, w_10000_2419, w_10000_2420, w_10000_2421, w_10000_2422, w_10000_2423, w_10000_2424, w_10000_2425, w_10000_2426, w_10000_2427, w_10000_2428, w_10000_2429, w_10000_2430, w_10000_2431, w_10000_2432, w_10000_2433, w_10000_2434, w_10000_2435, w_10000_2436, w_10000_2437, w_10000_2438, w_10000_2439, w_10000_2440, w_10000_2441, w_10000_2442, w_10000_2443, w_10000_2444, w_10000_2445, w_10000_2446, w_10000_2447, w_10000_2448, w_10000_2449, w_10000_2450, w_10000_2451, w_10000_2452, w_10000_2453, w_10000_2454, w_10000_2455, w_10000_2456, w_10000_2457, w_10000_2458, w_10000_2459, w_10000_2460, w_10000_2461, w_10000_2462, w_10000_2463, w_10000_2464, w_10000_2465, w_10000_2466, w_10000_2467, w_10000_2468, w_10000_2469, w_10000_2470, w_10000_2471, w_10000_2472, w_10000_2473, w_10000_2474, w_10000_2475, w_10000_2476, w_10000_2477, w_10000_2478, w_10000_2479, w_10000_2480, w_10000_2481, w_10000_2482, w_10000_2483, w_10000_2484, w_10000_2485, w_10000_2486, w_10000_2487, w_10000_2488, w_10000_2489, w_10000_2490, w_10000_2491, w_10000_2492, w_10000_2493, w_10000_2494, w_10000_2495, w_10000_2496, w_10000_2497, w_10000_2498, w_10000_2499, w_10000_2500, w_10000_2501, w_10000_2502, w_10000_2503, w_10000_2504, w_10000_2505, w_10000_2506, w_10000_2507, w_10000_2508, w_10000_2509, w_10000_2510, w_10000_2511, w_10000_2512, w_10000_2513, w_10000_2514, w_10000_2515, w_10000_2516, w_10000_2517, w_10000_2518, w_10000_2519, w_10000_2520, w_10000_2521, w_10000_2522, w_10000_2523, w_10000_2524, w_10000_2525, w_10000_2526, w_10000_2527, w_10000_2528, w_10000_2529, w_10000_2530, w_10000_2531, w_10000_2532, w_10000_2533, w_10000_2534, w_10000_2535, w_10000_2536, w_10000_2537, w_10000_2538, w_10000_2539, w_10000_2540, w_10000_2541, w_10000_2542, w_10000_2543, w_10000_2544, w_10000_2545, w_10000_2546, w_10000_2547, w_10000_2548, w_10000_2549, w_10000_2550, w_10000_2551, w_10000_2552, w_10000_2553, w_10000_2554, w_10000_2555, w_10000_2556, w_10000_2557, w_10000_2558, w_10000_2559, w_10000_2560, w_10000_2561, w_10000_2562, w_10000_2563, w_10000_2564, w_10000_2565, w_10000_2566, w_10000_2567, w_10000_2568, w_10000_2569, w_10000_2570, w_10000_2571, w_10000_2572, w_10000_2573, w_10000_2574, w_10000_2575, w_10000_2576, w_10000_2577, w_10000_2578, w_10000_2579, w_10000_2580, w_10000_2581, w_10000_2582, w_10000_2583, w_10000_2584, w_10000_2585, w_10000_2586, w_10000_2587, w_10000_2588, w_10000_2589, w_10000_2590, w_10000_2591, w_10000_2592, w_10000_2593, w_10000_2594, w_10000_2595, w_10000_2596, w_10000_2597, w_10000_2598, w_10000_2599, w_10000_2600, w_10000_2601, w_10000_2602, w_10000_2603, w_10000_2604, w_10000_2605, w_10000_2606, w_10000_2607, w_10000_2608, w_10000_2609, w_10000_2610, w_10000_2611, w_10000_2612, w_10000_2613, w_10000_2614, w_10000_2615, w_10000_2616, w_10000_2617, w_10000_2618, w_10000_2619, w_10000_2620, w_10000_2621, w_10000_2622, w_10000_2623, w_10000_2624, w_10000_2625, w_10000_2626, w_10000_2627, w_10000_2628, w_10000_2629, w_10000_2630, w_10000_2631, w_10000_2632, w_10000_2633, w_10000_2634, w_10000_2635, w_10000_2636, w_10000_2637, w_10000_2638, w_10000_2639, w_10000_2640, w_10000_2641, w_10000_2642, w_10000_2643, w_10000_2644, w_10000_2645, w_10000_2646, w_10000_2647, w_10000_2648, w_10000_2649, w_10000_2650, w_10000_2651, w_10000_2652, w_10000_2653, w_10000_2654, w_10000_2655, w_10000_2656, w_10000_2657, w_10000_2658, w_10000_2659, w_10000_2660, w_10000_2661, w_10000_2662, w_10000_2663, w_10000_2664, w_10000_2665, w_10000_2666, w_10000_2667, w_10000_2668, w_10000_2669, w_10000_2670, w_10000_2671, w_10000_2672, w_10000_2673, w_10000_2674, w_10000_2675, w_10000_2676, w_10000_2677, w_10000_2678, w_10000_2679, w_10000_2680, w_10000_2681, w_10000_2682, w_10000_2683, w_10000_2684, w_10000_2685, w_10000_2686, w_10000_2687, w_10000_2688, w_10000_2689, w_10000_2690, w_10000_2691, w_10000_2692, w_10000_2693, w_10000_2694, w_10000_2695, w_10000_2696, w_10000_2697, w_10000_2698, w_10000_2699, w_10000_2700, w_10000_2701, w_10000_2702, w_10000_2703, w_10000_2704, w_10000_2705, w_10000_2706, w_10000_2707, w_10000_2708, w_10000_2709, w_10000_2710, w_10000_2711, w_10000_2712, w_10000_2713, w_10000_2714, w_10000_2715, w_10000_2716, w_10000_2717, w_10000_2718, w_10000_2719, w_10000_2720, w_10000_2721, w_10000_2722, w_10000_2723, w_10000_2724, w_10000_2725, w_10000_2726, w_10000_2727, w_10000_2728, w_10000_2729, w_10000_2730, w_10000_2731, w_10000_2732, w_10000_2733, w_10000_2734, w_10000_2735, w_10000_2736, w_10000_2737, w_10000_2738, w_10000_2739, w_10000_2740, w_10000_2741, w_10000_2742, w_10000_2743, w_10000_2744, w_10000_2745, w_10000_2746, w_10000_2747, w_10000_2748, w_10000_2749, w_10000_2750, w_10000_2751, w_10000_2752, w_10000_2753, w_10000_2754, w_10000_2755, w_10000_2756, w_10000_2757, w_10000_2758, w_10000_2759, w_10000_2760, w_10000_2761, w_10000_2762, w_10000_2763, w_10000_2764, w_10000_2765, w_10000_2766, w_10000_2767, w_10000_2768, w_10000_2769, w_10000_2770, w_10000_2771, w_10000_2772, w_10000_2773, w_10000_2774, w_10000_2775, w_10000_2776, w_10000_2777, w_10000_2778, w_10000_2779, w_10000_2780, w_10000_2781, w_10000_2782, w_10000_2783, w_10000_2784, w_10000_2785, w_10000_2786, w_10000_2787, w_10000_2788, w_10000_2789, w_10000_2790, w_10000_2791, w_10000_2792, w_10000_2793, w_10000_2794, w_10000_2795, w_10000_2796, w_10000_2797, w_10000_2798, w_10000_2799, w_10000_2800, w_10000_2801, w_10000_2802, w_10000_2803, w_10000_2804, w_10000_2805, w_10000_2806, w_10000_2807, w_10000_2808, w_10000_2809, w_10000_2810, w_10000_2811, w_10000_2812, w_10000_2813, w_10000_2814, w_10000_2815, w_10000_2816, w_10000_2817, w_10000_2818, w_10000_2819, w_10000_2820, w_10000_2821, w_10000_2822, w_10000_2823, w_10000_2824, w_10000_2825, w_10000_2826, w_10000_2827, w_10000_2828, w_10000_2829, w_10000_2830, w_10000_2831, w_10000_2832, w_10000_2833, w_10000_2834, w_10000_2835, w_10000_2836, w_10000_2837, w_10000_2838, w_10000_2839, w_10000_2840, w_10000_2841, w_10000_2842, w_10000_2843, w_10000_2844, w_10000_2845, w_10000_2846, w_10000_2847, w_10000_2848, w_10000_2849, w_10000_2850, w_10000_2851, w_10000_2852, w_10000_2853, w_10000_2854, w_10000_2855, w_10000_2856, w_10000_2857, w_10000_2858, w_10000_2859, w_10000_2860, w_10000_2861, w_10000_2862, w_10000_2863, w_10000_2864, w_10000_2865, w_10000_2866, w_10000_2867, w_10000_2868, w_10000_2869, w_10000_2870, w_10000_2871, w_10000_2872, w_10000_2873, w_10000_2874, w_10000_2875, w_10000_2876, w_10000_2877, w_10000_2878, w_10000_2879, w_10000_2880, w_10000_2881, w_10000_2882, w_10000_2883, w_10000_2884, w_10000_2885, w_10000_2886, w_10000_2887, w_10000_2888, w_10000_2889, w_10000_2890, w_10000_2891, w_10000_2892, w_10000_2893, w_10000_2894, w_10000_2895, w_10000_2896, w_10000_2897, w_10000_2898, w_10000_2899, w_10000_2900, w_10000_2901, w_10000_2902, w_10000_2903, w_10000_2904, w_10000_2905, w_10000_2906, w_10000_2907, w_10000_2908, w_10000_2909, w_10000_2910, w_10000_2911, w_10000_2912, w_10000_2913, w_10000_2914, w_10000_2915, w_10000_2916, w_10000_2917, w_10000_2918, w_10000_2919, w_10000_2920, w_10000_2921, w_10000_2922, w_10000_2923, w_10000_2924, w_10000_2925, w_10000_2926, w_10000_2927, w_10000_2928, w_10000_2929, w_10000_2930, w_10000_2931, w_10000_2932, w_10000_2933, w_10000_2934, w_10000_2935, w_10000_2936, w_10000_2937, w_10000_2938, w_10000_2939, w_10000_2940, w_10000_2941, w_10000_2942, w_10000_2943, w_10000_2944, w_10000_2945, w_10000_2946, w_10000_2947, w_10000_2948, w_10000_2949, w_10000_2950, w_10000_2951, w_10000_2952, w_10000_2953, w_10000_2954, w_10000_2955, w_10000_2956, w_10000_2957, w_10000_2958, w_10000_2959, w_10000_2960, w_10000_2961, w_10000_2962, w_10000_2963, w_10000_2964, w_10000_2965, w_10000_2966, w_10000_2967, w_10000_2968, w_10000_2969, w_10000_2970, w_10000_2971, w_10000_2972, w_10000_2973, w_10000_2974, w_10000_2975, w_10000_2976, w_10000_2977, w_10000_2978, w_10000_2979, w_10000_2980, w_10000_2981, w_10000_2982, w_10000_2983, w_10000_2984, w_10000_2985, w_10000_2986, w_10000_2987, w_10000_2988, w_10000_2989, w_10000_2990, w_10000_2991, w_10000_2992, w_10000_2993, w_10000_2994, w_10000_2995, w_10000_2996, w_10000_2997, w_10000_2998, w_10000_2999, w_10000_3000, w_10000_3001, w_10000_3002, w_10000_3003, w_10000_3004, w_10000_3005, w_10000_3006, w_10000_3007, w_10000_3008, w_10000_3009, w_10000_3010, w_10000_3011, w_10000_3012, w_10000_3013, w_10000_3014, w_10000_3015, w_10000_3016, w_10000_3017, w_10000_3018, w_10000_3019, w_10000_3020, w_10000_3021, w_10000_3022, w_10000_3023, w_10000_3024, w_10000_3025, w_10000_3026, w_10000_3027, w_10000_3028, w_10000_3029, w_10000_3030, w_10000_3031, w_10000_3032, w_10000_3033, w_10000_3034, w_10000_3035, w_10000_3036, w_10000_3037, w_10000_3038, w_10000_3039, w_10000_3040, w_10000_3041, w_10000_3042, w_10000_3043, w_10000_3044, w_10000_3045, w_10000_3046, w_10000_3047, w_10000_3048, w_10000_3049, w_10000_3050, w_10000_3051, w_10000_3052, w_10000_3053, w_10000_3054, w_10000_3055, w_10000_3056, w_10000_3057, w_10000_3058, w_10000_3059, w_10000_3060, w_10000_3061, w_10000_3062, w_10000_3063, w_10000_3064, w_10000_3065, w_10000_3066, w_10000_3067, w_10000_3068, w_10000_3069, w_10000_3070, w_10000_3071, w_10000_3072, w_10000_3073, w_10000_3074, w_10000_3075, w_10000_3076, w_10000_3077, w_10000_3078, w_10000_3079, w_10000_3080, w_10000_3081, w_10000_3082, w_10000_3083, w_10000_3084, w_10000_3085, w_10000_3086, w_10000_3087, w_10000_3088, w_10000_3089, w_10000_3090, w_10000_3091, w_10000_3092, w_10000_3093, w_10000_3094, w_10000_3095, w_10000_3096, w_10000_3097, w_10000_3098, w_10000_3099, w_10000_3100, w_10000_3101, w_10000_3102, w_10000_3103, w_10000_3104, w_10000_3105, w_10000_3106, w_10000_3107, w_10000_3108, w_10000_3109, w_10000_3110, w_10000_3111, w_10000_3112, w_10000_3113, w_10000_3114, w_10000_3115, w_10000_3116, w_10000_3117, w_10000_3118, w_10000_3119, w_10000_3120, w_10000_3121, w_10000_3122, w_10000_3123, w_10000_3124, w_10000_3125, w_10000_3126, w_10000_3127, w_10000_3128, w_10000_3129, w_10000_3130, w_10000_3131, w_10000_3132, w_10000_3133, w_10000_3134, w_10000_3135, w_10000_3136, w_10000_3137, w_10000_3138, w_10000_3139, w_10000_3140, w_10000_3141, w_10000_3142, w_10000_3143, w_10000_3144, w_10000_3145, w_10000_3146, w_10000_3147, w_10000_3148, w_10000_3149, w_10000_3150, w_10000_3151, w_10000_3152, w_10000_3153, w_10000_3154, w_10000_3155, w_10000_3156, w_10000_3157, w_10000_3158, w_10000_3159, w_10000_3160, w_10000_3161, w_10000_3162, w_10000_3163, w_10000_3164, w_10000_3165, w_10000_3166, w_10000_3167, w_10000_3168, w_10000_3169, w_10000_3170, w_10000_3171, w_10000_3172, w_10000_3173, w_10000_3174, w_10000_3175, w_10000_3176, w_10000_3177, w_10000_3178, w_10000_3179, w_10000_3180, w_10000_3181, w_10000_3182, w_10000_3183, w_10000_3184, w_10000_3185, w_10000_3186, w_10000_3187, w_10000_3188, w_10000_3189, w_10000_3190, w_10000_3191, w_10000_3192, w_10000_3193, w_10000_3194, w_10000_3195, w_10000_3196, w_10000_3197, w_10000_3198, w_10000_3199, w_10000_3200, w_10000_3201, w_10000_3202, w_10000_3203, w_10000_3204, w_10000_3205, w_10000_3206, w_10000_3207, w_10000_3208, w_10000_3209, w_10000_3210, w_10000_3211, w_10000_3212, w_10000_3213, w_10000_3214, w_10000_3215, w_10000_3216, w_10000_3217, w_10000_3218, w_10000_3219, w_10000_3220, w_10000_3221, w_10000_3222, w_10000_3223, w_10000_3224, w_10000_3225, w_10000_3226, w_10000_3227, w_10000_3228, w_10000_3229, w_10000_3230, w_10000_3231, w_10000_3232, w_10000_3233, w_10000_3234, w_10000_3235, w_10000_3236, w_10000_3237, w_10000_3238, w_10000_3239, w_10000_3240, w_10000_3241, w_10000_3242, w_10000_3243, w_10000_3244, w_10000_3245, w_10000_3246, w_10000_3247, w_10000_3248, w_10000_3249, w_10000_3250, w_10000_3251, w_10000_3252, w_10000_3253, w_10000_3254, w_10000_3255, w_10000_3256, w_10000_3257, w_10000_3258, w_10000_3259, w_10000_3260, w_10000_3261, w_10000_3262, w_10000_3263, w_10000_3264, w_10000_3265, w_10000_3266, w_10000_3267, w_10000_3268, w_10000_3269, w_10000_3270, w_10000_3271, w_10000_3272, w_10000_3273, w_10000_3274, w_10000_3275, w_10000_3276, w_10000_3277, w_10000_3278, w_10000_3279, w_10000_3280, w_10000_3281, w_10000_3282, w_10000_3283, w_10000_3284, w_10000_3285, w_10000_3286, w_10000_3287, w_10000_3288, w_10000_3289, w_10000_3290, w_10000_3291, w_10000_3292, w_10000_3293, w_10000_3294, w_10000_3295, w_10000_3296, w_10000_3297, w_10000_3298, w_10000_3299, w_10000_3300, w_10000_3301, w_10000_3302, w_10000_3303, w_10000_3304, w_10000_3305, w_10000_3306, w_10000_3307, w_10000_3308, w_10000_3309, w_10000_3310, w_10000_3311, w_10000_3312, w_10000_3313, w_10000_3314, w_10000_3315, w_10000_3316, w_10000_3317, w_10000_3318, w_10000_3319, w_10000_3320, w_10000_3321, w_10000_3322, w_10000_3323, w_10000_3324, w_10000_3325, w_10000_3326, w_10000_3327, w_10000_3328, w_10000_3329, w_10000_3330, w_10000_3331, w_10000_3332, w_10000_3333, w_10000_3334, w_10000_3335, w_10000_3336, w_10000_3337, w_10000_3338, w_10000_3339, w_10000_3340, w_10000_3341, w_10000_3342, w_10000_3343, w_10000_3344, w_10000_3345, w_10000_3346, w_10000_3347, w_10000_3348, w_10000_3349, w_10000_3350, w_10000_3351, w_10000_3352, w_10000_3353, w_10000_3354, w_10000_3355, w_10000_3356, w_10000_3357, w_10000_3358, w_10000_3359, w_10000_3360, w_10000_3361, w_10000_3362, w_10000_3363, w_10000_3364, w_10000_3365, w_10000_3366, w_10000_3367, w_10000_3368, w_10000_3369, w_10000_3370, w_10000_3371, w_10000_3372, w_10000_3373, w_10000_3374, w_10000_3375, w_10000_3376, w_10000_3377, w_10000_3378, w_10000_3379, w_10000_3380, w_10000_3381, w_10000_3382, w_10000_3383, w_10000_3384, w_10000_3385, w_10000_3386, w_10000_3387, w_10000_3388, w_10000_3389, w_10000_3390, w_10000_3391, w_10000_3392, w_10000_3393, w_10000_3394, w_10000_3395, w_10000_3396, w_10000_3397, w_10000_3398, w_10000_3399, w_10000_3400, w_10000_3401, w_10000_3402, w_10000_3403, w_10000_3404, w_10000_3405, w_10000_3406, w_10000_3407, w_10000_3408, w_10000_3409, w_10000_3410, w_10000_3411, w_10000_3412, w_10000_3413, w_10000_3414, w_10000_3415, w_10000_3416, w_10000_3417, w_10000_3418, w_10000_3419, w_10000_3420, w_10000_3421, w_10000_3422, w_10000_3423, w_10000_3424, w_10000_3425, w_10000_3426, w_10000_3427, w_10000_3428, w_10000_3429, w_10000_3430, w_10000_3431, w_10000_3432, w_10000_3433, w_10000_3434, w_10000_3435, w_10000_3436, w_10000_3437, w_10000_3438, w_10000_3439, w_10000_3440, w_10000_3441, w_10000_3442, w_10000_3443, w_10000_3444, w_10000_3445, w_10000_3446, w_10000_3447, w_10000_3448, w_10000_3449, w_10000_3450, w_10000_3451, w_10000_3452, w_10000_3453, w_10000_3454, w_10000_3455, w_10000_3456, w_10000_3457, w_10000_3458, w_10000_3459, w_10000_3460, w_10000_3461, w_10000_3462, w_10000_3463, w_10000_3464, w_10000_3465, w_10000_3466, w_10000_3467, w_10000_3468, w_10000_3469, w_10000_3470, w_10000_3471, w_10000_3472, w_10000_3473, w_10000_3474, w_10000_3475, w_10000_3476, w_10000_3477, w_10000_3478, w_10000_3479, w_10000_3480, w_10000_3481, w_10000_3482, w_10000_3483, w_10000_3484, w_10000_3485, w_10000_3486, w_10000_3487, w_10000_3488, w_10000_3489, w_10000_3490, w_10000_3491, w_10000_3492, w_10000_3493, w_10000_3494, w_10000_3495, w_10000_3496, w_10000_3497, w_10000_3498, w_10000_3499, w_10000_3500, w_10000_3501, w_10000_3502, w_10000_3503, w_10000_3504, w_10000_3505, w_10000_3506, w_10000_3507, w_10000_3508, w_10000_3509, w_10000_3510, w_10000_3511, w_10000_3512, w_10000_3513, w_10000_3514, w_10000_3515, w_10000_3516, w_10000_3517, w_10000_3518, w_10000_3519, w_10000_3520, w_10000_3521, w_10000_3522, w_10000_3523, w_10000_3524, w_10000_3525, w_10000_3526, w_10000_3527, w_10000_3528, w_10000_3529, w_10000_3530, w_10000_3531, w_10000_3532, w_10000_3533, w_10000_3534, w_10000_3535, w_10000_3536, w_10000_3537, w_10000_3538, w_10000_3539, w_10000_3540, w_10000_3541, w_10000_3542, w_10000_3543, w_10000_3544, w_10000_3545, w_10000_3546, w_10000_3547, w_10000_3548, w_10000_3549, w_10000_3550, w_10000_3551, w_10000_3552, w_10000_3553, w_10000_3554, w_10000_3555, w_10000_3556, w_10000_3557, w_10000_3558, w_10000_3559, w_10000_3560, w_10000_3561, w_10000_3562, w_10000_3563, w_10000_3564, w_10000_3565, w_10000_3566, w_10000_3567, w_10000_3568, w_10000_3569, w_10000_3570, w_10000_3571, w_10000_3572, w_10000_3573, w_10000_3574, w_10000_3575, w_10000_3576, w_10000_3577, w_10000_3578, w_10000_3579, w_10000_3580, w_10000_3581, w_10000_3582, w_10000_3583, w_10000_3584, w_10000_3585, w_10000_3586, w_10000_3587, w_10000_3588, w_10000_3589, w_10000_3590, w_10000_3591, w_10000_3592, w_10000_3593, w_10000_3594, w_10000_3595, w_10000_3596, w_10000_3597, w_10000_3598, w_10000_3599, w_10000_3600, w_10000_3601, w_10000_3602, w_10000_3603, w_10000_3604, w_10000_3605, w_10000_3606, w_10000_3607, w_10000_3608, w_10000_3609, w_10000_3610, w_10000_3611, w_10000_3612, w_10000_3613, w_10000_3614, w_10000_3615, w_10000_3616, w_10000_3617, w_10000_3618, w_10000_3619, w_10000_3620, w_10000_3621, w_10000_3622, w_10000_3623, w_10000_3624, w_10000_3625, w_10000_3626, w_10000_3627, w_10000_3628, w_10000_3629, w_10000_3630, w_10000_3631, w_10000_3632, w_10000_3633, w_10000_3634, w_10000_3635, w_10000_3636, w_10000_3637, w_10000_3638, w_10000_3639, w_10000_3640, w_10000_3641, w_10000_3642, w_10000_3643, w_10000_3644, w_10000_3645, w_10000_3646, w_10000_3647, w_10000_3648, w_10000_3649, w_10000_3650, w_10000_3651, w_10000_3652, w_10000_3653, w_10000_3654, w_10000_3655, w_10000_3656, w_10000_3657, w_10000_3658, w_10000_3659, w_10000_3660, w_10000_3661, w_10000_3662, w_10000_3663, w_10000_3664, w_10000_3665, w_10000_3666, w_10000_3667, w_10000_3668, w_10000_3669, w_10000_3670, w_10000_3671, w_10000_3672, w_10000_3673, w_10000_3674, w_10000_3675, w_10000_3676, w_10000_3677, w_10000_3678, w_10000_3679, w_10000_3680, w_10000_3681, w_10000_3682, w_10000_3683, w_10000_3684, w_10000_3685, w_10000_3686, w_10000_3687, w_10000_3688, w_10000_3689, w_10000_3690, w_10000_3691, w_10000_3692, w_10000_3693, w_10000_3694, w_10000_3695, w_10000_3696, w_10000_3697, w_10000_3698, w_10000_3699, w_10000_3700, w_10000_3701, w_10000_3702, w_10000_3703, w_10000_3704, w_10000_3705, w_10000_3706, w_10000_3707, w_10000_3708, w_10000_3709, w_10000_3710, w_10000_3711, w_10000_3712, w_10000_3713, w_10000_3714, w_10000_3715, w_10000_3716, w_10000_3717, w_10000_3718, w_10000_3719, w_10000_3720, w_10000_3721, w_10000_3722, w_10000_3723, w_10000_3724, w_10000_3725, w_10000_3726, w_10000_3727, w_10000_3728, w_10000_3729, w_10000_3730, w_10000_3731, w_10000_3732, w_10000_3733, w_10000_3734, w_10000_3735, w_10000_3736, w_10000_3737, w_10000_3738, w_10000_3739, w_10000_3740, w_10000_3741, w_10000_3742, w_10000_3743, w_10000_3744, w_10000_3745, w_10000_3746, w_10000_3747, w_10000_3748, w_10000_3749, w_10000_3750, w_10000_3751, w_10000_3752, w_10000_3753, w_10000_3754, w_10000_3755, w_10000_3756, w_10000_3757, w_10000_3758, w_10000_3759, w_10000_3760, w_10000_3761, w_10000_3762, w_10000_3763, w_10000_3764, w_10000_3765, w_10000_3766, w_10000_3767, w_10000_3768, w_10000_3769, w_10000_3770, w_10000_3771, w_10000_3772, w_10000_3773, w_10000_3774, w_10000_3775, w_10000_3776, w_10000_3777, w_10000_3778, w_10000_3779, w_10000_3780, w_10000_3781, w_10000_3782, w_10000_3783, w_10000_3784, w_10000_3785, w_10000_3786, w_10000_3787, w_10000_3788, w_10000_3789, w_10000_3790, w_10000_3791, w_10000_3792, w_10000_3793, w_10000_3794, w_10000_3795, w_10000_3796, w_10000_3797, w_10000_3798, w_10000_3799, w_10000_3800, w_10000_3801, w_10000_3802, w_10000_3803, w_10000_3804, w_10000_3805, w_10000_3806, w_10000_3807, w_10000_3808, w_10000_3809, w_10000_3810, w_10000_3811, w_10000_3812, w_10000_3813, w_10000_3814, w_10000_3815, w_10000_3816, w_10000_3817, w_10000_3818, w_10000_3819, w_10000_3820, w_10000_3821, w_10000_3822, w_10000_3823, w_10000_3824, w_10000_3825, w_10000_3826, w_10000_3827, w_10000_3828, w_10000_3829, w_10000_3830, w_10000_3831, w_10000_3832, w_10000_3833, w_10000_3834, w_10000_3835, w_10000_3836, w_10000_3837, w_10000_3838, w_10000_3839, w_10000_3840, w_10000_3841, w_10000_3842, w_10000_3843, w_10000_3844, w_10000_3845, w_10000_3846, w_10000_3847, w_10000_3848, w_10000_3849, w_10000_3850, w_10000_3851, w_10000_3852, w_10000_3853, w_10000_3854, w_10000_3855, w_10000_3856, w_10000_3857, w_10000_3858, w_10000_3859, w_10000_3860, w_10000_3861, w_10000_3862, w_10000_3863, w_10000_3864, w_10000_3865, w_10000_3866, w_10000_3867, w_10000_3868, w_10000_3869, w_10000_3870, w_10000_3871, w_10000_3872, w_10000_3873, w_10000_3874, w_10000_3875, w_10000_3876, w_10000_3877, w_10000_3878, w_10000_3879, w_10000_3880, w_10000_3881, w_10000_3882, w_10000_3883, w_10000_3884, w_10000_3885, w_10000_3886, w_10000_3887, w_10000_3888, w_10000_3889, w_10000_3890, w_10000_3891, w_10000_3892, w_10000_3893, w_10000_3894, w_10000_3895, w_10000_3896, w_10000_3897, w_10000_3898, w_10000_3899, w_10000_3900, w_10000_3901, w_10000_3902, w_10000_3903, w_10000_3904, w_10000_3905, w_10000_3906, w_10000_3907, w_10000_3908, w_10000_3909, w_10000_3910, w_10000_3911, w_10000_3912, w_10000_3913, w_10000_3914, w_10000_3915, w_10000_3916, w_10000_3917, w_10000_3918, w_10000_3919, w_10000_3920, w_10000_3921, w_10000_3922, w_10000_3923, w_10000_3924, w_10000_3925, w_10000_3926, w_10000_3927, w_10000_3928, w_10000_3929, w_10000_3930, w_10000_3931, w_10000_3932, w_10000_3933, w_10000_3934, w_10000_3935, w_10000_3936, w_10000_3937, w_10000_3938, w_10000_3939, w_10000_3940, w_10000_3941, w_10000_3942, w_10000_3943, w_10000_3944, w_10000_3945, w_10000_3946, w_10000_3947, w_10000_3948, w_10000_3949, w_10000_3950, w_10000_3951, w_10000_3952, w_10000_3953, w_10000_3954, w_10000_3955, w_10000_3956, w_10000_3957, w_10000_3958, w_10000_3959, w_10000_3960, w_10000_3961, w_10000_3962, w_10000_3963, w_10000_3964, w_10000_3965, w_10000_3966, w_10000_3967, w_10000_3968, w_10000_3969, w_10000_3970, w_10000_3971, w_10000_3972, w_10000_3973, w_10000_3974, w_10000_3975, w_10000_3976, w_10000_3977, w_10000_3978, w_10000_3979, w_10000_3980, w_10000_3981, w_10000_3982, w_10000_3983, w_10000_3984, w_10000_3985, w_10000_3986, w_10000_3987, w_10000_3988, w_10000_3989, w_10000_3990, w_10000_3991, w_10000_3992, w_10000_3993, w_10000_3994, w_10000_3995, w_10000_3996, w_10000_3997, w_10000_3998, w_10000_3999, w_10000_4000, w_10000_4001, w_10000_4002, w_10000_4003, w_10000_4004, w_10000_4005, w_10000_4006, w_10000_4007, w_10000_4008, w_10000_4009, w_10000_4010, w_10000_4011, w_10000_4012, w_10000_4013, w_10000_4014, w_10000_4015, w_10000_4016, w_10000_4017, w_10000_4018, w_10000_4019, w_10000_4020, w_10000_4021, w_10000_4022, w_10000_4023, w_10000_4024, w_10000_4025, w_10000_4026, w_10000_4027, w_10000_4028, w_10000_4029, w_10000_4030, w_10000_4031, w_10000_4032, w_10000_4033, w_10000_4034, w_10000_4035, w_10000_4036, w_10000_4037, w_10000_4038, w_10000_4039, w_10000_4040, w_10000_4041, w_10000_4042, w_10000_4043, w_10000_4044, w_10000_4045, w_10000_4046, w_10000_4047, w_10000_4048, w_10000_4049, w_10000_4050, w_10000_4051, w_10000_4052, w_10000_4053, w_10000_4054, w_10000_4055, w_10000_4056, w_10000_4057, w_10000_4058, w_10000_4059, w_10000_4060, w_10000_4061, w_10000_4062, w_10000_4063, w_10000_4064, w_10000_4065, w_10000_4066, w_10000_4067, w_10000_4068, w_10000_4069, w_10000_4070, w_10000_4071, w_10000_4072, w_10000_4073, w_10000_4074, w_10000_4075, w_10000_4076, w_10000_4077, w_10000_4078, w_10000_4079, w_10000_4080, w_10000_4081, w_10000_4082, w_10000_4083, w_10000_4084, w_10000_4085, w_10000_4086, w_10000_4087, w_10000_4088, w_10000_4089, w_10000_4090, w_10000_4091, w_10000_4092, w_10000_4093, w_10000_4094, w_10000_4095, w_10000_4096, w_10000_4097, w_10000_4098, w_10000_4099, w_10000_4100, w_10000_4101, w_10000_4102, w_10000_4103, w_10000_4104, w_10000_4105, w_10000_4106, w_10000_4107, w_10000_4108, w_10000_4109, w_10000_4110, w_10000_4111, w_10000_4112, w_10000_4113, w_10000_4114, w_10000_4115, w_10000_4116, w_10000_4117, w_10000_4118, w_10000_4119, w_10000_4120, w_10000_4121, w_10000_4122, w_10000_4123, w_10000_4124, w_10000_4125, w_10000_4126, w_10000_4127, w_10000_4128, w_10000_4129, w_10000_4130, w_10000_4131, w_10000_4132, w_10000_4133, w_10000_4134, w_10000_4135, w_10000_4136, w_10000_4137, w_10000_4138, w_10000_4139, w_10000_4140, w_10000_4141, w_10000_4142, w_10000_4143, w_10000_4144, w_10000_4145, w_10000_4146, w_10000_4147, w_10000_4148, w_10000_4149, w_10000_4150, w_10000_4151, w_10000_4152, w_10000_4153, w_10000_4154, w_10000_4155, w_10000_4156, w_10000_4157, w_10000_4158, w_10000_4159, w_10000_4160, w_10000_4161, w_10000_4162, w_10000_4163, w_10000_4164, w_10000_4165, w_10000_4166, w_10000_4167, w_10000_4168, w_10000_4169, w_10000_4170, w_10000_4171, w_10000_4172, w_10000_4173, w_10000_4174, w_10000_4175, w_10000_4176, w_10000_4177, w_10000_4178, w_10000_4179, w_10000_4180, w_10000_4181, w_10000_4182, w_10000_4183, w_10000_4184, w_10000_4185, w_10000_4186, w_10000_4187, w_10000_4188, w_10000_4189, w_10000_4190, w_10000_4191, w_10000_4192, w_10000_4193, w_10000_4194, w_10000_4195, w_10000_4196, w_10000_4197, w_10000_4198, w_10000_4199, w_10000_4200, w_10000_4201, w_10000_4202, w_10000_4203, w_10000_4204, w_10000_4205, w_10000_4206, w_10000_4207, w_10000_4208, w_10000_4209, w_10000_4210, w_10000_4211, w_10000_4212, w_10000_4213, w_10000_4214, w_10000_4215, w_10000_4216, w_10000_4217, w_10000_4218, w_10000_4219, w_10000_4220, w_10000_4221, w_10000_4222, w_10000_4223, w_10000_4224, w_10000_4225, w_10000_4226, w_10000_4227, w_10000_4228, w_10000_4229, w_10000_4230, w_10000_4231, w_10000_4232, w_10000_4233, w_10000_4234, w_10000_4235, w_10000_4236, w_10000_4237, w_10000_4238, w_10000_4239, w_10000_4240, w_10000_4241, w_10000_4242, w_10000_4243, w_10000_4244, w_10000_4245, w_10000_4246, w_10000_4247, w_10000_4248, w_10000_4249, w_10000_4250, w_10000_4251, w_10000_4252, w_10000_4253, w_10000_4254, w_10000_4255, w_10000_4256, w_10000_4257, w_10000_4258, w_10000_4259, w_10000_4260, w_10000_4261, w_10000_4262, w_10000_4263, w_10000_4264, w_10000_4265, w_10000_4266, w_10000_4267, w_10000_4268, w_10000_4269, w_10000_4270, w_10000_4271, w_10000_4272, w_10000_4273, w_10000_4274, w_10000_4275, w_10000_4276, w_10000_4277, w_10000_4278, w_10000_4279, w_10000_4280, w_10000_4281, w_10000_4282, w_10000_4283, w_10000_4284, w_10000_4285, w_10000_4286, w_10000_4287, w_10000_4288, w_10000_4289, w_10000_4290, w_10000_4291, w_10000_4292, w_10000_4293, w_10000_4294, w_10000_4295, w_10000_4296, w_10000_4297, w_10000_4298, w_10000_4299, w_10000_4300, w_10000_4301, w_10000_4302, w_10000_4303, w_10000_4304, w_10000_4305, w_10000_4306, w_10000_4307, w_10000_4308, w_10000_4309, w_10000_4310, w_10000_4311, w_10000_4312, w_10000_4313, w_10000_4314, w_10000_4315, w_10000_4316, w_10000_4317, w_10000_4318, w_10000_4319, w_10000_4320, w_10000_4321, w_10000_4322, w_10000_4323, w_10000_4324, w_10000_4325, w_10000_4326, w_10000_4327, w_10000_4328, w_10000_4329, w_10000_4330, w_10000_4331, w_10000_4332, w_10000_4333, w_10000_4334, w_10000_4335, w_10000_4336, w_10000_4337, w_10000_4338, w_10000_4339, w_10000_4340, w_10000_4341, w_10000_4342, w_10000_4343, w_10000_4344, w_10000_4345, w_10000_4346, w_10000_4347, w_10000_4348, w_10000_4349, w_10000_4350, w_10000_4351, w_10000_4352, w_10000_4353, w_10000_4354, w_10000_4355, w_10000_4356, w_10000_4357, w_10000_4358, w_10000_4359, w_10000_4360, w_10000_4361, w_10000_4362, w_10000_4363, w_10000_4364, w_10000_4365, w_10000_4366, w_10000_4367, w_10000_4368, w_10000_4369, w_10000_4370, w_10000_4371, w_10000_4372, w_10000_4373, w_10000_4374, w_10000_4375, w_10000_4376, w_10000_4377, w_10000_4378, w_10000_4379, w_10000_4380, w_10000_4381, w_10000_4382, w_10000_4383, w_10000_4384, w_10000_4385, w_10000_4386, w_10000_4387, w_10000_4388, w_10000_4389, w_10000_4390, w_10000_4391, w_10000_4392, w_10000_4393, w_10000_4394, w_10000_4395, w_10000_4396, w_10000_4397, w_10000_4398, w_10000_4399, w_10000_4400, w_10000_4401, w_10000_4402, w_10000_4403, w_10000_4404, w_10000_4405, w_10000_4406, w_10000_4407, w_10000_4408, w_10000_4409, w_10000_4410, w_10000_4411, w_10000_4412, w_10000_4413, w_10000_4414, w_10000_4415, w_10000_4416, w_10000_4417, w_10000_4418, w_10000_4419, w_10000_4420, w_10000_4421, w_10000_4422, w_10000_4423, w_10000_4424, w_10000_4425, w_10000_4426, w_10000_4427, w_10000_4428, w_10000_4429, w_10000_4430, w_10000_4431, w_10000_4432, w_10000_4433, w_10000_4434, w_10000_4435, w_10000_4436, w_10000_4437, w_10000_4438, w_10000_4439, w_10000_4440, w_10000_4441, w_10000_4442, w_10000_4443, w_10000_4444, w_10000_4445, w_10000_4446, w_10000_4447, w_10000_4448, w_10000_4449, w_10000_4450, w_10000_4451, w_10000_4452, w_10000_4453, w_10000_4454, w_10000_4455, w_10000_4456, w_10000_4457, w_10000_4458, w_10000_4459, w_10000_4460, w_10000_4461, w_10000_4462, w_10000_4463, w_10000_4464, w_10000_4465, w_10000_4466, w_10000_4467, w_10000_4468, w_10000_4469, w_10000_4470, w_10000_4471, w_10000_4472, w_10000_4473, w_10000_4474, w_10000_4475, w_10000_4476, w_10000_4477, w_10000_4478, w_10000_4479, w_10000_4480, w_10000_4481, w_10000_4482, w_10000_4483, w_10000_4484, w_10000_4485, w_10000_4486, w_10000_4487, w_10000_4488, w_10000_4489, w_10000_4490, w_10000_4491, w_10000_4492, w_10000_4493, w_10000_4494, w_10000_4495, w_10000_4496, w_10000_4497, w_10000_4498, w_10000_4499, w_10000_4500, w_10000_4501, w_10000_4502, w_10000_4503, w_10000_4504, w_10000_4505, w_10000_4506, w_10000_4507, w_10000_4508, w_10000_4509, w_10000_4510, w_10000_4511, w_10000_4512, w_10000_4513, w_10000_4514, w_10000_4515, w_10000_4516, w_10000_4517, w_10000_4518, w_10000_4519, w_10000_4520, w_10000_4521, w_10000_4522, w_10000_4523, w_10000_4524, w_10000_4525, w_10000_4526, w_10000_4527, w_10000_4528, w_10000_4529, w_10000_4530, w_10000_4531, w_10000_4532, w_10000_4533, w_10000_4534, w_10000_4535, w_10000_4536, w_10000_4537, w_10000_4538, w_10000_4539, w_10000_4540, w_10000_4541, w_10000_4542, w_10000_4543, w_10000_4544, w_10000_4545, w_10000_4546, w_10000_4547, w_10000_4548, w_10000_4549, w_10000_4550, w_10000_4551, w_10000_4552, w_10000_4553, w_10000_4554, w_10000_4555, w_10000_4556, w_10000_4557, w_10000_4558, w_10000_4559, w_10000_4560, w_10000_4561, w_10000_4562, w_10000_4563, w_10000_4564, w_10000_4565, w_10000_4566, w_10000_4567, w_10000_4568, w_10000_4569, w_10000_4570, w_10000_4571, w_10000_4572, w_10000_4573, w_10000_4574, w_10000_4575, w_10000_4576, w_10000_4577, w_10000_4578, w_10000_4579, w_10000_4580, w_10000_4581, w_10000_4582, w_10000_4583, w_10000_4584, w_10000_4585, w_10000_4586, w_10000_4587, w_10000_4588, w_10000_4589, w_10000_4590, w_10000_4591, w_10000_4592, w_10000_4593, w_10000_4594, w_10000_4595, w_10000_4596, w_10000_4597, w_10000_4598, w_10000_4599, w_10000_4600, w_10000_4601, w_10000_4602, w_10000_4603, w_10000_4604, w_10000_4605, w_10000_4606, w_10000_4607, w_10000_4608, w_10000_4609, w_10000_4610, w_10000_4611, w_10000_4612, w_10000_4613, w_10000_4614, w_10000_4615, w_10000_4616, w_10000_4617, w_10000_4618, w_10000_4619, w_10000_4620, w_10000_4621, w_10000_4622, w_10000_4623, w_10000_4624, w_10000_4625, w_10000_4626, w_10000_4627, w_10000_4628, w_10000_4629, w_10000_4630, w_10000_4631, w_10000_4632, w_10000_4633, w_10000_4634, w_10000_4635, w_10000_4636, w_10000_4637, w_10000_4638, w_10000_4639, w_10000_4640, w_10000_4641, w_10000_4642, w_10000_4643, w_10000_4644, w_10000_4645, w_10000_4646, w_10000_4647, w_10000_4648, w_10000_4649, w_10000_4650, w_10000_4651, w_10000_4652, w_10000_4653, w_10000_4654, w_10000_4655, w_10000_4656, w_10000_4657, w_10000_4658, w_10000_4659, w_10000_4660, w_10000_4661, w_10000_4662, w_10000_4663, w_10000_4664, w_10000_4665, w_10000_4666, w_10000_4667, w_10000_4668, w_10000_4669, w_10000_4670, w_10000_4671, w_10000_4672, w_10000_4673, w_10000_4674, w_10000_4675, w_10000_4676, w_10000_4677, w_10000_4678, w_10000_4679, w_10000_4680, w_10000_4681, w_10000_4682, w_10000_4683, w_10000_4684, w_10000_4685, w_10000_4686, w_10000_4687, w_10000_4688, w_10000_4689, w_10000_4690, w_10000_4691, w_10000_4692, w_10000_4693, w_10000_4694, w_10000_4695, w_10000_4696, w_10000_4697, w_10000_4698, w_10000_4699, w_10000_4700, w_10000_4701, w_10000_4702, w_10000_4703, w_10000_4704, w_10000_4705, w_10000_4706, w_10000_4707, w_10000_4708, w_10000_4709, w_10000_4710, w_10000_4711, w_10000_4712, w_10000_4713, w_10000_4714, w_10000_4715, w_10000_4716, w_10000_4717, w_10000_4718, w_10000_4719, w_10000_4720, w_10000_4721, w_10000_4722, w_10000_4723, w_10000_4724, w_10000_4725, w_10000_4726, w_10000_4727, w_10000_4728, w_10000_4729, w_10000_4730, w_10000_4731, w_10000_4732, w_10000_4733, w_10000_4734, w_10000_4735, w_10000_4736, w_10000_4737, w_10000_4738, w_10000_4739, w_10000_4740, w_10000_4741, w_10000_4742, w_10000_4743, w_10000_4744, w_10000_4745, w_10000_4746, w_10000_4747, w_10000_4748, w_10000_4749, w_10000_4750, w_10000_4751, w_10000_4752, w_10000_4753, w_10000_4754, w_10000_4755, w_10000_4756, w_10000_4757, w_10000_4758, w_10000_4759, w_10000_4760, w_10000_4761, w_10000_4762, w_10000_4763, w_10000_4764, w_10000_4765, w_10000_4766, w_10000_4767, w_10000_4768, w_10000_4769, w_10000_4770, w_10000_4771, w_10000_4772, w_10000_4773, w_10000_4774, w_10000_4775, w_10000_4776, w_10000_4777, w_10000_4778, w_10000_4779, w_10000_4780, w_10000_4781, w_10000_4782, w_10000_4783, w_10000_4784, w_10000_4785, w_10000_4786, w_10000_4787, w_10000_4788, w_10000_4789, w_10000_4790, w_10000_4791, w_10000_4792, w_10000_4793, w_10000_4794, w_10000_4795, w_10000_4796, w_10000_4797, w_10000_4798, w_10000_4799, w_10000_4800, w_10000_4801, w_10000_4802, w_10000_4803, w_10000_4804, w_10000_4805, w_10000_4806, w_10000_4807, w_10000_4808, w_10000_4809, w_10000_4810, w_10000_4811, w_10000_4812, w_10000_4813, w_10000_4814, w_10000_4815, w_10000_4816, w_10000_4817, w_10000_4818, w_10000_4819, w_10000_4820, w_10000_4821, w_10000_4822, w_10000_4823, w_10000_4824, w_10000_4825, w_10000_4826, w_10000_4827, w_10000_4828, w_10000_4829, w_10000_4830, w_10000_4831, w_10000_4832, w_10000_4833, w_10000_4834, w_10000_4835, w_10000_4836, w_10000_4837, w_10000_4838, w_10000_4839, w_10000_4840, w_10000_4841, w_10000_4842, w_10000_4843, w_10000_4844, w_10000_4845, w_10000_4846, w_10000_4847, w_10000_4848, w_10000_4849, w_10000_4850, w_10000_4851, w_10000_4852, w_10000_4853, w_10000_4854, w_10000_4855, w_10000_4856, w_10000_4857, w_10000_4858, w_10000_4859, w_10000_4860, w_10000_4861, w_10000_4862, w_10000_4863, w_10000_4864, w_10000_4865, w_10000_4866, w_10000_4867, w_10000_4868, w_10000_4869, w_10000_4870, w_10000_4871, w_10000_4872, w_10000_4873, w_10000_4874, w_10000_4875, w_10000_4876, w_10000_4877, w_10000_4878, w_10000_4879, w_10000_4880, w_10000_4881, w_10000_4882, w_10000_4883, w_10000_4884, w_10000_4885, w_10000_4886, w_10000_4887, w_10000_4888, w_10000_4889, w_10000_4890, w_10000_4891, w_10000_4892, w_10000_4893, w_10000_4894, w_10000_4895, w_10000_4896, w_10000_4897, w_10000_4898, w_10000_4899, w_10000_4900, w_10000_4901, w_10000_4902, w_10000_4903, w_10000_4904, w_10000_4905, w_10000_4906, w_10000_4907, w_10000_4908, w_10000_4909, w_10000_4910, w_10000_4911, w_10000_4912, w_10000_4913, w_10000_4914, w_10000_4915, w_10000_4916, w_10000_4917, w_10000_4918, w_10000_4919, w_10000_4920, w_10000_4921, w_10000_4922, w_10000_4923, w_10000_4924, w_10000_4925, w_10000_4926, w_10000_4927, w_10000_4928, w_10000_4929, w_10000_4930, w_10000_4931, w_10000_4932, w_10000_4933, w_10000_4934, w_10000_4935, w_10000_4936, w_10000_4937, w_10000_4938, w_10000_4939, w_10000_4940, w_10000_4941, w_10000_4942, w_10000_4943, w_10000_4944, w_10000_4945, w_10000_4946, w_10000_4947, w_10000_4948, w_10000_4949, w_10000_4950, w_10000_4951, w_10000_4952, w_10000_4953, w_10000_4954, w_10000_4955, w_10000_4956, w_10000_4957, w_10000_4958, w_10000_4959, w_10000_4960, w_10000_4961, w_10000_4962, w_10000_4963, w_10000_4964, w_10000_4965, w_10000_4966, w_10000_4967, w_10000_4968, w_10000_4969, w_10000_4970, w_10000_4971, w_10000_4972, w_10000_4973, w_10000_4974, w_10000_4975, w_10000_4976, w_10000_4977, w_10000_4978, w_10000_4979, w_10000_4980, w_10000_4981, w_10000_4982, w_10000_4983, w_10000_4984, w_10000_4985, w_10000_4986, w_10000_4987, w_10000_4988, w_10000_4989, w_10000_4990, w_10000_4991, w_10000_4992, w_10000_4993, w_10000_4994, w_10000_4995, w_10000_4996, w_10000_4997, w_10000_4998, w_10000_4999, w_10000_5000, w_10000_5001, w_10000_5002, w_10000_5003, w_10000_5004, w_10000_5005, w_10000_5006, w_10000_5007, w_10000_5008, w_10000_5009, w_10000_5010, w_10000_5011, w_10000_5012, w_10000_5013, w_10000_5014, w_10000_5015, w_10000_5016, w_10000_5017, w_10000_5018, w_10000_5019, w_10000_5020, w_10000_5021, w_10000_5022, w_10000_5023, w_10000_5024, w_10000_5025, w_10000_5026, w_10000_5027, w_10000_5028, w_10000_5029, w_10000_5030, w_10000_5031, w_10000_5032, w_10000_5033, w_10000_5034, w_10000_5035, w_10000_5036, w_10000_5037, w_10000_5038, w_10000_5039, w_10000_5040, w_10000_5041, w_10000_5042, w_10000_5043, w_10000_5044, w_10000_5045, w_10000_5046, w_10000_5047, w_10000_5048, w_10000_5049, w_10000_5050, w_10000_5051, w_10000_5052, w_10000_5053, w_10000_5054, w_10000_5055, w_10000_5056, w_10000_5057, w_10000_5058, w_10000_5059, w_10000_5060, w_10000_5061, w_10000_5062, w_10000_5063, w_10000_5064, w_10000_5065, w_10000_5066, w_10000_5067, w_10000_5068, w_10000_5069, w_10000_5070, w_10000_5071, w_10000_5072, w_10000_5073, w_10000_5074, w_10000_5075, w_10000_5076, w_10000_5077, w_10000_5078, w_10000_5079, w_10000_5080, w_10000_5081, w_10000_5082, w_10000_5083, w_10000_5084, w_10000_5085, w_10000_5086, w_10000_5087, w_10000_5088, w_10000_5089, w_10000_5090, w_10000_5091, w_10000_5092, w_10000_5093, w_10000_5094, w_10000_5095, w_10000_5096, w_10000_5097, w_10000_5098, w_10000_5099, w_10000_5100, w_10000_5101, w_10000_5102, w_10000_5103, w_10000_5104, w_10000_5105, w_10000_5106, w_10000_5107, w_10000_5108, w_10000_5109, w_10000_5110, w_10000_5111, w_10000_5112, w_10000_5113, w_10000_5114, w_10000_5115, w_10000_5116, w_10000_5117, w_10000_5118, w_10000_5119, w_10000_5120, w_10000_5121, w_10000_5122, w_10000_5123, w_10000_5124, w_10000_5125, w_10000_5126, w_10000_5127, w_10000_5128, w_10000_5129, w_10000_5130, w_10000_5131, w_10000_5132, w_10000_5133, w_10000_5134, w_10000_5135, w_10000_5136, w_10000_5137, w_10000_5138, w_10000_5139, w_10000_5140, w_10000_5141, w_10000_5142, w_10000_5143, w_10000_5144, w_10000_5145, w_10000_5146, w_10000_5147, w_10000_5148, w_10000_5149, w_10000_5150, w_10000_5151, w_10000_5152, w_10000_5153, w_10000_5154, w_10000_5155, w_10000_5156, w_10000_5157, w_10000_5158, w_10000_5159, w_10000_5160, w_10000_5161, w_10000_5162, w_10000_5163, w_10000_5164, w_10000_5165, w_10000_5166, w_10000_5167, w_10000_5168, w_10000_5169, w_10000_5170, w_10000_5171, w_10000_5172, w_10000_5173, w_10000_5174, w_10000_5175, w_10000_5176, w_10000_5177, w_10000_5178, w_10000_5179, w_10000_5180, w_10000_5181, w_10000_5182, w_10000_5183, w_10000_5184, w_10000_5185, w_10000_5186, w_10000_5187, w_10000_5188, w_10000_5189, w_10000_5190, w_10000_5191, w_10000_5192, w_10000_5193, w_10000_5194, w_10000_5195, w_10000_5196, w_10000_5197, w_10000_5198, w_10000_5199, w_10000_5200, w_10000_5201, w_10000_5202, w_10000_5203, w_10000_5204, w_10000_5205, w_10000_5206, w_10000_5207, w_10000_5208, w_10000_5209, w_10000_5210, w_10000_5211, w_10000_5212, w_10000_5213, w_10000_5214, w_10000_5215, w_10000_5216, w_10000_5217, w_10000_5218, w_10000_5219, w_10000_5220, w_10000_5221, w_10000_5222, w_10000_5223, w_10000_5224, w_10000_5225, w_10000_5226, w_10000_5227, w_10000_5228, w_10000_5229, w_10000_5230, w_10000_5231, w_10000_5232, w_10000_5233, w_10000_5234, w_10000_5235, w_10000_5236, w_10000_5237, w_10000_5238, w_10000_5239, w_10000_5240, w_10000_5241, w_10000_5242, w_10000_5243, w_10000_5244, w_10000_5245, w_10000_5246, w_10000_5247, w_10000_5248, w_10000_5249, w_10000_5250, w_10000_5251, w_10000_5252, w_10000_5253, w_10000_5254, w_10000_5255, w_10000_5256, w_10000_5257, w_10000_5258, w_10000_5259, w_10000_5260, w_10000_5261, w_10000_5262, w_10000_5263, w_10000_5264, w_10000_5265, w_10000_5266, w_10000_5267, w_10000_5268, w_10000_5269, w_10000_5270, w_10000_5271, w_10000_5272, w_10000_5273, w_10000_5274, w_10000_5275, w_10000_5276, w_10000_5277, w_10000_5278, w_10000_5279, w_10000_5280, w_10000_5281, w_10000_5282, w_10000_5283, w_10000_5284, w_10000_5285, w_10000_5286, w_10000_5287, w_10000_5288, w_10000_5289, w_10000_5290, w_10000_5291, w_10000_5292, w_10000_5293, w_10000_5294, w_10000_5295, w_10000_5296, w_10000_5297, w_10000_5298, w_10000_5299, w_10000_5300, w_10000_5301, w_10000_5302, w_10000_5303, w_10000_5304, w_10000_5305, w_10000_5306, w_10000_5307, w_10000_5308, w_10000_5309, w_10000_5310, w_10000_5311, w_10000_5312, w_10000_5313, w_10000_5314, w_10000_5315, w_10000_5316, w_10000_5317, w_10000_5318, w_10000_5319, w_10000_5320, w_10000_5321, w_10000_5322, w_10000_5323, w_10000_5324, w_10000_5325, w_10000_5326, w_10000_5327, w_10000_5328, w_10000_5329, w_10000_5330, w_10000_5331, w_10000_5332, w_10000_5333, w_10000_5334, w_10000_5335, w_10000_5336, w_10000_5337, w_10000_5338, w_10000_5339, w_10000_5340, w_10000_5341, w_10000_5342, w_10000_5343, w_10000_5344, w_10000_5345, w_10000_5346, w_10000_5347, w_10000_5348, w_10000_5349, w_10000_5350, w_10000_5351, w_10000_5352, w_10000_5353, w_10000_5354, w_10000_5355, w_10000_5356, w_10000_5357, w_10000_5358, w_10000_5359, w_10000_5360, w_10000_5361, w_10000_5362, w_10000_5363, w_10000_5364, w_10000_5365, w_10000_5366, w_10000_5367, w_10000_5368, w_10000_5369, w_10000_5370, w_10000_5371, w_10000_5372, w_10000_5373, w_10000_5374, w_10000_5375, w_10000_5376, w_10000_5377, w_10000_5378, w_10000_5379, w_10000_5380, w_10000_5381, w_10000_5382, w_10000_5383, w_10000_5384, w_10000_5385, w_10000_5386, w_10000_5387, w_10000_5388, w_10000_5389, w_10000_5390, w_10000_5391, w_10000_5392, w_10000_5393, w_10000_5394, w_10000_5395, w_10000_5396, w_10000_5397, w_10000_5398, w_10000_5399, w_10000_5400, w_10000_5401, w_10000_5402, w_10000_5403, w_10000_5404, w_10000_5405, w_10000_5406, w_10000_5407, w_10000_5408, w_10000_5409, w_10000_5410, w_10000_5411, w_10000_5412, w_10000_5413, w_10000_5414, w_10000_5415, w_10000_5416, w_10000_5417, w_10000_5418, w_10000_5419, w_10000_5420, w_10000_5421, w_10000_5422, w_10000_5423, w_10000_5424, w_10000_5425, w_10000_5426, w_10000_5427, w_10000_5428, w_10000_5429, w_10000_5430, w_10000_5431, w_10000_5432, w_10000_5433, w_10000_5434, w_10000_5435, w_10000_5436, w_10000_5437, w_10000_5438, w_10000_5439, w_10000_5440, w_10000_5441, w_10000_5442, w_10000_5443, w_10000_5444, w_10000_5445, w_10000_5446, w_10000_5447, w_10000_5448, w_10000_5449, w_10000_5450, w_10000_5451, w_10000_5452, w_10000_5453, w_10000_5454, w_10000_5455, w_10000_5456, w_10000_5457, w_10000_5458, w_10000_5459, w_10000_5460, w_10000_5461, w_10000_5462, w_10000_5463, w_10000_5464, w_10000_5465, w_10000_5466, w_10000_5467, w_10000_5468, w_10000_5469, w_10000_5470, w_10000_5471, w_10000_5472, w_10000_5473, w_10000_5474, w_10000_5475, w_10000_5476, w_10000_5477, w_10000_5478, w_10000_5479, w_10000_5480, w_10000_5481, w_10000_5482, w_10000_5483, w_10000_5484, w_10000_5485, w_10000_5486, w_10000_5487, w_10000_5488, w_10000_5489, w_10000_5490, w_10000_5491, w_10000_5492, w_10000_5493, w_10000_5494, w_10000_5495, w_10000_5496, w_10000_5497, w_10000_5498, w_10000_5499, w_10000_5500, w_10000_5501, w_10000_5502, w_10000_5503, w_10000_5504, w_10000_5505, w_10000_5506, w_10000_5507, w_10000_5508, w_10000_5509, w_10000_5510, w_10000_5511, w_10000_5512, w_10000_5513, w_10000_5514, w_10000_5515, w_10000_5516, w_10000_5517, w_10000_5518, w_10000_5519, w_10000_5520, w_10000_5521, w_10000_5522, w_10000_5523, w_10000_5524, w_10000_5525, w_10000_5526, w_10000_5527, w_10000_5528, w_10000_5529, w_10000_5530, w_10000_5531, w_10000_5532, w_10000_5533, w_10000_5534, w_10000_5535, w_10000_5536, w_10000_5537, w_10000_5538, w_10000_5539, w_10000_5540, w_10000_5541, w_10000_5542, w_10000_5543, w_10000_5544, w_10000_5545, w_10000_5546, w_10000_5547, w_10000_5548, w_10000_5549, w_10000_5550, w_10000_5551, w_10000_5552, w_10000_5553, w_10000_5554, w_10000_5555, w_10000_5556, w_10000_5557, w_10000_5558, w_10000_5559, w_10000_5560, w_10000_5561, w_10000_5562, w_10000_5563, w_10000_5564, w_10000_5565, w_10000_5566, w_10000_5567, w_10000_5568, w_10000_5569, w_10000_5570, w_10000_5571, w_10000_5572, w_10000_5573, w_10000_5574, w_10000_5575, w_10000_5576, w_10000_5577, w_10000_5578, w_10000_5579, w_10000_5580, w_10000_5581, w_10000_5582, w_10000_5583, w_10000_5584, w_10000_5585, w_10000_5586, w_10000_5587, w_10000_5588, w_10000_5589, w_10000_5590, w_10000_5591, w_10000_5592, w_10000_5593, w_10000_5594, w_10000_5595, w_10000_5596, w_10000_5597, w_10000_5598, w_10000_5599, w_10000_5600, w_10000_5601, w_10000_5602, w_10000_5603, w_10000_5604, w_10000_5605, w_10000_5606, w_10000_5607, w_10000_5608, w_10000_5609, w_10000_5610, w_10000_5611, w_10000_5612, w_10000_5613, w_10000_5614, w_10000_5615, w_10000_5616, w_10000_5617, w_10000_5618, w_10000_5619, w_10000_5620, w_10000_5621, w_10000_5622, w_10000_5623, w_10000_5624, w_10000_5625, w_10000_5626, w_10000_5627, w_10000_5628, w_10000_5629, w_10000_5630, w_10000_5631, w_10000_5632, w_10000_5633, w_10000_5634, w_10000_5635, w_10000_5636, w_10000_5637, w_10000_5638, w_10000_5639, w_10000_5640, w_10000_5641, w_10000_5642, w_10000_5643, w_10000_5644, w_10000_5645, w_10000_5646, w_10000_5647, w_10000_5648, w_10000_5649, w_10000_5650, w_10000_5651, w_10000_5652, w_10000_5653, w_10000_5654, w_10000_5655, w_10000_5656, w_10000_5657, w_10000_5658, w_10000_5659, w_10000_5660, w_10000_5661, w_10000_5662, w_10000_5663, w_10000_5664, w_10000_5665, w_10000_5666, w_10000_5667, w_10000_5668, w_10000_5669, w_10000_5670, w_10000_5671, w_10000_5672, w_10000_5673, w_10000_5674, w_10000_5675, w_10000_5676, w_10000_5677, w_10000_5678, w_10000_5679, w_10000_5680, w_10000_5681, w_10000_5682, w_10000_5683, w_10000_5684, w_10000_5685, w_10000_5686, w_10000_5687, w_10000_5688, w_10000_5689, w_10000_5690, w_10000_5691, w_10000_5692, w_10000_5693, w_10000_5694, w_10000_5695, w_10000_5696, w_10000_5697, w_10000_5698, w_10000_5699, w_10000_5700, w_10000_5701, w_10000_5702, w_10000_5703, w_10000_5704, w_10000_5705, w_10000_5706, w_10000_5707, w_10000_5708, w_10000_5709, w_10000_5710, w_10000_5711, w_10000_5712, w_10000_5713, w_10000_5714, w_10000_5715, w_10000_5716, w_10000_5717, w_10000_5718, w_10000_5719, w_10000_5720, w_10000_5721, w_10000_5722, w_10000_5723, w_10000_5724, w_10000_5725, w_10000_5726, w_10000_5727, w_10000_5728, w_10000_5729, w_10000_5730, w_10000_5731, w_10000_5732, w_10000_5733, w_10000_5734, w_10000_5735, w_10000_5736, w_10000_5737, w_10000_5738, w_10000_5739, w_10000_5740, w_10000_5741, w_10000_5742, w_10000_5743, w_10000_5744, w_10000_5745, w_10000_5746, w_10000_5747, w_10000_5748, w_10000_5749, w_10000_5750, w_10000_5751, w_10000_5752, w_10000_5753, w_10000_5754, w_10000_5755, w_10000_5756, w_10000_5757, w_10000_5758, w_10000_5759, w_10000_5760, w_10000_5761, w_10000_5762, w_10000_5763, w_10000_5764, w_10000_5765, w_10000_5766, w_10000_5767, w_10000_5768, w_10000_5769, w_10000_5770, w_10000_5771, w_10000_5772, w_10000_5773, w_10000_5774, w_10000_5775, w_10000_5776, w_10000_5777, w_10000_5778, w_10000_5779, w_10000_5780, w_10000_5781, w_10000_5782, w_10000_5783, w_10000_5784, w_10000_5785, w_10000_5786, w_10000_5787, w_10000_5788, w_10000_5789, w_10000_5790, w_10000_5791, w_10000_5792, w_10000_5793, w_10000_5794, w_10000_5795, w_10000_5796, w_10000_5797, w_10000_5798, w_10000_5799, w_10000_5800, w_10000_5801, w_10000_5802, w_10000_5803, w_10000_5804, w_10000_5805, w_10000_5806, w_10000_5807, w_10000_5808, w_10000_5809, w_10000_5810, w_10000_5811, w_10000_5812, w_10000_5813, w_10000_5814, w_10000_5815, w_10000_5816, w_10000_5817, w_10000_5818, w_10000_5819, w_10000_5820, w_10000_5821, w_10000_5822, w_10000_5823, w_10000_5824, w_10000_5825, w_10000_5826, w_10000_5827, w_10000_5828, w_10000_5829, w_10000_5830, w_10000_5831, w_10000_5832, w_10000_5833, w_10000_5834, w_10000_5835, w_10000_5836, w_10000_5837, w_10000_5838, w_10000_5839, w_10000_5840, w_10000_5841, w_10000_5842, w_10000_5843, w_10000_5844, w_10000_5845, w_10000_5846, w_10000_5847, w_10000_5848, w_10000_5849, w_10000_5850, w_10000_5851, w_10000_5852, w_10000_5853, w_10000_5854, w_10000_5855, w_10000_5856, w_10000_5857, w_10000_5858, w_10000_5859, w_10000_5860, w_10000_5861, w_10000_5862, w_10000_5863, w_10000_5864, w_10000_5865, w_10000_5866, w_10000_5867, w_10000_5868, w_10000_5869, w_10000_5870, w_10000_5871, w_10000_5872, w_10000_5873, w_10000_5874, w_10000_5875, w_10000_5876, w_10000_5877, w_10000_5878, w_10000_5879, w_10000_5880, w_10000_5881, w_10000_5882, w_10000_5883, w_10000_5884, w_10000_5885, w_10000_5886, w_10000_5887, w_10000_5888, w_10000_5889, w_10000_5890, w_10000_5891, w_10000_5892, w_10000_5893, w_10000_5894, w_10000_5895, w_10000_5896, w_10000_5897, w_10000_5898, w_10000_5899, w_10000_5900, w_10000_5901, w_10000_5902, w_10000_5903, w_10000_5904, w_10000_5905, w_10000_5906, w_10000_5907, w_10000_5908, w_10000_5909, w_10000_5910, w_10000_5911, w_10000_5912, w_10000_5913, w_10000_5914, w_10000_5915, w_10000_5916, w_10000_5917, w_10000_5918, w_10000_5919, w_10000_5920, w_10000_5921, w_10000_5922, w_10000_5923, w_10000_5924, w_10000_5925, w_10000_5926, w_10000_5927, w_10000_5928, w_10000_5929, w_10000_5930, w_10000_5931, w_10000_5932, w_10000_5933, w_10000_5934, w_10000_5935, w_10000_5936, w_10000_5937, w_10000_5938, w_10000_5939, w_10000_5940, w_10000_5941, w_10000_5942, w_10000_5943, w_10000_5944, w_10000_5945, w_10000_5946, w_10000_5947, w_10000_5948, w_10000_5949, w_10000_5950, w_10000_5951, w_10000_5952, w_10000_5953, w_10000_5954, w_10000_5955, w_10000_5956, w_10000_5957, w_10000_5958, w_10000_5959, w_10000_5960, w_10000_5961, w_10000_5962, w_10000_5963, w_10000_5964, w_10000_5965, w_10000_5966, w_10000_5967, w_10000_5968, w_10000_5969, w_10000_5970, w_10000_5971, w_10000_5972, w_10000_5973, w_10000_5974, w_10000_5975, w_10000_5976, w_10000_5977, w_10000_5978, w_10000_5979, w_10000_5980, w_10000_5981, w_10000_5982, w_10000_5983, w_10000_5984, w_10000_5985, w_10000_5986, w_10000_5987, w_10000_5988, w_10000_5989, w_10000_5990, w_10000_5991, w_10000_5992, w_10000_5993, w_10000_5994, w_10000_5995, w_10000_5996, w_10000_5997, w_10000_5998, w_10000_5999, w_10000_6000, w_10000_6001, w_10000_6002, w_10000_6003, w_10000_6004, w_10000_6005, w_10000_6006, w_10000_6007, w_10000_6008, w_10000_6009, w_10000_6010, w_10000_6011, w_10000_6012, w_10000_6013, w_10000_6014, w_10000_6015, w_10000_6016, w_10000_6017, w_10000_6018, w_10000_6019, w_10000_6020, w_10000_6021, w_10000_6022, w_10000_6023, w_10000_6024, w_10000_6025, w_10000_6026, w_10000_6027, w_10000_6028, w_10000_6029, w_10000_6030, w_10000_6031, w_10000_6032, w_10000_6033, w_10000_6034, w_10000_6035, w_10000_6036, w_10000_6037, w_10000_6038, w_10000_6039, w_10000_6040, w_10000_6041, w_10000_6042, w_10000_6043, w_10000_6044, w_10000_6045, w_10000_6046, w_10000_6047, w_10000_6048, w_10000_6049, w_10000_6050, w_10000_6051, w_10000_6052, w_10000_6053, w_10000_6054, w_10000_6055, w_10000_6056, w_10000_6057, w_10000_6058, w_10000_6059, w_10000_6060, w_10000_6061, w_10000_6062, w_10000_6063, w_10000_6064, w_10000_6065, w_10000_6066, w_10000_6067, w_10000_6068, w_10000_6069, w_10000_6070, w_10000_6071, w_10000_6072, w_10000_6073, w_10000_6074, w_10000_6075, w_10000_6076, w_10000_6077, w_10000_6078, w_10000_6079, w_10000_6080, w_10000_6081, w_10000_6082, w_10000_6083, w_10000_6084, w_10000_6085, w_10000_6086, w_10000_6087, w_10000_6088, w_10000_6089, w_10000_6090, w_10000_6091, w_10000_6092, w_10000_6093, w_10000_6094, w_10000_6095, w_10000_6096, w_10000_6097, w_10000_6098, w_10000_6099, w_10000_6100, w_10000_6101, w_10000_6102, w_10000_6103, w_10000_6104, w_10000_6105, w_10000_6106, w_10000_6107, w_10000_6108, w_10000_6109, w_10000_6110, w_10000_6111, w_10000_6112, w_10000_6113, w_10000_6114, w_10000_6115, w_10000_6116, w_10000_6117, w_10000_6118, w_10000_6119, w_10000_6120, w_10000_6121, w_10000_6122, w_10000_6123, w_10000_6124, w_10000_6125, w_10000_6126, w_10000_6127, w_10000_6128, w_10000_6129, w_10000_6130, w_10000_6131, w_10000_6132, w_10000_6133, w_10000_6134, w_10000_6135, w_10000_6136, w_10000_6137, w_10000_6138, w_10000_6139, w_10000_6140, w_10000_6141, w_10000_6142, w_10000_6143, w_10000_6144, w_10000_6145, w_10000_6146, w_10000_6147, w_10000_6148, w_10000_6149, w_10000_6150, w_10000_6151, w_10000_6152, w_10000_6153, w_10000_6154, w_10000_6155, w_10000_6156, w_10000_6157, w_10000_6158, w_10000_6159, w_10000_6160, w_10000_6161, w_10000_6162, w_10000_6163, w_10000_6164, w_10000_6165, w_10000_6166, w_10000_6167, w_10000_6168, w_10000_6169, w_10000_6170, w_10000_6171, w_10000_6172, w_10000_6173, w_10000_6174, w_10000_6175, w_10000_6176, w_10000_6177, w_10000_6178, w_10000_6179, w_10000_6180, w_10000_6181, w_10000_6182, w_10000_6183, w_10000_6184, w_10000_6185, w_10000_6186, w_10000_6187, w_10000_6188, w_10000_6189, w_10000_6190, w_10000_6191, w_10000_6192, w_10000_6193, w_10000_6194, w_10000_6195, w_10000_6196, w_10000_6197, w_10000_6198, w_10000_6199, w_10000_6200, w_10000_6201, w_10000_6202, w_10000_6203, w_10000_6204, w_10000_6205, w_10000_6206, w_10000_6207, w_10000_6208, w_10000_6209, w_10000_6210, w_10000_6211, w_10000_6212, w_10000_6213, w_10000_6214, w_10000_6215, w_10000_6216, w_10000_6217, w_10000_6218, w_10000_6219, w_10000_6220, w_10000_6221, w_10000_6222, w_10000_6223, w_10000_6224, w_10000_6225, w_10000_6226, w_10000_6227, w_10000_6228, w_10000_6229, w_10000_6230, w_10000_6231, w_10000_6232, w_10000_6233, w_10000_6234, w_10000_6235, w_10000_6236, w_10000_6237, w_10000_6238, w_10000_6239, w_10000_6240, w_10000_6241, w_10000_6242, w_10000_6243, w_10000_6244, w_10000_6245, w_10000_6246, w_10000_6247, w_10000_6248, w_10000_6249, w_10000_6250, w_10000_6251, w_10000_6252, w_10000_6253, w_10000_6254, w_10000_6255, w_10000_6256, w_10000_6257, w_10000_6258, w_10000_6259, w_10000_6260, w_10000_6261, w_10000_6262, w_10000_6263, w_10000_6264, w_10000_6265, w_10000_6266, w_10000_6267, w_10000_6268, w_10000_6269, w_10000_6270, w_10000_6271, w_10000_6272, w_10000_6273, w_10000_6274, w_10000_6275, w_10000_6276, w_10000_6277, w_10000_6278, w_10000_6279, w_10000_6280, w_10000_6281, w_10000_6282, w_10000_6283, w_10000_6284, w_10000_6285, w_10000_6286, w_10000_6287, w_10000_6288, w_10000_6289, w_10000_6290, w_10000_6291, w_10000_6292, w_10000_6293, w_10000_6294, w_10000_6295, w_10000_6296, w_10000_6297, w_10000_6298, w_10000_6299, w_10000_6300, w_10000_6301, w_10000_6302, w_10000_6303, w_10000_6304, w_10000_6305, w_10000_6306, w_10000_6307, w_10000_6308, w_10000_6309, w_10000_6310, w_10000_6311, w_10000_6312, w_10000_6313, w_10000_6314, w_10000_6315, w_10000_6316, w_10000_6317, w_10000_6318, w_10000_6319, w_10000_6320, w_10000_6321, w_10000_6322, w_10000_6323, w_10000_6324, w_10000_6325, w_10000_6326, w_10000_6327, w_10000_6328, w_10000_6329, w_10000_6330, w_10000_6331, w_10000_6332, w_10000_6333, w_10000_6334, w_10000_6335, w_10000_6336, w_10000_6337, w_10000_6338, w_10000_6339, w_10000_6340, w_10000_6341, w_10000_6342, w_10000_6343, w_10000_6344, w_10000_6345, w_10000_6346, w_10000_6347, w_10000_6348, w_10000_6349, w_10000_6350, w_10000_6351, w_10000_6352, w_10000_6353, w_10000_6354, w_10000_6355, w_10000_6356, w_10000_6357, w_10000_6358, w_10000_6359, w_10000_6360, w_10000_6361, w_10000_6362, w_10000_6363, w_10000_6364, w_10000_6365, w_10000_6366, w_10000_6367, w_10000_6368, w_10000_6369, w_10000_6370, w_10000_6371, w_10000_6372, w_10000_6373, w_10000_6374, w_10000_6375, w_10000_6376, w_10000_6377, w_10000_6378, w_10000_6379, w_10000_6380, w_10000_6381, w_10000_6382, w_10000_6383, w_10000_6384, w_10000_6385, w_10000_6386, w_10000_6387, w_10000_6388, w_10000_6389, w_10000_6390, w_10000_6391, w_10000_6392, w_10000_6393, w_10000_6394, w_10000_6395, w_10000_6396, w_10000_6397, w_10000_6398, w_10000_6399, w_10000_6400, w_10000_6401, w_10000_6402, w_10000_6403, w_10000_6404, w_10000_6405, w_10000_6406, w_10000_6407, w_10000_6408, w_10000_6409, w_10000_6410, w_10000_6411, w_10000_6412, w_10000_6413, w_10000_6414, w_10000_6415, w_10000_6416, w_10000_6417, w_10000_6418, w_10000_6419, w_10000_6420, w_10000_6421, w_10000_6422, w_10000_6423, w_10000_6424, w_10000_6425, w_10000_6426, w_10000_6427, w_10000_6428, w_10000_6429, w_10000_6430, w_10000_6431, w_10000_6432, w_10000_6433, w_10000_6434, w_10000_6435, w_10000_6436, w_10000_6437, w_10000_6438, w_10000_6439, w_10000_6440, w_10000_6441, w_10000_6442, w_10000_6443, w_10000_6444, w_10000_6445, w_10000_6446, w_10000_6447, w_10000_6448, w_10000_6449, w_10000_6450, w_10000_6451, w_10000_6452, w_10000_6453, w_10000_6454, w_10000_6455, w_10000_6456, w_10000_6457, w_10000_6458, w_10000_6459, w_10000_6460, w_10000_6461, w_10000_6462, w_10000_6463, w_10000_6464, w_10000_6465, w_10000_6466, w_10000_6467, w_10000_6468, w_10000_6469, w_10000_6470, w_10000_6471, w_10000_6472, w_10000_6473, w_10000_6474, w_10000_6475, w_10000_6476, w_10000_6477, w_10000_6478, w_10000_6479, w_10000_6480, w_10000_6481, w_10000_6482, w_10000_6483, w_10000_6484, w_10000_6485, w_10000_6486, w_10000_6487, w_10000_6488, w_10000_6489, w_10000_6490, w_10000_6491, w_10000_6492, w_10000_6493, w_10000_6494, w_10000_6495, w_10000_6496, w_10000_6497, w_10000_6498, w_10000_6499, w_10000_6500, w_10000_6501, w_10000_6502, w_10000_6503, w_10000_6504, w_10000_6505, w_10000_6506, w_10000_6507, w_10000_6508, w_10000_6509, w_10000_6510, w_10000_6511, w_10000_6512, w_10000_6513, w_10000_6514, w_10000_6515, w_10000_6516, w_10000_6517, w_10000_6518, w_10000_6519, w_10000_6520, w_10000_6521, w_10000_6522, w_10000_6523, w_10000_6524, w_10000_6525, w_10000_6526, w_10000_6527, w_10000_6528, w_10000_6529, w_10000_6530, w_10000_6531, w_10000_6532, w_10000_6533, w_10000_6534, w_10000_6535, w_10000_6536, w_10000_6537, w_10000_6538, w_10000_6539, w_10000_6540, w_10000_6541, w_10000_6542, w_10000_6543, w_10000_6544, w_10000_6545, w_10000_6546, w_10000_6547, w_10000_6548, w_10000_6549, w_10000_6550, w_10000_6551, w_10000_6552, w_10000_6553, w_10000_6554, w_10000_6555, w_10000_6556, w_10000_6557, w_10000_6558, w_10000_6559, w_10000_6560, w_10000_6561, w_10000_6562, w_10000_6563, w_10000_6564, w_10000_6565, w_10000_6566, w_10000_6567, w_10000_6568, w_10000_6569, w_10000_6570, w_10000_6571, w_10000_6572, w_10000_6573, w_10000_6574, w_10000_6575, w_10000_6576, w_10000_6577, w_10000_6578, w_10000_6579, w_10000_6580, w_10000_6581, w_10000_6582, w_10000_6583, w_10000_6584, w_10000_6585, w_10000_6586, w_10000_6587, w_10000_6588, w_10000_6589, w_10000_6590, w_10000_6591, w_10000_6592, w_10000_6593, w_10000_6594, w_10000_6595, w_10000_6596, w_10000_6597, w_10000_6598, w_10000_6599, w_10000_6600, w_10000_6601, w_10000_6602, w_10000_6603, w_10000_6604, w_10000_6605, w_10000_6606, w_10000_6607, w_10000_6608, w_10000_6609, w_10000_6610, w_10000_6611, w_10000_6612, w_10000_6613, w_10000_6614, w_10000_6615, w_10000_6616, w_10000_6617, w_10000_6618, w_10000_6619, w_10000_6620, w_10000_6621, w_10000_6622, w_10000_6623, w_10000_6624, w_10000_6625, w_10000_6626, w_10000_6627, w_10000_6628, w_10000_6629, w_10000_6630, w_10000_6631, w_10000_6632, w_10000_6633, w_10000_6634, w_10000_6635, w_10000_6636, w_10000_6637, w_10000_6638, w_10000_6639, w_10000_6640, w_10000_6641, w_10000_6642, w_10000_6643, w_10000_6644, w_10000_6645, w_10000_6646, w_10000_6647, w_10000_6648, w_10000_6649, w_10000_6650, w_10000_6651, w_10000_6652, w_10000_6653, w_10000_6654, w_10000_6655, w_10000_6656, w_10000_6657, w_10000_6658, w_10000_6659, w_10000_6660, w_10000_6661, w_10000_6662, w_10000_6663, w_10000_6664, w_10000_6665, w_10000_6666, w_10000_6667, w_10000_6668, w_10000_6669, w_10000_6670, w_10000_6671, w_10000_6672, w_10000_6673, w_10000_6674, w_10000_6675, w_10000_6676, w_10000_6677, w_10000_6678, w_10000_6679, w_10000_6680, w_10000_6681, w_10000_6682, w_10000_6683, w_10000_6684, w_10000_6685, w_10000_6686, w_10000_6687, w_10000_6688, w_10000_6689, w_10000_6690, w_10000_6691, w_10000_6692, w_10000_6693, w_10000_6694, w_10000_6695, w_10000_6696, w_10000_6697, w_10000_6698, w_10000_6699, w_10000_6700, w_10000_6701, w_10000_6702, w_10000_6703, w_10000_6704, w_10000_6705, w_10000_6706, w_10000_6707, w_10000_6708, w_10000_6709, w_10000_6710, w_10000_6711, w_10000_6712, w_10000_6713, w_10000_6714, w_10000_6715, w_10000_6716, w_10000_6717, w_10000_6718, w_10000_6719, w_10000_6720, w_10000_6721, w_10000_6722, w_10000_6723, w_10000_6724, w_10000_6725, w_10000_6726, w_10000_6727, w_10000_6728, w_10000_6729, w_10000_6730, w_10000_6731, w_10000_6732, w_10000_6733, w_10000_6734, w_10000_6735, w_10000_6736, w_10000_6737, w_10000_6738, w_10000_6739, w_10000_6740, w_10000_6741, w_10000_6742, w_10000_6743, w_10000_6744, w_10000_6745, w_10000_6746, w_10000_6747, w_10000_6748, w_10000_6749, w_10000_6750, w_10000_6751, w_10000_6752, w_10000_6753, w_10000_6754, w_10000_6755, w_10000_6756, w_10000_6757, w_10000_6758, w_10000_6759, w_10000_6760, w_10000_6761, w_10000_6762, w_10000_6763, w_10000_6764, w_10000_6765, w_10000_6766, w_10000_6767, w_10000_6768, w_10000_6769, w_10000_6770, w_10000_6771, w_10000_6772, w_10000_6773, w_10000_6774, w_10000_6775, w_10000_6776, w_10000_6777, w_10000_6778, w_10000_6779, w_10000_6780, w_10000_6781, w_10000_6782, w_10000_6783, w_10000_6784, w_10000_6785, w_10000_6786, w_10000_6787, w_10000_6788, w_10000_6789, w_10000_6790, w_10000_6791, w_10000_6792, w_10000_6793, w_10000_6794, w_10000_6795, w_10000_6796, w_10000_6797, w_10000_6798, w_10000_6799, w_10000_6800, w_10000_6801, w_10000_6802, w_10000_6803, w_10000_6804, w_10000_6805, w_10000_6806, w_10000_6807, w_10000_6808, w_10000_6809, w_10000_6810, w_10000_6811, w_10000_6812, w_10000_6813, w_10000_6814, w_10000_6815, w_10000_6816, w_10000_6817, w_10000_6818, w_10000_6819, w_10000_6820, w_10000_6821, w_10000_6822, w_10000_6823, w_10000_6824, w_10000_6825, w_10000_6826, w_10000_6827, w_10000_6828, w_10000_6829, w_10000_6830, w_10000_6831, w_10000_6832, w_10000_6833, w_10000_6834, w_10000_6835, w_10000_6836, w_10000_6837, w_10000_6838, w_10000_6839, w_10000_6840, w_10000_6841, w_10000_6842, w_10000_6843, w_10000_6844, w_10000_6845, w_10000_6846, w_10000_6847, w_10000_6848, w_10000_6849, w_10000_6850, w_10000_6851, w_10000_6852, w_10000_6853, w_10000_6854, w_10000_6855, w_10000_6856, w_10000_6857, w_10000_6858, w_10000_6859, w_10000_6860, w_10000_6861, w_10000_6862, w_10000_6863, w_10000_6864, w_10000_6865, w_10000_6866, w_10000_6867, w_10000_6868, w_10000_6869, w_10000_6870, w_10000_6871, w_10000_6872, w_10000_6873, w_10000_6874, w_10000_6875, w_10000_6876, w_10000_6877, w_10000_6878, w_10000_6879, w_10000_6880, w_10000_6881, w_10000_6882, w_10000_6883, w_10000_6884, w_10000_6885, w_10000_6886, w_10000_6887, w_10000_6888, w_10000_6889, w_10000_6890, w_10000_6891, w_10000_6892, w_10000_6893, w_10000_6894, w_10000_6895, w_10000_6896, w_10000_6897, w_10000_6898, w_10000_6899, w_10000_6900, w_10000_6901, w_10000_6902, w_10000_6903, w_10000_6904, w_10000_6905, w_10000_6906, w_10000_6907, w_10000_6908, w_10000_6909, w_10000_6910, w_10000_6911, w_10000_6912, w_10000_6913, w_10000_6914, w_10000_6915, w_10000_6916, w_10000_6917, w_10000_6918, w_10000_6919, w_10000_6920, w_10000_6921, w_10000_6922, w_10000_6923, w_10000_6924, w_10000_6925, w_10000_6926, w_10000_6927, w_10000_6928, w_10000_6929, w_10000_6930, w_10000_6931, w_10000_6932, w_10000_6933, w_10000_6934, w_10000_6935, w_10000_6936, w_10000_6937, w_10000_6938, w_10000_6939, w_10000_6940, w_10000_6941, w_10000_6942, w_10000_6943, w_10000_6944, w_10000_6945, w_10000_6946, w_10000_6947, w_10000_6948, w_10000_6949, w_10000_6950, w_10000_6951, w_10000_6952, w_10000_6953, w_10000_6954, w_10000_6955, w_10000_6956, w_10000_6957, w_10000_6958, w_10000_6959, w_10000_6960, w_10000_6961, w_10000_6962, w_10000_6963, w_10000_6964, w_10000_6965, w_10000_6966, w_10000_6967, w_10000_6968, w_10000_6969, w_10000_6970, w_10000_6971, w_10000_6972, w_10000_6973, w_10000_6974, w_10000_6975, w_10000_6976, w_10000_6977, w_10000_6978, w_10000_6979, w_10000_6980, w_10000_6981, w_10000_6982, w_10000_6983, w_10000_6984, w_10000_6985, w_10000_6986, w_10000_6987, w_10000_6988, w_10000_6989, w_10000_6990, w_10000_6991, w_10000_6992, w_10000_6993, w_10000_6994, w_10000_6995, w_10000_6996, w_10000_6997, w_10000_6998, w_10000_6999, w_10000_7000, w_10000_7001, w_10000_7002, w_10000_7003, w_10000_7004, w_10000_7005, w_10000_7006, w_10000_7007, w_10000_7008, w_10000_7009, w_10000_7010, w_10000_7011, w_10000_7012, w_10000_7013, w_10000_7014, w_10000_7015, w_10000_7016, w_10000_7017, w_10000_7018, w_10000_7019, w_10000_7020, w_10000_7021, w_10000_7022, w_10000_7023, w_10000_7024, w_10000_7025, w_10000_7026, w_10000_7027, w_10000_7028, w_10000_7029, w_10000_7030, w_10000_7031, w_10000_7032, w_10000_7033, w_10000_7034, w_10000_7035, w_10000_7036, w_10000_7037, w_10000_7038, w_10000_7039, w_10000_7040, w_10000_7041, w_10000_7042, w_10000_7043, w_10000_7044, w_10000_7045, w_10000_7046, w_10000_7047, w_10000_7048, w_10000_7049, w_10000_7050, w_10000_7051, w_10000_7052, w_10000_7053, w_10000_7054, w_10000_7055, w_10000_7056, w_10000_7057, w_10000_7058, w_10000_7059, w_10000_7060, w_10000_7061, w_10000_7062, w_10000_7063, w_10000_7064, w_10000_7065, w_10000_7066, w_10000_7067, w_10000_7068, w_10000_7069, w_10000_7070, w_10000_7071, w_10000_7072, w_10000_7073, w_10000_7074, w_10000_7075, w_10000_7076, w_10000_7077, w_10000_7078, w_10000_7079, w_10000_7080, w_10000_7081, w_10000_7082, w_10000_7083, w_10000_7084, w_10000_7085, w_10000_7086, w_10000_7087, w_10000_7088, w_10000_7089, w_10000_7090, w_10000_7091, w_10000_7092, w_10000_7093, w_10000_7094, w_10000_7095, w_10000_7096, w_10000_7097, w_10000_7098, w_10000_7099, w_10000_7100, w_10000_7101, w_10000_7102, w_10000_7103, w_10000_7104, w_10000_7105, w_10000_7106, w_10000_7107, w_10000_7108, w_10000_7109, w_10000_7110, w_10000_7111, w_10000_7112, w_10000_7113, w_10000_7114, w_10000_7115, w_10000_7116, w_10000_7117, w_10000_7118, w_10000_7119, w_10000_7120, w_10000_7121, w_10000_7122, w_10000_7123, w_10000_7124, w_10000_7125, w_10000_7126, w_10000_7127, w_10000_7128, w_10000_7129, w_10000_7130, w_10000_7131, w_10000_7132, w_10000_7133, w_10000_7134, w_10000_7135, w_10000_7136, w_10000_7137, w_10000_7138, w_10000_7139, w_10000_7140, w_10000_7141, w_10000_7142, w_10000_7143, w_10000_7144, w_10000_7145, w_10000_7146, w_10000_7147, w_10000_7148, w_10000_7149, w_10000_7150, w_10000_7151, w_10000_7152, w_10000_7153, w_10000_7154, w_10000_7155, w_10000_7156, w_10000_7157, w_10000_7158, w_10000_7159, w_10000_7160, w_10000_7161, w_10000_7162, w_10000_7163, w_10000_7164, w_10000_7165, w_10000_7166, w_10000_7167, w_10000_7168, w_10000_7169, w_10000_7170, w_10000_7171, w_10000_7172, w_10000_7173, w_10000_7174, w_10000_7175, w_10000_7176, w_10000_7177, w_10000_7178, w_10000_7179, w_10000_7180, w_10000_7181, w_10000_7182, w_10000_7183, w_10000_7184, w_10000_7185, w_10000_7186, w_10000_7187, w_10000_7188, w_10000_7189, w_10000_7190, w_10000_7191, w_10000_7192, w_10000_7193, w_10000_7194, w_10000_7195, w_10000_7196, w_10000_7197, w_10000_7198, w_10000_7199, w_10000_7200, w_10000_7201, w_10000_7202, w_10000_7203, w_10000_7204, w_10000_7205, w_10000_7206, w_10000_7207, w_10000_7208, w_10000_7209, w_10000_7210, w_10000_7211, w_10000_7212, w_10000_7213, w_10000_7214, w_10000_7215, w_10000_7216, w_10000_7217, w_10000_7218, w_10000_7219, w_10000_7220, w_10000_7221, w_10000_7222, w_10000_7223, w_10000_7224, w_10000_7225, w_10000_7226, w_10000_7227, w_10000_7228, w_10000_7229, w_10000_7230, w_10000_7231, w_10000_7232, w_10000_7233, w_10000_7234, w_10000_7235, w_10000_7236, w_10000_7237, w_10000_7238, w_10000_7239, w_10000_7240, w_10000_7241, w_10000_7242, w_10000_7243, w_10000_7244, w_10000_7245, w_10000_7246, w_10000_7247, w_10000_7248, w_10000_7249, w_10000_7250, w_10000_7251, w_10000_7252, w_10000_7253, w_10000_7254, w_10000_7255, w_10000_7256, w_10000_7257, w_10000_7258, w_10000_7259, w_10000_7260, w_10000_7261, w_10000_7262, w_10000_7263, w_10000_7264, w_10000_7265, w_10000_7266, w_10000_7267, w_10000_7268, w_10000_7269, w_10000_7270, w_10000_7271, w_10000_7272, w_10000_7273, w_10000_7274, w_10000_7275, w_10000_7276, w_10000_7277, w_10000_7278, w_10000_7279, w_10000_7280, w_10000_7281, w_10000_7282, w_10000_7283, w_10000_7284, w_10000_7285, w_10000_7286, w_10000_7287, w_10000_7288;
  wire w_000_000, w_000_001, w_000_002, w_000_003, w_000_004, w_000_005, w_000_006, w_000_007, w_000_008, w_000_009, w_000_010, w_000_011, w_000_012, w_000_013, w_000_014, w_000_015, w_000_016, w_000_017, w_000_018, w_000_019, w_000_020, w_000_021, w_000_022, w_000_023, w_000_024, w_000_025, w_000_026, w_000_027, w_000_028, w_000_029, w_000_030, w_000_031, w_000_032, w_000_033, w_000_034, w_000_035, w_000_036, w_000_037, w_000_038, w_000_039, w_000_040, w_000_041, w_000_042, w_000_043, w_000_044, w_000_045, w_000_046, w_000_047, w_000_048, w_000_049, w_000_050, w_000_051, w_000_052, w_000_053, w_000_054, w_000_055, w_000_056, w_000_057, w_000_058, w_000_059, w_000_060, w_000_061, w_000_062, w_000_063, w_000_064, w_000_065, w_000_066, w_000_067, w_000_068, w_000_069, w_000_070, w_000_071, w_000_072, w_000_073, w_000_074, w_000_075, w_000_076, w_000_077, w_000_078, w_000_079, w_000_080, w_000_081, w_000_082, w_000_083, w_000_084, w_000_085, w_000_086, w_000_087, w_000_088, w_000_089, w_000_090, w_000_091, w_000_092, w_000_093, w_000_094, w_000_095, w_000_096, w_000_097, w_000_098, w_000_099, w_000_100, w_000_101, w_000_102, w_000_103, w_000_104, w_000_105, w_000_106, w_000_107, w_000_108, w_000_109, w_000_110, w_000_111, w_000_112, w_000_113, w_000_114, w_000_115, w_000_116, w_000_117, w_000_118, w_000_119, w_000_120, w_000_121, w_000_122, w_000_123, w_000_124, w_000_125, w_000_126, w_000_127, w_000_128, w_000_129, w_000_130, w_000_131, w_000_132, w_000_133, w_000_134, w_000_135, w_000_136, w_000_137, w_000_138, w_000_139, w_000_140, w_000_141, w_000_142, w_000_143, w_000_144, w_000_145, w_000_146, w_000_147, w_000_148, w_000_149, w_000_150, w_000_151, w_000_152, w_000_153, w_000_154, w_000_155, w_000_156, w_000_157, w_000_158, w_000_159, w_000_160, w_000_161, w_000_162, w_000_163, w_000_164, w_000_165, w_000_166, w_000_167, w_000_168, w_000_169, w_000_170, w_000_171, w_000_172, w_000_173, w_000_174, w_000_175, w_000_176, w_000_177, w_000_178, w_000_179, w_000_180, w_000_181, w_000_182, w_000_183, w_000_184, w_000_185, w_000_186, w_000_187, w_000_188, w_000_189, w_000_190, w_000_191, w_000_192, w_000_193, w_000_194, w_000_195, w_000_196, w_000_197, w_000_198, w_000_199, w_000_200, w_000_201, w_000_202, w_000_203, w_000_204, w_000_205, w_000_206, w_000_207, w_000_208, w_000_209, w_000_210, w_000_211, w_000_212, w_000_213, w_000_214, w_000_215, w_000_216, w_000_217, w_000_218, w_000_219, w_000_220, w_000_221, w_000_222, w_000_223, w_000_224, w_000_225, w_000_226, w_000_227, w_000_228, w_000_229, w_000_230, w_000_231, w_000_232, w_000_233, w_000_234, w_000_235, w_000_236, w_000_237, w_000_238, w_000_239, w_000_240, w_000_241, w_000_242, w_000_243, w_000_244, w_000_245, w_000_246, w_000_247, w_000_248, w_000_249, w_000_250, w_000_251, w_000_252, w_000_253, w_000_254, w_000_255, w_000_256, w_000_257, w_000_258, w_000_259, w_000_260, w_000_261, w_000_262, w_000_263, w_000_264, w_000_265, w_000_266, w_000_267, w_000_268, w_000_269, w_000_270, w_000_271, w_000_272, w_000_273, w_000_274, w_000_275, w_000_276, w_000_277, w_000_278, w_000_279, w_000_280, w_000_281, w_000_282, w_000_283, w_000_284, w_000_285, w_000_286, w_000_287, w_000_288, w_000_289, w_000_290, w_000_291, w_000_292, w_000_293, w_000_294, w_000_295, w_000_296, w_000_297, w_000_298, w_000_299, w_000_300, w_000_301, w_000_302, w_000_303, w_000_304, w_000_305, w_000_306, w_000_307, w_000_308, w_000_309, w_000_310, w_000_311, w_000_312, w_000_313, w_000_314, w_000_315, w_000_316, w_000_317, w_000_318, w_000_319, w_000_320, w_000_321, w_000_322, w_000_323, w_000_324, w_000_325, w_000_326, w_000_327, w_000_328, w_000_329, w_000_330, w_000_331, w_000_332, w_000_333, w_000_334, w_000_335, w_000_336, w_000_337, w_000_338, w_000_339, w_000_340, w_000_341, w_000_342, w_000_343, w_000_344, w_000_345, w_000_346, w_000_347, w_000_348, w_000_349, w_000_350, w_000_351, w_000_352, w_000_353, w_000_354, w_000_355, w_000_356, w_000_357, w_000_358, w_000_359, w_000_360, w_000_361, w_000_362, w_000_363, w_000_364, w_000_365, w_000_366, w_000_367, w_000_368, w_000_369, w_000_370, w_000_371, w_000_372, w_000_373, w_000_374, w_000_375, w_000_376, w_000_377, w_000_378, w_000_379, w_000_380, w_000_381, w_000_382, w_000_383, w_000_384, w_000_385, w_000_386, w_000_387, w_000_388, w_000_389, w_000_390, w_000_391, w_000_392, w_000_393, w_000_394, w_000_395, w_000_396, w_000_397, w_000_398, w_000_399, w_000_400, w_000_401, w_000_402, w_000_403, w_000_404, w_000_405, w_000_406, w_000_407, w_000_408, w_000_409, w_000_410, w_000_411, w_000_412, w_000_413, w_000_414, w_000_415, w_000_416, w_000_417, w_000_418, w_000_419, w_000_420, w_000_421, w_000_422, w_000_423, w_000_424, w_000_425, w_000_426, w_000_427, w_000_428, w_000_429, w_000_430, w_000_431, w_000_432, w_000_433, w_000_434, w_000_435, w_000_436, w_000_437, w_000_438, w_000_439, w_000_440, w_000_441, w_000_442, w_000_443, w_000_444, w_000_445, w_000_446, w_000_447, w_000_448, w_000_449, w_000_450, w_000_451, w_000_452, w_000_453, w_000_454, w_000_455, w_000_456, w_000_457, w_000_458, w_000_459, w_000_460, w_000_461, w_000_462, w_000_463, w_000_464, w_000_465, w_000_466, w_000_467, w_000_468, w_000_469, w_000_470, w_000_471, w_000_472, w_000_473, w_000_474, w_000_475, w_000_476, w_000_477, w_000_478, w_000_479, w_000_480, w_000_481, w_000_482, w_000_483, w_000_484, w_000_485, w_000_486, w_000_487, w_000_488, w_000_489, w_000_490, w_000_491, w_000_492, w_000_493, w_000_494, w_000_495, w_000_496, w_000_497, w_000_498, w_000_499, w_000_500, w_000_501, w_000_502, w_000_503, w_000_504, w_000_505, w_000_506, w_000_507, w_000_508, w_000_509, w_000_510, w_000_511, w_000_512, w_000_513, w_000_514, w_000_515, w_000_516, w_000_517, w_000_518, w_000_519, w_000_520, w_000_521, w_000_522, w_000_523, w_000_524, w_000_525, w_000_526, w_000_527, w_000_528, w_000_529, w_000_530, w_000_531, w_000_532, w_000_533, w_000_534, w_000_535, w_000_536, w_000_537, w_000_538, w_000_539, w_000_540, w_000_541, w_000_542, w_000_543, w_000_544, w_000_545, w_000_546, w_000_547, w_000_548, w_000_549, w_000_550, w_000_551, w_000_552, w_000_553, w_000_554, w_000_555, w_000_556, w_000_557, w_000_558, w_000_559, w_000_560, w_000_561, w_000_562, w_000_563, w_000_564, w_000_565, w_000_566, w_000_567, w_000_568, w_000_569, w_000_570, w_000_571, w_000_572, w_000_573, w_000_574, w_000_575, w_000_576, w_000_577, w_000_578, w_000_579, w_000_580, w_000_581, w_000_582, w_000_583, w_000_584, w_000_585, w_000_586, w_000_587, w_000_588, w_000_589, w_000_590, w_000_591, w_000_592, w_000_593, w_000_594, w_000_595, w_000_596, w_000_597, w_000_598, w_000_599, w_000_600, w_000_601, w_000_602, w_000_603, w_000_604, w_000_605, w_000_606, w_000_607, w_000_608, w_000_609, w_000_610, w_000_611, w_000_612, w_000_613, w_000_614, w_000_615, w_000_616, w_000_617, w_000_618, w_000_619, w_000_620, w_000_621, w_000_622, w_000_623, w_000_624, w_000_625, w_000_626, w_000_627, w_000_628, w_000_629, w_000_630, w_000_631, w_000_632, w_000_633, w_000_634, w_000_635, w_000_636, w_000_637, w_000_638, w_000_639, w_000_640, w_000_641, w_000_642, w_000_643, w_000_644, w_000_645, w_000_646, w_000_647, w_000_648, w_000_649, w_000_650, w_000_651, w_000_652, w_000_653, w_000_654, w_000_655, w_000_656, w_000_657, w_000_658, w_000_659, w_000_660, w_000_661, w_000_662, w_000_663, w_000_664, w_000_665, w_000_666, w_000_667, w_000_668, w_000_669, w_000_670, w_000_671, w_000_672, w_000_673, w_000_674, w_000_675, w_000_676, w_000_677, w_000_678, w_000_679, w_000_680, w_000_681, w_000_682, w_000_683, w_000_684, w_000_685, w_000_686, w_000_687, w_000_688, w_000_689, w_000_690, w_000_691, w_000_692, w_000_693, w_000_694, w_000_695, w_000_696, w_000_697, w_000_698, w_000_699, w_000_700, w_000_701, w_000_702, w_000_703, w_000_704, w_000_705, w_000_706, w_000_707, w_000_708, w_000_709, w_000_710, w_000_711, w_000_712, w_000_713, w_000_714, w_000_715, w_000_716, w_000_717, w_000_718, w_000_719, w_000_720, w_000_721, w_000_722, w_000_723, w_000_724, w_000_725, w_000_726, w_000_727, w_000_728, w_000_729, w_000_730, w_000_731, w_000_732, w_000_733, w_000_734, w_000_735, w_000_736, w_000_737, w_000_738, w_000_739, w_000_740, w_000_741, w_000_742, w_000_743, w_000_744, w_000_745, w_000_746, w_000_747, w_000_748, w_000_749, w_000_750, w_000_751, w_000_752, w_000_753, w_000_754, w_000_755, w_000_756, w_000_757, w_000_758, w_000_759, w_000_760, w_000_761, w_000_762, w_000_763, w_000_764, w_000_765, w_000_766, w_000_767, w_000_768, w_000_769, w_000_770, w_000_771, w_000_772, w_000_773, w_000_774, w_000_775, w_000_776, w_000_777, w_000_778, w_000_779, w_000_780, w_000_781, w_000_782, w_000_783, w_000_784, w_000_785, w_000_786, w_000_787, w_000_788, w_000_789, w_000_790, w_000_791, w_000_792, w_000_793, w_000_794, w_000_795, w_000_796, w_000_797, w_000_798, w_000_799, w_000_800, w_000_801, w_000_802, w_000_803, w_000_804, w_000_805, w_000_806, w_000_807, w_000_808, w_000_809, w_000_810, w_000_811, w_000_812, w_000_813, w_000_814, w_000_815, w_000_816, w_000_817, w_000_818, w_000_819, w_000_820, w_000_821, w_000_822, w_000_823, w_000_824, w_000_825, w_000_826, w_000_827, w_000_828, w_000_829, w_000_830, w_000_831, w_000_832, w_000_833, w_000_834, w_000_835, w_000_836, w_000_837, w_000_838, w_000_839, w_000_840, w_000_841, w_000_842, w_000_843, w_000_844, w_000_845, w_000_846, w_000_847, w_000_848, w_000_849, w_000_850, w_000_851, w_000_852, w_000_853, w_000_854, w_000_855, w_000_856, w_000_857, w_000_858, w_000_859, w_000_860, w_000_861, w_000_862, w_000_863, w_000_864, w_000_865, w_000_866, w_000_867, w_000_868, w_000_869, w_000_870, w_000_871, w_000_872, w_000_873, w_000_874, w_000_875, w_000_876, w_000_877, w_000_878, w_000_879, w_000_880, w_000_881, w_000_882, w_000_883, w_000_884, w_000_885, w_000_886, w_000_887, w_000_888, w_000_889, w_000_890, w_000_891, w_000_892, w_000_893, w_000_894, w_000_895, w_000_896, w_000_897, w_000_898, w_000_899, w_000_900, w_000_901, w_000_902, w_000_903, w_000_904, w_000_905, w_000_906, w_000_907, w_000_908, w_000_909, w_000_910, w_000_911, w_000_912, w_000_913, w_000_914, w_000_915, w_000_916, w_000_917, w_000_918, w_000_919, w_000_920, w_000_921, w_000_922, w_000_923, w_000_924, w_000_925, w_000_926, w_000_927, w_000_928, w_000_929, w_000_930, w_000_931, w_000_932, w_000_933, w_000_934, w_000_935, w_000_936, w_000_937, w_000_938, w_000_939, w_000_940, w_000_941, w_000_942, w_000_943, w_000_944, w_000_945, w_000_946, w_000_947, w_000_948, w_000_949, w_000_950, w_000_951, w_000_952, w_000_953, w_000_954, w_000_955, w_000_956, w_000_957, w_000_958, w_000_959, w_000_960, w_000_961, w_000_962, w_000_963, w_000_964, w_000_965, w_000_966, w_000_967, w_000_968, w_000_969, w_000_970, w_000_971, w_000_972, w_000_973, w_000_974, w_000_975, w_000_976, w_000_977, w_000_978, w_000_979, w_000_980, w_000_981, w_000_982, w_000_983, w_000_984, w_000_985, w_000_986, w_000_987, w_000_988, w_000_989, w_000_990, w_000_991, w_000_992, w_000_993, w_000_994, w_000_995, w_000_996, w_000_997, w_000_998, w_000_999, w_000_1000, w_000_1001, w_000_1002, w_000_1003, w_000_1004, w_000_1005, w_000_1006, w_000_1007, w_000_1008, w_000_1009, w_000_1010, w_000_1011, w_000_1012, w_000_1013, w_000_1014, w_000_1015, w_000_1016, w_000_1017, w_000_1018, w_000_1019, w_000_1020, w_000_1021, w_000_1022, w_000_1023, w_000_1024, w_000_1025, w_000_1026, w_000_1027, w_000_1028, w_000_1029, w_000_1030, w_000_1031, w_000_1032, w_000_1033, w_000_1034, w_000_1035, w_000_1036, w_000_1037, w_000_1038, w_000_1039, w_000_1040, w_000_1041, w_000_1042, w_000_1043, w_000_1044, w_000_1045, w_000_1046, w_000_1047, w_000_1048, w_000_1049, w_000_1050, w_000_1051, w_000_1052, w_000_1053, w_000_1054, w_000_1055, w_000_1056, w_000_1057, w_000_1058, w_000_1059, w_000_1060, w_000_1061, w_000_1062, w_000_1063, w_000_1064, w_000_1065, w_000_1066, w_000_1067, w_000_1068, w_000_1069, w_000_1070, w_000_1071, w_000_1072, w_000_1073, w_000_1074, w_000_1075, w_000_1076, w_000_1077, w_000_1078, w_000_1079, w_000_1080, w_000_1081, w_000_1082, w_000_1083, w_000_1084, w_000_1085, w_000_1086, w_000_1087, w_000_1088, w_000_1089, w_000_1090, w_000_1091, w_000_1092, w_000_1093, w_000_1094, w_000_1095, w_000_1096, w_000_1097, w_000_1098, w_000_1099, w_000_1100, w_000_1101, w_000_1102, w_000_1103, w_000_1104, w_000_1105, w_000_1106, w_000_1107, w_000_1108, w_000_1109, w_000_1110, w_000_1111, w_000_1112, w_000_1113, w_000_1114, w_000_1115, w_000_1116, w_000_1117, w_000_1118, w_000_1119, w_000_1120, w_000_1121, w_000_1122, w_000_1123, w_000_1124, w_000_1125, w_000_1126, w_000_1127, w_000_1128, w_000_1129, w_000_1130, w_000_1131, w_000_1132, w_000_1133, w_000_1134, w_000_1135, w_000_1136, w_000_1137, w_000_1138, w_000_1139, w_000_1140, w_000_1141, w_000_1142, w_000_1143, w_000_1144, w_000_1145, w_000_1146, w_000_1147, w_000_1148, w_000_1149, w_000_1150, w_000_1151, w_000_1152, w_000_1153, w_000_1154, w_000_1155, w_000_1156, w_000_1157, w_000_1158, w_000_1159, w_000_1160, w_000_1161, w_000_1162, w_000_1163, w_000_1164, w_000_1165, w_000_1166, w_000_1167, w_000_1168, w_000_1169, w_000_1170, w_000_1171, w_000_1172, w_000_1173, w_000_1174, w_000_1175, w_000_1176, w_000_1177, w_000_1178, w_000_1179, w_000_1180, w_000_1181, w_000_1182, w_000_1183, w_000_1184, w_000_1185, w_000_1186, w_000_1187, w_000_1188, w_000_1189, w_000_1190, w_000_1191, w_000_1192, w_000_1193, w_000_1194, w_000_1195, w_000_1196, w_000_1197, w_000_1198, w_000_1199, w_000_1200, w_000_1201, w_000_1202, w_000_1203, w_000_1204, w_000_1205, w_000_1206, w_000_1207, w_000_1208, w_000_1209, w_000_1210, w_000_1211, w_000_1212, w_000_1213, w_000_1214, w_000_1215, w_000_1216, w_000_1217, w_000_1218, w_000_1219, w_000_1220, w_000_1221, w_000_1222, w_000_1223, w_000_1224, w_000_1225, w_000_1226, w_000_1227, w_000_1228, w_000_1229, w_000_1230, w_000_1231, w_000_1232, w_000_1233, w_000_1234, w_000_1235, w_000_1236, w_000_1237, w_000_1238, w_000_1239, w_000_1240, w_000_1241, w_000_1242, w_000_1243, w_000_1244, w_000_1245, w_000_1246, w_000_1247, w_000_1248, w_000_1249, w_000_1250, w_000_1251, w_000_1252, w_000_1253, w_000_1254, w_000_1255, w_000_1256, w_000_1257, w_000_1258, w_000_1259, w_000_1260, w_000_1261, w_000_1262, w_000_1263, w_000_1264, w_000_1265, w_000_1266, w_000_1267, w_000_1268, w_000_1269, w_000_1270, w_000_1271, w_000_1272, w_000_1273, w_000_1274, w_000_1275, w_000_1276, w_000_1277, w_000_1278, w_000_1279, w_000_1280, w_000_1281, w_000_1282, w_000_1283, w_000_1284, w_000_1285, w_000_1286, w_000_1287, w_000_1288, w_000_1289, w_000_1290, w_000_1291, w_000_1292, w_000_1293, w_000_1294, w_000_1295, w_000_1296, w_000_1297, w_000_1298, w_000_1299, w_000_1300, w_000_1301, w_000_1302, w_000_1303, w_000_1304, w_000_1305, w_000_1306, w_000_1307, w_000_1308, w_000_1309, w_000_1310, w_000_1311, w_000_1312, w_000_1313, w_000_1314, w_000_1315, w_000_1316, w_000_1317, w_000_1318, w_000_1319, w_000_1320, w_000_1321, w_000_1322, w_000_1323, w_000_1324, w_000_1325, w_000_1326, w_000_1327, w_000_1328, w_000_1329, w_000_1330, w_000_1331, w_000_1332, w_000_1333, w_000_1334, w_000_1335, w_000_1336, w_000_1337, w_000_1338, w_000_1339, w_000_1340, w_000_1341, w_000_1342, w_000_1343, w_000_1344, w_000_1345, w_000_1346, w_000_1347, w_000_1348, w_000_1349, w_000_1350, w_000_1351, w_000_1352, w_000_1353, w_000_1354, w_000_1355, w_000_1356, w_000_1357, w_000_1358, w_000_1359, w_000_1360, w_000_1361, w_000_1362, w_000_1363, w_000_1364, w_000_1365, w_000_1366, w_000_1367, w_000_1368, w_000_1369, w_000_1370, w_000_1371, w_000_1372, w_000_1373, w_000_1374, w_000_1375, w_000_1376, w_000_1377, w_000_1378, w_000_1379, w_000_1380, w_000_1381, w_000_1382, w_000_1383, w_000_1384, w_000_1385, w_000_1386, w_000_1387, w_000_1388, w_000_1389, w_000_1390, w_000_1391, w_000_1392, w_000_1393, w_000_1394, w_000_1395, w_000_1396, w_000_1397, w_000_1398, w_000_1399, w_000_1400, w_000_1401, w_000_1402, w_000_1403, w_000_1404, w_000_1405, w_000_1406, w_000_1407, w_000_1408, w_000_1409, w_000_1410, w_000_1411, w_000_1412, w_000_1413, w_000_1414, w_000_1415, w_000_1416, w_000_1417, w_000_1418, w_000_1419, w_000_1420, w_000_1421, w_000_1422, w_000_1423, w_000_1424, w_000_1425, w_000_1426, w_000_1427, w_000_1428, w_000_1429, w_000_1430, w_000_1431, w_000_1432, w_000_1433, w_000_1434, w_000_1435, w_000_1436, w_000_1437, w_000_1438, w_000_1439, w_000_1440, w_000_1441, w_000_1442, w_000_1443, w_000_1444, w_000_1445, w_000_1446, w_000_1447, w_000_1448, w_000_1449, w_000_1450, w_000_1451, w_000_1452, w_000_1453, w_000_1454, w_000_1455, w_000_1456, w_000_1457, w_000_1458, w_000_1459, w_000_1460, w_000_1461, w_000_1462, w_000_1463, w_000_1464, w_000_1465, w_000_1466, w_000_1467, w_000_1468, w_000_1469, w_000_1470, w_000_1471, w_000_1472, w_000_1473, w_000_1474, w_000_1475, w_000_1476, w_000_1477, w_000_1478, w_000_1479, w_000_1480, w_000_1481, w_000_1482, w_000_1483, w_000_1484, w_000_1485, w_000_1486, w_000_1487, w_000_1488, w_000_1489, w_000_1490, w_000_1491, w_000_1492, w_000_1493, w_000_1494, w_000_1495, w_000_1496, w_000_1497, w_000_1498, w_000_1499, w_000_1500, w_000_1501, w_000_1502, w_000_1503, w_000_1504, w_000_1505, w_000_1506, w_000_1507, w_000_1508, w_000_1509, w_000_1510, w_000_1511, w_000_1512, w_000_1513, w_000_1514, w_000_1515, w_000_1516, w_000_1517, w_000_1518, w_000_1519, w_000_1520, w_000_1521, w_000_1522, w_000_1523, w_000_1524, w_000_1525, w_000_1526, w_000_1527, w_000_1528, w_000_1529, w_000_1530, w_000_1531, w_000_1532, w_000_1533, w_000_1534, w_000_1535, w_000_1536, w_000_1537, w_000_1538, w_000_1539, w_000_1540, w_000_1541, w_000_1542, w_000_1543, w_000_1544, w_000_1545, w_000_1546, w_000_1547, w_000_1548, w_000_1549, w_000_1550, w_000_1551, w_000_1552, w_000_1553, w_000_1554, w_000_1555, w_000_1556, w_000_1557, w_000_1558, w_000_1559, w_000_1560, w_000_1561, w_000_1562, w_000_1563, w_000_1564, w_000_1565, w_000_1566, w_000_1567, w_000_1568, w_000_1569, w_000_1570, w_000_1571, w_000_1572, w_000_1573, w_000_1574, w_000_1575, w_000_1576, w_000_1577, w_000_1578, w_000_1579, w_000_1580, w_000_1581, w_000_1582, w_000_1583, w_000_1584, w_000_1585, w_000_1586, w_000_1587, w_000_1588, w_000_1589, w_000_1590, w_000_1591, w_000_1592, w_000_1593, w_000_1594, w_000_1595, w_000_1596, w_000_1597, w_000_1598, w_000_1599, w_000_1600, w_000_1601, w_000_1602, w_000_1603, w_000_1604, w_000_1605, w_000_1606, w_000_1607, w_000_1608, w_000_1609, w_000_1610, w_000_1611, w_000_1612, w_000_1613, w_000_1614, w_000_1615, w_000_1616, w_000_1617, w_000_1618, w_000_1619, w_000_1620, w_000_1621, w_000_1622, w_000_1623, w_000_1624, w_000_1625, w_000_1626, w_000_1627, w_000_1628, w_000_1629, w_000_1630, w_000_1631, w_000_1632, w_000_1633, w_000_1634, w_000_1635, w_000_1636, w_000_1637, w_000_1638, w_000_1639, w_000_1640, w_000_1641, w_000_1642, w_000_1643, w_000_1644, w_000_1645, w_000_1646, w_000_1647, w_000_1648, w_000_1649, w_000_1650, w_000_1651, w_000_1652, w_000_1653, w_000_1654, w_000_1655, w_000_1656, w_000_1657, w_000_1658, w_000_1659, w_000_1660, w_000_1661, w_000_1662, w_000_1663, w_000_1664, w_000_1665, w_000_1666, w_000_1667, w_000_1668, w_000_1669, w_000_1670, w_000_1671, w_000_1672, w_000_1673, w_000_1674, w_000_1675, w_000_1676, w_000_1677, w_000_1678, w_000_1679, w_000_1680, w_000_1681, w_000_1682, w_000_1683, w_000_1684, w_000_1685, w_000_1686, w_000_1687, w_000_1688, w_000_1689, w_000_1690, w_000_1691, w_000_1692, w_000_1693, w_000_1694, w_000_1695, w_000_1696, w_000_1697, w_000_1698, w_000_1699, w_000_1700, w_000_1701, w_000_1702, w_000_1703, w_000_1704, w_000_1705, w_000_1706, w_000_1707, w_000_1708, w_000_1709, w_000_1710, w_000_1711, w_000_1712, w_000_1713, w_000_1714, w_000_1715, w_000_1716, w_000_1717, w_000_1718, w_000_1719, w_000_1720, w_000_1721, w_000_1722, w_000_1723, w_000_1724, w_000_1725, w_000_1726, w_000_1727, w_000_1728, w_000_1729, w_000_1730, w_000_1731, w_000_1732, w_000_1733, w_000_1734, w_000_1735, w_000_1736, w_000_1737, w_000_1738, w_000_1739, w_000_1740, w_000_1741, w_000_1742, w_000_1743, w_000_1744, w_000_1745, w_000_1746, w_000_1747, w_000_1748, w_000_1749, w_000_1750, w_000_1751, w_000_1752, w_000_1753, w_000_1754, w_000_1755, w_000_1756, w_000_1757, w_000_1758, w_000_1759, w_000_1760, w_000_1761, w_000_1762, w_000_1763, w_000_1764, w_000_1765, w_000_1766, w_000_1767, w_000_1768, w_000_1769, w_000_1770, w_000_1771, w_000_1772, w_000_1773, w_000_1774, w_000_1775, w_000_1776, w_000_1777, w_000_1778, w_000_1779, w_000_1780, w_000_1781, w_000_1782, w_000_1783, w_000_1784, w_000_1785, w_000_1786, w_000_1787, w_000_1788, w_000_1789, w_000_1790, w_000_1791, w_000_1792, w_000_1793, w_000_1794, w_000_1795, w_000_1796, w_000_1797, w_000_1798, w_000_1799, w_000_1800, w_000_1801, w_000_1802, w_000_1803, w_000_1804, w_000_1805, w_000_1806, w_000_1807, w_000_1808, w_000_1809, w_000_1810, w_000_1811, w_000_1812, w_000_1813, w_000_1814, w_000_1815, w_000_1816, w_000_1817, w_000_1818, w_000_1819, w_000_1820, w_000_1821, w_000_1822, w_000_1823, w_000_1824, w_000_1825, w_000_1826, w_000_1827, w_000_1828, w_000_1829, w_000_1830, w_000_1831, w_000_1832, w_000_1833, w_000_1834, w_000_1835, w_000_1836, w_000_1837, w_000_1838, w_000_1839, w_000_1840, w_000_1841, w_000_1842, w_000_1843, w_000_1844, w_000_1845, w_000_1846, w_000_1847, w_000_1848, w_000_1849, w_000_1850, w_000_1851, w_000_1852, w_000_1853, w_000_1854, w_000_1855, w_000_1856, w_000_1857, w_000_1858, w_000_1859, w_000_1860, w_000_1861, w_000_1862, w_000_1863, w_000_1864, w_000_1865, w_000_1866, w_000_1867, w_000_1868, w_000_1869, w_000_1870, w_000_1871, w_000_1872, w_000_1873, w_000_1874, w_000_1875, w_000_1876, w_000_1877, w_000_1878, w_000_1879, w_000_1880, w_000_1881, w_000_1882, w_000_1883, w_000_1884, w_000_1885, w_000_1886, w_000_1887, w_000_1888, w_000_1889, w_000_1890, w_000_1891, w_000_1892, w_000_1893, w_000_1894, w_000_1895, w_000_1896, w_000_1897, w_000_1898, w_000_1899, w_000_1900, w_000_1901, w_000_1902, w_000_1903, w_000_1904, w_000_1905, w_000_1906, w_000_1907, w_000_1908, w_000_1909, w_000_1910, w_000_1911, w_000_1912, w_000_1913, w_000_1914, w_000_1915, w_000_1916, w_000_1917, w_000_1918, w_000_1919, w_000_1920, w_000_1921, w_000_1922, w_000_1923, w_000_1924, w_000_1925, w_000_1926, w_000_1927, w_000_1928, w_000_1929, w_000_1930, w_000_1931, w_000_1932, w_000_1933, w_000_1934, w_000_1935, w_000_1936, w_000_1937, w_000_1938, w_000_1939, w_000_1940, w_000_1941, w_000_1942, w_000_1943, w_000_1944, w_000_1945, w_000_1946, w_000_1947, w_000_1948, w_000_1949, w_000_1950, w_000_1951, w_000_1952, w_000_1953, w_000_1954, w_000_1955, w_000_1956, w_000_1957, w_000_1958, w_000_1959, w_000_1960, w_000_1961, w_000_1962, w_000_1963, w_000_1964, w_000_1965, w_000_1966, w_000_1967, w_000_1968, w_000_1969, w_000_1970, w_000_1971, w_000_1972, w_000_1973, w_000_1974, w_000_1975, w_000_1976, w_000_1977, w_000_1978, w_000_1979, w_000_1980, w_000_1981, w_000_1982, w_000_1983, w_000_1984, w_000_1985, w_000_1986, w_000_1987, w_000_1988, w_000_1989, w_000_1990, w_000_1991, w_000_1992, w_000_1993, w_000_1994, w_000_1995, w_000_1996, w_000_1997, w_000_1998, w_000_1999, w_000_2000, w_000_2001, w_000_2002, w_000_2003, w_000_2004, w_000_2005, w_000_2006, w_000_2007, w_000_2008, w_000_2009, w_000_2010, w_000_2011, w_000_2012, w_000_2013, w_000_2014, w_000_2015, w_000_2016, w_000_2017, w_000_2018, w_000_2019, w_000_2020, w_000_2021, w_000_2022, w_000_2023, w_000_2024, w_000_2025, w_000_2026, w_000_2027, w_000_2028, w_000_2029, w_000_2030, w_000_2031, w_000_2032, w_000_2033, w_000_2034, w_000_2035, w_000_2036, w_000_2037, w_000_2038, w_000_2039, w_000_2040, w_000_2041, w_000_2042, w_000_2043, w_000_2044, w_000_2045, w_000_2046, w_000_2047, w_000_2048, w_000_2049, w_000_2050, w_000_2051, w_000_2052, w_000_2053, w_000_2054, w_000_2055, w_000_2056, w_000_2057, w_000_2058, w_000_2059, w_000_2060, w_000_2061, w_000_2062, w_000_2063, w_000_2064, w_000_2065, w_000_2066, w_000_2067, w_000_2068, w_000_2069, w_000_2070, w_000_2071, w_000_2072, w_000_2073, w_000_2074, w_000_2075, w_000_2076, w_000_2077, w_000_2078, w_000_2079, w_000_2080, w_000_2081, w_000_2082, w_000_2083, w_000_2084, w_000_2085, w_000_2086, w_000_2087, w_000_2088, w_000_2089, w_000_2090, w_000_2091, w_000_2092, w_000_2093, w_000_2094, w_000_2095, w_000_2096, w_000_2097, w_000_2098, w_000_2099, w_000_2100, w_000_2101, w_000_2102, w_000_2103, w_000_2104, w_000_2105, w_000_2106, w_000_2107, w_000_2108, w_000_2109, w_000_2110, w_000_2111, w_000_2112, w_000_2113, w_000_2114, w_000_2115, w_000_2116, w_000_2117, w_000_2118, w_000_2119, w_000_2120, w_000_2121, w_000_2122, w_000_2123, w_000_2124, w_000_2125, w_000_2126, w_000_2127, w_000_2128, w_000_2129, w_000_2130, w_000_2131, w_000_2132, w_000_2133, w_000_2134, w_000_2135, w_000_2136, w_000_2137, w_000_2138, w_000_2139, w_000_2140, w_000_2141, w_000_2142, w_000_2143, w_000_2144, w_000_2145, w_000_2146, w_000_2147, w_000_2148, w_000_2149, w_000_2150, w_000_2151, w_000_2152, w_000_2153, w_000_2154, w_000_2155, w_000_2156, w_000_2157, w_000_2158, w_000_2160, w_000_2161, w_000_2162, w_000_2163, w_000_2164, w_000_2165, w_000_2166, w_000_2167, w_000_2168, w_000_2169, w_000_2170, w_000_2171, w_000_2172, w_000_2173, w_000_2174, w_000_2175, w_000_2176, w_000_2177, w_000_2178, w_000_2179, w_000_2180, w_000_2181, w_000_2182, w_000_2183, w_000_2184, w_000_2185, w_000_2186, w_000_2187, w_000_2188, w_000_2189, w_000_2190, w_000_2191, w_000_2192, w_000_2193, w_000_2194, w_000_2195, w_000_2196, w_000_2197, w_000_2198, w_000_2199, w_000_2200, w_000_2201, w_000_2202, w_000_2203, w_000_2204, w_000_2205, w_000_2206, w_000_2207, w_000_2208, w_000_2209, w_000_2210, w_000_2211, w_000_2212, w_000_2213, w_000_2214, w_000_2215, w_000_2216, w_000_2217, w_000_2218, w_000_2219, w_000_2220, w_000_2221, w_000_2222, w_000_2223, w_000_2224, w_000_2225, w_000_2226, w_000_2227, w_000_2228, w_000_2229, w_000_2230, w_000_2231, w_000_2232, w_000_2233, w_000_2234, w_000_2235, w_000_2236, w_000_2237, w_000_2238, w_000_2239, w_000_2240, w_000_2241, w_000_2242, w_000_2243, w_000_2244, w_000_2245, w_000_2246, w_000_2247, w_000_2248, w_000_2249, w_000_2250, w_000_2251, w_000_2252, w_000_2253, w_000_2254, w_000_2255, w_000_2256, w_000_2257, w_000_2258, w_000_2259, w_000_2260, w_000_2261, w_000_2262, w_000_2263, w_000_2264, w_000_2265, w_000_2266, w_000_2267, w_000_2268, w_000_2269, w_000_2270, w_000_2271, w_000_2272, w_000_2273, w_000_2274, w_000_2275, w_000_2276, w_000_2277, w_000_2278, w_000_2279, w_000_2280, w_000_2281, w_000_2282, w_000_2283, w_000_2284, w_000_2285, w_000_2286, w_000_2287, w_000_2288, w_000_2289, w_000_2290, w_000_2291, w_000_2292, w_000_2293, w_000_2294, w_000_2295, w_000_2296, w_000_2297, w_000_2298, w_000_2299, w_000_2300, w_000_2301, w_000_2302, w_000_2303, w_000_2304, w_000_2305, w_000_2306, w_000_2307, w_000_2308, w_000_2309, w_000_2310, w_000_2311, w_000_2312, w_000_2313, w_000_2314, w_000_2315, w_000_2316, w_000_2317, w_000_2318, w_000_2319, w_000_2320, w_000_2321, w_000_2322, w_000_2323, w_000_2324, w_000_2325, w_000_2326, w_000_2327, w_000_2328, w_000_2329, w_000_2330, w_000_2331, w_000_2332, w_000_2333, w_000_2334, w_000_2335, w_000_2336, w_000_2337, w_000_2338, w_000_2339, w_000_2340, w_000_2341, w_000_2342, w_000_2343, w_000_2344, w_000_2345, w_000_2346, w_000_2347, w_000_2348, w_000_2349, w_000_2350, w_000_2351, w_000_2352, w_000_2353, w_000_2354, w_000_2355, w_000_2356, w_000_2357, w_000_2358, w_000_2359, w_000_2360, w_000_2361, w_000_2362, w_000_2363, w_000_2364, w_000_2365, w_000_2366, w_000_2367, w_000_2368, w_000_2369, w_000_2370, w_000_2371, w_000_2372, w_000_2373, w_000_2374, w_000_2375, w_000_2376, w_000_2377, w_000_2378, w_000_2379, w_000_2380, w_000_2381, w_000_2382, w_000_2383, w_000_2384, w_000_2385, w_000_2386, w_000_2387, w_000_2388, w_000_2389, w_000_2390, w_000_2391, w_000_2392, w_000_2393, w_000_2394, w_000_2395, w_000_2396, w_000_2397, w_000_2398, w_000_2399, w_000_2400, w_000_2401, w_000_2402, w_000_2403, w_000_2404, w_000_2405, w_000_2406, w_000_2407, w_000_2408, w_000_2410, w_000_2411, w_000_2412, w_000_2413, w_000_2414, w_000_2415, w_000_2416, w_000_2417, w_000_2418, w_000_2419, w_000_2420, w_000_2421, w_000_2422, w_000_2423, w_000_2424, w_000_2425, w_000_2426, w_000_2427, w_000_2428, w_000_2429, w_000_2430, w_000_2431, w_000_2432, w_000_2433, w_000_2434, w_000_2435, w_000_2436, w_000_2437, w_000_2438, w_000_2439, w_000_2440, w_000_2441, w_000_2442, w_000_2443, w_000_2444, w_000_2445, w_000_2446, w_000_2447, w_000_2448, w_000_2449, w_000_2450, w_000_2451, w_000_2452, w_000_2453, w_000_2454, w_000_2455, w_000_2456, w_000_2457, w_000_2458, w_000_2459, w_000_2460, w_000_2461, w_000_2462, w_000_2463, w_000_2464, w_000_2465, w_000_2466, w_000_2467, w_000_2468, w_000_2469, w_000_2470, w_000_2471, w_000_2472, w_000_2473, w_000_2474, w_000_2475, w_000_2476, w_000_2477, w_000_2478, w_000_2479, w_000_2480, w_000_2481, w_000_2482, w_000_2483, w_000_2484, w_000_2485, w_000_2486, w_000_2487, w_000_2488, w_000_2489, w_000_2490, w_000_2491, w_000_2492, w_000_2493, w_000_2494, w_000_2495, w_000_2496, w_000_2497, w_000_2498, w_000_2499, w_000_2500, w_000_2501, w_000_2502, w_000_2503, w_000_2504, w_000_2505, w_000_2506, w_000_2507, w_000_2508, w_000_2509, w_000_2510, w_000_2511, w_000_2512, w_000_2513, w_000_2514, w_000_2515, w_000_2516, w_000_2517, w_000_2518, w_000_2519, w_000_2520, w_000_2521, w_000_2522, w_000_2523, w_000_2524, w_000_2525, w_000_2526, w_000_2527, w_000_2528, w_000_2529, w_000_2530, w_000_2531, w_000_2532, w_000_2533, w_000_2534, w_000_2535, w_000_2536, w_000_2537, w_000_2538, w_000_2539, w_000_2540, w_000_2541, w_000_2542, w_000_2543, w_000_2544, w_000_2545, w_000_2546, w_000_2547, w_000_2548, w_000_2549, w_000_2550, w_000_2551, w_000_2552, w_000_2553, w_000_2554, w_000_2555, w_000_2556, w_000_2557, w_000_2558, w_000_2559, w_000_2560, w_000_2561, w_000_2562, w_000_2563, w_000_2564, w_000_2565, w_000_2566, w_000_2567, w_000_2568, w_000_2569, w_000_2570, w_000_2571, w_000_2572, w_000_2573, w_000_2574, w_000_2575, w_000_2576, w_000_2577, w_000_2578, w_000_2579, w_000_2580, w_000_2581, w_000_2582, w_000_2583, w_000_2584, w_000_2585, w_000_2586, w_000_2587, w_000_2588, w_000_2589, w_000_2590, w_000_2591, w_000_2592, w_000_2593, w_000_2594, w_000_2595, w_000_2596, w_000_2597, w_000_2598, w_000_2599, w_000_2600, w_000_2601, w_000_2602, w_000_2603, w_000_2604, w_000_2605, w_000_2606, w_000_2607, w_000_2608, w_000_2609, w_000_2610, w_000_2611, w_000_2612, w_000_2613, w_000_2614, w_000_2615, w_000_2616, w_000_2617, w_000_2618, w_000_2619, w_000_2620, w_000_2621, w_000_2622, w_000_2623, w_000_2624, w_000_2625, w_000_2626, w_000_2627, w_000_2628, w_000_2629, w_000_2630, w_000_2631, w_000_2632, w_000_2633, w_000_2634, w_000_2635, w_000_2636, w_000_2637, w_000_2638, w_000_2639, w_000_2640, w_000_2641, w_000_2642, w_000_2643, w_000_2644, w_000_2645, w_000_2646, w_000_2647, w_000_2648, w_000_2649, w_000_2650, w_000_2651, w_000_2652, w_000_2653, w_000_2654, w_000_2655, w_000_2656, w_000_2657, w_000_2658, w_000_2659, w_000_2660, w_000_2661, w_000_2662, w_000_2663, w_000_2664, w_000_2665, w_000_2666, w_000_2667, w_000_2668, w_000_2669, w_000_2670, w_000_2671, w_000_2672, w_000_2673, w_000_2674, w_000_2675, w_000_2676, w_000_2677, w_000_2678, w_000_2679, w_000_2680, w_000_2681, w_000_2682, w_000_2683, w_000_2684, w_000_2685, w_000_2686, w_000_2687, w_000_2688, w_000_2689, w_000_2690, w_000_2691, w_000_2692, w_000_2693, w_000_2694, w_000_2695, w_000_2696, w_000_2697, w_000_2698, w_000_2699, w_000_2700, w_000_2701, w_000_2702, w_000_2703, w_000_2704, w_000_2705, w_000_2706, w_000_2707, w_000_2708, w_000_2709, w_000_2710, w_000_2711, w_000_2712, w_000_2713, w_000_2714, w_000_2715, w_000_2716, w_000_2717, w_000_2718, w_000_2719, w_000_2720, w_000_2721, w_000_2722, w_000_2723, w_000_2724, w_000_2725, w_000_2726, w_000_2727, w_000_2728, w_000_2729, w_000_2730, w_000_2731, w_000_2732, w_000_2733, w_000_2734, w_000_2735, w_000_2736, w_000_2737, w_000_2738, w_000_2739, w_000_2740, w_000_2741, w_000_2742, w_000_2743, w_000_2744, w_000_2745, w_000_2746, w_000_2747, w_000_2748, w_000_2749, w_000_2750, w_000_2751, w_000_2752, w_000_2753, w_000_2754, w_000_2755, w_000_2756, w_000_2757, w_000_2758, w_000_2759, w_000_2760, w_000_2761, w_000_2762, w_000_2763, w_000_2764, w_000_2765, w_000_2766, w_000_2767, w_000_2768, w_000_2769, w_000_2770, w_000_2771, w_000_2772, w_000_2773, w_000_2774, w_000_2775, w_000_2776, w_000_2777, w_000_2778, w_000_2779, w_000_2780, w_000_2781, w_000_2782, w_000_2783, w_000_2784, w_000_2785, w_000_2786, w_000_2787, w_000_2788, w_000_2789, w_000_2790, w_000_2791, w_000_2792, w_000_2793, w_000_2794, w_000_2795, w_000_2796, w_000_2797, w_000_2798, w_000_2799, w_000_2800, w_000_2801, w_000_2802, w_000_2803, w_000_2804, w_000_2805, w_000_2806, w_000_2807, w_000_2808, w_000_2809, w_000_2810, w_000_2811, w_000_2812, w_000_2813, w_000_2814, w_000_2815, w_000_2816, w_000_2817, w_000_2818, w_000_2819, w_000_2820, w_000_2821, w_000_2822, w_000_2823, w_000_2824, w_000_2825, w_000_2826, w_000_2827, w_000_2828, w_000_2829, w_000_2830, w_000_2831, w_000_2832, w_000_2834, w_000_2835, w_000_2836, w_000_2837, w_000_2838, w_000_2839, w_000_2840, w_000_2841, w_000_2842, w_000_2843, w_000_2844, w_000_2845, w_000_2846, w_000_2847, w_000_2848, w_000_2849, w_000_2850, w_000_2851, w_000_2852, w_000_2853, w_000_2854, w_000_2855, w_000_2856, w_000_2857, w_000_2858, w_000_2859, w_000_2860, w_000_2861, w_000_2862, w_000_2863, w_000_2864, w_000_2865, w_000_2866, w_000_2867, w_000_2868, w_000_2869, w_000_2870, w_000_2871, w_000_2872, w_000_2873, w_000_2874, w_000_2875, w_000_2876, w_000_2877, w_000_2878, w_000_2879, w_000_2880, w_000_2881, w_000_2882, w_000_2883, w_000_2884, w_000_2885, w_000_2886, w_000_2887, w_000_2888, w_000_2889, w_000_2890, w_000_2891, w_000_2892, w_000_2893, w_000_2894, w_000_2895, w_000_2896, w_000_2897, w_000_2898, w_000_2899, w_000_2900, w_000_2901, w_000_2902, w_000_2903, w_000_2904, w_000_2905, w_000_2906, w_000_2907, w_000_2908, w_000_2909, w_000_2910, w_000_2911, w_000_2912, w_000_2913, w_000_2914, w_000_2915, w_000_2916, w_000_2917, w_000_2918, w_000_2919, w_000_2920, w_000_2921, w_000_2922, w_000_2923, w_000_2924, w_000_2925, w_000_2926, w_000_2927, w_000_2928, w_000_2929, w_000_2930, w_000_2931, w_000_2932, w_000_2933, w_000_2934, w_000_2935, w_000_2936, w_000_2937, w_000_2938, w_000_2939, w_000_2940, w_000_2941, w_000_2942, w_000_2943, w_000_2944, w_000_2945, w_000_2946, w_000_2947, w_000_2948, w_000_2949, w_000_2950, w_000_2951, w_000_2952, w_000_2953, w_000_2954, w_000_2955, w_000_2956, w_000_2957, w_000_2958, w_000_2959, w_000_2960, w_000_2961, w_000_2962, w_000_2963, w_000_2964, w_000_2965, w_000_2966, w_000_2967, w_000_2968, w_000_2969, w_000_2970, w_000_2971, w_000_2972, w_000_2973, w_000_2974, w_000_2975, w_000_2976, w_000_2977, w_000_2978, w_000_2979, w_000_2980, w_000_2981, w_000_2982, w_000_2983, w_000_2984, w_000_2985, w_000_2986, w_000_2987, w_000_2988, w_000_2989, w_000_2990, w_000_2991, w_000_2992, w_000_2993, w_000_2994, w_000_2995, w_000_2996, w_000_2997, w_000_2998, w_000_2999, w_000_3000, w_000_3001, w_000_3002, w_000_3003, w_000_3004, w_000_3005, w_000_3006, w_000_3007, w_000_3008, w_000_3009, w_000_3010, w_000_3011, w_000_3012, w_000_3013, w_000_3014, w_000_3015, w_000_3016, w_000_3017, w_000_3018, w_000_3019, w_000_3020, w_000_3021, w_000_3022, w_000_3023, w_000_3024, w_000_3025, w_000_3026, w_000_3027, w_000_3028, w_000_3029, w_000_3030, w_000_3031, w_000_3032, w_000_3033, w_000_3034, w_000_3035, w_000_3036, w_000_3037, w_000_3038, w_000_3039, w_000_3040, w_000_3041, w_000_3042, w_000_3043, w_000_3044, w_000_3045, w_000_3046, w_000_3047, w_000_3048, w_000_3049, w_000_3050, w_000_3051, w_000_3052, w_000_3053, w_000_3054, w_000_3055, w_000_3056, w_000_3057, w_000_3058, w_000_3059, w_000_3060, w_000_3061, w_000_3062, w_000_3063, w_000_3064, w_000_3065, w_000_3066, w_000_3067, w_000_3068, w_000_3069, w_000_3070, w_000_3071, w_000_3072, w_000_3073, w_000_3074, w_000_3075, w_000_3076, w_000_3077, w_000_3078, w_000_3079, w_000_3080, w_000_3081, w_000_3082, w_000_3083, w_000_3084, w_000_3085, w_000_3086, w_000_3087, w_000_3088, w_000_3089, w_000_3090, w_000_3091, w_000_3092, w_000_3093, w_000_3094, w_000_3095, w_000_3096, w_000_3097, w_000_3098, w_000_3099, w_000_3100, w_000_3101, w_000_3102, w_000_3103, w_000_3104, w_000_3105, w_000_3106, w_000_3107, w_000_3108, w_000_3109, w_000_3110, w_000_3111, w_000_3112, w_000_3113, w_000_3114, w_000_3115, w_000_3116, w_000_3117, w_000_3118, w_000_3119, w_000_3120, w_000_3121, w_000_3122, w_000_3123, w_000_3124, w_000_3125, w_000_3126, w_000_3127, w_000_3128, w_000_3129, w_000_3130, w_000_3131, w_000_3132, w_000_3133, w_000_3134, w_000_3135, w_000_3136, w_000_3137, w_000_3138, w_000_3139, w_000_3140, w_000_3141, w_000_3142, w_000_3143, w_000_3144, w_000_3145, w_000_3146, w_000_3147, w_000_3148, w_000_3149, w_000_3150, w_000_3151, w_000_3152, w_000_3153, w_000_3154, w_000_3155, w_000_3156, w_000_3157, w_000_3158, w_000_3159, w_000_3160, w_000_3161, w_000_3162, w_000_3163, w_000_3164, w_000_3165, w_000_3166, w_000_3167, w_000_3168, w_000_3169, w_000_3170, w_000_3171, w_000_3172, w_000_3173, w_000_3174, w_000_3175, w_000_3176, w_000_3177, w_000_3178, w_000_3179, w_000_3180, w_000_3181, w_000_3182, w_000_3183, w_000_3184, w_000_3185, w_000_3186, w_000_3187, w_000_3188, w_000_3189, w_000_3190, w_000_3191, w_000_3192, w_000_3193, w_000_3194, w_000_3195, w_000_3196, w_000_3197, w_000_3198, w_000_3199, w_000_3200, w_000_3201, w_000_3202, w_000_3203, w_000_3204, w_000_3205, w_000_3206, w_000_3207, w_000_3208, w_000_3209, w_000_3210, w_000_3211, w_000_3212, w_000_3213, w_000_3214, w_000_3215, w_000_3216, w_000_3217, w_000_3218, w_000_3219, w_000_3220, w_000_3221, w_000_3222, w_000_3223, w_000_3224, w_000_3225, w_000_3226, w_000_3227, w_000_3228, w_000_3229, w_000_3230, w_000_3231, w_000_3232, w_000_3233, w_000_3234, w_000_3235, w_000_3236, w_000_3237, w_000_3238, w_000_3239, w_000_3240, w_000_3241, w_000_3242, w_000_3243, w_000_3244, w_000_3245, w_000_3246, w_000_3247, w_000_3248, w_000_3249, w_000_3250, w_000_3251, w_000_3252, w_000_3253, w_000_3254, w_000_3255, w_000_3256, w_000_3257, w_000_3258, w_000_3259, w_000_3260, w_000_3261, w_000_3262, w_000_3263, w_000_3264, w_000_3265, w_000_3266, w_000_3267, w_000_3268, w_000_3269, w_000_3270, w_000_3271, w_000_3272, w_000_3273, w_000_3274, w_000_3275, w_000_3276, w_000_3277, w_000_3278, w_000_3279, w_000_3280, w_000_3281, w_000_3282, w_000_3283, w_000_3284, w_000_3285, w_000_3286, w_000_3287, w_000_3288, w_000_3289, w_000_3290, w_000_3291, w_000_3292, w_000_3293, w_000_3294, w_000_3295, w_000_3296, w_000_3297, w_000_3298, w_000_3299, w_000_3300, w_000_3301, w_000_3302, w_000_3303, w_000_3304, w_000_3305, w_000_3306, w_000_3307, w_000_3308, w_000_3309, w_000_3310, w_000_3311, w_000_3312, w_000_3313, w_000_3314, w_000_3315, w_000_3316, w_000_3317, w_000_3318, w_000_3319, w_000_3320, w_000_3321, w_000_3322, w_000_3323, w_000_3324, w_000_3325, w_000_3326, w_000_3327, w_000_3328, w_000_3329, w_000_3330, w_000_3331, w_000_3332, w_000_3333, w_000_3334, w_000_3335, w_000_3336, w_000_3337, w_000_3338, w_000_3339, w_000_3340, w_000_3341, w_000_3342, w_000_3343, w_000_3344, w_000_3345, w_000_3346, w_000_3347, w_000_3348, w_000_3349, w_000_3350, w_000_3351, w_000_3352, w_000_3353, w_000_3354, w_000_3355, w_000_3356, w_000_3357, w_000_3358, w_000_3359, w_000_3360, w_000_3361, w_000_3362, w_000_3363, w_000_3364, w_000_3365, w_000_3366, w_000_3367, w_000_3368, w_000_3369, w_000_3370, w_000_3371, w_000_3372, w_000_3373, w_000_3374, w_000_3375, w_000_3376, w_000_3377, w_000_3378, w_000_3379, w_000_3380, w_000_3381, w_000_3382, w_000_3383, w_000_3384, w_000_3385, w_000_3386, w_000_3387, w_000_3388, w_000_3389, w_000_3390, w_000_3391, w_000_3392, w_000_3393, w_000_3394, w_000_3395, w_000_3396, w_000_3397, w_000_3398, w_000_3399, w_000_3400, w_000_3401, w_000_3402, w_000_3403, w_000_3404, w_000_3405, w_000_3406, w_000_3407, w_000_3408, w_000_3409, w_000_3410, w_000_3411, w_000_3412, w_000_3413, w_000_3414, w_000_3415, w_000_3416, w_000_3417, w_000_3418, w_000_3419, w_000_3420, w_000_3421, w_000_3422, w_000_3423, w_000_3424, w_000_3425, w_000_3426, w_000_3427, w_000_3428, w_000_3429, w_000_3430, w_000_3431, w_000_3432, w_000_3433, w_000_3434, w_000_3435, w_000_3436, w_000_3437, w_000_3438, w_000_3439, w_000_3440, w_000_3441, w_000_3442, w_000_3443, w_000_3444, w_000_3445, w_000_3446, w_000_3447, w_000_3448, w_000_3449, w_000_3450, w_000_3451, w_000_3452, w_000_3453, w_000_3454, w_000_3455, w_000_3456, w_000_3457, w_000_3458, w_000_3459, w_000_3460, w_000_3461, w_000_3462, w_000_3463, w_000_3464, w_000_3465, w_000_3466, w_000_3467, w_000_3468, w_000_3469, w_000_3470, w_000_3471, w_000_3472, w_000_3473, w_000_3474, w_000_3475, w_000_3476, w_000_3477, w_000_3478, w_000_3479, w_000_3480, w_000_3481, w_000_3482, w_000_3483, w_000_3484, w_000_3485, w_000_3486, w_000_3487, w_000_3488, w_000_3489, w_000_3490, w_000_3491, w_000_3492, w_000_3493, w_000_3494, w_000_3495, w_000_3496, w_000_3497, w_000_3498, w_000_3499, w_000_3500, w_000_3501, w_000_3502, w_000_3503, w_000_3504, w_000_3505, w_000_3506, w_000_3507, w_000_3508, w_000_3509, w_000_3510, w_000_3511, w_000_3512, w_000_3513, w_000_3514, w_000_3515, w_000_3516, w_000_3517, w_000_3518, w_000_3519, w_000_3520, w_000_3521, w_000_3522, w_000_3523, w_000_3524, w_000_3525, w_000_3526, w_000_3527, w_000_3528, w_000_3529, w_000_3530, w_000_3531, w_000_3532, w_000_3533, w_000_3534, w_000_3535, w_000_3536, w_000_3537, w_000_3538, w_000_3539, w_000_3540, w_000_3541, w_000_3542, w_000_3543, w_000_3544, w_000_3545, w_000_3546, w_000_3547, w_000_3548, w_000_3549, w_000_3550, w_000_3551, w_000_3552, w_000_3553, w_000_3554, w_000_3555, w_000_3556, w_000_3557, w_000_3558, w_000_3559, w_000_3560, w_000_3561, w_000_3562, w_000_3563, w_000_3564, w_000_3565, w_000_3566, w_000_3567, w_000_3568, w_000_3569, w_000_3570, w_000_3571, w_000_3572, w_000_3573, w_000_3574, w_000_3575, w_000_3576, w_000_3577, w_000_3578, w_000_3579, w_000_3580, w_000_3581, w_000_3582, w_000_3583, w_000_3584, w_000_3585, w_000_3586, w_000_3587, w_000_3588, w_000_3589, w_000_3590, w_000_3591, w_000_3592, w_000_3593, w_000_3594, w_000_3595, w_000_3596, w_000_3597, w_000_3598, w_000_3599, w_000_3600, w_000_3601, w_000_3602, w_000_3603, w_000_3604, w_000_3605, w_000_3606, w_000_3607, w_000_3608, w_000_3609, w_000_3610, w_000_3611, w_000_3612, w_000_3613, w_000_3614, w_000_3615, w_000_3616, w_000_3617, w_000_3618, w_000_3619, w_000_3620, w_000_3621, w_000_3622, w_000_3623, w_000_3624, w_000_3625, w_000_3626, w_000_3627, w_000_3628, w_000_3629, w_000_3630, w_000_3631, w_000_3632, w_000_3633, w_000_3634, w_000_3635, w_000_3636, w_000_3637, w_000_3638, w_000_3639, w_000_3640, w_000_3641, w_000_3642, w_000_3643, w_000_3644, w_000_3645, w_000_3646, w_000_3647, w_000_3648, w_000_3649, w_000_3650, w_000_3651, w_000_3652, w_000_3653, w_000_3654, w_000_3655, w_000_3656, w_000_3657, w_000_3658, w_000_3659, w_000_3660, w_000_3661, w_000_3662, w_000_3663, w_000_3664, w_000_3665, w_000_3666, w_000_3667, w_000_3668, w_000_3669, w_000_3670, w_000_3671, w_000_3672, w_000_3673, w_000_3674, w_000_3675, w_000_3676, w_000_3677, w_000_3678, w_000_3679, w_000_3680, w_000_3681, w_000_3682, w_000_3683, w_000_3684, w_000_3685, w_000_3686, w_000_3687, w_000_3688, w_000_3689, w_000_3690, w_000_3691, w_000_3692, w_000_3693, w_000_3694, w_000_3695, w_000_3696, w_000_3697, w_000_3698, w_000_3699, w_000_3700, w_000_3701, w_000_3702, w_000_3703, w_000_3704, w_000_3705, w_000_3706, w_000_3707, w_000_3708, w_000_3709, w_000_3710, w_000_3711, w_000_3712, w_000_3713, w_000_3714, w_000_3715, w_000_3716, w_000_3717, w_000_3718, w_000_3719, w_000_3720, w_000_3721, w_000_3722, w_000_3723, w_000_3724, w_000_3725, w_000_3726, w_000_3727, w_000_3728, w_000_3729, w_000_3730, w_000_3731, w_000_3732, w_000_3733, w_000_3734, w_000_3735, w_000_3736, w_000_3737, w_000_3738, w_000_3739, w_000_3740, w_000_3741, w_000_3742, w_000_3743, w_000_3744, w_000_3745, w_000_3746, w_000_3747, w_000_3748, w_000_3749, w_000_3750, w_000_3751, w_000_3752, w_000_3753, w_000_3754, w_000_3755, w_000_3756, w_000_3757, w_000_3758, w_000_3759, w_000_3760, w_000_3761, w_000_3762, w_000_3763, w_000_3764, w_000_3765, w_000_3766, w_000_3767, w_000_3768, w_000_3769, w_000_3770, w_000_3771, w_000_3772, w_000_3773, w_000_3774, w_000_3775, w_000_3776, w_000_3777, w_000_3778, w_000_3779, w_000_3780, w_000_3781, w_000_3782, w_000_3783, w_000_3784, w_000_3785, w_000_3786, w_000_3787, w_000_3788, w_000_3789, w_000_3790, w_000_3791, w_000_3792, w_000_3793, w_000_3794, w_000_3795, w_000_3796, w_000_3797, w_000_3798, w_000_3799, w_000_3800, w_000_3801, w_000_3802, w_000_3803, w_000_3804, w_000_3805, w_000_3806, w_000_3807, w_000_3808, w_000_3809, w_000_3810, w_000_3811, w_000_3812, w_000_3813, w_000_3814, w_000_3815, w_000_3816, w_000_3817, w_000_3818, w_000_3819, w_000_3820, w_000_3821, w_000_3822, w_000_3823, w_000_3824, w_000_3825, w_000_3826, w_000_3827, w_000_3828, w_000_3829, w_000_3830, w_000_3831, w_000_3832, w_000_3833, w_000_3834, w_000_3835, w_000_3836, w_000_3837, w_000_3838, w_000_3839, w_000_3840, w_000_3841, w_000_3842, w_000_3843, w_000_3844, w_000_3845, w_000_3846, w_000_3847, w_000_3848, w_000_3849, w_000_3850, w_000_3851, w_000_3852, w_000_3853, w_000_3854, w_000_3855, w_000_3856, w_000_3857, w_000_3858, w_000_3859, w_000_3860, w_000_3861, w_000_3862, w_000_3863, w_000_3864, w_000_3865, w_000_3866, w_000_3867, w_000_3868, w_000_3869, w_000_3870, w_000_3871, w_000_3872, w_000_3873, w_000_3874, w_000_3875, w_000_3876, w_000_3877, w_000_3878, w_000_3879, w_000_3880, w_000_3881, w_000_3882, w_000_3883, w_000_3884, w_000_3885, w_000_3886, w_000_3887, w_000_3888, w_000_3889, w_000_3890, w_000_3891, w_000_3892, w_000_3893, w_000_3894, w_000_3895, w_000_3896, w_000_3897, w_000_3898, w_000_3899, w_000_3900, w_000_3901, w_000_3902, w_000_3903, w_000_3904, w_000_3905, w_000_3906, w_000_3907, w_000_3908, w_000_3909, w_000_3910, w_000_3911, w_000_3912, w_000_3913, w_000_3914, w_000_3915, w_000_3916, w_000_3917, w_000_3918, w_000_3919, w_000_3920, w_000_3921, w_000_3922, w_000_3923, w_000_3924, w_000_3925, w_000_3926, w_000_3927, w_000_3928, w_000_3929, w_000_3930, w_000_3931, w_000_3932, w_000_3933, w_000_3934, w_000_3935, w_000_3936, w_000_3937, w_000_3938, w_000_3939, w_000_3940, w_000_3941, w_000_3942, w_000_3943, w_000_3944, w_000_3945, w_000_3946, w_000_3947, w_000_3948, w_000_3949, w_000_3950, w_000_3951, w_000_3952, w_000_3953, w_000_3954, w_000_3955, w_000_3956, w_000_3957, w_000_3958, w_000_3959, w_000_3960, w_000_3961, w_000_3962, w_000_3963, w_000_3964, w_000_3965, w_000_3966, w_000_3967, w_000_3968, w_000_3969, w_000_3970, w_000_3971, w_000_3972, w_000_3973, w_000_3974, w_000_3975, w_000_3976, w_000_3977, w_000_3978, w_000_3979, w_000_3980, w_000_3981, w_000_3982, w_000_3983, w_000_3984, w_000_3985, w_000_3986, w_000_3987, w_000_3988, w_000_3989, w_000_3990, w_000_3991, w_000_3992, w_000_3993, w_000_3994, w_000_3995, w_000_3996, w_000_3997, w_000_3998, w_000_3999, w_000_4000, w_000_4001, w_000_4002, w_000_4003, w_000_4004, w_000_4005, w_000_4006, w_000_4007, w_000_4008, w_000_4009, w_000_4010, w_000_4011, w_000_4012, w_000_4013, w_000_4014, w_000_4015, w_000_4016, w_000_4017, w_000_4018, w_000_4019, w_000_4020, w_000_4022, w_000_4023, w_000_4024, w_000_4025, w_000_4026, w_000_4027, w_000_4028, w_000_4029, w_000_4030, w_000_4031, w_000_4032, w_000_4033, w_000_4034, w_000_4035, w_000_4036, w_000_4037, w_000_4038, w_000_4039, w_000_4040, w_000_4041, w_000_4042, w_000_4043, w_000_4044, w_000_4045, w_000_4046, w_000_4047, w_000_4048, w_000_4049, w_000_4050, w_000_4051, w_000_4052, w_000_4053, w_000_4054, w_000_4055, w_000_4056, w_000_4057, w_000_4058, w_000_4059, w_000_4060, w_000_4061, w_000_4062, w_000_4063, w_000_4064, w_000_4065, w_000_4066, w_000_4067, w_000_4068, w_000_4069, w_000_4070, w_000_4071, w_000_4072, w_000_4073, w_000_4074, w_000_4075, w_000_4076, w_000_4077, w_000_4078, w_000_4079, w_000_4080, w_000_4081, w_000_4082, w_000_4083, w_000_4084, w_000_4085, w_000_4086, w_000_4087, w_000_4088, w_000_4089, w_000_4090, w_000_4091, w_000_4092, w_000_4093, w_000_4094, w_000_4095, w_000_4096, w_000_4097, w_000_4098, w_000_4099, w_000_4100, w_000_4101, w_000_4102, w_000_4103, w_000_4104, w_000_4105, w_000_4106, w_000_4107, w_000_4108, w_000_4109, w_000_4110, w_000_4111, w_000_4112, w_000_4113, w_000_4114, w_000_4115, w_000_4116, w_000_4117, w_000_4118, w_000_4119, w_000_4120, w_000_4121, w_000_4122, w_000_4123, w_000_4124, w_000_4125, w_000_4126, w_000_4127, w_000_4128, w_000_4129, w_000_4130, w_000_4131, w_000_4132, w_000_4133, w_000_4134, w_000_4135, w_000_4136, w_000_4137, w_000_4138, w_000_4139, w_000_4140, w_000_4141, w_000_4142, w_000_4143, w_000_4144, w_000_4145, w_000_4146, w_000_4147, w_000_4148, w_000_4149, w_000_4150, w_000_4151, w_000_4152, w_000_4153, w_000_4154, w_000_4155, w_000_4156, w_000_4157, w_000_4158, w_000_4159, w_000_4160, w_000_4161, w_000_4162, w_000_4163, w_000_4164, w_000_4165, w_000_4166, w_000_4167, w_000_4168, w_000_4169, w_000_4170, w_000_4171, w_000_4172, w_000_4173, w_000_4174, w_000_4175, w_000_4176, w_000_4177, w_000_4178, w_000_4179, w_000_4180, w_000_4181, w_000_4182, w_000_4183, w_000_4184, w_000_4185, w_000_4186, w_000_4187, w_000_4188, w_000_4189, w_000_4190, w_000_4191, w_000_4192, w_000_4193, w_000_4194, w_000_4195, w_000_4196, w_000_4197, w_000_4198, w_000_4199, w_000_4200, w_000_4201, w_000_4202, w_000_4203, w_000_4204, w_000_4205, w_000_4206, w_000_4207, w_000_4208, w_000_4209, w_000_4210, w_000_4211, w_000_4212, w_000_4213, w_000_4214, w_000_4215, w_000_4216, w_000_4217, w_000_4218, w_000_4219, w_000_4220, w_000_4221, w_000_4222, w_000_4223, w_000_4224, w_000_4225, w_000_4226, w_000_4227, w_000_4228, w_000_4229, w_000_4230, w_000_4231, w_000_4232, w_000_4233, w_000_4234, w_000_4235, w_000_4236, w_000_4237, w_000_4238, w_000_4239, w_000_4240, w_000_4241, w_000_4242, w_000_4243, w_000_4245, w_000_4246, w_000_4247, w_000_4248, w_000_4249, w_000_4250, w_000_4251, w_000_4252, w_000_4253, w_000_4254, w_000_4255, w_000_4256, w_000_4257, w_000_4258, w_000_4259, w_000_4260, w_000_4261, w_000_4262, w_000_4263, w_000_4264, w_000_4265, w_000_4266, w_000_4267, w_000_4268, w_000_4269, w_000_4270, w_000_4271, w_000_4272, w_000_4273, w_000_4274, w_000_4275, w_000_4276, w_000_4277, w_000_4278, w_000_4279, w_000_4280, w_000_4281, w_000_4282, w_000_4283, w_000_4284, w_000_4285, w_000_4286, w_000_4287, w_000_4288, w_000_4289, w_000_4290, w_000_4291, w_000_4292, w_000_4293, w_000_4294, w_000_4295, w_000_4296, w_000_4297, w_000_4298, w_000_4299, w_000_4300, w_000_4301, w_000_4302, w_000_4303, w_000_4304, w_000_4305, w_000_4306, w_000_4307, w_000_4308, w_000_4309, w_000_4310, w_000_4311, w_000_4312, w_000_4313, w_000_4314, w_000_4315, w_000_4316, w_000_4317, w_000_4318, w_000_4319, w_000_4320, w_000_4321, w_000_4322, w_000_4323, w_000_4324, w_000_4325, w_000_4326, w_000_4327, w_000_4328, w_000_4329, w_000_4330, w_000_4331, w_000_4332, w_000_4333, w_000_4334, w_000_4335, w_000_4336, w_000_4337, w_000_4338, w_000_4339, w_000_4340, w_000_4341, w_000_4342, w_000_4343, w_000_4344, w_000_4345, w_000_4346, w_000_4347, w_000_4348, w_000_4349, w_000_4350, w_000_4351, w_000_4352, w_000_4353, w_000_4354, w_000_4355, w_000_4356, w_000_4357, w_000_4358, w_000_4359, w_000_4360, w_000_4361, w_000_4362, w_000_4363, w_000_4364, w_000_4365, w_000_4366, w_000_4367, w_000_4368, w_000_4369, w_000_4370, w_000_4371, w_000_4372, w_000_4373, w_000_4374, w_000_4375, w_000_4376, w_000_4377, w_000_4378, w_000_4379, w_000_4380, w_000_4381, w_000_4382, w_000_4383, w_000_4384, w_000_4385, w_000_4386, w_000_4387, w_000_4388, w_000_4389, w_000_4390, w_000_4391, w_000_4392, w_000_4393, w_000_4394, w_000_4395, w_000_4396, w_000_4397, w_000_4398, w_000_4399, w_000_4400, w_000_4401, w_000_4402, w_000_4403, w_000_4404, w_000_4405, w_000_4406, w_000_4407, w_000_4408, w_000_4409, w_000_4410, w_000_4411, w_000_4412, w_000_4413, w_000_4414, w_000_4415, w_000_4416, w_000_4417, w_000_4418, w_000_4419, w_000_4420, w_000_4421, w_000_4422, w_000_4423, w_000_4424, w_000_4425, w_000_4426, w_000_4427, w_000_4428, w_000_4429, w_000_4430, w_000_4431, w_000_4432, w_000_4433, w_000_4434, w_000_4435, w_000_4436, w_000_4437, w_000_4438, w_000_4439, w_000_4440, w_000_4441, w_000_4442, w_000_4443, w_000_4444, w_000_4445, w_000_4446, w_000_4447, w_000_4448, w_000_4449, w_000_4450, w_000_4451, w_000_4452, w_000_4453, w_000_4454, w_000_4455, w_000_4456, w_000_4457, w_000_4458, w_000_4459, w_000_4460, w_000_4461, w_000_4462, w_000_4463, w_000_4464, w_000_4465, w_000_4466, w_000_4467, w_000_4468, w_000_4469, w_000_4470, w_000_4471, w_000_4472, w_000_4473, w_000_4474, w_000_4475, w_000_4476, w_000_4477, w_000_4478, w_000_4479, w_000_4480, w_000_4481, w_000_4482, w_000_4483, w_000_4484, w_000_4485, w_000_4486, w_000_4487, w_000_4488, w_000_4489, w_000_4490, w_000_4491, w_000_4492, w_000_4493, w_000_4494, w_000_4495, w_000_4496, w_000_4497, w_000_4498, w_000_4499, w_000_4500, w_000_4501, w_000_4502, w_000_4503, w_000_4504, w_000_4505, w_000_4506, w_000_4507, w_000_4508, w_000_4509, w_000_4510, w_000_4511, w_000_4512, w_000_4513, w_000_4514, w_000_4515, w_000_4516, w_000_4517, w_000_4518, w_000_4519, w_000_4520, w_000_4521, w_000_4522, w_000_4523, w_000_4524, w_000_4525, w_000_4526, w_000_4527, w_000_4528, w_000_4529, w_000_4530, w_000_4531, w_000_4532, w_000_4533, w_000_4534, w_000_4535, w_000_4536, w_000_4537, w_000_4538, w_000_4539, w_000_4540, w_000_4541, w_000_4542, w_000_4543, w_000_4544, w_000_4545, w_000_4546, w_000_4547, w_000_4548, w_000_4549, w_000_4550, w_000_4551, w_000_4552, w_000_4553, w_000_4554, w_000_4555, w_000_4556, w_000_4557, w_000_4558, w_000_4559, w_000_4560, w_000_4561, w_000_4562, w_000_4563, w_000_4564, w_000_4565, w_000_4566, w_000_4567, w_000_4568, w_000_4569, w_000_4570, w_000_4571, w_000_4572, w_000_4573, w_000_4574, w_000_4575, w_000_4576, w_000_4577, w_000_4578, w_000_4579, w_000_4580, w_000_4581, w_000_4582, w_000_4583, w_000_4584, w_000_4585, w_000_4586, w_000_4588, w_000_4589, w_000_4590, w_000_4591, w_000_4592, w_000_4593, w_000_4594, w_000_4595, w_000_4596, w_000_4597, w_000_4598, w_000_4599, w_000_4600, w_000_4601, w_000_4602, w_000_4603, w_000_4604, w_000_4605, w_000_4606, w_000_4607, w_000_4608, w_000_4609, w_000_4610, w_000_4611, w_000_4612, w_000_4613, w_000_4614, w_000_4615, w_000_4616, w_000_4617, w_000_4618, w_000_4619, w_000_4620, w_000_4621, w_000_4622, w_000_4623, w_000_4624, w_000_4625, w_000_4626, w_000_4627, w_000_4628, w_000_4629, w_000_4630, w_000_4631, w_000_4632, w_000_4633, w_000_4634, w_000_4635, w_000_4636, w_000_4637, w_000_4638, w_000_4639, w_000_4640, w_000_4641, w_000_4642, w_000_4643, w_000_4644, w_000_4645, w_000_4646, w_000_4647, w_000_4648, w_000_4649, w_000_4650, w_000_4651, w_000_4652, w_000_4653, w_000_4654, w_000_4655, w_000_4656, w_000_4657, w_000_4658, w_000_4659, w_000_4660, w_000_4661, w_000_4662, w_000_4663, w_000_4664, w_000_4665, w_000_4666, w_000_4667, w_000_4668, w_000_4669, w_000_4670, w_000_4671, w_000_4672, w_000_4673, w_000_4674, w_000_4675, w_000_4676, w_000_4677, w_000_4678, w_000_4679, w_000_4680, w_000_4681, w_000_4682, w_000_4683, w_000_4684, w_000_4685, w_000_4686, w_000_4687, w_000_4688, w_000_4689, w_000_4690, w_000_4691, w_000_4692, w_000_4693, w_000_4694, w_000_4695, w_000_4696, w_000_4697, w_000_4698, w_000_4699, w_000_4700, w_000_4701, w_000_4702, w_000_4703, w_000_4704, w_000_4705, w_000_4706, w_000_4707, w_000_4708, w_000_4709, w_000_4710, w_000_4711, w_000_4712, w_000_4713, w_000_4714, w_000_4715, w_000_4716, w_000_4717, w_000_4718, w_000_4719, w_000_4720, w_000_4721, w_000_4722, w_000_4723, w_000_4724, w_000_4725, w_000_4726, w_000_4727, w_000_4728, w_000_4729, w_000_4730, w_000_4731, w_000_4732, w_000_4733, w_000_4734, w_000_4735, w_000_4736, w_000_4737, w_000_4738, w_000_4739, w_000_4740, w_000_4741, w_000_4742, w_000_4743, w_000_4744, w_000_4745, w_000_4746, w_000_4747, w_000_4748, w_000_4749, w_000_4750, w_000_4751, w_000_4752, w_000_4753, w_000_4754, w_000_4755, w_000_4756, w_000_4757, w_000_4758, w_000_4759, w_000_4760, w_000_4761, w_000_4762, w_000_4763, w_000_4764, w_000_4765, w_000_4766, w_000_4767, w_000_4768, w_000_4769, w_000_4770, w_000_4771, w_000_4772, w_000_4773, w_000_4774, w_000_4775, w_000_4776, w_000_4777, w_000_4778, w_000_4779, w_000_4780, w_000_4781, w_000_4782, w_000_4783, w_000_4784, w_000_4785, w_000_4786, w_000_4787, w_000_4788, w_000_4789, w_000_4790, w_000_4791, w_000_4792, w_000_4793, w_000_4794, w_000_4795, w_000_4796, w_000_4797, w_000_4798, w_000_4799, w_000_4800, w_000_4801, w_000_4802, w_000_4803, w_000_4804, w_000_4805, w_000_4806, w_000_4807, w_000_4808, w_000_4809, w_000_4810, w_000_4811, w_000_4812, w_000_4813, w_000_4814, w_000_4815, w_000_4816, w_000_4817, w_000_4818, w_000_4819, w_000_4820, w_000_4821, w_000_4822, w_000_4823, w_000_4824, w_000_4825, w_000_4826, w_000_4827, w_000_4828, w_000_4829, w_000_4830, w_000_4831, w_000_4832, w_000_4833, w_000_4834, w_000_4835, w_000_4836, w_000_4837, w_000_4838, w_000_4839, w_000_4840, w_000_4841, w_000_4842, w_000_4843, w_000_4844, w_000_4845, w_000_4846, w_000_4847, w_000_4848, w_000_4849, w_000_4850, w_000_4851, w_000_4852, w_000_4853, w_000_4854, w_000_4855, w_000_4856, w_000_4857, w_000_4858, w_000_4859, w_000_4860, w_000_4861, w_000_4862, w_000_4863, w_000_4864, w_000_4865, w_000_4866, w_000_4867, w_000_4868, w_000_4869, w_000_4870, w_000_4871, w_000_4872, w_000_4873, w_000_4874, w_000_4875, w_000_4876, w_000_4877, w_000_4878, w_000_4879, w_000_4880, w_000_4881, w_000_4882, w_000_4883, w_000_4884, w_000_4885, w_000_4886, w_000_4887, w_000_4888, w_000_4889, w_000_4890, w_000_4891, w_000_4892, w_000_4893, w_000_4894, w_000_4895, w_000_4896, w_000_4897, w_000_4898, w_000_4899, w_000_4900, w_000_4901, w_000_4902, w_000_4903, w_000_4904, w_000_4905, w_000_4906, w_000_4907, w_000_4908, w_000_4909, w_000_4910, w_000_4911, w_000_4912, w_000_4913, w_000_4914, w_000_4915, w_000_4916, w_000_4917, w_000_4918, w_000_4919, w_000_4920, w_000_4921, w_000_4922, w_000_4923, w_000_4924, w_000_4925, w_000_4926, w_000_4927, w_000_4928, w_000_4929, w_000_4930, w_000_4931, w_000_4932, w_000_4933, w_000_4934, w_000_4935, w_000_4936, w_000_4937, w_000_4938, w_000_4939, w_000_4940, w_000_4941, w_000_4942, w_000_4943, w_000_4944, w_000_4945, w_000_4946, w_000_4947, w_000_4948, w_000_4949, w_000_4950, w_000_4951, w_000_4952, w_000_4953, w_000_4954, w_000_4955, w_000_4956, w_000_4957, w_000_4958, w_000_4959, w_000_4960, w_000_4961, w_000_4962, w_000_4963, w_000_4964, w_000_4965, w_000_4966, w_000_4967, w_000_4968, w_000_4969, w_000_4970, w_000_4971, w_000_4972, w_000_4973, w_000_4974, w_000_4975, w_000_4976, w_000_4977, w_000_4978, w_000_4979, w_000_4980, w_000_4981, w_000_4982, w_000_4983, w_000_4984, w_000_4985, w_000_4986, w_000_4987, w_000_4988, w_000_4989, w_000_4990, w_000_4991, w_000_4992, w_000_4993, w_000_4994, w_000_4995, w_000_4996, w_000_4997, w_000_4998, w_000_4999, w_000_5000, w_000_5001, w_000_5002, w_000_5003, w_000_5004, w_000_5005, w_000_5006, w_000_5007, w_000_5008, w_000_5009, w_000_5010, w_000_5011, w_000_5012, w_000_5013, w_000_5014, w_000_5015, w_000_5016, w_000_5017, w_000_5018, w_000_5019, w_000_5020, w_000_5021, w_000_5022, w_000_5023, w_000_5024, w_000_5025, w_000_5026, w_000_5027, w_000_5028, w_000_5029, w_000_5030, w_000_5031, w_000_5032, w_000_5033, w_000_5034, w_000_5035, w_000_5036, w_000_5037, w_000_5038, w_000_5039, w_000_5040, w_000_5041, w_000_5042, w_000_5043, w_000_5044, w_000_5045, w_000_5046, w_000_5047, w_000_5048, w_000_5049, w_000_5050, w_000_5051, w_000_5052, w_000_5053, w_000_5054, w_000_5055, w_000_5056, w_000_5057, w_000_5058, w_000_5059, w_000_5060, w_000_5061, w_000_5062, w_000_5063, w_000_5064, w_000_5065, w_000_5066, w_000_5067, w_000_5068, w_000_5069, w_000_5070, w_000_5071, w_000_5072, w_000_5073, w_000_5074, w_000_5075, w_000_5076, w_000_5077, w_000_5078, w_000_5079, w_000_5080, w_000_5081, w_000_5082, w_000_5083, w_000_5084, w_000_5085, w_000_5086, w_000_5087, w_000_5088, w_000_5089, w_000_5090, w_000_5091, w_000_5092, w_000_5093, w_000_5094, w_000_5095, w_000_5096, w_000_5097, w_000_5098, w_000_5099, w_000_5100, w_000_5101, w_000_5102, w_000_5103, w_000_5104, w_000_5105, w_000_5106, w_000_5107, w_000_5108, w_000_5109, w_000_5110, w_000_5111, w_000_5112, w_000_5113, w_000_5114, w_000_5115, w_000_5116, w_000_5117, w_000_5118, w_000_5119, w_000_5120, w_000_5121, w_000_5122, w_000_5123, w_000_5124, w_000_5125, w_000_5126, w_000_5127, w_000_5128, w_000_5129, w_000_5130, w_000_5131, w_000_5132, w_000_5133, w_000_5134, w_000_5135, w_000_5136, w_000_5137, w_000_5138, w_000_5139, w_000_5140, w_000_5141, w_000_5142, w_000_5143, w_000_5144, w_000_5145, w_000_5146, w_000_5147, w_000_5148, w_000_5149, w_000_5150, w_000_5151, w_000_5152, w_000_5153, w_000_5154, w_000_5155, w_000_5156, w_000_5157, w_000_5158, w_000_5159, w_000_5160, w_000_5161, w_000_5162, w_000_5163, w_000_5164, w_000_5165, w_000_5166, w_000_5167, w_000_5168, w_000_5169, w_000_5170, w_000_5171, w_000_5172, w_000_5173, w_000_5174, w_000_5175, w_000_5176, w_000_5177, w_000_5178, w_000_5179, w_000_5180, w_000_5181, w_000_5182, w_000_5183, w_000_5184, w_000_5185, w_000_5186, w_000_5187, w_000_5188, w_000_5189, w_000_5190, w_000_5191, w_000_5192, w_000_5193, w_000_5194, w_000_5195, w_000_5196, w_000_5197, w_000_5198, w_000_5199, w_000_5200, w_000_5201, w_000_5202, w_000_5203, w_000_5204, w_000_5205, w_000_5206, w_000_5207, w_000_5208, w_000_5209, w_000_5210, w_000_5211, w_000_5212, w_000_5213, w_000_5214, w_000_5215, w_000_5216, w_000_5217, w_000_5218, w_000_5219, w_000_5220, w_000_5221, w_000_5222, w_000_5223, w_000_5224, w_000_5225, w_000_5226, w_000_5227, w_000_5228, w_000_5229, w_000_5230, w_000_5231, w_000_5232, w_000_5233, w_000_5234, w_000_5235, w_000_5236, w_000_5237, w_000_5238, w_000_5239, w_000_5240, w_000_5241, w_000_5242, w_000_5243, w_000_5244, w_000_5245, w_000_5246, w_000_5247, w_000_5248, w_000_5249, w_000_5250, w_000_5251, w_000_5252, w_000_5253, w_000_5254, w_000_5255, w_000_5256, w_000_5257, w_000_5258, w_000_5259, w_000_5260, w_000_5261, w_000_5262, w_000_5263, w_000_5264, w_000_5265, w_000_5266, w_000_5267, w_000_5268, w_000_5269, w_000_5270, w_000_5271, w_000_5272, w_000_5273, w_000_5274, w_000_5275, w_000_5276, w_000_5277, w_000_5278, w_000_5279, w_000_5280, w_000_5281, w_000_5282, w_000_5283, w_000_5284, w_000_5285, w_000_5286, w_000_5287, w_000_5288, w_000_5289, w_000_5290, w_000_5291, w_000_5292, w_000_5293, w_000_5294, w_000_5295, w_000_5296, w_000_5297, w_000_5298, w_000_5299, w_000_5300, w_000_5301, w_000_5302, w_000_5303, w_000_5304, w_000_5305, w_000_5306, w_000_5307, w_000_5308, w_000_5309, w_000_5310, w_000_5311, w_000_5312, w_000_5313, w_000_5314, w_000_5315, w_000_5316, w_000_5317, w_000_5318, w_000_5319, w_000_5320, w_000_5321, w_000_5322, w_000_5323, w_000_5324, w_000_5325, w_000_5326, w_000_5327, w_000_5328, w_000_5329, w_000_5330, w_000_5331, w_000_5332, w_000_5333, w_000_5334, w_000_5335, w_000_5336, w_000_5337, w_000_5338, w_000_5339, w_000_5340, w_000_5341, w_000_5342, w_000_5343, w_000_5344, w_000_5345, w_000_5346, w_000_5347, w_000_5348, w_000_5349, w_000_5350, w_000_5351, w_000_5352, w_000_5353, w_000_5354, w_000_5355, w_000_5356, w_000_5357, w_000_5358, w_000_5359, w_000_5360, w_000_5361, w_000_5362, w_000_5363, w_000_5364, w_000_5365, w_000_5366, w_000_5367, w_000_5368, w_000_5369, w_000_5370, w_000_5371, w_000_5372, w_000_5373, w_000_5374, w_000_5375, w_000_5376, w_000_5377, w_000_5378, w_000_5379, w_000_5380, w_000_5381, w_000_5382, w_000_5383, w_000_5384, w_000_5385, w_000_5386, w_000_5387, w_000_5388, w_000_5389, w_000_5390, w_000_5391, w_000_5392, w_000_5393, w_000_5394, w_000_5395, w_000_5396, w_000_5397, w_000_5398, w_000_5399, w_000_5400, w_000_5401, w_000_5402, w_000_5403, w_000_5404, w_000_5405, w_000_5406, w_000_5407, w_000_5408, w_000_5409, w_000_5410, w_000_5411, w_000_5412, w_000_5413, w_000_5414, w_000_5415, w_000_5416, w_000_5417, w_000_5418, w_000_5419, w_000_5420, w_000_5421, w_000_5422, w_000_5423, w_000_5424, w_000_5425, w_000_5426, w_000_5427, w_000_5428, w_000_5429, w_000_5430, w_000_5431, w_000_5432, w_000_5433, w_000_5434, w_000_5435, w_000_5436, w_000_5437, w_000_5438, w_000_5439, w_000_5440, w_000_5441, w_000_5442, w_000_5443, w_000_5444, w_000_5445, w_000_5446, w_000_5447, w_000_5448, w_000_5449, w_000_5450, w_000_5451, w_000_5452, w_000_5453, w_000_5454, w_000_5455, w_000_5456, w_000_5457, w_000_5458, w_000_5459, w_000_5460, w_000_5461, w_000_5462, w_000_5463, w_000_5464, w_000_5465, w_000_5466, w_000_5467, w_000_5468, w_000_5469, w_000_5470, w_000_5471, w_000_5472, w_000_5473, w_000_5474, w_000_5475, w_000_5476, w_000_5477, w_000_5478, w_000_5479, w_000_5480, w_000_5481, w_000_5482, w_000_5483, w_000_5484, w_000_5485, w_000_5486, w_000_5487, w_000_5488, w_000_5489, w_000_5490, w_000_5491, w_000_5492, w_000_5493, w_000_5494, w_000_5495, w_000_5496, w_000_5497, w_000_5498, w_000_5499, w_000_5500, w_000_5501, w_000_5502, w_000_5503, w_000_5504, w_000_5505, w_000_5506, w_000_5507, w_000_5508, w_000_5509, w_000_5510, w_000_5511, w_000_5512, w_000_5513, w_000_5514, w_000_5515, w_000_5516, w_000_5517, w_000_5518, w_000_5519, w_000_5520, w_000_5521, w_000_5522, w_000_5523, w_000_5524, w_000_5525, w_000_5526, w_000_5527, w_000_5528, w_000_5529, w_000_5530, w_000_5531, w_000_5532, w_000_5533, w_000_5534, w_000_5535, w_000_5536, w_000_5537, w_000_5538, w_000_5539, w_000_5540, w_000_5541, w_000_5542, w_000_5543, w_000_5544, w_000_5545, w_000_5546, w_000_5547, w_000_5548, w_000_5549, w_000_5550, w_000_5551, w_000_5552, w_000_5553, w_000_5554, w_000_5555, w_000_5556, w_000_5557, w_000_5558, w_000_5559, w_000_5560, w_000_5561, w_000_5562, w_000_5563, w_000_5564, w_000_5565, w_000_5566, w_000_5567, w_000_5568, w_000_5569, w_000_5570, w_000_5571, w_000_5572, w_000_5573, w_000_5574, w_000_5575, w_000_5576, w_000_5577, w_000_5578, w_000_5579, w_000_5580, w_000_5581, w_000_5582, w_000_5583, w_000_5584, w_000_5585, w_000_5586, w_000_5587, w_000_5588, w_000_5589, w_000_5590, w_000_5591, w_000_5592, w_000_5593, w_000_5594, w_000_5595, w_000_5596, w_000_5597, w_000_5598, w_000_5599, w_000_5600, w_000_5601, w_000_5602, w_000_5603, w_000_5604, w_000_5605, w_000_5606, w_000_5607, w_000_5608, w_000_5609, w_000_5610, w_000_5611, w_000_5612, w_000_5613, w_000_5614, w_000_5615, w_000_5616, w_000_5617, w_000_5618, w_000_5619, w_000_5620, w_000_5621, w_000_5622, w_000_5623, w_000_5624, w_000_5625, w_000_5626, w_000_5627, w_000_5628, w_000_5629, w_000_5630, w_000_5631, w_000_5632, w_000_5633, w_000_5634, w_000_5635, w_000_5636, w_000_5637, w_000_5638, w_000_5639, w_000_5640, w_000_5641, w_000_5642, w_000_5643, w_000_5644, w_000_5645, w_000_5646, w_000_5647, w_000_5648, w_000_5649, w_000_5650, w_000_5651, w_000_5652, w_000_5653, w_000_5654, w_000_5655, w_000_5656, w_000_5657, w_000_5658, w_000_5659, w_000_5660, w_000_5661, w_000_5662, w_000_5663, w_000_5664, w_000_5665, w_000_5666, w_000_5667, w_000_5668, w_000_5669, w_000_5670, w_000_5671, w_000_5672, w_000_5673, w_000_5674, w_000_5675, w_000_5676, w_000_5677, w_000_5678, w_000_5679, w_000_5680, w_000_5681, w_000_5682, w_000_5683, w_000_5684, w_000_5685, w_000_5686, w_000_5687, w_000_5688, w_000_5689, w_000_5690, w_000_5691, w_000_5692, w_000_5693, w_000_5694, w_000_5695, w_000_5696, w_000_5697, w_000_5698, w_000_5699, w_000_5700, w_000_5701, w_000_5702, w_000_5703, w_000_5704, w_000_5705, w_000_5706, w_000_5707, w_000_5708, w_000_5709, w_000_5710, w_000_5711, w_000_5712, w_000_5713, w_000_5714, w_000_5715, w_000_5716, w_000_5717, w_000_5718, w_000_5719, w_000_5720, w_000_5721, w_000_5722, w_000_5723, w_000_5724, w_000_5725, w_000_5726, w_000_5727, w_000_5728, w_000_5729, w_000_5730, w_000_5731, w_000_5732, w_000_5733, w_000_5734, w_000_5735, w_000_5736, w_000_5737, w_000_5738, w_000_5739, w_000_5740, w_000_5741, w_000_5742, w_000_5743, w_000_5744, w_000_5745, w_000_5746, w_000_5747, w_000_5748, w_000_5749, w_000_5750, w_000_5751, w_000_5752, w_000_5753, w_000_5754, w_000_5755, w_000_5756, w_000_5757, w_000_5758, w_000_5759, w_000_5760, w_000_5761, w_000_5762, w_000_5763, w_000_5764, w_000_5765, w_000_5766, w_000_5767, w_000_5768, w_000_5769, w_000_5770, w_000_5771, w_000_5772, w_000_5773, w_000_5774, w_000_5775, w_000_5776, w_000_5777, w_000_5778, w_000_5779, w_000_5780, w_000_5781, w_000_5782, w_000_5783, w_000_5784, w_000_5785, w_000_5786, w_000_5787, w_000_5788, w_000_5789, w_000_5790, w_000_5791, w_000_5792, w_000_5793, w_000_5794, w_000_5795, w_000_5796, w_000_5797, w_000_5798, w_000_5799, w_000_5800, w_000_5801, w_000_5802, w_000_5803, w_000_5804, w_000_5805, w_000_5806, w_000_5807, w_000_5808, w_000_5809, w_000_5810, w_000_5811, w_000_5812, w_000_5813, w_000_5814, w_000_5815, w_000_5816, w_000_5817, w_000_5818, w_000_5819, w_000_5820, w_000_5821, w_000_5822, w_000_5823, w_000_5824, w_000_5825, w_000_5826, w_000_5827, w_000_5828, w_000_5829, w_000_5830, w_000_5831, w_000_5832, w_000_5833, w_000_5834, w_000_5835, w_000_5836, w_000_5837, w_000_5838, w_000_5839, w_000_5840, w_000_5841, w_000_5842, w_000_5843, w_000_5844, w_000_5845, w_000_5846, w_000_5847, w_000_5848, w_000_5849, w_000_5850, w_000_5851, w_000_5852, w_000_5853, w_000_5854, w_000_5855, w_000_5856, w_000_5857, w_000_5858, w_000_5859, w_000_5860, w_000_5861, w_000_5862, w_000_5863, w_000_5864, w_000_5865, w_000_5866, w_000_5867, w_000_5868, w_000_5869, w_000_5870, w_000_5871, w_000_5872, w_000_5873, w_000_5874, w_000_5875, w_000_5876, w_000_5877, w_000_5878, w_000_5879, w_000_5880, w_000_5881, w_000_5882, w_000_5883, w_000_5884, w_000_5885, w_000_5886, w_000_5887, w_000_5888, w_000_5889, w_000_5890, w_000_5891, w_000_5892, w_000_5893, w_000_5894, w_000_5895, w_000_5896, w_000_5897, w_000_5898, w_000_5899, w_000_5900, w_000_5901, w_000_5902, w_000_5903, w_000_5904, w_000_5905, w_000_5906, w_000_5907, w_000_5908, w_000_5909, w_000_5910, w_000_5911, w_000_5912, w_000_5913, w_000_5914, w_000_5915, w_000_5916, w_000_5917, w_000_5918, w_000_5919, w_000_5920, w_000_5921, w_000_5922, w_000_5923, w_000_5924, w_000_5925, w_000_5926, w_000_5927, w_000_5928, w_000_5929, w_000_5930, w_000_5931, w_000_5932, w_000_5933, w_000_5934, w_000_5935, w_000_5936, w_000_5937, w_000_5938, w_000_5939, w_000_5940, w_000_5941, w_000_5942, w_000_5943, w_000_5944, w_000_5945, w_000_5946, w_000_5947, w_000_5948, w_000_5949, w_000_5950, w_000_5951, w_000_5952, w_000_5953, w_000_5954, w_000_5955, w_000_5956, w_000_5957, w_000_5958, w_000_5959, w_000_5960, w_000_5961, w_000_5962, w_000_5963, w_000_5964, w_000_5965, w_000_5966, w_000_5967, w_000_5968, w_000_5969, w_000_5970, w_000_5971, w_000_5972, w_000_5973, w_000_5974, w_000_5975, w_000_5976, w_000_5977, w_000_5978, w_000_5979, w_000_5980, w_000_5981, w_000_5982, w_000_5983, w_000_5984, w_000_5985, w_000_5986, w_000_5987, w_000_5988, w_000_5989, w_000_5990, w_000_5991, w_000_5992, w_000_5993, w_000_5994, w_000_5995, w_000_5996, w_000_5997, w_000_5998, w_000_5999, w_000_6000, w_000_6001, w_000_6002, w_000_6003, w_000_6004, w_000_6005, w_000_6006, w_000_6007, w_000_6008, w_000_6009, w_000_6010, w_000_6011, w_000_6012, w_000_6013, w_000_6014, w_000_6015, w_000_6016, w_000_6017, w_000_6018, w_000_6019, w_000_6020, w_000_6021, w_000_6022, w_000_6023, w_000_6024, w_000_6025, w_000_6026, w_000_6027, w_000_6028, w_000_6029, w_000_6030, w_000_6031, w_000_6032, w_000_6033, w_000_6034, w_000_6035, w_000_6036, w_000_6037, w_000_6038, w_000_6039, w_000_6040, w_000_6041, w_000_6042, w_000_6043, w_000_6044, w_000_6045, w_000_6046, w_000_6047, w_000_6048, w_000_6049, w_000_6050, w_000_6051, w_000_6052, w_000_6053, w_000_6054, w_000_6055, w_000_6056, w_000_6057, w_000_6058, w_000_6059, w_000_6060, w_000_6061, w_000_6062, w_000_6063, w_000_6064, w_000_6065, w_000_6066, w_000_6067, w_000_6068, w_000_6069, w_000_6070, w_000_6071, w_000_6072, w_000_6073, w_000_6074, w_000_6075, w_000_6076, w_000_6077, w_000_6078, w_000_6079, w_000_6080, w_000_6081, w_000_6082, w_000_6083, w_000_6084, w_000_6085, w_000_6086, w_000_6087, w_000_6088, w_000_6089, w_000_6090, w_000_6091, w_000_6092, w_000_6093, w_000_6094, w_000_6095, w_000_6096, w_000_6097, w_000_6098, w_000_6099, w_000_6100, w_000_6101, w_000_6102, w_000_6103, w_000_6104, w_000_6105, w_000_6106, w_000_6107, w_000_6108, w_000_6109, w_000_6110, w_000_6111, w_000_6112, w_000_6113, w_000_6114, w_000_6115, w_000_6116, w_000_6117, w_000_6118, w_000_6119, w_000_6120, w_000_6121, w_000_6122, w_000_6123, w_000_6124, w_000_6125, w_000_6126, w_000_6127, w_000_6128, w_000_6129, w_000_6130, w_000_6131, w_000_6132, w_000_6133, w_000_6134, w_000_6135, w_000_6136, w_000_6137, w_000_6138, w_000_6139, w_000_6140, w_000_6141, w_000_6142, w_000_6143, w_000_6144, w_000_6145, w_000_6146, w_000_6147, w_000_6148, w_000_6149, w_000_6150, w_000_6151, w_000_6152, w_000_6153, w_000_6154, w_000_6155, w_000_6156, w_000_6157, w_000_6158, w_000_6159, w_000_6160, w_000_6161, w_000_6162, w_000_6163, w_000_6164, w_000_6165, w_000_6166, w_000_6167, w_000_6168, w_000_6169, w_000_6170, w_000_6171, w_000_6172, w_000_6173, w_000_6174, w_000_6175, w_000_6176, w_000_6177, w_000_6178, w_000_6179, w_000_6180, w_000_6181, w_000_6182, w_000_6183, w_000_6184, w_000_6185, w_000_6186, w_000_6187, w_000_6188, w_000_6189, w_000_6190, w_000_6191, w_000_6192, w_000_6193, w_000_6194, w_000_6195, w_000_6196, w_000_6197, w_000_6198, w_000_6199, w_000_6200, w_000_6201, w_000_6202, w_000_6203, w_000_6204, w_000_6205, w_000_6206, w_000_6207, w_000_6208, w_000_6209, w_000_6210, w_000_6211, w_000_6212, w_000_6213, w_000_6214, w_000_6215, w_000_6216, w_000_6217, w_000_6218, w_000_6219, w_000_6220, w_000_6221, w_000_6222, w_000_6223, w_000_6224, w_000_6225, w_000_6226, w_000_6227, w_000_6228, w_000_6229, w_000_6230, w_000_6231, w_000_6232, w_000_6233, w_000_6234, w_000_6235, w_000_6236, w_000_6237, w_000_6238, w_000_6239, w_000_6240, w_000_6241, w_000_6242, w_000_6243, w_000_6244, w_000_6245, w_000_6246, w_000_6247, w_000_6248, w_000_6249, w_000_6250, w_000_6251, w_000_6252, w_000_6253, w_000_6254, w_000_6255, w_000_6256, w_000_6257, w_000_6258, w_000_6259, w_000_6260, w_000_6261, w_000_6262, w_000_6263, w_000_6264, w_000_6265, w_000_6266, w_000_6267, w_000_6268, w_000_6269, w_000_6270, w_000_6271, w_000_6272, w_000_6273, w_000_6274, w_000_6275, w_000_6276, w_000_6277, w_000_6278, w_000_6279, w_000_6280, w_000_6281, w_000_6282, w_000_6283, w_000_6284, w_000_6285, w_000_6286, w_000_6287, w_000_6288, w_000_6289, w_000_6290, w_000_6291, w_000_6293, w_000_6294, w_000_6295, w_000_6296, w_000_6297, w_000_6298, w_000_6299, w_000_6300, w_000_6301, w_000_6302, w_000_6303, w_000_6304, w_000_6305, w_000_6306, w_000_6307, w_000_6308, w_000_6309, w_000_6310, w_000_6311, w_000_6312, w_000_6313, w_000_6314, w_000_6315, w_000_6316, w_000_6317, w_000_6318, w_000_6319, w_000_6320, w_000_6321, w_000_6322, w_000_6323, w_000_6324, w_000_6325, w_000_6326, w_000_6327, w_000_6328, w_000_6329, w_000_6330, w_000_6331, w_000_6332, w_000_6333, w_000_6334, w_000_6335, w_000_6336, w_000_6337, w_000_6338, w_000_6339, w_000_6340, w_000_6341, w_000_6342, w_000_6343, w_000_6344, w_000_6345, w_000_6346, w_000_6347, w_000_6348, w_000_6349, w_000_6350, w_000_6351, w_000_6352, w_000_6353, w_000_6354, w_000_6355, w_000_6356, w_000_6357, w_000_6358, w_000_6359, w_000_6360, w_000_6361, w_000_6362, w_000_6363, w_000_6364, w_000_6365, w_000_6366, w_000_6367, w_000_6368, w_000_6369, w_000_6370, w_000_6371, w_000_6372, w_000_6373, w_000_6374, w_000_6375, w_000_6376, w_000_6377, w_000_6378, w_000_6379, w_000_6380, w_000_6381, w_000_6382, w_000_6383, w_000_6384, w_000_6385, w_000_6386, w_000_6387, w_000_6388, w_000_6389, w_000_6390, w_000_6391, w_000_6392, w_000_6393, w_000_6394, w_000_6395, w_000_6396, w_000_6397, w_000_6398, w_000_6399, w_000_6400, w_000_6401, w_000_6402, w_000_6403, w_000_6404, w_000_6405, w_000_6406, w_000_6407, w_000_6408, w_000_6409, w_000_6410, w_000_6411, w_000_6412, w_000_6413, w_000_6414, w_000_6415, w_000_6416, w_000_6417, w_000_6418, w_000_6419, w_000_6420, w_000_6421, w_000_6422, w_000_6423, w_000_6424, w_000_6425, w_000_6426, w_000_6427, w_000_6428, w_000_6429, w_000_6430, w_000_6431, w_000_6432, w_000_6433, w_000_6434, w_000_6435, w_000_6436, w_000_6437, w_000_6438, w_000_6439, w_000_6440, w_000_6441, w_000_6442, w_000_6443, w_000_6444, w_000_6445, w_000_6446, w_000_6447, w_000_6448, w_000_6449, w_000_6450, w_000_6451, w_000_6452, w_000_6453, w_000_6454, w_000_6455, w_000_6456, w_000_6457, w_000_6458, w_000_6459, w_000_6460, w_000_6461, w_000_6462, w_000_6463, w_000_6464, w_000_6465, w_000_6466, w_000_6467, w_000_6468, w_000_6469, w_000_6470, w_000_6471, w_000_6472, w_000_6473, w_000_6474, w_000_6475, w_000_6476, w_000_6477, w_000_6478, w_000_6479, w_000_6480, w_000_6481, w_000_6482, w_000_6483, w_000_6484, w_000_6485, w_000_6486, w_000_6487, w_000_6488, w_000_6489, w_000_6490, w_000_6491, w_000_6492, w_000_6493, w_000_6494, w_000_6495, w_000_6496, w_000_6497, w_000_6498, w_000_6499, w_000_6500, w_000_6501, w_000_6502, w_000_6503, w_000_6504, w_000_6505, w_000_6506, w_000_6507, w_000_6508, w_000_6509, w_000_6510, w_000_6511, w_000_6512, w_000_6513, w_000_6514, w_000_6515, w_000_6516, w_000_6517, w_000_6518, w_000_6519, w_000_6520, w_000_6521, w_000_6522, w_000_6523, w_000_6524, w_000_6525, w_000_6526, w_000_6527, w_000_6528, w_000_6529, w_000_6530, w_000_6531, w_000_6532, w_000_6533, w_000_6534, w_000_6535, w_000_6536, w_000_6537, w_000_6538, w_000_6539, w_000_6540, w_000_6541, w_000_6542, w_000_6543, w_000_6544, w_000_6545, w_000_6546, w_000_6547, w_000_6548, w_000_6549, w_000_6550, w_000_6551, w_000_6552, w_000_6553, w_000_6554, w_000_6555, w_000_6556, w_000_6557, w_000_6558, w_000_6559, w_000_6560, w_000_6561, w_000_6562, w_000_6563, w_000_6564, w_000_6565, w_000_6566, w_000_6567, w_000_6568, w_000_6569, w_000_6570, w_000_6571, w_000_6572, w_000_6573, w_000_6574, w_000_6575, w_000_6576, w_000_6577, w_000_6578, w_000_6579, w_000_6580, w_000_6581, w_000_6582, w_000_6583, w_000_6584, w_000_6585, w_000_6586, w_000_6587, w_000_6588, w_000_6589, w_000_6590, w_000_6591, w_000_6592, w_000_6593, w_000_6594, w_000_6595, w_000_6596, w_000_6597, w_000_6598, w_000_6599, w_000_6600, w_000_6601, w_000_6602, w_000_6603, w_000_6604, w_000_6605, w_000_6606, w_000_6607, w_000_6608, w_000_6609, w_000_6610, w_000_6611, w_000_6612, w_000_6613, w_000_6614, w_000_6615, w_000_6616, w_000_6617, w_000_6618, w_000_6619, w_000_6620, w_000_6621, w_000_6622, w_000_6623, w_000_6624, w_000_6625, w_000_6626, w_000_6627, w_000_6628, w_000_6629, w_000_6630, w_000_6631, w_000_6632, w_000_6633, w_000_6634, w_000_6635, w_000_6636, w_000_6637, w_000_6638, w_000_6639, w_000_6640, w_000_6641, w_000_6642, w_000_6643, w_000_6644, w_000_6645, w_000_6646, w_000_6647, w_000_6648, w_000_6649, w_000_6650, w_000_6651, w_000_6652, w_000_6653, w_000_6654, w_000_6655, w_000_6656, w_000_6657, w_000_6658, w_000_6659, w_000_6660, w_000_6661, w_000_6662, w_000_6663, w_000_6664, w_000_6665, w_000_6666, w_000_6667, w_000_6668, w_000_6669, w_000_6670, w_000_6671, w_000_6672, w_000_6673, w_000_6674, w_000_6675, w_000_6676, w_000_6677, w_000_6678, w_000_6679, w_000_6680, w_000_6681, w_000_6682, w_000_6683, w_000_6684, w_000_6685, w_000_6686, w_000_6687, w_000_6688, w_000_6689, w_000_6690, w_000_6691, w_000_6692, w_000_6693, w_000_6694, w_000_6695, w_000_6696, w_000_6697, w_000_6698, w_000_6699, w_000_6700, w_000_6701, w_000_6702, w_000_6703, w_000_6704, w_000_6705, w_000_6706, w_000_6707, w_000_6708, w_000_6709, w_000_6710, w_000_6711, w_000_6712, w_000_6714, w_000_6715, w_000_6716, w_000_6717, w_000_6718, w_000_6719, w_000_6720, w_000_6721, w_000_6722, w_000_6723, w_000_6724, w_000_6725, w_000_6726, w_000_6727, w_000_6728, w_000_6729, w_000_6730, w_000_6731, w_000_6732, w_000_6733, w_000_6734, w_000_6735, w_000_6736, w_000_6737, w_000_6738, w_000_6739, w_000_6740, w_000_6741, w_000_6742, w_000_6743, w_000_6744, w_000_6745, w_000_6746, w_000_6747, w_000_6748, w_000_6749, w_000_6750, w_000_6751, w_000_6752, w_000_6753, w_000_6754, w_000_6755, w_000_6756, w_000_6757, w_000_6758, w_000_6759, w_000_6760, w_000_6761, w_000_6762, w_000_6763, w_000_6764, w_000_6765, w_000_6766, w_000_6767, w_000_6768, w_000_6769, w_000_6770, w_000_6771, w_000_6772, w_000_6773, w_000_6774, w_000_6775, w_000_6776, w_000_6777, w_000_6778, w_000_6779, w_000_6780, w_000_6781, w_000_6782, w_000_6783, w_000_6784, w_000_6785, w_000_6786, w_000_6787, w_000_6788, w_000_6789, w_000_6790, w_000_6791, w_000_6792, w_000_6793, w_000_6794, w_000_6795, w_000_6796, w_000_6797, w_000_6798, w_000_6799, w_000_6800, w_000_6801, w_000_6802, w_000_6803, w_000_6804, w_000_6805, w_000_6806, w_000_6807, w_000_6808, w_000_6809, w_000_6810, w_000_6811, w_000_6812, w_000_6813, w_000_6814, w_000_6815, w_000_6816, w_000_6817, w_000_6818, w_000_6819, w_000_6820, w_000_6821, w_000_6822, w_000_6823, w_000_6824, w_000_6825, w_000_6826, w_000_6827, w_000_6828, w_000_6829, w_000_6830, w_000_6831, w_000_6832, w_000_6833, w_000_6834, w_000_6835, w_000_6836, w_000_6837, w_000_6838, w_000_6839, w_000_6840, w_000_6841, w_000_6842, w_000_6843, w_000_6844, w_000_6845, w_000_6846, w_000_6847, w_000_6848, w_000_6849, w_000_6850, w_000_6851, w_000_6852, w_000_6853, w_000_6854, w_000_6855, w_000_6856, w_000_6857, w_000_6858, w_000_6859, w_000_6860, w_000_6861, w_000_6862, w_000_6863, w_000_6864, w_000_6865, w_000_6866, w_000_6867, w_000_6868, w_000_6869, w_000_6870, w_000_6871, w_000_6872, w_000_6873, w_000_6874, w_000_6875, w_000_6876, w_000_6877, w_000_6878, w_000_6879, w_000_6880, w_000_6881, w_000_6882, w_000_6883, w_000_6884, w_000_6885, w_000_6886, w_000_6887, w_000_6888, w_000_6889, w_000_6890, w_000_6891, w_000_6892, w_000_6893, w_000_6894, w_000_6895, w_000_6896, w_000_6897, w_000_6898, w_000_6899, w_000_6900, w_000_6901, w_000_6902, w_000_6903, w_000_6904, w_000_6905, w_000_6906, w_000_6907, w_000_6908, w_000_6909, w_000_6910, w_000_6911, w_000_6912, w_000_6913, w_000_6914, w_000_6915, w_000_6916, w_000_6917, w_000_6918, w_000_6919, w_000_6920, w_000_6921, w_000_6922, w_000_6923, w_000_6924, w_000_6925, w_000_6926, w_000_6927, w_000_6928, w_000_6929, w_000_6930, w_000_6931, w_000_6932, w_000_6933, w_000_6934, w_000_6935, w_000_6936, w_000_6937, w_000_6938, w_000_6939, w_000_6940, w_000_6941, w_000_6942, w_000_6943, w_000_6944, w_000_6945, w_000_6946, w_000_6947, w_000_6948, w_000_6949, w_000_6950, w_000_6951, w_000_6952, w_000_6953, w_000_6954, w_000_6955, w_000_6956, w_000_6957, w_000_6958, w_000_6959, w_000_6960, w_000_6961, w_000_6962, w_000_6963, w_000_6964, w_000_6965, w_000_6966, w_000_6967, w_000_6968, w_000_6969, w_000_6970, w_000_6971, w_000_6972, w_000_6973, w_000_6974, w_000_6975, w_000_6976, w_000_6977, w_000_6978, w_000_6979, w_000_6980, w_000_6981, w_000_6982, w_000_6983, w_000_6984, w_000_6985, w_000_6986, w_000_6987, w_000_6988, w_000_6989, w_000_6990, w_000_6991, w_000_6992, w_000_6993, w_000_6994, w_000_6995, w_000_6996, w_000_6997, w_000_6998, w_000_6999, w_000_7000, w_000_7001, w_000_7002, w_000_7003, w_000_7004, w_000_7005, w_000_7006, w_000_7007, w_000_7008, w_000_7009, w_000_7010, w_000_7011, w_000_7012, w_000_7013, w_000_7014, w_000_7015, w_000_7016, w_000_7017, w_000_7018, w_000_7019, w_000_7020, w_000_7021, w_000_7022, w_000_7023, w_000_7024, w_000_7025, w_000_7026, w_000_7027, w_000_7028, w_000_7029, w_000_7030, w_000_7031, w_000_7032, w_000_7033, w_000_7034, w_000_7035, w_000_7036, w_000_7037, w_000_7038, w_000_7039, w_000_7040, w_000_7041, w_000_7042, w_000_7043, w_000_7044, w_000_7045, w_000_7046, w_000_7047, w_000_7048, w_000_7049, w_000_7050, w_000_7051, w_000_7052, w_000_7053, w_000_7054, w_000_7055, w_000_7056, w_000_7057, w_000_7058, w_000_7059, w_000_7060, w_000_7061, w_000_7062, w_000_7063, w_000_7064, w_000_7065, w_000_7066, w_000_7067, w_000_7068, w_000_7069, w_000_7070, w_000_7071, w_000_7072, w_000_7073, w_000_7074, w_000_7075, w_000_7076, w_000_7077, w_000_7078, w_000_7079, w_000_7080, w_000_7081, w_000_7082, w_000_7083, w_000_7084, w_000_7085, w_000_7086, w_000_7087, w_000_7088, w_000_7089, w_000_7090, w_000_7091, w_000_7092, w_000_7093, w_000_7094, w_000_7095, w_000_7096, w_000_7097, w_000_7098, w_000_7099, w_000_7100, w_000_7101, w_000_7102, w_000_7103, w_000_7104, w_000_7105, w_000_7106, w_000_7107, w_000_7108, w_000_7109, w_000_7110, w_000_7111, w_000_7112, w_000_7113, w_000_7114, w_000_7115, w_000_7116, w_000_7117, w_000_7118, w_000_7119, w_000_7120, w_000_7121, w_000_7122, w_000_7123, w_000_7124, w_000_7125, w_000_7126, w_000_7127, w_000_7128, w_000_7129, w_000_7130, w_000_7131, w_000_7132, w_000_7133, w_000_7134, w_000_7135, w_000_7136, w_000_7137, w_000_7138, w_000_7139, w_000_7140, w_000_7141, w_000_7142, w_000_7143, w_000_7144, w_000_7145, w_000_7146, w_000_7147, w_000_7148, w_000_7149, w_000_7150, w_000_7151, w_000_7152, w_000_7153, w_000_7154, w_000_7155, w_000_7156, w_000_7157, w_000_7158, w_000_7159, w_000_7160, w_000_7161, w_000_7162, w_000_7163, w_000_7164, w_000_7165, w_000_7166, w_000_7167, w_000_7168, w_000_7169, w_000_7170, w_000_7171, w_000_7172, w_000_7173, w_000_7174, w_000_7175, w_000_7176, w_000_7177, w_000_7178, w_000_7179, w_000_7180, w_000_7181, w_000_7182, w_000_7183, w_000_7184, w_000_7185, w_000_7186, w_000_7187, w_000_7188, w_000_7189, w_000_7190, w_000_7191, w_000_7192, w_000_7193, w_000_7194, w_000_7195, w_000_7196, w_000_7197, w_000_7198, w_000_7199, w_000_7200, w_000_7201, w_000_7202, w_000_7203, w_000_7204, w_000_7205, w_000_7206, w_000_7207, w_000_7208, w_000_7209, w_000_7210, w_000_7211, w_000_7212, w_000_7213, w_000_7214, w_000_7215, w_000_7216, w_000_7217, w_000_7218, w_000_7219, w_000_7220, w_000_7221, w_000_7222, w_000_7223, w_000_7224, w_000_7225, w_000_7226, w_000_7227, w_000_7228, w_000_7229, w_000_7230, w_000_7231, w_000_7232, w_000_7233, w_000_7234, w_000_7235, w_000_7236, w_000_7237, w_000_7238, w_000_7239, w_000_7240, w_000_7241, w_000_7242, w_000_7243, w_000_7244, w_000_7245, w_000_7246, w_000_7247, w_000_7248, w_000_7249, w_000_7250, w_000_7251, w_000_7252, w_000_7253, w_000_7254, w_000_7255, w_000_7256, w_000_7257, w_000_7258, w_000_7259, w_000_7260, w_000_7261, w_000_7262, w_000_7263, w_000_7264, w_000_7265, w_000_7266, w_000_7267, w_000_7268, w_000_7269, w_000_7270, w_000_7271, w_000_7272, w_000_7273, w_000_7274, w_000_7275, w_000_7276, w_000_7277, w_000_7278, w_000_7279, w_000_7280, w_000_7281, w_000_7282, w_000_7283, w_000_7284, w_000_7285, w_000_7286, w_000_7287, w_000_7288, w_000_7289, w_000_7290, w_000_7291, w_000_7292, w_000_7293, w_000_7294, w_000_7295, w_000_7296, w_000_7297, w_000_7298, w_000_7299, w_000_7300, w_000_7301, w_000_7302, w_000_7303, w_000_7304, w_000_7305, w_000_7306, w_000_7307, w_000_7308, w_000_7309, w_000_7310, w_000_7311, w_000_7312, w_000_7313, w_000_7314, w_000_7315, w_000_7316, w_000_7317, w_000_7318, w_000_7319, w_000_7320, w_000_7321, w_000_7322, w_000_7323, w_000_7324, w_000_7325, w_000_7326, w_000_7327, w_000_7328, w_000_7329, w_000_7330, w_000_7331, w_000_7332, w_000_7333, w_000_7334, w_000_7335, w_000_7336, w_000_7337, w_000_7338, w_000_7339, w_000_7340, w_000_7341, w_000_7342, w_000_7343, w_000_7344, w_000_7345, w_000_7346, w_000_7347, w_000_7348, w_000_7349, w_000_7350, w_000_7351, w_000_7352, w_000_7353, w_000_7354, w_000_7355, w_000_7356, w_000_7357, w_000_7358, w_000_7359, w_000_7360, w_000_7361, w_000_7362, w_000_7363, w_000_7364, w_000_7365, w_000_7366, w_000_7367, w_000_7368, w_000_7369, w_000_7370, w_000_7371, w_000_7372, w_000_7373, w_000_7374, w_000_7375, w_000_7376, w_000_7377, w_000_7378, w_000_7379, w_000_7380, w_000_7381, w_000_7382, w_000_7383, w_000_7384, w_000_7385, w_000_7386, w_000_7387, w_000_7388, w_000_7389, w_000_7390, w_000_7391, w_000_7392, w_000_7393, w_000_7394, w_000_7395, w_000_7396, w_000_7397, w_000_7398, w_000_7399, w_000_7400, w_000_7401, w_000_7402, w_000_7403, w_000_7404, w_000_7405, w_000_7406, w_000_7407, w_000_7408, w_000_7409, w_000_7410, w_000_7411, w_000_7412, w_000_7413, w_000_7414, w_000_7415, w_000_7416, w_000_7417, w_000_7418, w_000_7419, w_000_7420, w_000_7421, w_000_7422, w_000_7423, w_000_7424, w_000_7425, w_000_7426, w_000_7427, w_000_7428, w_000_7429, w_000_7430, w_000_7431, w_000_7432, w_000_7433, w_000_7434, w_000_7435, w_000_7436, w_000_7437, w_000_7438, w_000_7439, w_000_7440, w_000_7441, w_000_7442, w_000_7443, w_000_7444, w_000_7445, w_000_7446, w_000_7447, w_000_7448, w_000_7449, w_000_7450, w_000_7451, w_000_7452, w_000_7453, w_000_7454, w_000_7455, w_000_7456, w_000_7457, w_000_7458, w_000_7459, w_000_7460, w_000_7461, w_000_7462, w_000_7463, w_000_7464, w_000_7465, w_000_7466, w_000_7467, w_000_7468, w_000_7469, w_000_7470, w_000_7471, w_000_7472, w_000_7473, w_000_7474, w_000_7475, w_000_7476, w_000_7477, w_000_7478, w_000_7479, w_000_7480, w_000_7481, w_000_7482, w_000_7483, w_000_7484, w_000_7485, w_000_7486, w_000_7487, w_000_7488, w_000_7489, w_000_7490, w_000_7491, w_000_7492, w_000_7493, w_000_7494, w_000_7495, w_000_7496, w_000_7497, w_000_7498, w_000_7499, w_000_7500, w_000_7501, w_000_7502, w_000_7503, w_000_7504, w_000_7505, w_000_7506, w_000_7507, w_000_7508, w_000_7509, w_000_7510, w_000_7511, w_000_7512, w_000_7513, w_000_7514, w_000_7515, w_000_7516, w_000_7517, w_000_7518, w_000_7519, w_000_7520, w_000_7521, w_000_7522, w_000_7523, w_000_7524, w_000_7525, w_000_7526, w_000_7527, w_000_7528, w_000_7529, w_000_7530, w_000_7531, w_000_7532, w_000_7533, w_000_7534, w_000_7535, w_000_7536, w_000_7537, w_000_7538, w_000_7539, w_000_7540, w_000_7541, w_000_7542, w_000_7543, w_000_7544, w_000_7545, w_000_7546, w_000_7547, w_000_7548, w_000_7549, w_000_7550, w_000_7551, w_000_7552, w_000_7553, w_000_7554, w_000_7555, w_000_7556, w_000_7557, w_000_7558, w_000_7559, w_000_7560, w_000_7561, w_000_7562, w_000_7563, w_000_7564, w_000_7565, w_000_7566, w_000_7567, w_000_7568, w_000_7569, w_000_7570, w_000_7571, w_000_7572, w_000_7573, w_000_7574, w_000_7575, w_000_7576, w_000_7577, w_000_7578, w_000_7579, w_000_7580, w_000_7581, w_000_7582, w_000_7583, w_000_7584, w_000_7585, w_000_7586, w_000_7587, w_000_7588, w_000_7589, w_000_7590, w_000_7591, w_000_7592, w_000_7593, w_000_7594, w_000_7595, w_000_7596, w_000_7597, w_000_7598, w_000_7599, w_000_7600, w_000_7601, w_000_7602, w_000_7603, w_000_7604, w_000_7605, w_000_7606, w_000_7607, w_000_7608, w_000_7610, w_000_7611, w_000_7612, w_000_7613, w_000_7614, w_000_7615, w_000_7616, w_000_7617, w_000_7618, w_000_7619, w_000_7620, w_000_7621, w_000_7622, w_000_7623, w_000_7624, w_000_7625, w_000_7626, w_000_7627, w_000_7628, w_000_7629, w_000_7630, w_000_7631, w_000_7632, w_000_7633, w_000_7634, w_000_7635, w_000_7636, w_000_7637, w_000_7638, w_000_7639, w_000_7640, w_000_7641, w_000_7642, w_000_7643, w_000_7644, w_000_7645, w_000_7646, w_000_7647, w_000_7648, w_000_7649, w_000_7650, w_000_7651, w_000_7652, w_000_7653, w_000_7654, w_000_7655, w_000_7656, w_000_7657, w_000_7658, w_000_7659, w_000_7660, w_000_7661, w_000_7662, w_000_7663, w_000_7664, w_000_7665, w_000_7666, w_000_7667, w_000_7668, w_000_7669, w_000_7670, w_000_7671, w_000_7672, w_000_7673, w_000_7674, w_000_7675, w_000_7676, w_000_7677, w_000_7678, w_000_7679, w_000_7680, w_000_7681, w_000_7682, w_000_7683, w_000_7684, w_000_7685, w_000_7686, w_000_7687, w_000_7688, w_000_7689, w_000_7690, w_000_7692, w_000_7693, w_000_7694, w_000_7695, w_000_7696, w_000_7697, w_000_7698, w_000_7699, w_000_7700, w_000_7701, w_000_7702, w_000_7703, w_000_7704, w_000_7705, w_000_7706, w_000_7707, w_000_7708, w_000_7709, w_000_7710, w_000_7711, w_000_7712, w_000_7713, w_000_7714, w_000_7715, w_000_7716, w_000_7717, w_000_7718, w_000_7719, w_000_7720, w_000_7721, w_000_7722, w_000_7723, w_000_7724, w_000_7725, w_000_7726, w_000_7727, w_000_7728, w_000_7729, w_000_7730, w_000_7731, w_000_7732, w_000_7733, w_000_7734, w_000_7735, w_000_7736, w_000_7737, w_000_7738, w_000_7739, w_000_7740, w_000_7741, w_000_7742, w_000_7743, w_000_7744, w_000_7745, w_000_7746, w_000_7747, w_000_7748, w_000_7749, w_000_7750, w_000_7751, w_000_7752, w_000_7753, w_000_7754, w_000_7755, w_000_7756, w_000_7757, w_000_7758, w_000_7759, w_000_7760, w_000_7761, w_000_7762, w_000_7763, w_000_7764, w_000_7765, w_000_7766, w_000_7767, w_000_7768, w_000_7769, w_000_7770, w_000_7771, w_000_7772, w_000_7773, w_000_7774, w_000_7775, w_000_7776, w_000_7777, w_000_7778, w_000_7779, w_000_7780, w_000_7781, w_000_7782, w_000_7784, w_000_7785, w_000_7786, w_000_7787, w_000_7788, w_000_7789, w_000_7790, w_000_7791, w_000_7792, w_000_7793, w_000_7794, w_000_7795, w_000_7796, w_000_7797, w_000_7799, w_000_7800, w_000_7801, w_000_7802, w_000_7803, w_000_7804, w_000_7805, w_000_7806, w_000_7807, w_000_7808, w_000_7809, w_000_7810, w_000_7811, w_000_7812, w_000_7813, w_000_7814, w_000_7815, w_000_7816, w_000_7817, w_000_7818, w_000_7819, w_000_7820, w_000_7821, w_000_7822, w_000_7823, w_000_7824, w_000_7825, w_000_7826, w_000_7827, w_000_7828, w_000_7829, w_000_7830, w_000_7831, w_000_7832, w_000_7833, w_000_7834, w_000_7835, w_000_7836, w_000_7837, w_000_7838, w_000_7839, w_000_7840, w_000_7841, w_000_7842, w_000_7843, w_000_7844, w_000_7845, w_000_7846, w_000_7847, w_000_7848, w_000_7849, w_000_7850, w_000_7851, w_000_7852, w_000_7853, w_000_7854, w_000_7855, w_000_7856, w_000_7857, w_000_7858, w_000_7859, w_000_7860, w_000_7861, w_000_7862, w_000_7863, w_000_7864, w_000_7865, w_000_7866, w_000_7867, w_000_7868, w_000_7869, w_000_7870, w_000_7871, w_000_7872, w_000_7874, w_000_7875, w_000_7876, w_000_7877, w_000_7878, w_000_7879, w_000_7880, w_000_7881, w_000_7882, w_000_7883, w_000_7884, w_000_7885, w_000_7886, w_000_7887, w_000_7888, w_000_7889, w_000_7890, w_000_7891, w_000_7892, w_000_7893, w_000_7894, w_000_7895, w_000_7896, w_000_7897, w_000_7898, w_000_7899, w_000_7900, w_000_7901, w_000_7902, w_000_7903, w_000_7904, w_000_7905, w_000_7906, w_000_7907, w_000_7908, w_000_7909, w_000_7910, w_000_7911, w_000_7912, w_000_7913, w_000_7914, w_000_7915, w_000_7916, w_000_7917, w_000_7918, w_000_7919, w_000_7920, w_000_7921, w_000_7922, w_000_7923, w_000_7924, w_000_7925, w_000_7926, w_000_7927, w_000_7928, w_000_7929, w_000_7930, w_000_7931, w_000_7932, w_000_7933, w_000_7934, w_000_7935, w_000_7936, w_000_7937, w_000_7938, w_000_7939, w_000_7940, w_000_7941, w_000_7942, w_000_7943, w_000_7944, w_000_7945, w_000_7946, w_000_7947, w_000_7948, w_000_7949, w_000_7950, w_000_7951, w_000_7952, w_000_7953, w_000_7954, w_000_7955, w_000_7956, w_000_7957, w_000_7958, w_000_7959, w_000_7960, w_000_7961, w_000_7962, w_000_7963, w_000_7964, w_000_7965, w_000_7966, w_000_7967, w_000_7968, w_000_7969, w_000_7970, w_000_7971, w_000_7972, w_000_7973, w_000_7974, w_000_7975, w_000_7976, w_000_7977, w_000_7978, w_000_7979, w_000_7980, w_000_7981, w_000_7982, w_000_7983, w_000_7984, w_000_7985, w_000_7986, w_000_7987, w_000_7988, w_000_7989, w_000_7990, w_000_7991, w_000_7992, w_000_7993, w_000_7994, w_000_7995, w_000_7996, w_000_7997, w_000_7998, w_000_7999, w_000_8000, w_000_8001, w_000_8002, w_000_8003, w_000_8004, w_000_8005, w_000_8006, w_000_8007, w_000_8008, w_000_8009, w_000_8010, w_000_8011, w_000_8012, w_000_8013, w_000_8014, w_000_8015, w_000_8016, w_000_8017, w_000_8018, w_000_8019, w_000_8020, w_000_8021, w_000_8022, w_000_8023, w_000_8024, w_000_8025, w_000_8026, w_000_8027, w_000_8028, w_000_8029, w_000_8030, w_000_8031, w_000_8032, w_000_8033, w_000_8034, w_000_8035, w_000_8036, w_000_8037, w_000_8038, w_000_8039, w_000_8040, w_000_8041, w_000_8042, w_000_8043, w_000_8044, w_000_8045, w_000_8046, w_000_8047, w_000_8048, w_000_8049, w_000_8050, w_000_8051, w_000_8052, w_000_8053, w_000_8054, w_000_8055, w_000_8056, w_000_8057, w_000_8058, w_000_8059, w_000_8060, w_000_8061, w_000_8062, w_000_8063, w_000_8064, w_000_8065, w_000_8066, w_000_8067, w_000_8068, w_000_8069, w_000_8070, w_000_8071, w_000_8072, w_000_8073, w_000_8074, w_000_8075, w_000_8076, w_000_8077, w_000_8078, w_000_8079, w_000_8080, w_000_8081, w_000_8082, w_000_8083, w_000_8084, w_000_8085, w_000_8086, w_000_8087, w_000_8088, w_000_8089, w_000_8090, w_000_8091, w_000_8092, w_000_8093, w_000_8094, w_000_8095, w_000_8096, w_000_8097, w_000_8098, w_000_8099, w_000_8100, w_000_8101, w_000_8102, w_000_8103, w_000_8104, w_000_8105, w_000_8106, w_000_8107, w_000_8108, w_000_8109, w_000_8110, w_000_8111, w_000_8112, w_000_8113, w_000_8114, w_000_8115, w_000_8116, w_000_8117, w_000_8118, w_000_8119, w_000_8120, w_000_8121, w_000_8122, w_000_8123, w_000_8124, w_000_8125, w_000_8126, w_000_8127, w_000_8128, w_000_8129, w_000_8130, w_000_8131, w_000_8132, w_000_8133, w_000_8134, w_000_8135, w_000_8136, w_000_8137, w_000_8138, w_000_8139, w_000_8140, w_000_8141, w_000_8142, w_000_8143, w_000_8144, w_000_8145, w_000_8146, w_000_8147, w_000_8148, w_000_8149, w_000_8150, w_000_8151, w_000_8152, w_000_8153, w_000_8154, w_000_8155, w_000_8156, w_000_8157, w_000_8158, w_000_8159, w_000_8160, w_000_8161, w_000_8162, w_000_8163, w_000_8164, w_000_8165, w_000_8166, w_000_8167, w_000_8168, w_000_8169, w_000_8170, w_000_8171, w_000_8172, w_000_8173, w_000_8174, w_000_8175, w_000_8176, w_000_8177, w_000_8178, w_000_8179, w_000_8180, w_000_8181, w_000_8182, w_000_8183, w_000_8184, w_000_8185, w_000_8186, w_000_8187, w_000_8188, w_000_8189, w_000_8190, w_000_8191, w_000_8192, w_000_8193, w_000_8194, w_000_8195, w_000_8196, w_000_8197, w_000_8198, w_000_8199, w_000_8200, w_000_8201, w_000_8202, w_000_8203, w_000_8204, w_000_8205, w_000_8206, w_000_8207, w_000_8208, w_000_8209, w_000_8210, w_000_8211, w_000_8212, w_000_8213, w_000_8214, w_000_8215, w_000_8216, w_000_8217, w_000_8218, w_000_8219, w_000_8220, w_000_8221, w_000_8222, w_000_8223, w_000_8224, w_000_8225, w_000_8226, w_000_8227, w_000_8228, w_000_8229, w_000_8230, w_000_8231, w_000_8232, w_000_8233, w_000_8234, w_000_8235, w_000_8236, w_000_8237, w_000_8238, w_000_8239, w_000_8240, w_000_8241, w_000_8242, w_000_8243, w_000_8244, w_000_8245, w_000_8246, w_000_8247, w_000_8248, w_000_8249, w_000_8250, w_000_8251, w_000_8252, w_000_8253, w_000_8254, w_000_8255, w_000_8256, w_000_8257, w_000_8258, w_000_8259, w_000_8260, w_000_8261, w_000_8262, w_000_8263, w_000_8264, w_000_8265, w_000_8266, w_000_8267, w_000_8268, w_000_8269, w_000_8270, w_000_8271, w_000_8272, w_000_8273, w_000_8274, w_000_8275, w_000_8276, w_000_8277, w_000_8278, w_000_8279, w_000_8280, w_000_8281, w_000_8282, w_000_8283, w_000_8284, w_000_8285, w_000_8286, w_000_8287, w_000_8288, w_000_8289, w_000_8290, w_000_8291, w_000_8292, w_000_8293, w_000_8294, w_000_8295, w_000_8296, w_000_8297, w_000_8298, w_000_8299, w_000_8300, w_000_8301, w_000_8302, w_000_8303, w_000_8304, w_000_8305, w_000_8306, w_000_8307, w_000_8308, w_000_8309, w_000_8310, w_000_8311, w_000_8312, w_000_8313, w_000_8314, w_000_8315, w_000_8316, w_000_8317, w_000_8318, w_000_8319, w_000_8320, w_000_8321, w_000_8322, w_000_8323, w_000_8324, w_000_8325, w_000_8326, w_000_8327, w_000_8328, w_000_8329, w_000_8330, w_000_8331, w_000_8332, w_000_8333, w_000_8334, w_000_8335, w_000_8336, w_000_8337, w_000_8338, w_000_8339, w_000_8340, w_000_8341, w_000_8342, w_000_8343, w_000_8344, w_000_8345, w_000_8346, w_000_8347, w_000_8348, w_000_8349, w_000_8350, w_000_8351, w_000_8352, w_000_8353, w_000_8354, w_000_8355, w_000_8356, w_000_8357, w_000_8358, w_000_8359, w_000_8360, w_000_8361, w_000_8362, w_000_8363, w_000_8364, w_000_8365, w_000_8366, w_000_8367, w_000_8368, w_000_8369, w_000_8370, w_000_8371, w_000_8372, w_000_8373, w_000_8374, w_000_8375, w_000_8376, w_000_8377, w_000_8378, w_000_8379, w_000_8380, w_000_8381, w_000_8382, w_000_8383, w_000_8384, w_000_8385, w_000_8386, w_000_8387, w_000_8388, w_000_8389, w_000_8390, w_000_8391, w_000_8392, w_000_8393, w_000_8394, w_000_8395, w_000_8396, w_000_8397, w_000_8398, w_000_8399, w_000_8400, w_000_8401, w_000_8402, w_000_8403, w_000_8404, w_000_8405, w_000_8406, w_000_8407, w_000_8408, w_000_8409, w_000_8410, w_000_8411, w_000_8412, w_000_8413, w_000_8414, w_000_8415, w_000_8416, w_000_8417, w_000_8418, w_000_8419, w_000_8420, w_000_8421, w_000_8422, w_000_8423, w_000_8424, w_000_8425, w_000_8426, w_000_8427, w_000_8428, w_000_8429, w_000_8430, w_000_8431, w_000_8432, w_000_8433, w_000_8434, w_000_8435, w_000_8436, w_000_8437, w_000_8438, w_000_8439, w_000_8440, w_000_8441, w_000_8442, w_000_8443, w_000_8444, w_000_8445, w_000_8446, w_000_8447, w_000_8448, w_000_8449, w_000_8450, w_000_8451, w_000_8452, w_000_8453, w_000_8454, w_000_8455, w_000_8456, w_000_8457, w_000_8458, w_000_8459, w_000_8460, w_000_8461, w_000_8462, w_000_8463, w_000_8464, w_000_8465, w_000_8466, w_000_8467, w_000_8468, w_000_8469, w_000_8470, w_000_8471, w_000_8472, w_000_8473, w_000_8474, w_000_8475, w_000_8476, w_000_8477, w_000_8478, w_000_8479, w_000_8480, w_000_8481, w_000_8482, w_000_8483, w_000_8484, w_000_8485, w_000_8486, w_000_8487, w_000_8488, w_000_8489, w_000_8490, w_000_8491, w_000_8492, w_000_8493, w_000_8494, w_000_8495, w_000_8496, w_000_8497, w_000_8498, w_000_8499, w_000_8500, w_000_8501, w_000_8502, w_000_8503, w_000_8504, w_000_8505, w_000_8506, w_000_8507, w_000_8508, w_000_8509, w_000_8510, w_000_8511, w_000_8512, w_000_8513, w_000_8514, w_000_8515, w_000_8516, w_000_8517, w_000_8518, w_000_8519, w_000_8520, w_000_8521, w_000_8522, w_000_8523, w_000_8524, w_000_8525, w_000_8526, w_000_8527, w_000_8528, w_000_8529, w_000_8530, w_000_8531, w_000_8532, w_000_8533, w_000_8534, w_000_8535, w_000_8536, w_000_8537, w_000_8538, w_000_8539, w_000_8540, w_000_8541, w_000_8542, w_000_8543, w_000_8544, w_000_8545, w_000_8546, w_000_8547, w_000_8548, w_000_8549, w_000_8550, w_000_8551, w_000_8552, w_000_8553, w_000_8554, w_000_8555, w_000_8556, w_000_8557, w_000_8558, w_000_8559, w_000_8560, w_000_8561, w_000_8562, w_000_8563, w_000_8564, w_000_8565, w_000_8566, w_000_8567, w_000_8568, w_000_8569, w_000_8570, w_000_8571, w_000_8572, w_000_8573, w_000_8574, w_000_8575, w_000_8576, w_000_8577, w_000_8578, w_000_8579, w_000_8580, w_000_8581, w_000_8582, w_000_8583, w_000_8584, w_000_8585, w_000_8586, w_000_8587, w_000_8588, w_000_8589, w_000_8590, w_000_8591, w_000_8592, w_000_8593, w_000_8594, w_000_8595, w_000_8596, w_000_8597, w_000_8598, w_000_8599, w_000_8600, w_000_8601, w_000_8602, w_000_8603, w_000_8604, w_000_8605, w_000_8606, w_000_8607, w_000_8608, w_000_8609, w_000_8610, w_000_8611, w_000_8612, w_000_8613, w_000_8614, w_000_8615, w_000_8616, w_000_8617, w_000_8618, w_000_8619, w_000_8620, w_000_8621, w_000_8622, w_000_8623, w_000_8624, w_000_8625, w_000_8626, w_000_8627, w_000_8628, w_000_8629, w_000_8630, w_000_8631, w_000_8632, w_000_8633, w_000_8634, w_000_8635, w_000_8636, w_000_8637, w_000_8638, w_000_8639, w_000_8640, w_000_8641, w_000_8642, w_000_8643, w_000_8644, w_000_8645, w_000_8646, w_000_8647, w_000_8648, w_000_8649, w_000_8650, w_000_8651, w_000_8652, w_000_8653, w_000_8654, w_000_8655, w_000_8656, w_000_8657, w_000_8658, w_000_8659, w_000_8660, w_000_8661, w_000_8662, w_000_8663, w_000_8664, w_000_8665, w_000_8666, w_000_8667, w_000_8668, w_000_8669, w_000_8670, w_000_8671, w_000_8672, w_000_8673, w_000_8674, w_000_8675, w_000_8676, w_000_8677, w_000_8678, w_000_8679, w_000_8680, w_000_8681, w_000_8682, w_000_8683, w_000_8684, w_000_8685, w_000_8686, w_000_8687, w_000_8688, w_000_8689, w_000_8690, w_000_8691, w_000_8692, w_000_8693, w_000_8694, w_000_8695, w_000_8696, w_000_8697, w_000_8698, w_000_8699, w_000_8700, w_000_8701, w_000_8702, w_000_8703, w_000_8704, w_000_8705, w_000_8706, w_000_8707, w_000_8708, w_000_8709, w_000_8710, w_000_8711, w_000_8712, w_000_8713, w_000_8714, w_000_8715, w_000_8716, w_000_8717, w_000_8718, w_000_8719, w_000_8720, w_000_8721, w_000_8722, w_000_8723, w_000_8724, w_000_8725, w_000_8726, w_000_8728, w_000_8729, w_000_8730, w_000_8731, w_000_8732, w_000_8733, w_000_8734, w_000_8735, w_000_8736, w_000_8737, w_000_8738, w_000_8739, w_000_8740, w_000_8741, w_000_8742, w_000_8743, w_000_8744, w_000_8745, w_000_8746, w_000_8747, w_000_8748, w_000_8749, w_000_8751, w_000_8752, w_000_8753, w_000_8754, w_000_8755, w_000_8756, w_000_8757, w_000_8758, w_000_8759, w_000_8760, w_000_8761, w_000_8762, w_000_8763, w_000_8764, w_000_8765, w_000_8766, w_000_8767, w_000_8768, w_000_8769, w_000_8770, w_000_8771, w_000_8772, w_000_8773, w_000_8774, w_000_8775, w_000_8776, w_000_8777, w_000_8778, w_000_8779, w_000_8780, w_000_8781, w_000_8782, w_000_8783, w_000_8784, w_000_8785, w_000_8786, w_000_8787, w_000_8788, w_000_8789, w_000_8790, w_000_8791, w_000_8792, w_000_8793, w_000_8794, w_000_8795, w_000_8796, w_000_8797, w_000_8798, w_000_8799, w_000_8800, w_000_8801, w_000_8802, w_000_8803, w_000_8804, w_000_8805, w_000_8806, w_000_8807, w_000_8808, w_000_8809, w_000_8810, w_000_8811, w_000_8812, w_000_8813, w_000_8814, w_000_8815, w_000_8816, w_000_8817, w_000_8818, w_000_8819, w_000_8820, w_000_8821, w_000_8822, w_000_8823, w_000_8824, w_000_8825, w_000_8826, w_000_8827, w_000_8828, w_000_8829, w_000_8830, w_000_8831, w_000_8832, w_000_8833, w_000_8834, w_000_8835, w_000_8836, w_000_8837, w_000_8838, w_000_8839, w_000_8840, w_000_8841, w_000_8842, w_000_8843, w_000_8844, w_000_8845, w_000_8846, w_000_8848, w_000_8849, w_000_8850, w_000_8851, w_000_8852, w_000_8853, w_000_8854, w_000_8855, w_000_8856, w_000_8857, w_000_8858, w_000_8859, w_000_8860, w_000_8861, w_000_8862, w_000_8863, w_000_8864, w_000_8865, w_000_8866, w_000_8867, w_000_8868, w_000_8869, w_000_8870, w_000_8871, w_000_8872, w_000_8873, w_000_8874, w_000_8875, w_000_8876, w_000_8877, w_000_8878, w_000_8879, w_000_8880, w_000_8881, w_000_8882, w_000_8883, w_000_8884, w_000_8885, w_000_8886, w_000_8887, w_000_8888, w_000_8889, w_000_8891, w_000_8892, w_000_8893, w_000_8894, w_000_8895, w_000_8896, w_000_8897, w_000_8898, w_000_8899, w_000_8900, w_000_8901, w_000_8902, w_000_8903, w_000_8904, w_000_8905, w_000_8906, w_000_8907, w_000_8908, w_000_8909, w_000_8910, w_000_8911, w_000_8912, w_000_8913, w_000_8914, w_000_8916, w_000_8917, w_000_8918, w_000_8919, w_000_8920, w_000_8921, w_000_8922, w_000_8923, w_000_8924, w_000_8925, w_000_8926, w_000_8927, w_000_8928, w_000_8929, w_000_8930, w_000_8931, w_000_8932, w_000_8933, w_000_8934, w_000_8935, w_000_8936, w_000_8937, w_000_8938, w_000_8939, w_000_8940, w_000_8941, w_000_8942, w_000_8943, w_000_8944, w_000_8945, w_000_8946, w_000_8947, w_000_8948, w_000_8949, w_000_8950, w_000_8951, w_000_8952, w_000_8953, w_000_8954, w_000_8955, w_000_8956, w_000_8957, w_000_8958, w_000_8959, w_000_8960, w_000_8961, w_000_8962, w_000_8963, w_000_8964, w_000_8965, w_000_8966, w_000_8967, w_000_8968, w_000_8969, w_000_8970, w_000_8971, w_000_8972, w_000_8973, w_000_8974, w_000_8975, w_000_8976, w_000_8977, w_000_8978, w_000_8979, w_000_8980, w_000_8981, w_000_8982, w_000_8983, w_000_8984, w_000_8985, w_000_8986, w_000_8987, w_000_8988, w_000_8989, w_000_8990, w_000_8991, w_000_8992, w_000_8993, w_000_8994, w_000_8995, w_000_8996, w_000_8997, w_000_8998, w_000_8999, w_000_9000, w_000_9001, w_000_9002, w_000_9003, w_000_9004, w_000_9005, w_000_9006, w_000_9007, w_000_9008, w_000_9009, w_000_9010, w_000_9011, w_000_9012, w_000_9013, w_000_9014, w_000_9015, w_000_9016, w_000_9017, w_000_9018, w_000_9019, w_000_9020, w_000_9021, w_000_9022, w_000_9023, w_000_9024, w_000_9025, w_000_9026, w_000_9027, w_000_9028, w_000_9029, w_000_9030, w_000_9031, w_000_9032, w_000_9033, w_000_9034, w_000_9035, w_000_9036, w_000_9037, w_000_9038, w_000_9039, w_000_9040, w_000_9041, w_000_9042, w_000_9043, w_000_9044, w_000_9045, w_000_9046, w_000_9047, w_000_9048, w_000_9049, w_000_9050, w_000_9051, w_000_9052, w_000_9053, w_000_9054, w_000_9055, w_000_9056, w_000_9057, w_000_9058, w_000_9059, w_000_9060, w_000_9061, w_000_9062, w_000_9063, w_000_9064, w_000_9065, w_000_9066, w_000_9067, w_000_9068, w_000_9069, w_000_9070, w_000_9071, w_000_9072, w_000_9073, w_000_9074, w_000_9075, w_000_9076, w_000_9077, w_000_9078, w_000_9079, w_000_9080, w_000_9081, w_000_9082, w_000_9083, w_000_9084, w_000_9085, w_000_9086, w_000_9087, w_000_9088, w_000_9089, w_000_9090, w_000_9091, w_000_9092, w_000_9093, w_000_9094, w_000_9095, w_000_9096, w_000_9097, w_000_9098, w_000_9099, w_000_9100, w_000_9101, w_000_9102, w_000_9103, w_000_9104, w_000_9105, w_000_9106, w_000_9107, w_000_9108, w_000_9109, w_000_9110, w_000_9111, w_000_9112, w_000_9113, w_000_9114, w_000_9115, w_000_9116, w_000_9117, w_000_9118, w_000_9119, w_000_9120, w_000_9121, w_000_9122, w_000_9123, w_000_9124, w_000_9125, w_000_9126, w_000_9127, w_000_9128, w_000_9129, w_000_9130, w_000_9131, w_000_9132, w_000_9133, w_000_9134, w_000_9135, w_000_9136, w_000_9137, w_000_9138, w_000_9139, w_000_9140, w_000_9141, w_000_9142, w_000_9143, w_000_9144, w_000_9145, w_000_9146, w_000_9147, w_000_9148, w_000_9149, w_000_9150, w_000_9151, w_000_9152, w_000_9153, w_000_9154, w_000_9155, w_000_9156, w_000_9157, w_000_9158, w_000_9159, w_000_9160, w_000_9161, w_000_9162, w_000_9163, w_000_9164, w_000_9165, w_000_9166, w_000_9167, w_000_9168, w_000_9169, w_000_9170, w_000_9171, w_000_9172, w_000_9173, w_000_9174, w_000_9175, w_000_9176, w_000_9177, w_000_9178, w_000_9179, w_000_9180, w_000_9181, w_000_9182, w_000_9183, w_000_9184, w_000_9185, w_000_9186, w_000_9187, w_000_9188, w_000_9189, w_000_9190, w_000_9191, w_000_9192, w_000_9193, w_000_9194, w_000_9195, w_000_9196, w_000_9197, w_000_9198, w_000_9199, w_000_9200, w_000_9201, w_000_9202, w_000_9203, w_000_9204, w_000_9205, w_000_9206, w_000_9207, w_000_9208, w_000_9209, w_000_9210, w_000_9211, w_000_9212, w_000_9213, w_000_9214, w_000_9215, w_000_9216, w_000_9217, w_000_9218, w_000_9219, w_000_9220, w_000_9221, w_000_9222, w_000_9223, w_000_9224, w_000_9225, w_000_9226, w_000_9227, w_000_9228, w_000_9229, w_000_9230, w_000_9231, w_000_9232, w_000_9233, w_000_9234, w_000_9235, w_000_9236, w_000_9237, w_000_9238, w_000_9239, w_000_9240, w_000_9241, w_000_9242, w_000_9243, w_000_9244, w_000_9245, w_000_9246, w_000_9247, w_000_9248, w_000_9249, w_000_9250, w_000_9251, w_000_9252, w_000_9253, w_000_9254, w_000_9255, w_000_9256, w_000_9257, w_000_9258, w_000_9259, w_000_9260, w_000_9261, w_000_9262, w_000_9263, w_000_9264, w_000_9265, w_000_9266, w_000_9267, w_000_9268, w_000_9269, w_000_9270, w_000_9271, w_000_9272, w_000_9273, w_000_9274, w_000_9275, w_000_9276, w_000_9277, w_000_9278, w_000_9279, w_000_9280, w_000_9281, w_000_9282, w_000_9283, w_000_9284, w_000_9285, w_000_9286, w_000_9287, w_000_9288, w_000_9289, w_000_9290, w_000_9291, w_000_9292, w_000_9293, w_000_9294, w_000_9295, w_000_9296, w_000_9297, w_000_9298, w_000_9299, w_000_9300, w_000_9301, w_000_9302, w_000_9303, w_000_9304, w_000_9305, w_000_9306, w_000_9307, w_000_9308, w_000_9309, w_000_9310, w_000_9311, w_000_9312, w_000_9313, w_000_9314, w_000_9315, w_000_9316, w_000_9317, w_000_9318, w_000_9319, w_000_9320, w_000_9321, w_000_9322, w_000_9323, w_000_9324, w_000_9325, w_000_9326, w_000_9327, w_000_9328, w_000_9329, w_000_9330, w_000_9331, w_000_9332, w_000_9333, w_000_9334, w_000_9335, w_000_9336, w_000_9337, w_000_9338, w_000_9339, w_000_9340, w_000_9341, w_000_9342, w_000_9343, w_000_9344, w_000_9345, w_000_9346, w_000_9347, w_000_9348, w_000_9349, w_000_9350, w_000_9351, w_000_9352, w_000_9353, w_000_9354, w_000_9355, w_000_9356, w_000_9357, w_000_9358, w_000_9359, w_000_9360, w_000_9361, w_000_9362, w_000_9363, w_000_9364, w_000_9365, w_000_9366, w_000_9367, w_000_9368, w_000_9369, w_000_9370, w_000_9371, w_000_9372, w_000_9373, w_000_9374, w_000_9375, w_000_9376, w_000_9377, w_000_9378, w_000_9379, w_000_9380, w_000_9381, w_000_9382, w_000_9383, w_000_9384, w_000_9385, w_000_9386, w_000_9387, w_000_9388, w_000_9389, w_000_9390, w_000_9391, w_000_9392, w_000_9393, w_000_9394, w_000_9395, w_000_9396, w_000_9397, w_000_9398, w_000_9399, w_000_9400, w_000_9401, w_000_9402, w_000_9403, w_000_9404, w_000_9405, w_000_9406, w_000_9407, w_000_9408, w_000_9409, w_000_9410, w_000_9411, w_000_9412, w_000_9413, w_000_9414, w_000_9415, w_000_9416, w_000_9417, w_000_9418, w_000_9419, w_000_9420, w_000_9421, w_000_9422, w_000_9423, w_000_9424, w_000_9425, w_000_9426, w_000_9427, w_000_9428, w_000_9429, w_000_9430, w_000_9431, w_000_9432, w_000_9433, w_000_9434, w_000_9435, w_000_9436, w_000_9437, w_000_9438, w_000_9439, w_000_9440, w_000_9441, w_000_9442, w_000_9443, w_000_9444, w_000_9445, w_000_9446, w_000_9447, w_000_9448, w_000_9449, w_000_9450, w_000_9451, w_000_9452, w_000_9453, w_000_9454, w_000_9455, w_000_9456, w_000_9457, w_000_9458, w_000_9459, w_000_9460, w_000_9461, w_000_9462, w_000_9463, w_000_9464, w_000_9465, w_000_9466, w_000_9467, w_000_9468, w_000_9469, w_000_9470, w_000_9471, w_000_9472, w_000_9473, w_000_9474, w_000_9475, w_000_9476, w_000_9477, w_000_9478, w_000_9479, w_000_9480, w_000_9481, w_000_9482, w_000_9483, w_000_9484, w_000_9485, w_000_9486, w_000_9487, w_000_9488, w_000_9489, w_000_9490, w_000_9491, w_000_9492, w_000_9493, w_000_9494, w_000_9495, w_000_9496, w_000_9497, w_000_9498, w_000_9499, w_000_9500, w_000_9501, w_000_9502, w_000_9504, w_000_9505, w_000_9506, w_000_9507, w_000_9508, w_000_9509, w_000_9510, w_000_9511, w_000_9512, w_000_9513, w_000_9514, w_000_9515, w_000_9516, w_000_9517, w_000_9518, w_000_9519, w_000_9520, w_000_9521, w_000_9522, w_000_9523, w_000_9524, w_000_9525, w_000_9526, w_000_9527, w_000_9528, w_000_9529, w_000_9530, w_000_9531, w_000_9532, w_000_9533, w_000_9534, w_000_9535, w_000_9536, w_000_9537, w_000_9538, w_000_9539, w_000_9540, w_000_9541, w_000_9542, w_000_9543, w_000_9544, w_000_9545, w_000_9547, w_000_9548, w_000_9549, w_000_9550, w_000_9551, w_000_9552, w_000_9554, w_000_9555, w_000_9556, w_000_9557, w_000_9558, w_000_9559, w_000_9560, w_000_9561, w_000_9563, w_000_9564, w_000_9565, w_000_9566, w_000_9567, w_000_9569, w_000_9570, w_000_9571, w_000_9572, w_000_9573, w_000_9574, w_000_9575, w_000_9576, w_000_9577, w_000_9578, w_000_9579, w_000_9580, w_000_9581, w_000_9582, w_000_9583, w_000_9584, w_000_9585, w_000_9586, w_000_9587, w_000_9588, w_000_9589, w_000_9590, w_000_9591, w_000_9592, w_000_9593, w_000_9594, w_000_9595, w_000_9596, w_000_9597, w_000_9598, w_000_9599, w_000_9600, w_000_9601, w_000_9602, w_000_9603, w_000_9604, w_000_9605, w_000_9606, w_000_9607, w_000_9608, w_000_9609, w_000_9610, w_000_9611, w_000_9612, w_000_9613, w_000_9614, w_000_9615, w_000_9616, w_000_9617, w_000_9618, w_000_9619, w_000_9620, w_000_9621, w_000_9622, w_000_9623, w_000_9624, w_000_9625, w_000_9626, w_000_9627, w_000_9628, w_000_9629, w_000_9630, w_000_9632, w_000_9633, w_000_9634, w_000_9635, w_000_9636, w_000_9637, w_000_9639, w_000_9640, w_000_9641, w_000_9642, w_000_9643, w_000_9644, w_000_9646, w_000_9647, w_000_9648, w_000_9649, w_000_9650, w_000_9651, w_000_9652, w_000_9653, w_000_9654, w_000_9655, w_000_9656, w_000_9657, w_000_9658, w_000_9659, w_000_9660, w_000_9661, w_000_9662, w_000_9663, w_000_9664, w_000_9666, w_000_9667, w_000_9668, w_000_9669, w_000_9670, w_000_9671, w_000_9672, w_000_9673, w_000_9674, w_000_9675, w_000_9676, w_000_9677, w_000_9678, w_000_9679, w_000_9682, w_000_9683, w_000_9684, w_000_9685, w_000_9686, w_000_9687, w_000_9688, w_000_9689, w_000_9690, w_000_9691, w_000_9692, w_000_9693, w_000_9694, w_000_9695, w_000_9696, w_000_9697, w_000_9698, w_000_9699, w_000_9701, w_000_9702, w_000_9704, w_000_9706, w_000_9708, w_000_9709, w_000_9710, w_000_9711, w_000_9713, w_000_9715, w_000_9716, w_000_9717, w_000_9719, w_000_9720, w_000_9721, w_000_9723, w_000_9725, w_000_9727, w_000_9728, w_000_9729, w_000_9730, w_000_9731, w_000_9732, w_000_9733, w_000_9734, w_000_9735, w_000_9736, w_000_9737, w_000_9738, w_000_9739, w_000_9740, w_000_9741, w_000_9742, w_000_9743, w_000_9744, w_000_9745, w_000_9747, w_000_9748, w_000_9749, w_000_9750, w_000_9752, w_000_9753, w_000_9754, w_000_9755, w_000_9756, w_000_9757, w_000_9758, w_000_9759, w_000_9760, w_000_9761, w_000_9765, w_000_9766, w_000_9767, w_000_9769, w_000_9770, w_000_9771, w_000_9772, w_000_9774, w_000_9776, w_000_9777, w_000_9778, w_000_9779, w_000_9780, w_000_9781, w_000_9782, w_000_9783, w_000_9785, w_000_9786, w_000_9788, w_000_9789, w_000_9790, w_000_9791, w_000_9792, w_000_9793, w_000_9794, w_000_9795, w_000_9796, w_000_9797, w_000_9798, w_000_9799, w_000_9800, w_000_9801, w_000_9802, w_000_9803, w_000_9804, w_000_9805, w_000_9806, w_000_9807, w_000_9808, w_000_9809, w_000_9810, w_000_9811, w_000_9812, w_000_9813, w_000_9814, w_000_9815, w_000_9816, w_000_9817, w_000_9819, w_000_9820, w_000_9821, w_000_9822, w_000_9823, w_000_9824, w_000_9825, w_000_9826, w_000_9827, w_000_9828, w_000_9829, w_000_9830, w_000_9831, w_000_9832, w_000_9833, w_000_9834, w_000_9835, w_000_9837, w_000_9838, w_000_9841, w_000_9842, w_000_9843, w_000_9844, w_000_9846, w_000_9847, w_000_9848, w_000_9849, w_000_9851, w_000_9853, w_000_9854, w_000_9855, w_000_9856, w_000_9857, w_000_9858, w_000_9859, w_000_9860, w_000_9861, w_000_9862, w_000_9864, w_000_9865, w_000_9866, w_000_9867, w_000_9871, w_000_9872, w_000_9874, w_000_9875, w_000_9877, w_000_9878, w_000_9879, w_000_9880, w_000_9882, w_000_9884, w_000_9887, w_000_9889, w_000_9890, w_000_9892, w_000_9893, w_000_9894, w_000_9895, w_000_9896, w_000_9897, w_000_9898, w_000_9899, w_000_9900, w_000_9902, w_000_9904, w_000_9905, w_000_9907, w_000_9908, w_000_9910, w_000_9914, w_000_9920, w_000_9922, w_000_9925, w_000_9926, w_000_9929, w_000_9930, w_000_9934, w_000_9936, w_000_9937, w_000_9938, w_000_9941, w_000_9949, w_000_9951, w_000_9958, w_000_9970, w_000_9978, w_000_9985, w_000_9996;
  wire w_001_000, w_001_001, w_001_002, w_001_003, w_001_004, w_001_005, w_001_006, w_001_007, w_001_008, w_001_009, w_001_010, w_001_011, w_001_012, w_001_013, w_001_014, w_001_015, w_001_016, w_001_017, w_001_018, w_001_019, w_001_020, w_001_021, w_001_022, w_001_023, w_001_024, w_001_025, w_001_026, w_001_027, w_001_028, w_001_029, w_001_030, w_001_031, w_001_032, w_001_033, w_001_034, w_001_035, w_001_036, w_001_037, w_001_038, w_001_039, w_001_040, w_001_041, w_001_042, w_001_043, w_001_044, w_001_045, w_001_046, w_001_047, w_001_048, w_001_049, w_001_050, w_001_051, w_001_052, w_001_053, w_001_054, w_001_055, w_001_056, w_001_057, w_001_058, w_001_059, w_001_060, w_001_061, w_001_062, w_001_063, w_001_064, w_001_065, w_001_066, w_001_067, w_001_068, w_001_069, w_001_070, w_001_071, w_001_072, w_001_073, w_001_074, w_001_075, w_001_076, w_001_077, w_001_078, w_001_079, w_001_080, w_001_081, w_001_082, w_001_083, w_001_084, w_001_085, w_001_086, w_001_087, w_001_088, w_001_089, w_001_090, w_001_091, w_001_092, w_001_093, w_001_094, w_001_095, w_001_096, w_001_097, w_001_098, w_001_099, w_001_100, w_001_101, w_001_102, w_001_103, w_001_104, w_001_105, w_001_106, w_001_107, w_001_108, w_001_109, w_001_110, w_001_111, w_001_112, w_001_113, w_001_114, w_001_115, w_001_116, w_001_117, w_001_118, w_001_119, w_001_120, w_001_121, w_001_122, w_001_123, w_001_124, w_001_125, w_001_126, w_001_127, w_001_128, w_001_129, w_001_130, w_001_131, w_001_132, w_001_133, w_001_134, w_001_135, w_001_136, w_001_137, w_001_138, w_001_139, w_001_140, w_001_141, w_001_142, w_001_143, w_001_144, w_001_145, w_001_146, w_001_147, w_001_148, w_001_149, w_001_150, w_001_151, w_001_152, w_001_153, w_001_154, w_001_155, w_001_156, w_001_157, w_001_158, w_001_159, w_001_160, w_001_161, w_001_162, w_001_163, w_001_164, w_001_165, w_001_166, w_001_167, w_001_168, w_001_169, w_001_170, w_001_171, w_001_172, w_001_173, w_001_174, w_001_175, w_001_176, w_001_177, w_001_178, w_001_179, w_001_180, w_001_181, w_001_182, w_001_183, w_001_184, w_001_185, w_001_186, w_001_187, w_001_188, w_001_189, w_001_190, w_001_191, w_001_192, w_001_193, w_001_194, w_001_195, w_001_196, w_001_197, w_001_198, w_001_199, w_001_200, w_001_201, w_001_202, w_001_203, w_001_204, w_001_205, w_001_206, w_001_207, w_001_208, w_001_209, w_001_210, w_001_211, w_001_212, w_001_213, w_001_214, w_001_215, w_001_216, w_001_217, w_001_218, w_001_219, w_001_220, w_001_221, w_001_222, w_001_223, w_001_224, w_001_225, w_001_226, w_001_227, w_001_228, w_001_229, w_001_230, w_001_231, w_001_232, w_001_233, w_001_234, w_001_235, w_001_236, w_001_237, w_001_238, w_001_239, w_001_240, w_001_241, w_001_242, w_001_243, w_001_244, w_001_245, w_001_246, w_001_247, w_001_248, w_001_249, w_001_250, w_001_251, w_001_252, w_001_253, w_001_254, w_001_255, w_001_256, w_001_257, w_001_258, w_001_259, w_001_260, w_001_261, w_001_262, w_001_263, w_001_264, w_001_265, w_001_266, w_001_267, w_001_268, w_001_269, w_001_270, w_001_271, w_001_272, w_001_273, w_001_274, w_001_275, w_001_276, w_001_277, w_001_278, w_001_279, w_001_280, w_001_281, w_001_282, w_001_283, w_001_284, w_001_285, w_001_286, w_001_287, w_001_288, w_001_289, w_001_290, w_001_291, w_001_292, w_001_293, w_001_294, w_001_295, w_001_296, w_001_297, w_001_298, w_001_299, w_001_300, w_001_301, w_001_302, w_001_303, w_001_304, w_001_305, w_001_306, w_001_307, w_001_308, w_001_309, w_001_310, w_001_311, w_001_312, w_001_313, w_001_314, w_001_315, w_001_316, w_001_317, w_001_318, w_001_319, w_001_320, w_001_321, w_001_322, w_001_323, w_001_324, w_001_325, w_001_326, w_001_327, w_001_328, w_001_329, w_001_330, w_001_331, w_001_332, w_001_333, w_001_334, w_001_335, w_001_336, w_001_337, w_001_338, w_001_339, w_001_340, w_001_341, w_001_342, w_001_343, w_001_344, w_001_345, w_001_346, w_001_347, w_001_348, w_001_349, w_001_350, w_001_351, w_001_352, w_001_353, w_001_354, w_001_355, w_001_356, w_001_357, w_001_358, w_001_359, w_001_360, w_001_361, w_001_362, w_001_363, w_001_364, w_001_365, w_001_366, w_001_367, w_001_368, w_001_369, w_001_370, w_001_371, w_001_372, w_001_373, w_001_374, w_001_375, w_001_376, w_001_377, w_001_378, w_001_379, w_001_380, w_001_381, w_001_382, w_001_383, w_001_384, w_001_385, w_001_386, w_001_387, w_001_388, w_001_389, w_001_390, w_001_391, w_001_392, w_001_393, w_001_394, w_001_395, w_001_396, w_001_397, w_001_398, w_001_399, w_001_400, w_001_401, w_001_402, w_001_403, w_001_404, w_001_405, w_001_406, w_001_407, w_001_408, w_001_409, w_001_410, w_001_411, w_001_412, w_001_413, w_001_414, w_001_415, w_001_416, w_001_417, w_001_418, w_001_419, w_001_420, w_001_421, w_001_422, w_001_423, w_001_424, w_001_425, w_001_426, w_001_427, w_001_428, w_001_429, w_001_430, w_001_431, w_001_432, w_001_433, w_001_434, w_001_435, w_001_436, w_001_437, w_001_438, w_001_439, w_001_440, w_001_441, w_001_442, w_001_443, w_001_444, w_001_445, w_001_446, w_001_447, w_001_448, w_001_449, w_001_450, w_001_451, w_001_452, w_001_453, w_001_454, w_001_455, w_001_456, w_001_457, w_001_458, w_001_459, w_001_460, w_001_461, w_001_462, w_001_463, w_001_464, w_001_465, w_001_466, w_001_467, w_001_468, w_001_469, w_001_470, w_001_471, w_001_472, w_001_473, w_001_474, w_001_475, w_001_476, w_001_477, w_001_478, w_001_479, w_001_480, w_001_481, w_001_482, w_001_483, w_001_484, w_001_485, w_001_486, w_001_487, w_001_488, w_001_489, w_001_490, w_001_491, w_001_492, w_001_493, w_001_494, w_001_495, w_001_496, w_001_497, w_001_498, w_001_499, w_001_500, w_001_501, w_001_502, w_001_503, w_001_504, w_001_505, w_001_506, w_001_507, w_001_508, w_001_509, w_001_510, w_001_511, w_001_512, w_001_513, w_001_514, w_001_515, w_001_516, w_001_517, w_001_518, w_001_519, w_001_520, w_001_521, w_001_522, w_001_523, w_001_524, w_001_525, w_001_526, w_001_527, w_001_528, w_001_529, w_001_530, w_001_531, w_001_532, w_001_533, w_001_534, w_001_535, w_001_536, w_001_537, w_001_538, w_001_539, w_001_540, w_001_541, w_001_542, w_001_543, w_001_544, w_001_545, w_001_546, w_001_547, w_001_548, w_001_549, w_001_550, w_001_551, w_001_552, w_001_553, w_001_554, w_001_555, w_001_556, w_001_557, w_001_558, w_001_559, w_001_560, w_001_561, w_001_562, w_001_563, w_001_564, w_001_565, w_001_566, w_001_567, w_001_568, w_001_569, w_001_570, w_001_571, w_001_572, w_001_573, w_001_574, w_001_575, w_001_576, w_001_577, w_001_578, w_001_579, w_001_580, w_001_581, w_001_582, w_001_583, w_001_584, w_001_585, w_001_586, w_001_587, w_001_588, w_001_589, w_001_590, w_001_591, w_001_592, w_001_593, w_001_594, w_001_595, w_001_596, w_001_597, w_001_598, w_001_599, w_001_600, w_001_601, w_001_602, w_001_603, w_001_604, w_001_605, w_001_606, w_001_607, w_001_608, w_001_609, w_001_610, w_001_611, w_001_612, w_001_613, w_001_614, w_001_615, w_001_616, w_001_617, w_001_618, w_001_619, w_001_620, w_001_621, w_001_622, w_001_623, w_001_624, w_001_625, w_001_626, w_001_627, w_001_628, w_001_629, w_001_630, w_001_631, w_001_632, w_001_633, w_001_634, w_001_635, w_001_636, w_001_637, w_001_638, w_001_639, w_001_640, w_001_641, w_001_642, w_001_643, w_001_644, w_001_645, w_001_646, w_001_647, w_001_648, w_001_649, w_001_650, w_001_651, w_001_652, w_001_653, w_001_654, w_001_655, w_001_656, w_001_657, w_001_658, w_001_659, w_001_660, w_001_661, w_001_662, w_001_663, w_001_664, w_001_665, w_001_667, w_001_668, w_001_669, w_001_670, w_001_671, w_001_672, w_001_673, w_001_674, w_001_675, w_001_676, w_001_677, w_001_678, w_001_679, w_001_680, w_001_681, w_001_682, w_001_683, w_001_684, w_001_685, w_001_686, w_001_687, w_001_688, w_001_689, w_001_690, w_001_691, w_001_692, w_001_693, w_001_694, w_001_695, w_001_696, w_001_697, w_001_698, w_001_699, w_001_700, w_001_701, w_001_702, w_001_703, w_001_704, w_001_705, w_001_706, w_001_707, w_001_708, w_001_709, w_001_710, w_001_711, w_001_712, w_001_713, w_001_714, w_001_715, w_001_716, w_001_717, w_001_718, w_001_719, w_001_720, w_001_721, w_001_722, w_001_723, w_001_724, w_001_725, w_001_726, w_001_727, w_001_728, w_001_729, w_001_730, w_001_731, w_001_732, w_001_733, w_001_734, w_001_735, w_001_736, w_001_737, w_001_738, w_001_739, w_001_740, w_001_741, w_001_742, w_001_743, w_001_744, w_001_745, w_001_746, w_001_747, w_001_748, w_001_749, w_001_750, w_001_751, w_001_752, w_001_753, w_001_754, w_001_755, w_001_756, w_001_757, w_001_758, w_001_759, w_001_760, w_001_761, w_001_762, w_001_763, w_001_764, w_001_765, w_001_766, w_001_767, w_001_768, w_001_769, w_001_770, w_001_771, w_001_772, w_001_773, w_001_774, w_001_775, w_001_776, w_001_777, w_001_778, w_001_779, w_001_780, w_001_781, w_001_782, w_001_783, w_001_784, w_001_785, w_001_786, w_001_787, w_001_788, w_001_789, w_001_790, w_001_791, w_001_792, w_001_793, w_001_794, w_001_795, w_001_796, w_001_797, w_001_798, w_001_799, w_001_800, w_001_801, w_001_802, w_001_803, w_001_804, w_001_805, w_001_806, w_001_807, w_001_808, w_001_809, w_001_810, w_001_811, w_001_812, w_001_813, w_001_814, w_001_815, w_001_816, w_001_817, w_001_818, w_001_819, w_001_820, w_001_821, w_001_822, w_001_823, w_001_824, w_001_825, w_001_826, w_001_827, w_001_828, w_001_829, w_001_830, w_001_831, w_001_832, w_001_833, w_001_834, w_001_835, w_001_836, w_001_837, w_001_838, w_001_839, w_001_840, w_001_841, w_001_842, w_001_843, w_001_844, w_001_845, w_001_846, w_001_847, w_001_848, w_001_849, w_001_850, w_001_851, w_001_852, w_001_853, w_001_854, w_001_855, w_001_856, w_001_857, w_001_858, w_001_859, w_001_860, w_001_861, w_001_862, w_001_863, w_001_864, w_001_865, w_001_866, w_001_867, w_001_868, w_001_869, w_001_870, w_001_871, w_001_872, w_001_873, w_001_874, w_001_875, w_001_876, w_001_877, w_001_878, w_001_879, w_001_880, w_001_881, w_001_882, w_001_883, w_001_884, w_001_885, w_001_886, w_001_887, w_001_888, w_001_889, w_001_890, w_001_891, w_001_892, w_001_893, w_001_894, w_001_895, w_001_896, w_001_897, w_001_898, w_001_899, w_001_900, w_001_901, w_001_902, w_001_903, w_001_904, w_001_905, w_001_906, w_001_907, w_001_908, w_001_909, w_001_910, w_001_912, w_001_913, w_001_914, w_001_915, w_001_916, w_001_917, w_001_918, w_001_919, w_001_920, w_001_921, w_001_922, w_001_923, w_001_924, w_001_925, w_001_926, w_001_927, w_001_928, w_001_930, w_001_931, w_001_932, w_001_933, w_001_934, w_001_935, w_001_936, w_001_937, w_001_938, w_001_939, w_001_940, w_001_941, w_001_942, w_001_943, w_001_944, w_001_945, w_001_946, w_001_947, w_001_948, w_001_949, w_001_950, w_001_951, w_001_952, w_001_953, w_001_954, w_001_955, w_001_956, w_001_957, w_001_958, w_001_959, w_001_960, w_001_961, w_001_962, w_001_963, w_001_964, w_001_965, w_001_966, w_001_967, w_001_968, w_001_969, w_001_970, w_001_971, w_001_972, w_001_973, w_001_974, w_001_975, w_001_976, w_001_977, w_001_978, w_001_979, w_001_980, w_001_981, w_001_982, w_001_983, w_001_984, w_001_985, w_001_986, w_001_987, w_001_988, w_001_989, w_001_990, w_001_991, w_001_992, w_001_993, w_001_994, w_001_995, w_001_996, w_001_997, w_001_998, w_001_999, w_001_1000, w_001_1001, w_001_1002, w_001_1003, w_001_1004, w_001_1005, w_001_1006, w_001_1007, w_001_1008, w_001_1009, w_001_1010, w_001_1011, w_001_1012, w_001_1013, w_001_1014, w_001_1015, w_001_1016, w_001_1017, w_001_1018, w_001_1019, w_001_1020, w_001_1021, w_001_1022, w_001_1023, w_001_1024, w_001_1025, w_001_1026, w_001_1027, w_001_1028, w_001_1029, w_001_1030, w_001_1031, w_001_1032, w_001_1033, w_001_1034, w_001_1035, w_001_1036, w_001_1037, w_001_1038, w_001_1039, w_001_1040, w_001_1041, w_001_1042, w_001_1043, w_001_1044, w_001_1045, w_001_1046, w_001_1047, w_001_1048, w_001_1049, w_001_1050, w_001_1051, w_001_1052, w_001_1053, w_001_1054, w_001_1055, w_001_1056, w_001_1057, w_001_1058, w_001_1059, w_001_1060, w_001_1061, w_001_1062, w_001_1063, w_001_1064, w_001_1065, w_001_1066, w_001_1067, w_001_1068, w_001_1069, w_001_1070, w_001_1071, w_001_1072, w_001_1073, w_001_1074, w_001_1075, w_001_1077, w_001_1078, w_001_1079, w_001_1082, w_001_1083, w_001_1084, w_001_1085, w_001_1086, w_001_1087, w_001_1088, w_001_1089, w_001_1090, w_001_1091, w_001_1092, w_001_1093, w_001_1095, w_001_1097, w_001_1098, w_001_1099, w_001_1100, w_001_1101, w_001_1102, w_001_1103, w_001_1104, w_001_1106, w_001_1107, w_001_1108, w_001_1109, w_001_1110, w_001_1111, w_001_1112, w_001_1113, w_001_1114, w_001_1115, w_001_1117, w_001_1118, w_001_1119, w_001_1120, w_001_1121, w_001_1122, w_001_1123, w_001_1124, w_001_1125, w_001_1127, w_001_1128, w_001_1129, w_001_1130, w_001_1131, w_001_1132, w_001_1133, w_001_1134, w_001_1135, w_001_1136, w_001_1137, w_001_1138, w_001_1139, w_001_1140, w_001_1141, w_001_1142, w_001_1143, w_001_1144, w_001_1145, w_001_1146, w_001_1147, w_001_1148, w_001_1149, w_001_1152, w_001_1153, w_001_1154, w_001_1155, w_001_1156, w_001_1157, w_001_1158, w_001_1159, w_001_1160, w_001_1161, w_001_1162, w_001_1163, w_001_1164, w_001_1165, w_001_1166, w_001_1167, w_001_1168, w_001_1169, w_001_1170, w_001_1171, w_001_1172, w_001_1173, w_001_1174, w_001_1175, w_001_1176, w_001_1177, w_001_1178, w_001_1179, w_001_1180, w_001_1181, w_001_1182, w_001_1183, w_001_1184, w_001_1185, w_001_1186, w_001_1187, w_001_1188, w_001_1189, w_001_1190, w_001_1191, w_001_1192, w_001_1193, w_001_1194, w_001_1195, w_001_1196, w_001_1198, w_001_1199, w_001_1200, w_001_1201, w_001_1202, w_001_1203, w_001_1204, w_001_1206, w_001_1207, w_001_1208, w_001_1209, w_001_1210, w_001_1211, w_001_1212, w_001_1213, w_001_1214, w_001_1216, w_001_1218, w_001_1219, w_001_1220, w_001_1221, w_001_1222, w_001_1223, w_001_1224, w_001_1225, w_001_1226, w_001_1227, w_001_1228, w_001_1229, w_001_1230, w_001_1232, w_001_1233, w_001_1234, w_001_1235, w_001_1236, w_001_1237, w_001_1238, w_001_1240, w_001_1241, w_001_1242, w_001_1243, w_001_1244, w_001_1245, w_001_1246, w_001_1247, w_001_1249, w_001_1250, w_001_1251, w_001_1252, w_001_1253, w_001_1254, w_001_1256, w_001_1257, w_001_1258, w_001_1259, w_001_1260, w_001_1261, w_001_1262, w_001_1263, w_001_1264, w_001_1265, w_001_1266, w_001_1268, w_001_1269, w_001_1270, w_001_1271, w_001_1272, w_001_1273, w_001_1274, w_001_1275, w_001_1276, w_001_1277, w_001_1278, w_001_1279, w_001_1280, w_001_1281, w_001_1282, w_001_1283, w_001_1284, w_001_1285, w_001_1286, w_001_1287, w_001_1288, w_001_1289, w_001_1290, w_001_1291, w_001_1292, w_001_1293, w_001_1295, w_001_1296, w_001_1297, w_001_1299, w_001_1300, w_001_1301, w_001_1302, w_001_1303, w_001_1304, w_001_1305, w_001_1306, w_001_1307, w_001_1308, w_001_1309, w_001_1310, w_001_1311, w_001_1313, w_001_1314, w_001_1315, w_001_1316, w_001_1317, w_001_1318, w_001_1319, w_001_1320, w_001_1321, w_001_1322, w_001_1323, w_001_1324, w_001_1325, w_001_1327, w_001_1328, w_001_1329, w_001_1330, w_001_1331, w_001_1333, w_001_1334, w_001_1335, w_001_1336, w_001_1337, w_001_1338, w_001_1339, w_001_1341, w_001_1342, w_001_1343, w_001_1344, w_001_1345, w_001_1346, w_001_1347, w_001_1348, w_001_1349, w_001_1350, w_001_1351, w_001_1352, w_001_1353, w_001_1354, w_001_1355, w_001_1356, w_001_1357, w_001_1358, w_001_1359, w_001_1360, w_001_1361, w_001_1362, w_001_1363, w_001_1364, w_001_1365, w_001_1366, w_001_1368, w_001_1369, w_001_1370, w_001_1371, w_001_1372, w_001_1373, w_001_1374, w_001_1375, w_001_1376, w_001_1377, w_001_1378, w_001_1379, w_001_1380, w_001_1381, w_001_1382, w_001_1383, w_001_1384, w_001_1385, w_001_1386, w_001_1388, w_001_1389, w_001_1390, w_001_1391, w_001_1392, w_001_1393, w_001_1394, w_001_1395, w_001_1396, w_001_1397, w_001_1398, w_001_1399, w_001_1400, w_001_1402, w_001_1403, w_001_1404, w_001_1405, w_001_1406, w_001_1408, w_001_1409, w_001_1410, w_001_1411, w_001_1412, w_001_1413, w_001_1414, w_001_1415, w_001_1416, w_001_1417, w_001_1418, w_001_1419, w_001_1420, w_001_1421, w_001_1422, w_001_1423, w_001_1424, w_001_1425, w_001_1426, w_001_1427, w_001_1428, w_001_1429, w_001_1430, w_001_1431, w_001_1432, w_001_1433, w_001_1434, w_001_1435, w_001_1436, w_001_1437, w_001_1438, w_001_1439, w_001_1440, w_001_1441, w_001_1443, w_001_1444, w_001_1445, w_001_1446, w_001_1447, w_001_1448, w_001_1449, w_001_1450, w_001_1451, w_001_1452, w_001_1453, w_001_1454, w_001_1455, w_001_1457, w_001_1459, w_001_1460, w_001_1461, w_001_1462, w_001_1463, w_001_1464, w_001_1465, w_001_1466, w_001_1467, w_001_1469, w_001_1470, w_001_1471, w_001_1472, w_001_1473, w_001_1474, w_001_1475, w_001_1476, w_001_1478, w_001_1479, w_001_1480, w_001_1481, w_001_1482, w_001_1483, w_001_1484, w_001_1485, w_001_1486, w_001_1487, w_001_1488, w_001_1489, w_001_1490, w_001_1492, w_001_1493, w_001_1494, w_001_1495, w_001_1496, w_001_1498, w_001_1499, w_001_1500, w_001_1501, w_001_1502, w_001_1503, w_001_1504, w_001_1505, w_001_1506, w_001_1507, w_001_1508, w_001_1509, w_001_1510, w_001_1511, w_001_1512, w_001_1513, w_001_1515, w_001_1516, w_001_1517, w_001_1518, w_001_1519, w_001_1520, w_001_1521, w_001_1522, w_001_1523, w_001_1524, w_001_1525, w_001_1526, w_001_1527, w_001_1528, w_001_1529, w_001_1530, w_001_1531, w_001_1532, w_001_1533, w_001_1534, w_001_1535, w_001_1536, w_001_1537, w_001_1538, w_001_1539, w_001_1540, w_001_1541, w_001_1542, w_001_1543, w_001_1544, w_001_1545, w_001_1546, w_001_1547, w_001_1548, w_001_1549, w_001_1550, w_001_1551, w_001_1552, w_001_1553, w_001_1554, w_001_1555, w_001_1556, w_001_1557, w_001_1558, w_001_1559, w_001_1560, w_001_1561, w_001_1562, w_001_1563, w_001_1564, w_001_1565, w_001_1566, w_001_1567, w_001_1568, w_001_1569, w_001_1570, w_001_1571, w_001_1572, w_001_1573, w_001_1574, w_001_1575, w_001_1576, w_001_1577, w_001_1578, w_001_1579, w_001_1580, w_001_1581, w_001_1582, w_001_1583, w_001_1584, w_001_1585, w_001_1586, w_001_1587, w_001_1588, w_001_1589, w_001_1590, w_001_1591, w_001_1592, w_001_1593, w_001_1595, w_001_1596, w_001_1597, w_001_1598, w_001_1599, w_001_1601, w_001_1602, w_001_1603, w_001_1604, w_001_1605, w_001_1606, w_001_1607, w_001_1608, w_001_1609, w_001_1610, w_001_1611, w_001_1612, w_001_1613, w_001_1614, w_001_1615, w_001_1616, w_001_1617, w_001_1618, w_001_1619, w_001_1620, w_001_1621, w_001_1622, w_001_1623, w_001_1624, w_001_1625, w_001_1626, w_001_1627, w_001_1628, w_001_1629, w_001_1630, w_001_1631, w_001_1632, w_001_1633, w_001_1634, w_001_1635, w_001_1636, w_001_1637, w_001_1638, w_001_1639, w_001_1640, w_001_1641, w_001_1642, w_001_1643, w_001_1644, w_001_1645, w_001_1646, w_001_1647, w_001_1648, w_001_1649, w_001_1650, w_001_1651, w_001_1652, w_001_1653, w_001_1654, w_001_1655, w_001_1656, w_001_1657, w_001_1658, w_001_1659, w_001_1660, w_001_1661, w_001_1662, w_001_1663, w_001_1664, w_001_1665, w_001_1666, w_001_1667, w_001_1668, w_001_1669, w_001_1670, w_001_1671, w_001_1672, w_001_1673, w_001_1674, w_001_1675, w_001_1676, w_001_1677, w_001_1678, w_001_1679, w_001_1681, w_001_1682, w_001_1683, w_001_1684, w_001_1685, w_001_1686, w_001_1687, w_001_1688, w_001_1689, w_001_1690, w_001_1691, w_001_1692, w_001_1693, w_001_1694, w_001_1696, w_001_1697, w_001_1698, w_001_1699, w_001_1700, w_001_1701, w_001_1702, w_001_1703, w_001_1704, w_001_1705, w_001_1706, w_001_1707, w_001_1708, w_001_1709, w_001_1710, w_001_1711, w_001_1712, w_001_1713, w_001_1714, w_001_1715, w_001_1716, w_001_1717, w_001_1718, w_001_1719, w_001_1720, w_001_1721, w_001_1722, w_001_1723, w_001_1724, w_001_1725, w_001_1726, w_001_1727, w_001_1728, w_001_1729, w_001_1730, w_001_1731, w_001_1732, w_001_1733, w_001_1734, w_001_1735, w_001_1736, w_001_1737, w_001_1738, w_001_1740, w_001_1742, w_001_1743, w_001_1745, w_001_1746, w_001_1747, w_001_1748, w_001_1749, w_001_1750, w_001_1751, w_001_1753, w_001_1754, w_001_1755, w_001_1756, w_001_1757, w_001_1758, w_001_1759, w_001_1760, w_001_1761, w_001_1762, w_001_1763, w_001_1764, w_001_1765, w_001_1766, w_001_1767, w_001_1768, w_001_1769, w_001_1770, w_001_1771, w_001_1772, w_001_1773, w_001_1774, w_001_1775, w_001_1776, w_001_1777, w_001_1778, w_001_1779, w_001_1780, w_001_1781, w_001_1782, w_001_1783, w_001_1784, w_001_1785, w_001_1786, w_001_1787, w_001_1788, w_001_1789, w_001_1790, w_001_1791, w_001_1792, w_001_1793, w_001_1795, w_001_1797, w_001_1799, w_001_1800, w_001_1801, w_001_1802, w_001_1803, w_001_1804, w_001_1805, w_001_1806, w_001_1807, w_001_1808, w_001_1809, w_001_1810, w_001_1811, w_001_1812, w_001_1813, w_001_1814, w_001_1815, w_001_1816, w_001_1818, w_001_1819, w_001_1820, w_001_1821, w_001_1822, w_001_1823, w_001_1825, w_001_1826, w_001_1827, w_001_1828, w_001_1829, w_001_1830, w_001_1831, w_001_1832, w_001_1833, w_001_1834, w_001_1835, w_001_1836, w_001_1837, w_001_1839, w_001_1840, w_001_1841, w_001_1843, w_001_1844, w_001_1845, w_001_1846, w_001_1847, w_001_1848, w_001_1849, w_001_1850, w_001_1851, w_001_1852, w_001_1853, w_001_1855, w_001_1856, w_001_1857, w_001_1858, w_001_1859, w_001_1860, w_001_1861, w_001_1862, w_001_1863, w_001_1864, w_001_1865, w_001_1866, w_001_1867, w_001_1868, w_001_1869, w_001_1870, w_001_1872, w_001_1873, w_001_1874, w_001_1875, w_001_1876, w_001_1877, w_001_1878, w_001_1879, w_001_1880, w_001_1881, w_001_1882, w_001_1883, w_001_1884, w_001_1885, w_001_1886, w_001_1888, w_001_1890, w_001_1891, w_001_1892, w_001_1893, w_001_1894, w_001_1895, w_001_1896, w_001_1898, w_001_1899, w_001_1900, w_001_1901, w_001_1902, w_001_1903, w_001_1904, w_001_1905, w_001_1906, w_001_1907, w_001_1909, w_001_1910, w_001_1911, w_001_1912, w_001_1913, w_001_1914, w_001_1915, w_001_1916, w_001_1917, w_001_1918, w_001_1920, w_001_1921, w_001_1922, w_001_1923, w_001_1924, w_001_1925, w_001_1926, w_001_1927, w_001_1928, w_001_1929, w_001_1930, w_001_1931, w_001_1932, w_001_1933, w_001_1934, w_001_1935, w_001_1936, w_001_1937, w_001_1938, w_001_1939, w_001_1940, w_001_1941, w_001_1942, w_001_1943, w_001_1944, w_001_1945, w_001_1947, w_001_1948, w_001_1949, w_001_1950, w_001_1951, w_001_1952, w_001_1953, w_001_1954, w_001_1955, w_001_1956, w_001_1957, w_001_1958, w_001_1959, w_001_1960, w_001_1961, w_001_1962, w_001_1963, w_001_1964, w_001_1965, w_001_1966, w_001_1967, w_001_1968, w_001_1969, w_001_1970, w_001_1971, w_001_1972, w_001_1973, w_001_1974, w_001_1975, w_001_1976, w_001_1977, w_001_1978, w_001_1979, w_001_1980, w_001_1981, w_001_1982, w_001_1983, w_001_1984, w_001_1985, w_001_1986, w_001_1987, w_001_1988, w_001_1989, w_001_1990, w_001_1991, w_001_1992, w_001_1993, w_001_1994, w_001_1995, w_001_1996, w_001_1997, w_001_1998, w_001_1999, w_001_2000, w_001_2001, w_001_2002, w_001_2003, w_001_2004, w_001_2005, w_001_2006, w_001_2007, w_001_2008, w_001_2009, w_001_2010, w_001_2012, w_001_2013, w_001_2014, w_001_2015, w_001_2016, w_001_2017, w_001_2018, w_001_2019, w_001_2020, w_001_2021, w_001_2022, w_001_2023, w_001_2024, w_001_2025, w_001_2026, w_001_2027, w_001_2028, w_001_2029, w_001_2030, w_001_2031, w_001_2032, w_001_2033, w_001_2034, w_001_2035, w_001_2036, w_001_2037, w_001_2038, w_001_2039, w_001_2040, w_001_2041, w_001_2042, w_001_2043, w_001_2044, w_001_2045, w_001_2046, w_001_2047, w_001_2048, w_001_2049, w_001_2050, w_001_2051, w_001_2052, w_001_2053, w_001_2054, w_001_2055, w_001_2056, w_001_2057, w_001_2058, w_001_2060, w_001_2061, w_001_2062, w_001_2064, w_001_2065, w_001_2066, w_001_2068, w_001_2070, w_001_2071, w_001_2072, w_001_2073, w_001_2074, w_001_2075, w_001_2076, w_001_2077, w_001_2078, w_001_2079, w_001_2080, w_001_2081, w_001_2082, w_001_2083, w_001_2084, w_001_2085, w_001_2086, w_001_2087, w_001_2088, w_001_2089, w_001_2090, w_001_2091, w_001_2092, w_001_2093, w_001_2094, w_001_2095, w_001_2096, w_001_2097, w_001_2098, w_001_2099, w_001_2100, w_001_2102, w_001_2103, w_001_2105, w_001_2106, w_001_2107, w_001_2108, w_001_2109, w_001_2110, w_001_2111, w_001_2112, w_001_2113, w_001_2114, w_001_2115, w_001_2116, w_001_2117, w_001_2118, w_001_2121, w_001_2122, w_001_2123, w_001_2124, w_001_2125, w_001_2126, w_001_2127, w_001_2128, w_001_2130, w_001_2131, w_001_2132, w_001_2133, w_001_2134, w_001_2135, w_001_2136, w_001_2137, w_001_2138, w_001_2139, w_001_2140, w_001_2141, w_001_2142, w_001_2143, w_001_2144, w_001_2145, w_001_2146, w_001_2147, w_001_2148, w_001_2149, w_001_2151, w_001_2152, w_001_2153, w_001_2154, w_001_2155, w_001_2156, w_001_2157, w_001_2158, w_001_2159, w_001_2160, w_001_2161, w_001_2162, w_001_2163, w_001_2164, w_001_2165, w_001_2166, w_001_2167, w_001_2168, w_001_2169, w_001_2170, w_001_2171, w_001_2172, w_001_2173, w_001_2174, w_001_2175, w_001_2176, w_001_2177, w_001_2179, w_001_2180, w_001_2181, w_001_2182, w_001_2183, w_001_2184, w_001_2185, w_001_2186, w_001_2187, w_001_2188, w_001_2189, w_001_2190, w_001_2192, w_001_2193, w_001_2194, w_001_2195, w_001_2196, w_001_2197, w_001_2198, w_001_2199, w_001_2200, w_001_2201, w_001_2205, w_001_2206, w_001_2207, w_001_2208, w_001_2209, w_001_2210, w_001_2211, w_001_2212, w_001_2213, w_001_2214, w_001_2215, w_001_2216, w_001_2217, w_001_2218, w_001_2219, w_001_2220, w_001_2221, w_001_2222, w_001_2223, w_001_2224, w_001_2225, w_001_2226, w_001_2227, w_001_2228, w_001_2229, w_001_2230, w_001_2231, w_001_2232, w_001_2233, w_001_2234, w_001_2235, w_001_2236, w_001_2237, w_001_2238, w_001_2239, w_001_2240, w_001_2241, w_001_2242, w_001_2243, w_001_2244, w_001_2245, w_001_2246, w_001_2247, w_001_2248, w_001_2250, w_001_2252, w_001_2253, w_001_2254, w_001_2256, w_001_2257, w_001_2258, w_001_2259, w_001_2260, w_001_2261, w_001_2262, w_001_2263, w_001_2264, w_001_2265, w_001_2266, w_001_2268, w_001_2269, w_001_2270, w_001_2272, w_001_2273, w_001_2274, w_001_2275, w_001_2276, w_001_2277, w_001_2279, w_001_2280, w_001_2281, w_001_2282, w_001_2283, w_001_2284, w_001_2286, w_001_2287, w_001_2288, w_001_2289, w_001_2290, w_001_2291, w_001_2293, w_001_2295, w_001_2296, w_001_2297, w_001_2298, w_001_2299, w_001_2300, w_001_2301, w_001_2302, w_001_2303, w_001_2304, w_001_2305, w_001_2306, w_001_2307, w_001_2309, w_001_2310, w_001_2311, w_001_2312, w_001_2313, w_001_2314, w_001_2315, w_001_2316, w_001_2317, w_001_2318, w_001_2319, w_001_2320, w_001_2321, w_001_2322, w_001_2323, w_001_2324, w_001_2325, w_001_2326, w_001_2327, w_001_2328, w_001_2330, w_001_2331, w_001_2332, w_001_2333, w_001_2334, w_001_2335, w_001_2336, w_001_2337, w_001_2338, w_001_2339, w_001_2340, w_001_2341, w_001_2342, w_001_2343, w_001_2345, w_001_2346, w_001_2347, w_001_2348, w_001_2349, w_001_2350, w_001_2351, w_001_2352, w_001_2353, w_001_2354, w_001_2356, w_001_2357, w_001_2358, w_001_2359, w_001_2360, w_001_2361, w_001_2362, w_001_2363, w_001_2364, w_001_2365, w_001_2366, w_001_2367, w_001_2368, w_001_2369, w_001_2370, w_001_2371, w_001_2372, w_001_2373, w_001_2374, w_001_2375, w_001_2376, w_001_2377, w_001_2378, w_001_2379, w_001_2380, w_001_2381, w_001_2382, w_001_2383, w_001_2384, w_001_2385, w_001_2386, w_001_2387, w_001_2388, w_001_2389, w_001_2390, w_001_2391, w_001_2392, w_001_2393, w_001_2394, w_001_2395, w_001_2396, w_001_2398, w_001_2399, w_001_2401, w_001_2402, w_001_2403, w_001_2405, w_001_2406, w_001_2407, w_001_2408, w_001_2409, w_001_2410, w_001_2411, w_001_2412, w_001_2413, w_001_2414, w_001_2415, w_001_2416, w_001_2418, w_001_2420, w_001_2421, w_001_2422, w_001_2424, w_001_2425, w_001_2426, w_001_2427, w_001_2428, w_001_2429, w_001_2430, w_001_2431, w_001_2432, w_001_2433, w_001_2434, w_001_2435, w_001_2436, w_001_2437, w_001_2438, w_001_2439, w_001_2440, w_001_2441, w_001_2442, w_001_2443, w_001_2444, w_001_2445, w_001_2446, w_001_2447, w_001_2448, w_001_2449, w_001_2450, w_001_2451, w_001_2452, w_001_2453, w_001_2454, w_001_2455, w_001_2456, w_001_2457, w_001_2458, w_001_2459, w_001_2460, w_001_2461, w_001_2462, w_001_2463, w_001_2464, w_001_2465, w_001_2466, w_001_2467, w_001_2468, w_001_2470, w_001_2471, w_001_2472, w_001_2473, w_001_2474, w_001_2476, w_001_2477, w_001_2478, w_001_2479, w_001_2480, w_001_2481, w_001_2482, w_001_2483, w_001_2484, w_001_2485, w_001_2486, w_001_2487, w_001_2488, w_001_2489, w_001_2490, w_001_2491, w_001_2492, w_001_2493, w_001_2494, w_001_2495, w_001_2496, w_001_2497, w_001_2498, w_001_2499, w_001_2500, w_001_2501, w_001_2502, w_001_2503, w_001_2504, w_001_2505, w_001_2506, w_001_2507, w_001_2508, w_001_2509, w_001_2510, w_001_2512, w_001_2513, w_001_2514, w_001_2515, w_001_2516, w_001_2517, w_001_2518, w_001_2519, w_001_2520, w_001_2521, w_001_2522, w_001_2523, w_001_2524, w_001_2525, w_001_2526, w_001_2527, w_001_2528, w_001_2529, w_001_2530, w_001_2531, w_001_2532, w_001_2533, w_001_2535, w_001_2536, w_001_2537, w_001_2538, w_001_2539, w_001_2540, w_001_2541, w_001_2542, w_001_2543, w_001_2544, w_001_2545, w_001_2547, w_001_2548, w_001_2549, w_001_2550, w_001_2551, w_001_2552, w_001_2553, w_001_2554, w_001_2555, w_001_2557, w_001_2558, w_001_2559, w_001_2560, w_001_2561, w_001_2562, w_001_2563, w_001_2564, w_001_2565, w_001_2566, w_001_2567, w_001_2568, w_001_2569, w_001_2570, w_001_2571, w_001_2573, w_001_2575, w_001_2576, w_001_2577, w_001_2578, w_001_2580, w_001_2581, w_001_2583, w_001_2584, w_001_2585, w_001_2586, w_001_2587, w_001_2588, w_001_2589, w_001_2590, w_001_2591, w_001_2592, w_001_2593, w_001_2594, w_001_2595, w_001_2596, w_001_2597, w_001_2598, w_001_2599, w_001_2600, w_001_2601, w_001_2602, w_001_2603, w_001_2604, w_001_2605, w_001_2607, w_001_2608, w_001_2609, w_001_2610, w_001_2611, w_001_2612, w_001_2614, w_001_2615, w_001_2616, w_001_2617, w_001_2618, w_001_2619, w_001_2620, w_001_2621, w_001_2622, w_001_2623, w_001_2624, w_001_2625, w_001_2626, w_001_2627, w_001_2628, w_001_2629, w_001_2630, w_001_2632, w_001_2633, w_001_2634, w_001_2635, w_001_2636, w_001_2637, w_001_2638, w_001_2639, w_001_2640, w_001_2641, w_001_2642, w_001_2643, w_001_2644, w_001_2645, w_001_2646, w_001_2647, w_001_2648, w_001_2649, w_001_2650, w_001_2651, w_001_2652, w_001_2653, w_001_2654, w_001_2655, w_001_2656, w_001_2657, w_001_2658, w_001_2659, w_001_2660, w_001_2661, w_001_2662, w_001_2663, w_001_2664, w_001_2665, w_001_2666, w_001_2667, w_001_2668, w_001_2670, w_001_2671, w_001_2672, w_001_2673, w_001_2674, w_001_2675, w_001_2676, w_001_2677, w_001_2678, w_001_2680, w_001_2681, w_001_2682, w_001_2684, w_001_2685, w_001_2687, w_001_2688, w_001_2689, w_001_2690, w_001_2691, w_001_2692, w_001_2693, w_001_2694, w_001_2696, w_001_2697, w_001_2698, w_001_2699, w_001_2700, w_001_2701, w_001_2702, w_001_2703, w_001_2704, w_001_2705, w_001_2706, w_001_2707, w_001_2708, w_001_2709, w_001_2710, w_001_2711, w_001_2712, w_001_2713, w_001_2714, w_001_2715, w_001_2716, w_001_2717, w_001_2718, w_001_2719, w_001_2720, w_001_2722, w_001_2723, w_001_2724, w_001_2725, w_001_2726, w_001_2727, w_001_2728, w_001_2729, w_001_2730, w_001_2731, w_001_2732, w_001_2733, w_001_2734, w_001_2735, w_001_2736, w_001_2738, w_001_2739, w_001_2741, w_001_2742, w_001_2743, w_001_2744, w_001_2745, w_001_2746, w_001_2747, w_001_2748, w_001_2749, w_001_2750, w_001_2751, w_001_2752, w_001_2753, w_001_2754, w_001_2755, w_001_2756, w_001_2757, w_001_2758, w_001_2759, w_001_2760, w_001_2761, w_001_2762, w_001_2763, w_001_2764, w_001_2765, w_001_2766, w_001_2768, w_001_2769, w_001_2770, w_001_2772, w_001_2773, w_001_2774, w_001_2775, w_001_2776, w_001_2777, w_001_2778, w_001_2779, w_001_2780, w_001_2781, w_001_2782, w_001_2783, w_001_2784, w_001_2785, w_001_2786, w_001_2787, w_001_2788, w_001_2789, w_001_2790, w_001_2792, w_001_2793, w_001_2794, w_001_2795, w_001_2796, w_001_2797, w_001_2798, w_001_2799, w_001_2800, w_001_2801, w_001_2802, w_001_2803, w_001_2804, w_001_2805, w_001_2806, w_001_2807, w_001_2808, w_001_2809, w_001_2810, w_001_2811, w_001_2812, w_001_2813, w_001_2814, w_001_2815, w_001_2816, w_001_2817, w_001_2818, w_001_2819, w_001_2820, w_001_2821, w_001_2822, w_001_2823, w_001_2825, w_001_2827, w_001_2828, w_001_2829, w_001_2830, w_001_2831, w_001_2832, w_001_2833, w_001_2834, w_001_2835, w_001_2836, w_001_2837, w_001_2838, w_001_2839, w_001_2840, w_001_2841, w_001_2842, w_001_2843, w_001_2844, w_001_2845, w_001_2846, w_001_2847, w_001_2848, w_001_2850, w_001_2851, w_001_2852, w_001_2853, w_001_2854, w_001_2856, w_001_2857, w_001_2859, w_001_2860, w_001_2861, w_001_2862, w_001_2864, w_001_2865, w_001_2866, w_001_2867, w_001_2868, w_001_2869, w_001_2870, w_001_2871, w_001_2872, w_001_2873, w_001_2874, w_001_2875, w_001_2876, w_001_2877, w_001_2878, w_001_2879, w_001_2880, w_001_2881, w_001_2882, w_001_2884, w_001_2885, w_001_2886, w_001_2887, w_001_2888, w_001_2889, w_001_2890, w_001_2891, w_001_2892, w_001_2893, w_001_2894, w_001_2895, w_001_2896, w_001_2897, w_001_2898, w_001_2899, w_001_2900, w_001_2901, w_001_2902, w_001_2903, w_001_2904, w_001_2905, w_001_2906, w_001_2907, w_001_2908, w_001_2909, w_001_2910, w_001_2911, w_001_2912, w_001_2913, w_001_2914, w_001_2915, w_001_2916, w_001_2917, w_001_2918, w_001_2919, w_001_2920, w_001_2921, w_001_2922, w_001_2924, w_001_2925, w_001_2927, w_001_2928, w_001_2929, w_001_2931, w_001_2932, w_001_2933, w_001_2934, w_001_2935, w_001_2936, w_001_2937, w_001_2938, w_001_2939, w_001_2940, w_001_2941, w_001_2942, w_001_2943, w_001_2944, w_001_2945, w_001_2946, w_001_2947, w_001_2948, w_001_2949, w_001_2950, w_001_2951, w_001_2952, w_001_2953, w_001_2954, w_001_2955, w_001_2956, w_001_2957, w_001_2958, w_001_2959, w_001_2960, w_001_2961, w_001_2962, w_001_2965, w_001_2967, w_001_2968, w_001_2969, w_001_2970, w_001_2971, w_001_2972, w_001_2973, w_001_2974, w_001_2975, w_001_2976, w_001_2977, w_001_2978, w_001_2979, w_001_2980, w_001_2982, w_001_2983, w_001_2984, w_001_2985, w_001_2986, w_001_2987, w_001_2988, w_001_2989, w_001_2990, w_001_2991, w_001_2992, w_001_2993, w_001_2994, w_001_2995, w_001_2996, w_001_2997, w_001_2998, w_001_2999, w_001_3000, w_001_3001, w_001_3002, w_001_3003, w_001_3004, w_001_3005, w_001_3006, w_001_3007, w_001_3008, w_001_3009, w_001_3010, w_001_3011, w_001_3012, w_001_3013, w_001_3014, w_001_3015, w_001_3016, w_001_3018, w_001_3019, w_001_3020, w_001_3021, w_001_3022, w_001_3023, w_001_3024, w_001_3025, w_001_3026, w_001_3027, w_001_3028, w_001_3029, w_001_3031, w_001_3032, w_001_3033, w_001_3035, w_001_3036, w_001_3037, w_001_3038, w_001_3039, w_001_3040, w_001_3041, w_001_3042, w_001_3043, w_001_3044, w_001_3045, w_001_3046, w_001_3047, w_001_3048, w_001_3049, w_001_3050, w_001_3051, w_001_3052, w_001_3054, w_001_3055, w_001_3056, w_001_3057, w_001_3058, w_001_3059, w_001_3060, w_001_3061, w_001_3062, w_001_3063, w_001_3064, w_001_3065, w_001_3066, w_001_3067, w_001_3068, w_001_3069, w_001_3070, w_001_3071, w_001_3072, w_001_3073, w_001_3074, w_001_3075, w_001_3076, w_001_3077, w_001_3078, w_001_3079, w_001_3081, w_001_3082, w_001_3083, w_001_3084, w_001_3085, w_001_3086, w_001_3087, w_001_3089, w_001_3090, w_001_3091, w_001_3092, w_001_3093, w_001_3094, w_001_3095, w_001_3096, w_001_3097, w_001_3098, w_001_3099, w_001_3101, w_001_3102, w_001_3103, w_001_3104, w_001_3107, w_001_3108, w_001_3109, w_001_3110, w_001_3111, w_001_3112, w_001_3113, w_001_3114, w_001_3115, w_001_3116, w_001_3117, w_001_3118, w_001_3119, w_001_3120, w_001_3121, w_001_3122, w_001_3123, w_001_3124, w_001_3125, w_001_3126, w_001_3127, w_001_3128, w_001_3129, w_001_3130, w_001_3131, w_001_3132, w_001_3133, w_001_3134, w_001_3135, w_001_3136, w_001_3137, w_001_3139, w_001_3140, w_001_3141, w_001_3142, w_001_3143, w_001_3144, w_001_3146, w_001_3147, w_001_3148, w_001_3149, w_001_3150, w_001_3151, w_001_3152, w_001_3154, w_001_3155, w_001_3156, w_001_3157, w_001_3158, w_001_3159, w_001_3160, w_001_3161, w_001_3162, w_001_3163, w_001_3164, w_001_3165, w_001_3166, w_001_3167, w_001_3168, w_001_3169, w_001_3170, w_001_3171, w_001_3173, w_001_3174, w_001_3175, w_001_3176, w_001_3177, w_001_3178, w_001_3179, w_001_3180, w_001_3181, w_001_3182, w_001_3183, w_001_3186, w_001_3187, w_001_3188, w_001_3189, w_001_3190, w_001_3191, w_001_3192, w_001_3193, w_001_3195, w_001_3196, w_001_3197, w_001_3198, w_001_3199, w_001_3200, w_001_3201, w_001_3202, w_001_3203, w_001_3204, w_001_3205, w_001_3206, w_001_3207, w_001_3208, w_001_3209, w_001_3210, w_001_3211, w_001_3212, w_001_3214, w_001_3215, w_001_3216, w_001_3217, w_001_3218, w_001_3219, w_001_3220, w_001_3221, w_001_3222, w_001_3223, w_001_3224, w_001_3225, w_001_3226, w_001_3227, w_001_3228, w_001_3229, w_001_3230, w_001_3231, w_001_3232, w_001_3233, w_001_3234, w_001_3235, w_001_3236, w_001_3237, w_001_3238, w_001_3239, w_001_3240, w_001_3241, w_001_3242, w_001_3243, w_001_3244, w_001_3245, w_001_3246, w_001_3247, w_001_3249, w_001_3250, w_001_3251, w_001_3252, w_001_3253, w_001_3254, w_001_3255, w_001_3256, w_001_3257, w_001_3258, w_001_3259, w_001_3260, w_001_3261, w_001_3262, w_001_3263, w_001_3264, w_001_3265, w_001_3266, w_001_3267, w_001_3268, w_001_3269, w_001_3270, w_001_3271, w_001_3272, w_001_3273, w_001_3274, w_001_3275, w_001_3276, w_001_3277, w_001_3278, w_001_3280, w_001_3282, w_001_3283, w_001_3284, w_001_3285, w_001_3286, w_001_3287, w_001_3288, w_001_3289, w_001_3290, w_001_3291, w_001_3292, w_001_3293, w_001_3294, w_001_3295, w_001_3296, w_001_3297, w_001_3298, w_001_3299, w_001_3300, w_001_3301, w_001_3303, w_001_3305, w_001_3306, w_001_3307, w_001_3308, w_001_3309, w_001_3310, w_001_3311, w_001_3312, w_001_3313, w_001_3314, w_001_3315, w_001_3316, w_001_3317, w_001_3318, w_001_3319, w_001_3320, w_001_3321, w_001_3322, w_001_3323, w_001_3324, w_001_3326, w_001_3327, w_001_3328, w_001_3329, w_001_3330, w_001_3331, w_001_3332, w_001_3333, w_001_3334, w_001_3335, w_001_3336, w_001_3338, w_001_3339, w_001_3340, w_001_3341, w_001_3342, w_001_3343, w_001_3344, w_001_3345, w_001_3347, w_001_3348, w_001_3349, w_001_3350, w_001_3351, w_001_3353, w_001_3354, w_001_3355, w_001_3357, w_001_3358, w_001_3360, w_001_3361, w_001_3363, w_001_3364, w_001_3366, w_001_3367, w_001_3368, w_001_3369, w_001_3371, w_001_3372, w_001_3373, w_001_3374, w_001_3375, w_001_3376, w_001_3377, w_001_3378, w_001_3379, w_001_3380, w_001_3381, w_001_3382, w_001_3383, w_001_3384, w_001_3385, w_001_3386, w_001_3388, w_001_3389, w_001_3390, w_001_3392, w_001_3393, w_001_3394, w_001_3395, w_001_3396, w_001_3397, w_001_3398, w_001_3399, w_001_3400, w_001_3401, w_001_3402, w_001_3403, w_001_3404, w_001_3405, w_001_3406, w_001_3408, w_001_3409, w_001_3410, w_001_3411, w_001_3412, w_001_3413, w_001_3414, w_001_3415, w_001_3416, w_001_3417, w_001_3418, w_001_3419, w_001_3420, w_001_3422, w_001_3423, w_001_3424, w_001_3425, w_001_3426, w_001_3427, w_001_3428, w_001_3429, w_001_3430, w_001_3431, w_001_3432, w_001_3433, w_001_3434, w_001_3435, w_001_3436, w_001_3437, w_001_3438, w_001_3439, w_001_3440, w_001_3441, w_001_3442, w_001_3443, w_001_3444, w_001_3445, w_001_3446, w_001_3447, w_001_3448, w_001_3449, w_001_3450, w_001_3451, w_001_3452, w_001_3453, w_001_3454, w_001_3455, w_001_3456, w_001_3457, w_001_3458, w_001_3459, w_001_3460, w_001_3461, w_001_3462, w_001_3463, w_001_3464, w_001_3465, w_001_3467, w_001_3468, w_001_3469, w_001_3470, w_001_3471, w_001_3472, w_001_3473, w_001_3474, w_001_3475, w_001_3476, w_001_3477, w_001_3478, w_001_3479, w_001_3480, w_001_3481, w_001_3482, w_001_3483, w_001_3485, w_001_3486, w_001_3487, w_001_3488, w_001_3489, w_001_3490, w_001_3491, w_001_3492, w_001_3493, w_001_3494, w_001_3495, w_001_3496, w_001_3497, w_001_3498, w_001_3499, w_001_3500, w_001_3501, w_001_3502, w_001_3503, w_001_3504, w_001_3505, w_001_3506, w_001_3507, w_001_3508, w_001_3509, w_001_3510, w_001_3511, w_001_3512, w_001_3513, w_001_3514, w_001_3515, w_001_3516, w_001_3517, w_001_3518, w_001_3520, w_001_3521, w_001_3522, w_001_3523, w_001_3524, w_001_3525, w_001_3526, w_001_3527, w_001_3529, w_001_3530, w_001_3531, w_001_3532, w_001_3533, w_001_3534, w_001_3535, w_001_3536, w_001_3537, w_001_3538, w_001_3539, w_001_3540, w_001_3541, w_001_3544, w_001_3545, w_001_3546, w_001_3547, w_001_3548, w_001_3549, w_001_3550, w_001_3551, w_001_3552, w_001_3553, w_001_3554, w_001_3555, w_001_3556, w_001_3557, w_001_3558, w_001_3559, w_001_3560, w_001_3562, w_001_3563, w_001_3564, w_001_3566, w_001_3567, w_001_3568, w_001_3569, w_001_3570, w_001_3571, w_001_3572, w_001_3573, w_001_3574, w_001_3575, w_001_3576, w_001_3577, w_001_3578, w_001_3579, w_001_3580, w_001_3581, w_001_3582, w_001_3583, w_001_3584, w_001_3585, w_001_3586, w_001_3587, w_001_3588, w_001_3589, w_001_3590, w_001_3591, w_001_3592, w_001_3593, w_001_3594, w_001_3595, w_001_3596, w_001_3597, w_001_3598, w_001_3599, w_001_3600, w_001_3601, w_001_3602, w_001_3603, w_001_3604, w_001_3605, w_001_3606, w_001_3607, w_001_3608, w_001_3609, w_001_3610, w_001_3611, w_001_3612, w_001_3613, w_001_3614, w_001_3615, w_001_3616, w_001_3617, w_001_3618, w_001_3619, w_001_3620, w_001_3621, w_001_3622, w_001_3623, w_001_3624, w_001_3625, w_001_3626, w_001_3628, w_001_3629, w_001_3630, w_001_3631, w_001_3632, w_001_3633, w_001_3634, w_001_3635, w_001_3636, w_001_3637, w_001_3638, w_001_3639, w_001_3640, w_001_3641, w_001_3642, w_001_3643, w_001_3644, w_001_3645, w_001_3646, w_001_3648, w_001_3649, w_001_3650, w_001_3651, w_001_3652, w_001_3653, w_001_3654, w_001_3655, w_001_3656, w_001_3657, w_001_3658, w_001_3660, w_001_3661, w_001_3663, w_001_3665, w_001_3666, w_001_3667, w_001_3668, w_001_3669, w_001_3670, w_001_3671, w_001_3672, w_001_3673, w_001_3675, w_001_3677, w_001_3678, w_001_3679, w_001_3680, w_001_3681, w_001_3682, w_001_3683, w_001_3684, w_001_3685, w_001_3686, w_001_3687, w_001_3688, w_001_3689, w_001_3690, w_001_3691, w_001_3692, w_001_3693, w_001_3694, w_001_3696, w_001_3697, w_001_3698, w_001_3699, w_001_3700, w_001_3701, w_001_3702, w_001_3703, w_001_3704, w_001_3705, w_001_3706, w_001_3707, w_001_3708, w_001_3709, w_001_3710, w_001_3711, w_001_3712, w_001_3713, w_001_3714, w_001_3715, w_001_3716, w_001_3717, w_001_3718, w_001_3719, w_001_3720, w_001_3721, w_001_3722, w_001_3723, w_001_3724, w_001_3725, w_001_3726, w_001_3727, w_001_3728, w_001_3729, w_001_3730, w_001_3731, w_001_3733, w_001_3734, w_001_3735, w_001_3736, w_001_3738, w_001_3739, w_001_3740, w_001_3742, w_001_3743, w_001_3744, w_001_3745, w_001_3746, w_001_3747, w_001_3749, w_001_3750, w_001_3751, w_001_3752, w_001_3753, w_001_3754, w_001_3755, w_001_3756, w_001_3757, w_001_3758, w_001_3759, w_001_3760, w_001_3761, w_001_3762, w_001_3763, w_001_3764, w_001_3765, w_001_3766, w_001_3768, w_001_3769, w_001_3770, w_001_3771, w_001_3772, w_001_3773, w_001_3774, w_001_3775, w_001_3776, w_001_3777, w_001_3778, w_001_3780, w_001_3781, w_001_3782, w_001_3783, w_001_3784, w_001_3785, w_001_3786, w_001_3787, w_001_3788, w_001_3789, w_001_3790, w_001_3791, w_001_3793, w_001_3794, w_001_3795, w_001_3796, w_001_3797, w_001_3798, w_001_3800, w_001_3801, w_001_3802, w_001_3803, w_001_3804, w_001_3805, w_001_3807, w_001_3808, w_001_3809, w_001_3810, w_001_3811, w_001_3812, w_001_3813, w_001_3814, w_001_3815, w_001_3816, w_001_3818, w_001_3819, w_001_3820, w_001_3821, w_001_3822, w_001_3823, w_001_3824, w_001_3825, w_001_3826, w_001_3827, w_001_3828, w_001_3829, w_001_3830, w_001_3831, w_001_3832, w_001_3833, w_001_3835, w_001_3836, w_001_3837, w_001_3838, w_001_3839, w_001_3840, w_001_3841, w_001_3842, w_001_3843, w_001_3844, w_001_3845, w_001_3846, w_001_3847, w_001_3848, w_001_3849, w_001_3850, w_001_3851, w_001_3852, w_001_3853, w_001_3854, w_001_3855, w_001_3856, w_001_3857, w_001_3858, w_001_3859, w_001_3860, w_001_3861, w_001_3862, w_001_3863, w_001_3864, w_001_3865, w_001_3866, w_001_3867, w_001_3869, w_001_3870, w_001_3871, w_001_3872, w_001_3873, w_001_3874, w_001_3875, w_001_3876, w_001_3877, w_001_3878, w_001_3879, w_001_3880, w_001_3881, w_001_3882, w_001_3883, w_001_3884, w_001_3885, w_001_3886, w_001_3887, w_001_3888, w_001_3889, w_001_3890, w_001_3891, w_001_3892, w_001_3893, w_001_3894, w_001_3895, w_001_3896, w_001_3897, w_001_3899, w_001_3900, w_001_3901, w_001_3902, w_001_3903, w_001_3904, w_001_3905, w_001_3906, w_001_3907, w_001_3908, w_001_3909, w_001_3910, w_001_3911, w_001_3912, w_001_3913, w_001_3914, w_001_3915, w_001_3916, w_001_3917, w_001_3918, w_001_3919, w_001_3920, w_001_3921, w_001_3922, w_001_3923, w_001_3924, w_001_3925, w_001_3926, w_001_3927, w_001_3928, w_001_3929, w_001_3930, w_001_3932, w_001_3933, w_001_3934, w_001_3935, w_001_3936, w_001_3937, w_001_3938, w_001_3939, w_001_3940, w_001_3941, w_001_3942, w_001_3943, w_001_3944, w_001_3945, w_001_3947, w_001_3948, w_001_3949, w_001_3951, w_001_3952, w_001_3953, w_001_3955, w_001_3956, w_001_3957, w_001_3958, w_001_3959, w_001_3960, w_001_3961, w_001_3962, w_001_3963, w_001_3965, w_001_3966, w_001_3968, w_001_3969, w_001_3970, w_001_3971, w_001_3972, w_001_3973, w_001_3974, w_001_3975, w_001_3976, w_001_3977, w_001_3978, w_001_3979, w_001_3981, w_001_3982, w_001_3983, w_001_3984, w_001_3985, w_001_3986, w_001_3987, w_001_3988, w_001_3989, w_001_3991, w_001_3992, w_001_3993, w_001_3994, w_001_3995, w_001_3996, w_001_3997, w_001_3998, w_001_3999, w_001_4000, w_001_4001, w_001_4002, w_001_4003, w_001_4004, w_001_4005, w_001_4006, w_001_4007, w_001_4008, w_001_4010, w_001_4011, w_001_4012, w_001_4013, w_001_4014, w_001_4015, w_001_4016, w_001_4017, w_001_4018, w_001_4020, w_001_4021, w_001_4022, w_001_4023, w_001_4024, w_001_4025, w_001_4026, w_001_4027, w_001_4028, w_001_4029, w_001_4030, w_001_4031, w_001_4032, w_001_4033, w_001_4034, w_001_4035, w_001_4036, w_001_4037, w_001_4038, w_001_4039, w_001_4040, w_001_4041, w_001_4042, w_001_4043, w_001_4044, w_001_4046, w_001_4047, w_001_4049, w_001_4050, w_001_4051, w_001_4052, w_001_4053, w_001_4054, w_001_4055, w_001_4056, w_001_4057, w_001_4058, w_001_4059, w_001_4060, w_001_4062, w_001_4063, w_001_4064, w_001_4065, w_001_4066, w_001_4067, w_001_4068, w_001_4069, w_001_4070, w_001_4071, w_001_4072, w_001_4073, w_001_4074, w_001_4075, w_001_4076, w_001_4077, w_001_4078, w_001_4079, w_001_4080, w_001_4081, w_001_4082, w_001_4083, w_001_4084, w_001_4085, w_001_4087, w_001_4088, w_001_4089, w_001_4090, w_001_4091, w_001_4092, w_001_4093, w_001_4094, w_001_4095, w_001_4096, w_001_4097, w_001_4099, w_001_4100, w_001_4101, w_001_4102, w_001_4103, w_001_4104, w_001_4105, w_001_4107, w_001_4109, w_001_4110, w_001_4111, w_001_4112, w_001_4113, w_001_4114, w_001_4115, w_001_4116, w_001_4117, w_001_4118, w_001_4119, w_001_4120, w_001_4121, w_001_4123, w_001_4124, w_001_4125, w_001_4127, w_001_4128, w_001_4129, w_001_4130, w_001_4131, w_001_4132, w_001_4133, w_001_4134, w_001_4135, w_001_4136, w_001_4137, w_001_4139, w_001_4140, w_001_4141, w_001_4142, w_001_4143, w_001_4144, w_001_4145, w_001_4146, w_001_4147, w_001_4148, w_001_4149, w_001_4150, w_001_4151, w_001_4152, w_001_4153, w_001_4154, w_001_4156, w_001_4157, w_001_4158, w_001_4159, w_001_4160, w_001_4161, w_001_4162, w_001_4163, w_001_4164, w_001_4165, w_001_4166, w_001_4167, w_001_4168, w_001_4169, w_001_4170, w_001_4171, w_001_4172, w_001_4173, w_001_4174, w_001_4175, w_001_4176, w_001_4177, w_001_4178, w_001_4179, w_001_4180, w_001_4181, w_001_4182, w_001_4183, w_001_4184, w_001_4186, w_001_4188, w_001_4189, w_001_4190, w_001_4191, w_001_4192, w_001_4193, w_001_4194, w_001_4195, w_001_4196, w_001_4197, w_001_4198, w_001_4199, w_001_4200, w_001_4201, w_001_4202, w_001_4203, w_001_4204, w_001_4205, w_001_4207, w_001_4208, w_001_4209, w_001_4210, w_001_4211, w_001_4212, w_001_4213, w_001_4214, w_001_4215, w_001_4216, w_001_4217, w_001_4218, w_001_4219, w_001_4220, w_001_4222, w_001_4223, w_001_4224, w_001_4225, w_001_4226, w_001_4227, w_001_4228, w_001_4229, w_001_4230, w_001_4231, w_001_4232, w_001_4233, w_001_4234, w_001_4235, w_001_4236, w_001_4238, w_001_4239, w_001_4240, w_001_4241, w_001_4242, w_001_4243, w_001_4244, w_001_4245, w_001_4246, w_001_4247, w_001_4248, w_001_4249, w_001_4250, w_001_4251, w_001_4252, w_001_4253, w_001_4254, w_001_4255, w_001_4256, w_001_4257, w_001_4258, w_001_4259, w_001_4260, w_001_4261, w_001_4262, w_001_4263, w_001_4264, w_001_4265, w_001_4266, w_001_4267, w_001_4268, w_001_4269, w_001_4270, w_001_4271, w_001_4272, w_001_4273, w_001_4274, w_001_4275, w_001_4276, w_001_4277, w_001_4278, w_001_4279, w_001_4280, w_001_4281, w_001_4282, w_001_4283, w_001_4284, w_001_4285, w_001_4286, w_001_4287, w_001_4288, w_001_4289, w_001_4290, w_001_4291, w_001_4292, w_001_4293, w_001_4294, w_001_4295, w_001_4296, w_001_4297, w_001_4298, w_001_4299, w_001_4300, w_001_4301, w_001_4302, w_001_4303, w_001_4304, w_001_4305, w_001_4307, w_001_4308, w_001_4309, w_001_4310, w_001_4311, w_001_4312, w_001_4313, w_001_4314, w_001_4315, w_001_4316, w_001_4317, w_001_4318, w_001_4319, w_001_4320, w_001_4321, w_001_4322, w_001_4323, w_001_4324, w_001_4325, w_001_4326, w_001_4327, w_001_4328, w_001_4329, w_001_4330, w_001_4331, w_001_4332, w_001_4333, w_001_4335, w_001_4336, w_001_4337, w_001_4338, w_001_4339, w_001_4340, w_001_4341, w_001_4342, w_001_4343, w_001_4345, w_001_4346, w_001_4347, w_001_4348, w_001_4349, w_001_4351, w_001_4353, w_001_4354, w_001_4355, w_001_4356, w_001_4357, w_001_4358, w_001_4359, w_001_4361, w_001_4362, w_001_4363, w_001_4364, w_001_4365, w_001_4366, w_001_4367, w_001_4368, w_001_4369, w_001_4370, w_001_4371, w_001_4372, w_001_4373, w_001_4374, w_001_4375, w_001_4376, w_001_4377, w_001_4378, w_001_4379, w_001_4380, w_001_4381, w_001_4383, w_001_4384, w_001_4385, w_001_4386, w_001_4387, w_001_4389, w_001_4390, w_001_4391, w_001_4392, w_001_4394, w_001_4396, w_001_4397, w_001_4398, w_001_4399, w_001_4400, w_001_4402, w_001_4403, w_001_4404, w_001_4405, w_001_4406, w_001_4407, w_001_4408, w_001_4409, w_001_4411, w_001_4413, w_001_4414, w_001_4416, w_001_4417, w_001_4418, w_001_4420, w_001_4421, w_001_4422, w_001_4423, w_001_4424, w_001_4425, w_001_4426, w_001_4427, w_001_4428, w_001_4429, w_001_4430, w_001_4431, w_001_4432, w_001_4433, w_001_4434, w_001_4436, w_001_4437, w_001_4438, w_001_4439, w_001_4440, w_001_4441, w_001_4442, w_001_4443, w_001_4444, w_001_4445, w_001_4446, w_001_4447, w_001_4448, w_001_4450, w_001_4451, w_001_4452, w_001_4453, w_001_4454, w_001_4455, w_001_4456, w_001_4457, w_001_4458, w_001_4460, w_001_4461, w_001_4462, w_001_4463, w_001_4464, w_001_4465, w_001_4466, w_001_4467, w_001_4468, w_001_4469, w_001_4470, w_001_4471, w_001_4472, w_001_4473, w_001_4474, w_001_4475, w_001_4476, w_001_4477, w_001_4478, w_001_4479, w_001_4480, w_001_4481, w_001_4482, w_001_4483, w_001_4484, w_001_4485, w_001_4486, w_001_4487, w_001_4489, w_001_4490, w_001_4491, w_001_4492, w_001_4493, w_001_4494, w_001_4495, w_001_4496, w_001_4497, w_001_4498, w_001_4499, w_001_4500, w_001_4501, w_001_4502, w_001_4503, w_001_4504, w_001_4505, w_001_4506, w_001_4507, w_001_4508, w_001_4509, w_001_4510, w_001_4511, w_001_4512, w_001_4513, w_001_4514, w_001_4515, w_001_4516, w_001_4517, w_001_4518, w_001_4519, w_001_4520, w_001_4521, w_001_4522, w_001_4523, w_001_4524, w_001_4525, w_001_4526, w_001_4527, w_001_4528, w_001_4529, w_001_4530, w_001_4531, w_001_4532, w_001_4533, w_001_4534, w_001_4535, w_001_4536, w_001_4537, w_001_4538, w_001_4539, w_001_4540, w_001_4541, w_001_4542, w_001_4543, w_001_4544, w_001_4545, w_001_4546, w_001_4547, w_001_4548, w_001_4549, w_001_4551, w_001_4552, w_001_4553, w_001_4554, w_001_4555, w_001_4556, w_001_4557, w_001_4558, w_001_4559, w_001_4560, w_001_4561, w_001_4562, w_001_4563, w_001_4564, w_001_4565, w_001_4566, w_001_4567, w_001_4568, w_001_4569, w_001_4570, w_001_4571, w_001_4572, w_001_4573, w_001_4574, w_001_4575, w_001_4576, w_001_4577, w_001_4578, w_001_4579, w_001_4580, w_001_4581, w_001_4582, w_001_4583, w_001_4584, w_001_4585, w_001_4586, w_001_4587, w_001_4588, w_001_4589, w_001_4590, w_001_4591, w_001_4592, w_001_4593, w_001_4594, w_001_4597, w_001_4598, w_001_4600, w_001_4601, w_001_4602, w_001_4603, w_001_4604, w_001_4605, w_001_4607, w_001_4608, w_001_4609, w_001_4610, w_001_4611, w_001_4612, w_001_4613, w_001_4614, w_001_4615, w_001_4616, w_001_4617, w_001_4618, w_001_4619, w_001_4620, w_001_4621, w_001_4622, w_001_4623, w_001_4624, w_001_4625, w_001_4626, w_001_4627, w_001_4628, w_001_4629, w_001_4630, w_001_4631, w_001_4632, w_001_4633, w_001_4634, w_001_4635, w_001_4636, w_001_4637, w_001_4638, w_001_4639, w_001_4640, w_001_4641, w_001_4642, w_001_4643, w_001_4644, w_001_4645, w_001_4646, w_001_4647, w_001_4648, w_001_4649, w_001_4650, w_001_4651, w_001_4652, w_001_4653, w_001_4655, w_001_4656, w_001_4657, w_001_4658, w_001_4659, w_001_4660, w_001_4661, w_001_4662, w_001_4663, w_001_4664, w_001_4665, w_001_4666, w_001_4668, w_001_4669, w_001_4670, w_001_4671, w_001_4672, w_001_4673, w_001_4674, w_001_4675, w_001_4676, w_001_4677, w_001_4679, w_001_4680, w_001_4681, w_001_4682, w_001_4683, w_001_4684, w_001_4685, w_001_4686, w_001_4687, w_001_4688, w_001_4689, w_001_4690, w_001_4691, w_001_4693, w_001_4695, w_001_4696, w_001_4697, w_001_4698, w_001_4699, w_001_4700, w_001_4701, w_001_4702, w_001_4703, w_001_4704, w_001_4705, w_001_4706, w_001_4707, w_001_4708, w_001_4709, w_001_4710, w_001_4711, w_001_4712, w_001_4713, w_001_4714, w_001_4716, w_001_4717, w_001_4718, w_001_4719, w_001_4720, w_001_4721, w_001_4722, w_001_4723, w_001_4724, w_001_4725, w_001_4726, w_001_4727, w_001_4728, w_001_4729, w_001_4730, w_001_4731, w_001_4732, w_001_4733, w_001_4734, w_001_4735, w_001_4736, w_001_4737, w_001_4738, w_001_4739, w_001_4740, w_001_4741, w_001_4742, w_001_4743, w_001_4744, w_001_4745, w_001_4746, w_001_4747, w_001_4748, w_001_4749, w_001_4750, w_001_4753, w_001_4754, w_001_4755, w_001_4756, w_001_4757, w_001_4758, w_001_4759, w_001_4760, w_001_4761, w_001_4762, w_001_4763, w_001_4764, w_001_4765, w_001_4766, w_001_4767, w_001_4768, w_001_4769, w_001_4770, w_001_4771, w_001_4772, w_001_4773, w_001_4774, w_001_4775, w_001_4776, w_001_4777, w_001_4778, w_001_4779, w_001_4780, w_001_4781, w_001_4782, w_001_4783, w_001_4784, w_001_4785, w_001_4786, w_001_4787, w_001_4788, w_001_4790, w_001_4792, w_001_4793, w_001_4794, w_001_4795, w_001_4796, w_001_4798, w_001_4799, w_001_4800, w_001_4801, w_001_4802, w_001_4803, w_001_4804, w_001_4805, w_001_4806, w_001_4807, w_001_4808, w_001_4809, w_001_4810, w_001_4811, w_001_4812, w_001_4813, w_001_4814, w_001_4815, w_001_4816, w_001_4817, w_001_4818, w_001_4819, w_001_4820, w_001_4821, w_001_4822, w_001_4823, w_001_4824, w_001_4825, w_001_4826, w_001_4827, w_001_4828, w_001_4829, w_001_4830, w_001_4831, w_001_4832, w_001_4833, w_001_4834, w_001_4835, w_001_4836, w_001_4837, w_001_4839, w_001_4840, w_001_4841, w_001_4842, w_001_4843, w_001_4844, w_001_4845, w_001_4846, w_001_4847, w_001_4848, w_001_4850, w_001_4851, w_001_4852, w_001_4853, w_001_4854, w_001_4856, w_001_4857, w_001_4858, w_001_4859, w_001_4860, w_001_4862, w_001_4863, w_001_4864, w_001_4865, w_001_4866, w_001_4867, w_001_4868, w_001_4869, w_001_4870, w_001_4871, w_001_4872, w_001_4873, w_001_4874, w_001_4875, w_001_4876, w_001_4877, w_001_4879, w_001_4880, w_001_4881, w_001_4882, w_001_4884, w_001_4885, w_001_4886, w_001_4887, w_001_4888, w_001_4889, w_001_4890, w_001_4891, w_001_4892, w_001_4893, w_001_4894, w_001_4895, w_001_4896, w_001_4897, w_001_4898, w_001_4899, w_001_4900, w_001_4901, w_001_4902, w_001_4903, w_001_4904, w_001_4905, w_001_4906, w_001_4907, w_001_4909, w_001_4910, w_001_4911, w_001_4912, w_001_4913, w_001_4914, w_001_4915, w_001_4916, w_001_4917, w_001_4918, w_001_4919, w_001_4920, w_001_4921, w_001_4922, w_001_4923, w_001_4925, w_001_4927, w_001_4928, w_001_4929, w_001_4930, w_001_4931, w_001_4932, w_001_4933, w_001_4934, w_001_4936, w_001_4937, w_001_4938, w_001_4939, w_001_4940, w_001_4941, w_001_4943, w_001_4944, w_001_4946, w_001_4947, w_001_4948, w_001_4949, w_001_4951, w_001_4952, w_001_4953, w_001_4954, w_001_4955, w_001_4956, w_001_4957, w_001_4958, w_001_4960, w_001_4961, w_001_4962, w_001_4963, w_001_4964, w_001_4965, w_001_4966, w_001_4967, w_001_4968, w_001_4969, w_001_4970, w_001_4971, w_001_4972, w_001_4973, w_001_4974, w_001_4975, w_001_4976, w_001_4977, w_001_4978, w_001_4979, w_001_4980, w_001_4981, w_001_4982, w_001_4983, w_001_4984, w_001_4985, w_001_4986, w_001_4987, w_001_4988, w_001_4990, w_001_4991, w_001_4992, w_001_4993, w_001_4994, w_001_4995, w_001_4996, w_001_4997, w_001_4998, w_001_4999, w_001_5000, w_001_5001, w_001_5002, w_001_5003, w_001_5004, w_001_5005, w_001_5006, w_001_5007, w_001_5008, w_001_5009, w_001_5010, w_001_5012, w_001_5013, w_001_5014, w_001_5015, w_001_5016, w_001_5017, w_001_5018, w_001_5019, w_001_5020, w_001_5021, w_001_5022, w_001_5023, w_001_5024, w_001_5025, w_001_5026, w_001_5027, w_001_5028, w_001_5029, w_001_5030, w_001_5031, w_001_5032, w_001_5033, w_001_5034, w_001_5036, w_001_5037, w_001_5038, w_001_5039, w_001_5040, w_001_5041, w_001_5043, w_001_5044, w_001_5045, w_001_5046, w_001_5047, w_001_5048, w_001_5049, w_001_5050, w_001_5051, w_001_5052, w_001_5053, w_001_5054, w_001_5055, w_001_5056, w_001_5057, w_001_5058, w_001_5059, w_001_5060, w_001_5062, w_001_5063, w_001_5064, w_001_5065, w_001_5066, w_001_5067, w_001_5068, w_001_5069, w_001_5070, w_001_5071, w_001_5072, w_001_5073, w_001_5074, w_001_5075, w_001_5076, w_001_5077, w_001_5078, w_001_5080, w_001_5082, w_001_5083, w_001_5084, w_001_5085, w_001_5086, w_001_5087, w_001_5088, w_001_5089, w_001_5090, w_001_5091, w_001_5092, w_001_5093, w_001_5094, w_001_5095, w_001_5096, w_001_5098, w_001_5099, w_001_5100, w_001_5101, w_001_5102, w_001_5103, w_001_5106, w_001_5107, w_001_5108, w_001_5109, w_001_5110, w_001_5111, w_001_5112, w_001_5114, w_001_5115, w_001_5116, w_001_5117, w_001_5118, w_001_5119, w_001_5120, w_001_5121, w_001_5122, w_001_5123, w_001_5124, w_001_5125, w_001_5126, w_001_5127, w_001_5128, w_001_5129, w_001_5130, w_001_5131, w_001_5132, w_001_5133, w_001_5134, w_001_5135, w_001_5136, w_001_5137, w_001_5138, w_001_5140, w_001_5141, w_001_5142, w_001_5143, w_001_5144, w_001_5145, w_001_5146, w_001_5147, w_001_5148, w_001_5149, w_001_5150, w_001_5151, w_001_5152, w_001_5153, w_001_5154, w_001_5155, w_001_5157, w_001_5158, w_001_5159, w_001_5160, w_001_5161, w_001_5163, w_001_5164, w_001_5165, w_001_5167, w_001_5168, w_001_5169, w_001_5170, w_001_5171, w_001_5172, w_001_5173, w_001_5174, w_001_5175, w_001_5176, w_001_5177, w_001_5178, w_001_5179, w_001_5180, w_001_5181, w_001_5182, w_001_5183, w_001_5184, w_001_5185, w_001_5186, w_001_5187, w_001_5188, w_001_5189, w_001_5190, w_001_5191, w_001_5192, w_001_5194, w_001_5195, w_001_5196, w_001_5197, w_001_5198, w_001_5199, w_001_5200, w_001_5201, w_001_5202, w_001_5203, w_001_5204, w_001_5205, w_001_5206, w_001_5207, w_001_5208, w_001_5209, w_001_5210, w_001_5211, w_001_5212, w_001_5213, w_001_5214, w_001_5215, w_001_5216, w_001_5217, w_001_5218, w_001_5219, w_001_5220, w_001_5221, w_001_5222, w_001_5223, w_001_5224, w_001_5226, w_001_5227, w_001_5228, w_001_5229, w_001_5230, w_001_5231, w_001_5232, w_001_5233, w_001_5234, w_001_5235, w_001_5236, w_001_5237, w_001_5238, w_001_5239, w_001_5240, w_001_5241, w_001_5242, w_001_5243, w_001_5245, w_001_5246, w_001_5247, w_001_5248, w_001_5249, w_001_5250, w_001_5251, w_001_5253, w_001_5254, w_001_5255, w_001_5256, w_001_5257, w_001_5258, w_001_5259, w_001_5260, w_001_5261, w_001_5262, w_001_5263, w_001_5264, w_001_5265, w_001_5266, w_001_5267, w_001_5268, w_001_5269, w_001_5270, w_001_5271, w_001_5272, w_001_5273, w_001_5274, w_001_5275, w_001_5276, w_001_5278, w_001_5279, w_001_5280, w_001_5281, w_001_5282, w_001_5283, w_001_5284, w_001_5285, w_001_5286, w_001_5287, w_001_5288, w_001_5290, w_001_5291, w_001_5292, w_001_5293, w_001_5294, w_001_5295, w_001_5297, w_001_5299, w_001_5301, w_001_5303, w_001_5304, w_001_5305, w_001_5306, w_001_5307, w_001_5308, w_001_5309, w_001_5310, w_001_5311, w_001_5312, w_001_5313, w_001_5314, w_001_5315, w_001_5316, w_001_5318, w_001_5319, w_001_5320, w_001_5321, w_001_5322, w_001_5323, w_001_5324, w_001_5325, w_001_5326, w_001_5327, w_001_5328, w_001_5330, w_001_5331, w_001_5332, w_001_5333, w_001_5335, w_001_5336, w_001_5337, w_001_5338, w_001_5339, w_001_5340, w_001_5341, w_001_5342, w_001_5343, w_001_5344, w_001_5345, w_001_5346, w_001_5347, w_001_5348, w_001_5349, w_001_5350, w_001_5351, w_001_5352, w_001_5353, w_001_5354, w_001_5355, w_001_5356, w_001_5357, w_001_5358, w_001_5359, w_001_5360, w_001_5361, w_001_5362, w_001_5363, w_001_5365, w_001_5366, w_001_5367, w_001_5368, w_001_5369, w_001_5370, w_001_5371, w_001_5372, w_001_5373, w_001_5374, w_001_5375, w_001_5376, w_001_5377, w_001_5378, w_001_5379, w_001_5380, w_001_5381, w_001_5382, w_001_5383, w_001_5384, w_001_5385, w_001_5386, w_001_5387, w_001_5388, w_001_5389, w_001_5390, w_001_5392, w_001_5393, w_001_5394, w_001_5395, w_001_5396, w_001_5397, w_001_5398, w_001_5399, w_001_5400, w_001_5401, w_001_5402, w_001_5403, w_001_5404, w_001_5405, w_001_5406, w_001_5408, w_001_5409, w_001_5410, w_001_5411, w_001_5412, w_001_5413, w_001_5414, w_001_5415, w_001_5416, w_001_5417, w_001_5418, w_001_5419, w_001_5420, w_001_5422, w_001_5423, w_001_5424, w_001_5425, w_001_5426, w_001_5427, w_001_5428, w_001_5429, w_001_5430, w_001_5431, w_001_5432, w_001_5433, w_001_5434, w_001_5435, w_001_5436, w_001_5437, w_001_5438, w_001_5439, w_001_5440, w_001_5441, w_001_5443, w_001_5444, w_001_5445, w_001_5446, w_001_5447, w_001_5448, w_001_5449, w_001_5450, w_001_5451, w_001_5452, w_001_5453, w_001_5454, w_001_5455, w_001_5456, w_001_5457, w_001_5458, w_001_5459, w_001_5460, w_001_5461, w_001_5462, w_001_5463, w_001_5464, w_001_5465, w_001_5466, w_001_5467, w_001_5468, w_001_5469, w_001_5470, w_001_5471, w_001_5472, w_001_5473, w_001_5474, w_001_5475, w_001_5476, w_001_5477, w_001_5478, w_001_5479, w_001_5480, w_001_5481, w_001_5482, w_001_5483, w_001_5485, w_001_5486, w_001_5487, w_001_5488, w_001_5489, w_001_5490, w_001_5491, w_001_5492, w_001_5494, w_001_5495, w_001_5496, w_001_5497, w_001_5498, w_001_5499, w_001_5500, w_001_5501, w_001_5502, w_001_5503, w_001_5504, w_001_5505, w_001_5507, w_001_5508, w_001_5509, w_001_5510, w_001_5511, w_001_5512, w_001_5514, w_001_5515, w_001_5516, w_001_5517, w_001_5518, w_001_5519, w_001_5520, w_001_5521, w_001_5522, w_001_5523, w_001_5524, w_001_5525, w_001_5526, w_001_5527, w_001_5528, w_001_5529, w_001_5530, w_001_5531, w_001_5532, w_001_5533, w_001_5534, w_001_5535, w_001_5536, w_001_5538, w_001_5540, w_001_5541, w_001_5542, w_001_5543, w_001_5544, w_001_5545, w_001_5546, w_001_5547, w_001_5548, w_001_5549, w_001_5550, w_001_5552, w_001_5553, w_001_5554, w_001_5555, w_001_5556, w_001_5557, w_001_5558, w_001_5559, w_001_5560, w_001_5561, w_001_5562, w_001_5564, w_001_5565, w_001_5566, w_001_5567, w_001_5568, w_001_5570, w_001_5571, w_001_5572, w_001_5573, w_001_5574, w_001_5575, w_001_5576, w_001_5577, w_001_5578, w_001_5579, w_001_5580, w_001_5584, w_001_5585, w_001_5586, w_001_5588, w_001_5589, w_001_5590, w_001_5591, w_001_5592, w_001_5593, w_001_5594, w_001_5596, w_001_5597, w_001_5598, w_001_5599, w_001_5600, w_001_5601, w_001_5602, w_001_5603, w_001_5604, w_001_5605, w_001_5606, w_001_5607, w_001_5608, w_001_5609, w_001_5610, w_001_5611, w_001_5612, w_001_5613, w_001_5614, w_001_5615, w_001_5616, w_001_5617, w_001_5618, w_001_5619, w_001_5620, w_001_5621, w_001_5622, w_001_5623, w_001_5624, w_001_5625, w_001_5626, w_001_5627, w_001_5628, w_001_5630, w_001_5631, w_001_5633, w_001_5634, w_001_5635, w_001_5637, w_001_5638, w_001_5639, w_001_5640, w_001_5641, w_001_5642, w_001_5643, w_001_5644, w_001_5645, w_001_5646, w_001_5647, w_001_5648, w_001_5649, w_001_5650, w_001_5651, w_001_5652, w_001_5653, w_001_5654, w_001_5655, w_001_5656, w_001_5657, w_001_5658, w_001_5659, w_001_5660, w_001_5661, w_001_5662, w_001_5663, w_001_5664, w_001_5665, w_001_5666, w_001_5667, w_001_5668, w_001_5669, w_001_5671, w_001_5672, w_001_5673, w_001_5674, w_001_5675, w_001_5676, w_001_5677, w_001_5678, w_001_5679, w_001_5680, w_001_5681, w_001_5682, w_001_5684, w_001_5686, w_001_5687, w_001_5688, w_001_5689, w_001_5690, w_001_5691, w_001_5692, w_001_5693, w_001_5694, w_001_5695, w_001_5696, w_001_5697, w_001_5698, w_001_5699, w_001_5700, w_001_5701, w_001_5702, w_001_5703, w_001_5704, w_001_5705, w_001_5707, w_001_5708, w_001_5709, w_001_5710, w_001_5711, w_001_5712, w_001_5713, w_001_5714, w_001_5715, w_001_5716, w_001_5717, w_001_5720, w_001_5721, w_001_5722, w_001_5723, w_001_5724, w_001_5725, w_001_5726, w_001_5727, w_001_5728, w_001_5729, w_001_5730, w_001_5731, w_001_5732, w_001_5733, w_001_5734, w_001_5735, w_001_5736, w_001_5737, w_001_5738, w_001_5739, w_001_5740, w_001_5742, w_001_5743, w_001_5744, w_001_5745, w_001_5746, w_001_5747, w_001_5748, w_001_5749, w_001_5750, w_001_5751, w_001_5752, w_001_5753, w_001_5754, w_001_5755, w_001_5756, w_001_5757, w_001_5758, w_001_5759, w_001_5760, w_001_5761, w_001_5762, w_001_5763, w_001_5764, w_001_5765, w_001_5766, w_001_5767, w_001_5768, w_001_5769, w_001_5770, w_001_5771, w_001_5772, w_001_5773, w_001_5775, w_001_5776, w_001_5777, w_001_5778, w_001_5779, w_001_5780, w_001_5781, w_001_5782, w_001_5783, w_001_5784, w_001_5785, w_001_5786, w_001_5787, w_001_5788, w_001_5789, w_001_5790, w_001_5791, w_001_5792, w_001_5793, w_001_5794, w_001_5796, w_001_5797, w_001_5798, w_001_5799, w_001_5800, w_001_5801, w_001_5802, w_001_5803, w_001_5804, w_001_5805, w_001_5806, w_001_5807, w_001_5808, w_001_5810, w_001_5811, w_001_5812, w_001_5813, w_001_5814, w_001_5815, w_001_5816, w_001_5817, w_001_5818, w_001_5819, w_001_5820, w_001_5821, w_001_5822, w_001_5823, w_001_5824, w_001_5825, w_001_5826, w_001_5827, w_001_5828, w_001_5829, w_001_5831, w_001_5833, w_001_5834, w_001_5835, w_001_5836, w_001_5837, w_001_5838, w_001_5839, w_001_5840, w_001_5841, w_001_5842, w_001_5844, w_001_5845, w_001_5846, w_001_5847, w_001_5848, w_001_5849, w_001_5850, w_001_5851, w_001_5852, w_001_5853, w_001_5854, w_001_5855, w_001_5857, w_001_5858, w_001_5859, w_001_5861, w_001_5862, w_001_5863, w_001_5864, w_001_5865, w_001_5866, w_001_5867, w_001_5868, w_001_5869, w_001_5870, w_001_5871, w_001_5872, w_001_5873, w_001_5874, w_001_5875, w_001_5876, w_001_5877, w_001_5878, w_001_5879, w_001_5880, w_001_5881, w_001_5882, w_001_5883, w_001_5884, w_001_5885, w_001_5886, w_001_5887, w_001_5888, w_001_5889, w_001_5890, w_001_5891, w_001_5893, w_001_5895, w_001_5896, w_001_5898, w_001_5899, w_001_5900, w_001_5901, w_001_5902, w_001_5903, w_001_5904, w_001_5905, w_001_5906, w_001_5907, w_001_5908, w_001_5909, w_001_5911, w_001_5912, w_001_5913, w_001_5914, w_001_5915, w_001_5916, w_001_5917, w_001_5918, w_001_5919, w_001_5920, w_001_5921, w_001_5922, w_001_5925, w_001_5926, w_001_5927, w_001_5928, w_001_5929, w_001_5930, w_001_5931, w_001_5932, w_001_5933, w_001_5934, w_001_5935, w_001_5936, w_001_5937, w_001_5938, w_001_5939, w_001_5940, w_001_5941, w_001_5942, w_001_5943, w_001_5944, w_001_5945, w_001_5946, w_001_5947, w_001_5948, w_001_5949, w_001_5950, w_001_5952, w_001_5954, w_001_5955, w_001_5956, w_001_5957, w_001_5958, w_001_5959, w_001_5960, w_001_5961, w_001_5962, w_001_5963, w_001_5964, w_001_5965, w_001_5967, w_001_5968, w_001_5969, w_001_5970, w_001_5971, w_001_5972, w_001_5973, w_001_5975, w_001_5976, w_001_5977, w_001_5978, w_001_5979, w_001_5980, w_001_5981, w_001_5982, w_001_5983, w_001_5985, w_001_5986, w_001_5987, w_001_5988, w_001_5989, w_001_5990, w_001_5991, w_001_5992, w_001_5993, w_001_5994, w_001_5995, w_001_5996, w_001_5997, w_001_5998, w_001_5999, w_001_6000, w_001_6001, w_001_6002, w_001_6003, w_001_6004, w_001_6005, w_001_6006, w_001_6007, w_001_6008, w_001_6009, w_001_6010, w_001_6011, w_001_6012, w_001_6013, w_001_6014, w_001_6015, w_001_6016, w_001_6017, w_001_6018, w_001_6019, w_001_6020, w_001_6021, w_001_6022, w_001_6023, w_001_6024, w_001_6025, w_001_6026, w_001_6027, w_001_6028, w_001_6029, w_001_6030, w_001_6031, w_001_6032, w_001_6033, w_001_6034, w_001_6035, w_001_6036, w_001_6037, w_001_6038, w_001_6039, w_001_6040, w_001_6042, w_001_6043, w_001_6044, w_001_6045, w_001_6046, w_001_6047, w_001_6049, w_001_6050, w_001_6051, w_001_6052, w_001_6053, w_001_6054, w_001_6055, w_001_6057, w_001_6059, w_001_6060, w_001_6061, w_001_6062, w_001_6063, w_001_6064, w_001_6065, w_001_6066, w_001_6068, w_001_6069, w_001_6070, w_001_6071, w_001_6072, w_001_6073, w_001_6074, w_001_6075, w_001_6078, w_001_6079, w_001_6080, w_001_6081, w_001_6082, w_001_6083, w_001_6084, w_001_6085, w_001_6086, w_001_6087, w_001_6088, w_001_6089, w_001_6090, w_001_6091, w_001_6092, w_001_6093, w_001_6094, w_001_6095, w_001_6096, w_001_6098, w_001_6099, w_001_6100, w_001_6101, w_001_6102, w_001_6103, w_001_6104, w_001_6105, w_001_6106, w_001_6107, w_001_6108, w_001_6109, w_001_6110, w_001_6111, w_001_6112, w_001_6113, w_001_6114, w_001_6115, w_001_6117, w_001_6118, w_001_6119, w_001_6120, w_001_6121, w_001_6122, w_001_6123, w_001_6124, w_001_6125, w_001_6126, w_001_6127, w_001_6128, w_001_6129, w_001_6130, w_001_6131, w_001_6132, w_001_6133, w_001_6134, w_001_6135, w_001_6136, w_001_6137, w_001_6138, w_001_6139, w_001_6140, w_001_6141, w_001_6142, w_001_6143, w_001_6144, w_001_6145, w_001_6146, w_001_6147, w_001_6148, w_001_6149, w_001_6150, w_001_6151, w_001_6152, w_001_6153, w_001_6154, w_001_6155, w_001_6156, w_001_6157, w_001_6158, w_001_6159, w_001_6160, w_001_6161, w_001_6162, w_001_6163, w_001_6164, w_001_6165, w_001_6166, w_001_6167, w_001_6168, w_001_6169, w_001_6170, w_001_6171, w_001_6172, w_001_6173, w_001_6174, w_001_6175, w_001_6176, w_001_6177, w_001_6179, w_001_6180, w_001_6181, w_001_6182, w_001_6184, w_001_6185, w_001_6186, w_001_6187, w_001_6188, w_001_6189, w_001_6190, w_001_6191, w_001_6192, w_001_6193, w_001_6194, w_001_6195, w_001_6196, w_001_6197, w_001_6198, w_001_6199, w_001_6200, w_001_6201, w_001_6202, w_001_6203, w_001_6204, w_001_6205, w_001_6206, w_001_6207, w_001_6208, w_001_6209, w_001_6210, w_001_6211, w_001_6212, w_001_6213, w_001_6214, w_001_6215, w_001_6217, w_001_6218, w_001_6219, w_001_6220, w_001_6221, w_001_6222, w_001_6223, w_001_6224, w_001_6225, w_001_6226, w_001_6227, w_001_6228, w_001_6229, w_001_6230, w_001_6231, w_001_6232, w_001_6233, w_001_6234, w_001_6235, w_001_6236, w_001_6237, w_001_6238, w_001_6239, w_001_6240, w_001_6243, w_001_6244, w_001_6246, w_001_6247, w_001_6248, w_001_6249, w_001_6250, w_001_6251, w_001_6252, w_001_6253, w_001_6254, w_001_6255, w_001_6256, w_001_6258, w_001_6259, w_001_6260, w_001_6261, w_001_6262, w_001_6263, w_001_6265, w_001_6266, w_001_6267, w_001_6268, w_001_6269, w_001_6270, w_001_6271, w_001_6272, w_001_6273, w_001_6274, w_001_6275, w_001_6276, w_001_6277, w_001_6278, w_001_6279, w_001_6280, w_001_6281, w_001_6282, w_001_6283, w_001_6284, w_001_6285, w_001_6286, w_001_6287, w_001_6288, w_001_6289, w_001_6290, w_001_6291, w_001_6292, w_001_6293, w_001_6294, w_001_6295, w_001_6296, w_001_6297, w_001_6298, w_001_6299, w_001_6300, w_001_6301, w_001_6302, w_001_6303, w_001_6304, w_001_6305, w_001_6306, w_001_6307, w_001_6308, w_001_6309, w_001_6310, w_001_6311, w_001_6312, w_001_6313, w_001_6314, w_001_6315, w_001_6316, w_001_6317, w_001_6318, w_001_6319, w_001_6320, w_001_6321, w_001_6322, w_001_6323, w_001_6324, w_001_6325, w_001_6326, w_001_6327, w_001_6328, w_001_6329, w_001_6330, w_001_6332, w_001_6333, w_001_6334, w_001_6337, w_001_6338, w_001_6339, w_001_6340, w_001_6341, w_001_6342, w_001_6344, w_001_6345, w_001_6346, w_001_6347, w_001_6348, w_001_6349, w_001_6351, w_001_6352, w_001_6353, w_001_6354, w_001_6355, w_001_6356, w_001_6357, w_001_6358, w_001_6359, w_001_6360, w_001_6361, w_001_6362, w_001_6363, w_001_6364, w_001_6365, w_001_6366, w_001_6367, w_001_6368, w_001_6369, w_001_6370, w_001_6371, w_001_6372, w_001_6373, w_001_6375, w_001_6376, w_001_6377, w_001_6378, w_001_6379, w_001_6380, w_001_6381, w_001_6382, w_001_6383, w_001_6384, w_001_6385, w_001_6386, w_001_6387, w_001_6388, w_001_6389, w_001_6390, w_001_6391, w_001_6392, w_001_6393, w_001_6394, w_001_6395, w_001_6396, w_001_6397, w_001_6398, w_001_6399, w_001_6400, w_001_6401, w_001_6402, w_001_6403, w_001_6404, w_001_6405, w_001_6406, w_001_6407, w_001_6408, w_001_6409, w_001_6410, w_001_6411, w_001_6412, w_001_6413, w_001_6414, w_001_6416, w_001_6417, w_001_6419, w_001_6420, w_001_6421, w_001_6422, w_001_6423, w_001_6424, w_001_6425, w_001_6426, w_001_6427, w_001_6428, w_001_6429, w_001_6431, w_001_6432, w_001_6433, w_001_6434, w_001_6435, w_001_6436, w_001_6437, w_001_6438, w_001_6439, w_001_6440, w_001_6441, w_001_6442, w_001_6443, w_001_6444, w_001_6445, w_001_6446, w_001_6447, w_001_6448, w_001_6449, w_001_6450, w_001_6451, w_001_6452, w_001_6453, w_001_6454, w_001_6455, w_001_6456, w_001_6457, w_001_6458, w_001_6460, w_001_6461, w_001_6463, w_001_6464, w_001_6465, w_001_6466, w_001_6467, w_001_6468, w_001_6469, w_001_6470, w_001_6471, w_001_6472, w_001_6473, w_001_6474, w_001_6475, w_001_6476, w_001_6477, w_001_6478, w_001_6479, w_001_6480, w_001_6481, w_001_6482, w_001_6483, w_001_6484, w_001_6485, w_001_6486, w_001_6487, w_001_6488, w_001_6489, w_001_6490, w_001_6491, w_001_6492, w_001_6493, w_001_6494, w_001_6495, w_001_6496, w_001_6498, w_001_6499, w_001_6500, w_001_6501, w_001_6502, w_001_6503, w_001_6504, w_001_6505, w_001_6506, w_001_6509, w_001_6510, w_001_6511, w_001_6512, w_001_6513, w_001_6514, w_001_6515, w_001_6516, w_001_6517, w_001_6518, w_001_6519, w_001_6520, w_001_6521, w_001_6522, w_001_6523, w_001_6524, w_001_6525, w_001_6526, w_001_6527, w_001_6528, w_001_6529, w_001_6530, w_001_6531, w_001_6532, w_001_6533, w_001_6534, w_001_6535, w_001_6536, w_001_6537, w_001_6538, w_001_6539, w_001_6540, w_001_6541, w_001_6543, w_001_6544, w_001_6545, w_001_6546, w_001_6547, w_001_6548, w_001_6549, w_001_6550, w_001_6551, w_001_6552, w_001_6553, w_001_6554, w_001_6555, w_001_6556, w_001_6557, w_001_6558, w_001_6559, w_001_6560, w_001_6561, w_001_6562, w_001_6563, w_001_6564, w_001_6565, w_001_6566, w_001_6567, w_001_6568, w_001_6569, w_001_6570, w_001_6571, w_001_6572, w_001_6573, w_001_6574, w_001_6575, w_001_6576, w_001_6577, w_001_6579, w_001_6580, w_001_6581, w_001_6582, w_001_6583, w_001_6584, w_001_6585, w_001_6586, w_001_6587, w_001_6588, w_001_6590, w_001_6591, w_001_6592, w_001_6593, w_001_6594, w_001_6595, w_001_6596, w_001_6597, w_001_6598, w_001_6599, w_001_6600, w_001_6601, w_001_6602, w_001_6603, w_001_6604, w_001_6605, w_001_6606, w_001_6607, w_001_6608, w_001_6609, w_001_6610, w_001_6611, w_001_6613, w_001_6614, w_001_6615, w_001_6616, w_001_6617, w_001_6620, w_001_6621, w_001_6622, w_001_6623, w_001_6624, w_001_6626, w_001_6627, w_001_6628, w_001_6629, w_001_6630, w_001_6631, w_001_6632, w_001_6633, w_001_6634, w_001_6635, w_001_6636, w_001_6637, w_001_6638, w_001_6639, w_001_6640, w_001_6641, w_001_6642, w_001_6643, w_001_6644, w_001_6645, w_001_6646, w_001_6647, w_001_6649, w_001_6650, w_001_6651, w_001_6652, w_001_6653, w_001_6654, w_001_6655, w_001_6656, w_001_6657, w_001_6658, w_001_6659, w_001_6660, w_001_6663, w_001_6664, w_001_6665, w_001_6666, w_001_6667, w_001_6668, w_001_6669, w_001_6670, w_001_6671, w_001_6672, w_001_6673, w_001_6674, w_001_6676, w_001_6677, w_001_6678, w_001_6679, w_001_6680, w_001_6681, w_001_6682, w_001_6683, w_001_6684, w_001_6685, w_001_6686, w_001_6687, w_001_6688, w_001_6689, w_001_6690, w_001_6691, w_001_6692, w_001_6693, w_001_6694, w_001_6695, w_001_6696, w_001_6698, w_001_6699, w_001_6700, w_001_6701, w_001_6702, w_001_6703, w_001_6704, w_001_6705, w_001_6706, w_001_6707, w_001_6708, w_001_6709, w_001_6710, w_001_6711, w_001_6714, w_001_6715, w_001_6716, w_001_6717, w_001_6719, w_001_6720, w_001_6721, w_001_6722, w_001_6723, w_001_6724, w_001_6725, w_001_6727, w_001_6728, w_001_6729, w_001_6731, w_001_6732, w_001_6733, w_001_6734, w_001_6735, w_001_6736, w_001_6737, w_001_6738, w_001_6739, w_001_6740, w_001_6741, w_001_6742, w_001_6743, w_001_6744, w_001_6745, w_001_6746, w_001_6747, w_001_6748, w_001_6749, w_001_6750, w_001_6751, w_001_6752, w_001_6753, w_001_6754, w_001_6755, w_001_6756, w_001_6757, w_001_6759, w_001_6760, w_001_6761, w_001_6762, w_001_6763, w_001_6764, w_001_6765, w_001_6766, w_001_6767, w_001_6768, w_001_6770, w_001_6771, w_001_6772, w_001_6773, w_001_6774, w_001_6775, w_001_6776, w_001_6777, w_001_6778, w_001_6779, w_001_6780, w_001_6781, w_001_6782, w_001_6783, w_001_6784, w_001_6785, w_001_6786, w_001_6787, w_001_6788, w_001_6789, w_001_6790, w_001_6791, w_001_6792, w_001_6793, w_001_6794, w_001_6795, w_001_6796, w_001_6797, w_001_6798, w_001_6799, w_001_6800, w_001_6801, w_001_6802, w_001_6803, w_001_6804, w_001_6807, w_001_6808, w_001_6809, w_001_6810, w_001_6811, w_001_6812, w_001_6813, w_001_6814, w_001_6815, w_001_6816, w_001_6817, w_001_6818, w_001_6819, w_001_6820, w_001_6821, w_001_6822, w_001_6823, w_001_6824, w_001_6825, w_001_6826, w_001_6827, w_001_6828, w_001_6829, w_001_6830, w_001_6831, w_001_6832, w_001_6833, w_001_6835, w_001_6836, w_001_6837, w_001_6838, w_001_6839, w_001_6840, w_001_6841, w_001_6842, w_001_6843, w_001_6844, w_001_6845, w_001_6846, w_001_6847, w_001_6848, w_001_6849, w_001_6850, w_001_6851, w_001_6852, w_001_6853, w_001_6854, w_001_6855, w_001_6856, w_001_6857, w_001_6858, w_001_6859, w_001_6860, w_001_6861, w_001_6862, w_001_6863, w_001_6864, w_001_6865, w_001_6866, w_001_6867, w_001_6868, w_001_6869, w_001_6870, w_001_6871, w_001_6872, w_001_6873, w_001_6874, w_001_6875, w_001_6876, w_001_6877, w_001_6878, w_001_6879, w_001_6880, w_001_6881, w_001_6882, w_001_6884, w_001_6885, w_001_6886, w_001_6887, w_001_6888, w_001_6889, w_001_6890, w_001_6891, w_001_6892, w_001_6893, w_001_6894, w_001_6895, w_001_6896, w_001_6897, w_001_6898, w_001_6899, w_001_6900, w_001_6901, w_001_6903, w_001_6904, w_001_6905, w_001_6906, w_001_6907, w_001_6908, w_001_6909, w_001_6910, w_001_6911, w_001_6912, w_001_6913, w_001_6914, w_001_6915, w_001_6916, w_001_6917, w_001_6918, w_001_6919, w_001_6920, w_001_6921, w_001_6922, w_001_6923, w_001_6924, w_001_6925, w_001_6927, w_001_6928, w_001_6929, w_001_6930, w_001_6931, w_001_6932, w_001_6933, w_001_6935, w_001_6936, w_001_6937, w_001_6938, w_001_6939, w_001_6940, w_001_6941, w_001_6942, w_001_6943, w_001_6944, w_001_6945, w_001_6946, w_001_6947, w_001_6948, w_001_6949, w_001_6950, w_001_6951, w_001_6952, w_001_6953, w_001_6954, w_001_6955, w_001_6956, w_001_6957, w_001_6958, w_001_6959, w_001_6960, w_001_6961, w_001_6962, w_001_6963, w_001_6964, w_001_6965, w_001_6966, w_001_6967, w_001_6968, w_001_6969, w_001_6970, w_001_6971, w_001_6972, w_001_6973, w_001_6974, w_001_6975, w_001_6976, w_001_6977, w_001_6978, w_001_6979, w_001_6980, w_001_6981, w_001_6982, w_001_6983, w_001_6984, w_001_6985, w_001_6986, w_001_6987, w_001_6989, w_001_6990, w_001_6991, w_001_6992, w_001_6993, w_001_6994, w_001_6995, w_001_6996, w_001_6997, w_001_6999, w_001_7001, w_001_7002, w_001_7003, w_001_7004, w_001_7005, w_001_7006, w_001_7007, w_001_7008, w_001_7009, w_001_7011, w_001_7012, w_001_7013, w_001_7014, w_001_7015, w_001_7016, w_001_7017, w_001_7018, w_001_7019, w_001_7020, w_001_7021, w_001_7022, w_001_7024, w_001_7025, w_001_7026, w_001_7027, w_001_7028, w_001_7029, w_001_7030, w_001_7032, w_001_7033, w_001_7034, w_001_7035, w_001_7036, w_001_7037, w_001_7038, w_001_7039, w_001_7040, w_001_7041, w_001_7042, w_001_7043, w_001_7044, w_001_7045, w_001_7046, w_001_7047, w_001_7048, w_001_7049, w_001_7050, w_001_7051, w_001_7052, w_001_7053, w_001_7055, w_001_7056, w_001_7057, w_001_7058, w_001_7059, w_001_7060, w_001_7061, w_001_7062, w_001_7063, w_001_7064, w_001_7065, w_001_7066, w_001_7067, w_001_7068, w_001_7069, w_001_7070, w_001_7071, w_001_7072, w_001_7074, w_001_7075, w_001_7077, w_001_7078, w_001_7079, w_001_7080, w_001_7081, w_001_7082, w_001_7083, w_001_7084, w_001_7085, w_001_7086, w_001_7087, w_001_7088, w_001_7089, w_001_7090, w_001_7091, w_001_7092, w_001_7093, w_001_7094, w_001_7095, w_001_7096, w_001_7097, w_001_7098, w_001_7099, w_001_7100, w_001_7101, w_001_7102, w_001_7103, w_001_7104, w_001_7105, w_001_7107, w_001_7108, w_001_7109, w_001_7110, w_001_7111, w_001_7112, w_001_7113, w_001_7114, w_001_7115, w_001_7116, w_001_7117, w_001_7118, w_001_7119, w_001_7120, w_001_7121, w_001_7122, w_001_7123, w_001_7124, w_001_7125, w_001_7126, w_001_7127, w_001_7128, w_001_7129, w_001_7130, w_001_7131, w_001_7132, w_001_7133, w_001_7134, w_001_7135, w_001_7136, w_001_7137, w_001_7139, w_001_7140, w_001_7141, w_001_7142, w_001_7143, w_001_7144, w_001_7145, w_001_7146, w_001_7147, w_001_7148, w_001_7149, w_001_7150, w_001_7151, w_001_7152, w_001_7153, w_001_7154, w_001_7156, w_001_7157, w_001_7158, w_001_7159, w_001_7160, w_001_7161, w_001_7162, w_001_7163, w_001_7164, w_001_7165, w_001_7166, w_001_7167, w_001_7168, w_001_7169, w_001_7170, w_001_7171, w_001_7172, w_001_7173, w_001_7174, w_001_7175, w_001_7176, w_001_7177, w_001_7178, w_001_7180, w_001_7181, w_001_7182, w_001_7183, w_001_7184, w_001_7185, w_001_7186, w_001_7187, w_001_7188, w_001_7189, w_001_7190, w_001_7192, w_001_7193, w_001_7194, w_001_7195, w_001_7196, w_001_7197, w_001_7198, w_001_7199, w_001_7200, w_001_7201, w_001_7202, w_001_7203, w_001_7204, w_001_7205, w_001_7206, w_001_7207, w_001_7208, w_001_7209, w_001_7210, w_001_7211, w_001_7213, w_001_7214, w_001_7215, w_001_7216, w_001_7217, w_001_7218, w_001_7219, w_001_7220, w_001_7221, w_001_7222, w_001_7223, w_001_7224, w_001_7225, w_001_7226, w_001_7227, w_001_7228, w_001_7230, w_001_7231, w_001_7232, w_001_7233, w_001_7234, w_001_7235, w_001_7236, w_001_7237, w_001_7238, w_001_7239, w_001_7240, w_001_7241, w_001_7242, w_001_7244, w_001_7245, w_001_7246, w_001_7247, w_001_7248, w_001_7249, w_001_7250, w_001_7251, w_001_7253, w_001_7254, w_001_7255, w_001_7256, w_001_7257, w_001_7258, w_001_7259, w_001_7260, w_001_7261, w_001_7262, w_001_7263, w_001_7264, w_001_7265, w_001_7267, w_001_7268, w_001_7269, w_001_7270, w_001_7271, w_001_7272, w_001_7273, w_001_7274, w_001_7275, w_001_7276, w_001_7277, w_001_7278, w_001_7279, w_001_7280, w_001_7281, w_001_7282, w_001_7283, w_001_7284, w_001_7285, w_001_7286, w_001_7287, w_001_7288, w_001_7289, w_001_7290, w_001_7292, w_001_7293, w_001_7294, w_001_7295, w_001_7296, w_001_7297, w_001_7298, w_001_7299, w_001_7300, w_001_7301, w_001_7302, w_001_7303, w_001_7304, w_001_7305, w_001_7306, w_001_7307, w_001_7308, w_001_7309, w_001_7310, w_001_7311, w_001_7312, w_001_7313, w_001_7314, w_001_7315, w_001_7316, w_001_7317, w_001_7318, w_001_7319, w_001_7320, w_001_7321, w_001_7322, w_001_7323, w_001_7324, w_001_7325, w_001_7326, w_001_7327, w_001_7328, w_001_7329, w_001_7330, w_001_7331, w_001_7332, w_001_7333, w_001_7334, w_001_7335, w_001_7336, w_001_7337, w_001_7338, w_001_7339, w_001_7340, w_001_7341, w_001_7342, w_001_7343, w_001_7344, w_001_7345, w_001_7346, w_001_7347, w_001_7348, w_001_7349, w_001_7350, w_001_7351, w_001_7352, w_001_7353, w_001_7354, w_001_7355, w_001_7356, w_001_7358, w_001_7359, w_001_7360, w_001_7361, w_001_7362, w_001_7364, w_001_7365, w_001_7366, w_001_7367, w_001_7368, w_001_7369, w_001_7370, w_001_7371, w_001_7372, w_001_7373, w_001_7374, w_001_7375, w_001_7376, w_001_7377, w_001_7378, w_001_7379, w_001_7380, w_001_7381, w_001_7382, w_001_7383, w_001_7384, w_001_7385, w_001_7386, w_001_7387, w_001_7388, w_001_7389, w_001_7390, w_001_7391, w_001_7392, w_001_7393, w_001_7394, w_001_7395, w_001_7396, w_001_7397, w_001_7398, w_001_7399, w_001_7401, w_001_7402, w_001_7403, w_001_7404, w_001_7405, w_001_7406, w_001_7407, w_001_7408, w_001_7409, w_001_7410, w_001_7411, w_001_7412, w_001_7413, w_001_7414, w_001_7416, w_001_7417, w_001_7418, w_001_7419, w_001_7420, w_001_7421, w_001_7422, w_001_7423, w_001_7424, w_001_7425, w_001_7426, w_001_7427, w_001_7428, w_001_7430, w_001_7431, w_001_7432, w_001_7433, w_001_7434, w_001_7435, w_001_7436, w_001_7437, w_001_7438, w_001_7439, w_001_7440, w_001_7442, w_001_7443, w_001_7444, w_001_7445, w_001_7446, w_001_7447, w_001_7448, w_001_7449, w_001_7450, w_001_7451, w_001_7452, w_001_7453, w_001_7454, w_001_7455, w_001_7456, w_001_7457, w_001_7458, w_001_7459, w_001_7460, w_001_7461, w_001_7462, w_001_7463, w_001_7464, w_001_7465, w_001_7467, w_001_7468, w_001_7469, w_001_7470, w_001_7471, w_001_7472, w_001_7473, w_001_7474, w_001_7475, w_001_7476, w_001_7477, w_001_7478, w_001_7479, w_001_7480, w_001_7481, w_001_7482, w_001_7483, w_001_7484, w_001_7485, w_001_7486, w_001_7487, w_001_7488, w_001_7489, w_001_7490, w_001_7491, w_001_7492, w_001_7493, w_001_7494, w_001_7495, w_001_7496, w_001_7497, w_001_7498, w_001_7499, w_001_7500, w_001_7501, w_001_7502, w_001_7503, w_001_7504, w_001_7505, w_001_7506, w_001_7507, w_001_7508, w_001_7509, w_001_7510, w_001_7511, w_001_7512, w_001_7513, w_001_7514, w_001_7515, w_001_7516, w_001_7517, w_001_7518, w_001_7520, w_001_7521, w_001_7522, w_001_7523, w_001_7524, w_001_7525, w_001_7526, w_001_7528, w_001_7529, w_001_7530, w_001_7531, w_001_7532, w_001_7533, w_001_7534, w_001_7535, w_001_7537, w_001_7538, w_001_7539, w_001_7540, w_001_7541, w_001_7542, w_001_7543, w_001_7544, w_001_7545, w_001_7546, w_001_7547, w_001_7548, w_001_7549, w_001_7550, w_001_7551, w_001_7552, w_001_7553, w_001_7554, w_001_7555, w_001_7556, w_001_7557, w_001_7558, w_001_7559, w_001_7560, w_001_7561, w_001_7562, w_001_7563, w_001_7564, w_001_7565, w_001_7566, w_001_7567, w_001_7568, w_001_7569, w_001_7570, w_001_7571, w_001_7572, w_001_7573, w_001_7574, w_001_7575, w_001_7576, w_001_7577, w_001_7580, w_001_7581, w_001_7582, w_001_7583, w_001_7584, w_001_7585, w_001_7586, w_001_7587, w_001_7588, w_001_7589, w_001_7590, w_001_7591, w_001_7593, w_001_7594, w_001_7595, w_001_7596, w_001_7597, w_001_7598, w_001_7599, w_001_7600, w_001_7601, w_001_7602, w_001_7603, w_001_7604, w_001_7605, w_001_7606, w_001_7607, w_001_7608, w_001_7609, w_001_7610, w_001_7611, w_001_7612, w_001_7613, w_001_7615, w_001_7616, w_001_7617, w_001_7618, w_001_7619, w_001_7620, w_001_7621, w_001_7622, w_001_7623, w_001_7624, w_001_7625, w_001_7626, w_001_7627, w_001_7628, w_001_7629, w_001_7630, w_001_7631, w_001_7632, w_001_7633, w_001_7634, w_001_7635, w_001_7636, w_001_7637, w_001_7638, w_001_7639, w_001_7640, w_001_7641, w_001_7642, w_001_7643, w_001_7644, w_001_7645, w_001_7646, w_001_7647, w_001_7648, w_001_7649, w_001_7650, w_001_7651, w_001_7652, w_001_7653, w_001_7654, w_001_7655, w_001_7656, w_001_7657, w_001_7658, w_001_7659, w_001_7660, w_001_7661, w_001_7662, w_001_7663, w_001_7664, w_001_7665, w_001_7666, w_001_7667, w_001_7668, w_001_7669, w_001_7670, w_001_7671, w_001_7673, w_001_7674, w_001_7675, w_001_7676, w_001_7677, w_001_7678, w_001_7679, w_001_7680, w_001_7681, w_001_7682, w_001_7683, w_001_7684, w_001_7685, w_001_7686, w_001_7687, w_001_7688, w_001_7689, w_001_7690, w_001_7691, w_001_7693, w_001_7694, w_001_7695, w_001_7696, w_001_7697, w_001_7698, w_001_7699, w_001_7700, w_001_7701, w_001_7703, w_001_7704, w_001_7705, w_001_7706, w_001_7707, w_001_7708, w_001_7709, w_001_7710, w_001_7711, w_001_7712, w_001_7713, w_001_7715, w_001_7716, w_001_7717, w_001_7718, w_001_7719, w_001_7720, w_001_7721, w_001_7722, w_001_7723, w_001_7724, w_001_7725, w_001_7728, w_001_7729, w_001_7730, w_001_7731, w_001_7732, w_001_7733, w_001_7734, w_001_7735, w_001_7736, w_001_7737, w_001_7738, w_001_7739, w_001_7740, w_001_7741, w_001_7742, w_001_7743, w_001_7744, w_001_7745, w_001_7746, w_001_7747, w_001_7748, w_001_7749, w_001_7750, w_001_7752, w_001_7753, w_001_7754, w_001_7755, w_001_7756, w_001_7757, w_001_7758, w_001_7759, w_001_7760, w_001_7761, w_001_7762, w_001_7763, w_001_7764, w_001_7765, w_001_7766, w_001_7767, w_001_7768, w_001_7769, w_001_7770, w_001_7771, w_001_7772, w_001_7773, w_001_7774, w_001_7775, w_001_7776, w_001_7777, w_001_7778, w_001_7779, w_001_7781, w_001_7782, w_001_7783, w_001_7784, w_001_7785, w_001_7786, w_001_7787, w_001_7788, w_001_7789, w_001_7790, w_001_7792, w_001_7793, w_001_7794, w_001_7795, w_001_7796, w_001_7797, w_001_7798, w_001_7799, w_001_7801, w_001_7802, w_001_7803, w_001_7804, w_001_7805, w_001_7806, w_001_7807, w_001_7808, w_001_7809, w_001_7810, w_001_7811, w_001_7812, w_001_7813, w_001_7814, w_001_7816, w_001_7817, w_001_7818, w_001_7819, w_001_7820, w_001_7821, w_001_7822, w_001_7823, w_001_7824, w_001_7825, w_001_7826, w_001_7827, w_001_7828, w_001_7829, w_001_7830, w_001_7831, w_001_7832, w_001_7833, w_001_7834, w_001_7835, w_001_7836, w_001_7837, w_001_7838, w_001_7839, w_001_7840, w_001_7841, w_001_7842, w_001_7844, w_001_7845, w_001_7846, w_001_7847, w_001_7848, w_001_7849, w_001_7850, w_001_7851, w_001_7852, w_001_7853, w_001_7854, w_001_7855, w_001_7856, w_001_7857, w_001_7858, w_001_7859, w_001_7860, w_001_7861, w_001_7862, w_001_7863, w_001_7864, w_001_7865, w_001_7866, w_001_7867, w_001_7868, w_001_7870, w_001_7871, w_001_7872, w_001_7873, w_001_7874, w_001_7876, w_001_7878, w_001_7879, w_001_7880, w_001_7881, w_001_7884, w_001_7885, w_001_7886, w_001_7887, w_001_7888, w_001_7889, w_001_7890, w_001_7892, w_001_7894, w_001_7895, w_001_7896, w_001_7897, w_001_7898, w_001_7899, w_001_7900, w_001_7901, w_001_7902, w_001_7903, w_001_7906, w_001_7907, w_001_7908, w_001_7909, w_001_7910, w_001_7911, w_001_7912, w_001_7913, w_001_7914, w_001_7915, w_001_7917, w_001_7918, w_001_7919, w_001_7920, w_001_7921, w_001_7922, w_001_7923, w_001_7924, w_001_7925, w_001_7926, w_001_7927, w_001_7928, w_001_7929, w_001_7930, w_001_7931, w_001_7932, w_001_7933, w_001_7934, w_001_7935, w_001_7936, w_001_7938, w_001_7939, w_001_7940, w_001_7942, w_001_7943, w_001_7944, w_001_7945, w_001_7946, w_001_7947, w_001_7948, w_001_7950, w_001_7951, w_001_7952, w_001_7953, w_001_7954, w_001_7955, w_001_7956, w_001_7957, w_001_7958, w_001_7959, w_001_7960, w_001_7961, w_001_7962, w_001_7963, w_001_7964, w_001_7965, w_001_7966, w_001_7967, w_001_7968, w_001_7969, w_001_7970, w_001_7971, w_001_7972, w_001_7973, w_001_7974, w_001_7975, w_001_7976, w_001_7977, w_001_7978, w_001_7979, w_001_7980, w_001_7981, w_001_7982, w_001_7983, w_001_7984, w_001_7985, w_001_7986, w_001_7987, w_001_7988, w_001_7989, w_001_7990, w_001_7991, w_001_7992, w_001_7993, w_001_7994, w_001_7995, w_001_7996, w_001_7997, w_001_7998, w_001_7999, w_001_8000, w_001_8001, w_001_8002, w_001_8003, w_001_8004, w_001_8006, w_001_8007, w_001_8008, w_001_8009, w_001_8010, w_001_8011, w_001_8012, w_001_8013, w_001_8014, w_001_8015, w_001_8016, w_001_8017, w_001_8018, w_001_8019, w_001_8020, w_001_8021, w_001_8022, w_001_8023, w_001_8024, w_001_8025, w_001_8026, w_001_8027, w_001_8028, w_001_8029, w_001_8030, w_001_8031, w_001_8032, w_001_8033, w_001_8034, w_001_8036, w_001_8037, w_001_8038, w_001_8039, w_001_8040, w_001_8042, w_001_8043, w_001_8044, w_001_8045, w_001_8046, w_001_8047, w_001_8048, w_001_8049, w_001_8050, w_001_8051, w_001_8052, w_001_8054, w_001_8055, w_001_8056, w_001_8057, w_001_8058, w_001_8059, w_001_8061, w_001_8062, w_001_8063, w_001_8064, w_001_8065, w_001_8066, w_001_8067, w_001_8068, w_001_8069, w_001_8070, w_001_8072, w_001_8073, w_001_8074, w_001_8075, w_001_8078, w_001_8079, w_001_8080, w_001_8081, w_001_8082, w_001_8083, w_001_8084, w_001_8085, w_001_8086, w_001_8087, w_001_8088, w_001_8089, w_001_8090, w_001_8091, w_001_8092, w_001_8093, w_001_8094, w_001_8095, w_001_8096, w_001_8097, w_001_8098, w_001_8099, w_001_8100, w_001_8101, w_001_8102, w_001_8104, w_001_8105, w_001_8106, w_001_8107, w_001_8108, w_001_8109, w_001_8110, w_001_8111, w_001_8112, w_001_8113, w_001_8114, w_001_8115, w_001_8116, w_001_8117, w_001_8118, w_001_8119, w_001_8120, w_001_8121, w_001_8122, w_001_8123, w_001_8124, w_001_8125, w_001_8126, w_001_8127, w_001_8128, w_001_8129, w_001_8130, w_001_8131, w_001_8132, w_001_8133, w_001_8134, w_001_8135, w_001_8136, w_001_8138, w_001_8139, w_001_8140, w_001_8141, w_001_8142, w_001_8143, w_001_8144, w_001_8145, w_001_8146, w_001_8147, w_001_8148, w_001_8149, w_001_8150, w_001_8151, w_001_8152, w_001_8153, w_001_8155, w_001_8156, w_001_8157, w_001_8158, w_001_8159, w_001_8160, w_001_8161, w_001_8162, w_001_8163, w_001_8164, w_001_8165, w_001_8166, w_001_8167, w_001_8168, w_001_8169, w_001_8170, w_001_8171, w_001_8172, w_001_8173, w_001_8174, w_001_8175, w_001_8176, w_001_8177, w_001_8178, w_001_8179, w_001_8180, w_001_8181, w_001_8182, w_001_8183, w_001_8185, w_001_8186, w_001_8187, w_001_8188, w_001_8189, w_001_8190, w_001_8191, w_001_8193, w_001_8194, w_001_8195, w_001_8196, w_001_8197, w_001_8198, w_001_8199, w_001_8201, w_001_8202, w_001_8203, w_001_8204, w_001_8206, w_001_8207, w_001_8208, w_001_8209, w_001_8210, w_001_8211, w_001_8212, w_001_8213, w_001_8214, w_001_8215, w_001_8216, w_001_8217, w_001_8218, w_001_8219, w_001_8220, w_001_8221, w_001_8222, w_001_8223, w_001_8224, w_001_8225, w_001_8226, w_001_8227, w_001_8228, w_001_8229, w_001_8230, w_001_8231, w_001_8232, w_001_8233, w_001_8234, w_001_8235, w_001_8236, w_001_8237, w_001_8238, w_001_8239, w_001_8240, w_001_8241, w_001_8242, w_001_8243, w_001_8244, w_001_8246, w_001_8247, w_001_8248, w_001_8249, w_001_8250, w_001_8252, w_001_8253, w_001_8255, w_001_8256, w_001_8257, w_001_8258, w_001_8259, w_001_8260, w_001_8261, w_001_8262, w_001_8263, w_001_8264, w_001_8266, w_001_8267, w_001_8268, w_001_8269, w_001_8270, w_001_8271, w_001_8272, w_001_8273, w_001_8274, w_001_8275, w_001_8276, w_001_8277, w_001_8278, w_001_8279, w_001_8280, w_001_8281, w_001_8282, w_001_8283, w_001_8284, w_001_8285, w_001_8286, w_001_8287, w_001_8288, w_001_8289, w_001_8290, w_001_8291, w_001_8292, w_001_8293, w_001_8294, w_001_8295, w_001_8296, w_001_8297, w_001_8298, w_001_8299, w_001_8300, w_001_8301, w_001_8302, w_001_8303, w_001_8304, w_001_8305, w_001_8306, w_001_8307, w_001_8308, w_001_8309, w_001_8310, w_001_8311, w_001_8313, w_001_8314, w_001_8315, w_001_8316, w_001_8317, w_001_8318, w_001_8319, w_001_8320, w_001_8321, w_001_8322, w_001_8323, w_001_8324, w_001_8325, w_001_8326, w_001_8327, w_001_8328, w_001_8329, w_001_8330, w_001_8331, w_001_8332, w_001_8334, w_001_8335, w_001_8336, w_001_8337, w_001_8338, w_001_8339, w_001_8340, w_001_8341, w_001_8342, w_001_8343, w_001_8345, w_001_8346, w_001_8347, w_001_8348, w_001_8350, w_001_8351, w_001_8352, w_001_8353, w_001_8354, w_001_8356, w_001_8357, w_001_8359, w_001_8360, w_001_8361, w_001_8362, w_001_8363, w_001_8364, w_001_8365, w_001_8366, w_001_8367, w_001_8368, w_001_8369, w_001_8370, w_001_8371, w_001_8372, w_001_8373, w_001_8374, w_001_8375, w_001_8376, w_001_8377, w_001_8378, w_001_8379, w_001_8380, w_001_8381, w_001_8382, w_001_8383, w_001_8384, w_001_8385, w_001_8386, w_001_8387, w_001_8388, w_001_8389, w_001_8391, w_001_8392, w_001_8393, w_001_8394, w_001_8395, w_001_8396, w_001_8397, w_001_8398, w_001_8400, w_001_8401, w_001_8402, w_001_8403, w_001_8404, w_001_8405, w_001_8406, w_001_8407, w_001_8408, w_001_8409, w_001_8410, w_001_8411, w_001_8412, w_001_8413, w_001_8414, w_001_8415, w_001_8416, w_001_8417, w_001_8419, w_001_8420, w_001_8421, w_001_8422, w_001_8423, w_001_8424, w_001_8425, w_001_8426, w_001_8427, w_001_8428, w_001_8429, w_001_8430, w_001_8431, w_001_8432, w_001_8433, w_001_8434, w_001_8435, w_001_8436, w_001_8437, w_001_8438, w_001_8439, w_001_8440, w_001_8441, w_001_8442, w_001_8443, w_001_8444, w_001_8445, w_001_8446, w_001_8447, w_001_8448, w_001_8449, w_001_8450, w_001_8451, w_001_8452, w_001_8453, w_001_8454, w_001_8455, w_001_8456, w_001_8457, w_001_8458, w_001_8459, w_001_8460, w_001_8461, w_001_8462, w_001_8463, w_001_8464, w_001_8465, w_001_8466, w_001_8467, w_001_8468, w_001_8470, w_001_8471, w_001_8472, w_001_8473, w_001_8474, w_001_8475, w_001_8477, w_001_8478, w_001_8479, w_001_8480, w_001_8481, w_001_8482, w_001_8483, w_001_8484, w_001_8485, w_001_8486, w_001_8488, w_001_8489, w_001_8490, w_001_8491, w_001_8492, w_001_8493, w_001_8494, w_001_8495, w_001_8496, w_001_8497, w_001_8498, w_001_8500, w_001_8501, w_001_8502, w_001_8503, w_001_8504, w_001_8506, w_001_8507, w_001_8508, w_001_8509, w_001_8510, w_001_8511, w_001_8512, w_001_8513, w_001_8514, w_001_8517, w_001_8518, w_001_8519, w_001_8520, w_001_8521, w_001_8522, w_001_8523, w_001_8524, w_001_8525, w_001_8526, w_001_8527, w_001_8528, w_001_8529, w_001_8530, w_001_8531, w_001_8532, w_001_8533, w_001_8534, w_001_8535, w_001_8536, w_001_8537, w_001_8538, w_001_8539, w_001_8540, w_001_8541, w_001_8542, w_001_8544, w_001_8545, w_001_8546, w_001_8548, w_001_8549, w_001_8550, w_001_8551, w_001_8552, w_001_8553, w_001_8554, w_001_8555, w_001_8556, w_001_8557, w_001_8558, w_001_8559, w_001_8560, w_001_8561, w_001_8562, w_001_8563, w_001_8564, w_001_8565, w_001_8566, w_001_8567, w_001_8568, w_001_8569, w_001_8570, w_001_8571, w_001_8572, w_001_8573, w_001_8574, w_001_8575, w_001_8576, w_001_8577, w_001_8578, w_001_8579, w_001_8580, w_001_8581, w_001_8582, w_001_8583, w_001_8584, w_001_8585, w_001_8586, w_001_8587, w_001_8588, w_001_8589, w_001_8590, w_001_8591, w_001_8592, w_001_8593, w_001_8594, w_001_8598, w_001_8599, w_001_8600, w_001_8601, w_001_8602, w_001_8603, w_001_8604, w_001_8605, w_001_8606, w_001_8607, w_001_8608, w_001_8609, w_001_8610, w_001_8611, w_001_8612, w_001_8614, w_001_8615, w_001_8616, w_001_8617, w_001_8618, w_001_8619, w_001_8620, w_001_8621, w_001_8622, w_001_8623, w_001_8625, w_001_8626, w_001_8627, w_001_8628, w_001_8630, w_001_8631, w_001_8632, w_001_8633, w_001_8634, w_001_8635, w_001_8637, w_001_8638, w_001_8639, w_001_8640, w_001_8641, w_001_8643, w_001_8644, w_001_8645, w_001_8646, w_001_8647, w_001_8648, w_001_8649, w_001_8650, w_001_8652, w_001_8653, w_001_8654, w_001_8655, w_001_8656, w_001_8657, w_001_8658, w_001_8659, w_001_8660, w_001_8661, w_001_8662, w_001_8663, w_001_8664, w_001_8665, w_001_8666, w_001_8668, w_001_8669, w_001_8670, w_001_8671, w_001_8672, w_001_8673, w_001_8674, w_001_8675, w_001_8676, w_001_8677, w_001_8678, w_001_8679, w_001_8680, w_001_8682, w_001_8683, w_001_8684, w_001_8685, w_001_8686, w_001_8687, w_001_8689, w_001_8690, w_001_8691, w_001_8692, w_001_8693, w_001_8694, w_001_8696, w_001_8697, w_001_8699, w_001_8700, w_001_8701, w_001_8703, w_001_8704, w_001_8705, w_001_8706, w_001_8707, w_001_8708, w_001_8709, w_001_8710, w_001_8711, w_001_8712, w_001_8716, w_001_8717, w_001_8718, w_001_8719, w_001_8720, w_001_8721, w_001_8722, w_001_8723, w_001_8724, w_001_8725, w_001_8726, w_001_8727, w_001_8729, w_001_8730, w_001_8731, w_001_8732, w_001_8734, w_001_8735, w_001_8736, w_001_8737, w_001_8738, w_001_8739, w_001_8740, w_001_8741, w_001_8743, w_001_8744, w_001_8745, w_001_8746, w_001_8747, w_001_8748, w_001_8749, w_001_8750, w_001_8751, w_001_8752, w_001_8753, w_001_8754, w_001_8755, w_001_8756, w_001_8757, w_001_8758, w_001_8759, w_001_8760, w_001_8761, w_001_8762, w_001_8763, w_001_8764, w_001_8765, w_001_8766, w_001_8767, w_001_8768, w_001_8769, w_001_8770, w_001_8771, w_001_8772, w_001_8773, w_001_8774, w_001_8775, w_001_8776, w_001_8777, w_001_8778, w_001_8779, w_001_8780, w_001_8781, w_001_8782, w_001_8783, w_001_8784, w_001_8785, w_001_8786, w_001_8787, w_001_8788, w_001_8789, w_001_8790, w_001_8791, w_001_8792, w_001_8793, w_001_8794, w_001_8795, w_001_8797, w_001_8798, w_001_8799, w_001_8800, w_001_8801, w_001_8802, w_001_8804, w_001_8805, w_001_8807, w_001_8808, w_001_8809, w_001_8810, w_001_8811, w_001_8812, w_001_8813, w_001_8814, w_001_8815, w_001_8816, w_001_8817, w_001_8819, w_001_8820, w_001_8821, w_001_8822, w_001_8823, w_001_8824, w_001_8826, w_001_8827, w_001_8829, w_001_8830, w_001_8831, w_001_8832, w_001_8833, w_001_8835, w_001_8836, w_001_8837, w_001_8838, w_001_8839, w_001_8840, w_001_8841, w_001_8842, w_001_8843, w_001_8844, w_001_8845, w_001_8846, w_001_8847, w_001_8849, w_001_8851, w_001_8852, w_001_8853, w_001_8855, w_001_8856, w_001_8857, w_001_8858, w_001_8859, w_001_8860, w_001_8861, w_001_8862, w_001_8863, w_001_8864, w_001_8865, w_001_8866, w_001_8867, w_001_8868, w_001_8869, w_001_8870, w_001_8871, w_001_8872, w_001_8873, w_001_8874, w_001_8875, w_001_8876, w_001_8877, w_001_8878, w_001_8879, w_001_8880, w_001_8881, w_001_8882, w_001_8883, w_001_8884, w_001_8886, w_001_8887, w_001_8889, w_001_8890, w_001_8891, w_001_8892, w_001_8893, w_001_8894, w_001_8895, w_001_8896, w_001_8897, w_001_8898, w_001_8899, w_001_8900, w_001_8901, w_001_8902, w_001_8903, w_001_8904, w_001_8905, w_001_8906, w_001_8907, w_001_8908, w_001_8909, w_001_8910, w_001_8911, w_001_8912, w_001_8913, w_001_8914, w_001_8915, w_001_8916, w_001_8917, w_001_8918, w_001_8919, w_001_8920, w_001_8921, w_001_8922, w_001_8923, w_001_8924, w_001_8925, w_001_8926, w_001_8927, w_001_8928, w_001_8929, w_001_8930, w_001_8931, w_001_8932, w_001_8933, w_001_8934, w_001_8935, w_001_8936, w_001_8937, w_001_8939, w_001_8940, w_001_8941, w_001_8942, w_001_8943, w_001_8944, w_001_8945, w_001_8947, w_001_8948, w_001_8949, w_001_8950, w_001_8952, w_001_8953, w_001_8954, w_001_8955, w_001_8956, w_001_8957, w_001_8958, w_001_8959, w_001_8960, w_001_8962, w_001_8963, w_001_8964, w_001_8965, w_001_8966, w_001_8967, w_001_8968, w_001_8970, w_001_8971, w_001_8972;
  wire w_002_000, w_002_001, w_002_002, w_002_003, w_002_004, w_002_005, w_002_006, w_002_007, w_002_008, w_002_009, w_002_010, w_002_011, w_002_012, w_002_013, w_002_014, w_002_015, w_002_016, w_002_017, w_002_018, w_002_019, w_002_020, w_002_021, w_002_022, w_002_023, w_002_024, w_002_025, w_002_026, w_002_027, w_002_028, w_002_029, w_002_030, w_002_031, w_002_032, w_002_033, w_002_034, w_002_035, w_002_036, w_002_037, w_002_038, w_002_039, w_002_040, w_002_041, w_002_042, w_002_043, w_002_044, w_002_045, w_002_046, w_002_047, w_002_048, w_002_049, w_002_050, w_002_051, w_002_052, w_002_053, w_002_054, w_002_055, w_002_056, w_002_057, w_002_058, w_002_059, w_002_060, w_002_061, w_002_062, w_002_063, w_002_064, w_002_065, w_002_066, w_002_067, w_002_068, w_002_069, w_002_070, w_002_071, w_002_072, w_002_073, w_002_074, w_002_075, w_002_076, w_002_077, w_002_078, w_002_079, w_002_080, w_002_081, w_002_082, w_002_083, w_002_084, w_002_085, w_002_086, w_002_087, w_002_088, w_002_089, w_002_090, w_002_091, w_002_092, w_002_093, w_002_094, w_002_095, w_002_096, w_002_097, w_002_098, w_002_099, w_002_100, w_002_101, w_002_102, w_002_103, w_002_104, w_002_105, w_002_106, w_002_107, w_002_108, w_002_109, w_002_110, w_002_111, w_002_112, w_002_113, w_002_114, w_002_115, w_002_116, w_002_117, w_002_118, w_002_119, w_002_120, w_002_121, w_002_122, w_002_123, w_002_124, w_002_125, w_002_126, w_002_127, w_002_128, w_002_129, w_002_130, w_002_131, w_002_132, w_002_133, w_002_134, w_002_135, w_002_136, w_002_137, w_002_138, w_002_139, w_002_140, w_002_141, w_002_142, w_002_143, w_002_144, w_002_145, w_002_146, w_002_147, w_002_148, w_002_149, w_002_150, w_002_151, w_002_152, w_002_153, w_002_154, w_002_155, w_002_156, w_002_157, w_002_158, w_002_159, w_002_160, w_002_161, w_002_162, w_002_163, w_002_164, w_002_165, w_002_166, w_002_167, w_002_168, w_002_169, w_002_170, w_002_171, w_002_172, w_002_173, w_002_174, w_002_175, w_002_176, w_002_177, w_002_178, w_002_179, w_002_180, w_002_181, w_002_182, w_002_183, w_002_184, w_002_185, w_002_186, w_002_187, w_002_188, w_002_189, w_002_190, w_002_191, w_002_192, w_002_193, w_002_194, w_002_195, w_002_196, w_002_197, w_002_198, w_002_199, w_002_200, w_002_201, w_002_202, w_002_203, w_002_204, w_002_205, w_002_206, w_002_207, w_002_208, w_002_209, w_002_210, w_002_211, w_002_212, w_002_213, w_002_214, w_002_215, w_002_216, w_002_217, w_002_218, w_002_219, w_002_220, w_002_221, w_002_222, w_002_223, w_002_224, w_002_225, w_002_226, w_002_227, w_002_228, w_002_229, w_002_230, w_002_231, w_002_232, w_002_233, w_002_234, w_002_235, w_002_236, w_002_237, w_002_238, w_002_239, w_002_240, w_002_241, w_002_242, w_002_243, w_002_244, w_002_245, w_002_246, w_002_247, w_002_248, w_002_249, w_002_250, w_002_251, w_002_252, w_002_253, w_002_254, w_002_255, w_002_256, w_002_257, w_002_258, w_002_259, w_002_260, w_002_261, w_002_262, w_002_263, w_002_264, w_002_265, w_002_266, w_002_267, w_002_268, w_002_269, w_002_270, w_002_271, w_002_272, w_002_273, w_002_274, w_002_275, w_002_276, w_002_277, w_002_278, w_002_279, w_002_280, w_002_281, w_002_282, w_002_283, w_002_284, w_002_285, w_002_286, w_002_287, w_002_288, w_002_289, w_002_290, w_002_291, w_002_292, w_002_293, w_002_294, w_002_295, w_002_296, w_002_297, w_002_298, w_002_299, w_002_300, w_002_301, w_002_302, w_002_303, w_002_304, w_002_305, w_002_306, w_002_307, w_002_308, w_002_309, w_002_310, w_002_311, w_002_312, w_002_313, w_002_314, w_002_315, w_002_316, w_002_317, w_002_318, w_002_319, w_002_320, w_002_321, w_002_322, w_002_323, w_002_324, w_002_325, w_002_326, w_002_327, w_002_328, w_002_329, w_002_330, w_002_331, w_002_332, w_002_333, w_002_334, w_002_335, w_002_336, w_002_337, w_002_338, w_002_339, w_002_340, w_002_341, w_002_342, w_002_343, w_002_344, w_002_345, w_002_346, w_002_347, w_002_348, w_002_349, w_002_350, w_002_351, w_002_352, w_002_353, w_002_354, w_002_355, w_002_356, w_002_357, w_002_358, w_002_359, w_002_360, w_002_361, w_002_362, w_002_363, w_002_364, w_002_365, w_002_366, w_002_367, w_002_368, w_002_369, w_002_370, w_002_371, w_002_372, w_002_373, w_002_374, w_002_375, w_002_376, w_002_377, w_002_378, w_002_379, w_002_380, w_002_381, w_002_382, w_002_383, w_002_384, w_002_385, w_002_386, w_002_387, w_002_388, w_002_389, w_002_390, w_002_391, w_002_392, w_002_393, w_002_394, w_002_395, w_002_396, w_002_397, w_002_398, w_002_399, w_002_400, w_002_401, w_002_402, w_002_403, w_002_404, w_002_405, w_002_406, w_002_407, w_002_408, w_002_409, w_002_410, w_002_411, w_002_412, w_002_413, w_002_414, w_002_415, w_002_416, w_002_417, w_002_418, w_002_419, w_002_420, w_002_421, w_002_422, w_002_423, w_002_424, w_002_425, w_002_426, w_002_427, w_002_428, w_002_429, w_002_430, w_002_431, w_002_432, w_002_433, w_002_434, w_002_435, w_002_436, w_002_437, w_002_438, w_002_439, w_002_440, w_002_441, w_002_442, w_002_443, w_002_444, w_002_445, w_002_446, w_002_447, w_002_448, w_002_449, w_002_450, w_002_451, w_002_452, w_002_453, w_002_454, w_002_455, w_002_456, w_002_457, w_002_458, w_002_459, w_002_460, w_002_461, w_002_462, w_002_463, w_002_464, w_002_465, w_002_466, w_002_467, w_002_468, w_002_469, w_002_470, w_002_471, w_002_472, w_002_473, w_002_474, w_002_475, w_002_476, w_002_477, w_002_478, w_002_479, w_002_480, w_002_481, w_002_482, w_002_483, w_002_484, w_002_485, w_002_486, w_002_487, w_002_488, w_002_489, w_002_490, w_002_491, w_002_492, w_002_493, w_002_494, w_002_495, w_002_496, w_002_497, w_002_498, w_002_499, w_002_500, w_002_501, w_002_502, w_002_503, w_002_504, w_002_505, w_002_506, w_002_507, w_002_508, w_002_509, w_002_510, w_002_511, w_002_512, w_002_513, w_002_514, w_002_515, w_002_516, w_002_517, w_002_518, w_002_519, w_002_520, w_002_521, w_002_522, w_002_523, w_002_524, w_002_525, w_002_526, w_002_527, w_002_528, w_002_529, w_002_530, w_002_531, w_002_532, w_002_533, w_002_534, w_002_535, w_002_536, w_002_537, w_002_538, w_002_539, w_002_540, w_002_541, w_002_542, w_002_543, w_002_544, w_002_545, w_002_546, w_002_547, w_002_548, w_002_549, w_002_550, w_002_551, w_002_552, w_002_553, w_002_554, w_002_555, w_002_556, w_002_557, w_002_558, w_002_559, w_002_560, w_002_561, w_002_562, w_002_563, w_002_564, w_002_565, w_002_566, w_002_567, w_002_568, w_002_569, w_002_570, w_002_571, w_002_572, w_002_573, w_002_574, w_002_575, w_002_576, w_002_577, w_002_578, w_002_579, w_002_580, w_002_581, w_002_582, w_002_583, w_002_584, w_002_585, w_002_586, w_002_587, w_002_588, w_002_589, w_002_590, w_002_591, w_002_592, w_002_593, w_002_594, w_002_595, w_002_596, w_002_597, w_002_598, w_002_599, w_002_600, w_002_601, w_002_602, w_002_603, w_002_604, w_002_605, w_002_606, w_002_607, w_002_608, w_002_609, w_002_610, w_002_611, w_002_612, w_002_613, w_002_614, w_002_615, w_002_616, w_002_617, w_002_618, w_002_619, w_002_620, w_002_621, w_002_622, w_002_623, w_002_624, w_002_625, w_002_626, w_002_627, w_002_628, w_002_629, w_002_630, w_002_631, w_002_632, w_002_633, w_002_634, w_002_635, w_002_636, w_002_637, w_002_638, w_002_639, w_002_640, w_002_641, w_002_642, w_002_643, w_002_644, w_002_645, w_002_646, w_002_647, w_002_648, w_002_649, w_002_650, w_002_651, w_002_652, w_002_653, w_002_654, w_002_655, w_002_656, w_002_657, w_002_658, w_002_659, w_002_660, w_002_661, w_002_662, w_002_663, w_002_664, w_002_665, w_002_666, w_002_667, w_002_668, w_002_669, w_002_670, w_002_671, w_002_672, w_002_673, w_002_674, w_002_675, w_002_676, w_002_677, w_002_678, w_002_679, w_002_680, w_002_681, w_002_682, w_002_683, w_002_684, w_002_685, w_002_686, w_002_687, w_002_688, w_002_689, w_002_690, w_002_691, w_002_692, w_002_693, w_002_694, w_002_695, w_002_696, w_002_697, w_002_698, w_002_699, w_002_700, w_002_701, w_002_702, w_002_703, w_002_704, w_002_705, w_002_706, w_002_707, w_002_708, w_002_709, w_002_710, w_002_711, w_002_712, w_002_713, w_002_714, w_002_715, w_002_716, w_002_717, w_002_718, w_002_719, w_002_720, w_002_721, w_002_722, w_002_723, w_002_724, w_002_725, w_002_726, w_002_727, w_002_728, w_002_729, w_002_730, w_002_731, w_002_732, w_002_733, w_002_734, w_002_735, w_002_736, w_002_737, w_002_738, w_002_739, w_002_740, w_002_741, w_002_742, w_002_743, w_002_744, w_002_745, w_002_746, w_002_747, w_002_748, w_002_749, w_002_750, w_002_751, w_002_752, w_002_753, w_002_754, w_002_755, w_002_756, w_002_757, w_002_758, w_002_759, w_002_760, w_002_761, w_002_762, w_002_763, w_002_764, w_002_765, w_002_766, w_002_767, w_002_768, w_002_769, w_002_770, w_002_771, w_002_772, w_002_773, w_002_774, w_002_775, w_002_776, w_002_777, w_002_778, w_002_779, w_002_780, w_002_781, w_002_782, w_002_783, w_002_784, w_002_785, w_002_786, w_002_787, w_002_788, w_002_789, w_002_790, w_002_791, w_002_792, w_002_793, w_002_794, w_002_795, w_002_796, w_002_797, w_002_798, w_002_799, w_002_800, w_002_801, w_002_802, w_002_803, w_002_804, w_002_805, w_002_806, w_002_807, w_002_808, w_002_809, w_002_810, w_002_811, w_002_812, w_002_813, w_002_814, w_002_815, w_002_816, w_002_817, w_002_818, w_002_819, w_002_820, w_002_821, w_002_822, w_002_823, w_002_824, w_002_825, w_002_826, w_002_827, w_002_828, w_002_829, w_002_830, w_002_831, w_002_832, w_002_833, w_002_834, w_002_835, w_002_836, w_002_837, w_002_838, w_002_839, w_002_840, w_002_841, w_002_842, w_002_843, w_002_844, w_002_845, w_002_846, w_002_847, w_002_848, w_002_849, w_002_850, w_002_851, w_002_852, w_002_853, w_002_854, w_002_855, w_002_856, w_002_857, w_002_858, w_002_859, w_002_860, w_002_861, w_002_862, w_002_863, w_002_864, w_002_865, w_002_866, w_002_867, w_002_868, w_002_869, w_002_870, w_002_871, w_002_872, w_002_873, w_002_874, w_002_875, w_002_876, w_002_877, w_002_878, w_002_879, w_002_880, w_002_881, w_002_882, w_002_883, w_002_884, w_002_885, w_002_886, w_002_887, w_002_888, w_002_889, w_002_890, w_002_891, w_002_892, w_002_893, w_002_894, w_002_895, w_002_896, w_002_897, w_002_898, w_002_899, w_002_900, w_002_901, w_002_902, w_002_903, w_002_904, w_002_905, w_002_906, w_002_907, w_002_908, w_002_909, w_002_910, w_002_911, w_002_912, w_002_913, w_002_914, w_002_915, w_002_916, w_002_917, w_002_918, w_002_919, w_002_920, w_002_921, w_002_922, w_002_923, w_002_924, w_002_925, w_002_926, w_002_927, w_002_928, w_002_929, w_002_930, w_002_931, w_002_932, w_002_933, w_002_934, w_002_935, w_002_936, w_002_937, w_002_938, w_002_939, w_002_940, w_002_941, w_002_942, w_002_943, w_002_944, w_002_945, w_002_946, w_002_947, w_002_948, w_002_949, w_002_950, w_002_951, w_002_952, w_002_953, w_002_954, w_002_955, w_002_956, w_002_957, w_002_958, w_002_959, w_002_960, w_002_961, w_002_962, w_002_963, w_002_964, w_002_965, w_002_966, w_002_967, w_002_968, w_002_969, w_002_970, w_002_971, w_002_972, w_002_973, w_002_974, w_002_975, w_002_976, w_002_977, w_002_978, w_002_979, w_002_980, w_002_981, w_002_982, w_002_983, w_002_984, w_002_985, w_002_986, w_002_987, w_002_988, w_002_989, w_002_990, w_002_991, w_002_992, w_002_993, w_002_994, w_002_995, w_002_996, w_002_997, w_002_998, w_002_999, w_002_1000, w_002_1001, w_002_1002, w_002_1003, w_002_1004, w_002_1005, w_002_1006, w_002_1007, w_002_1008, w_002_1009, w_002_1010, w_002_1011, w_002_1012, w_002_1013, w_002_1014, w_002_1015, w_002_1016, w_002_1017, w_002_1018, w_002_1019, w_002_1020, w_002_1021, w_002_1022, w_002_1023, w_002_1024, w_002_1025, w_002_1026, w_002_1027, w_002_1028, w_002_1029, w_002_1030, w_002_1031, w_002_1032, w_002_1033, w_002_1034, w_002_1035, w_002_1036, w_002_1037, w_002_1038, w_002_1039, w_002_1040, w_002_1041, w_002_1042, w_002_1043, w_002_1044, w_002_1045, w_002_1046, w_002_1047, w_002_1048, w_002_1049, w_002_1050, w_002_1051, w_002_1052, w_002_1053, w_002_1054, w_002_1055, w_002_1056, w_002_1057, w_002_1058, w_002_1059, w_002_1060, w_002_1061, w_002_1062, w_002_1063, w_002_1064, w_002_1065, w_002_1066, w_002_1067, w_002_1068, w_002_1069, w_002_1070, w_002_1071, w_002_1072, w_002_1073, w_002_1074, w_002_1075, w_002_1076, w_002_1077, w_002_1078, w_002_1079, w_002_1080, w_002_1081, w_002_1082, w_002_1083, w_002_1084, w_002_1085, w_002_1086, w_002_1087, w_002_1088, w_002_1089, w_002_1090, w_002_1091, w_002_1092, w_002_1093, w_002_1094, w_002_1095, w_002_1096, w_002_1097, w_002_1098, w_002_1099, w_002_1101, w_002_1102, w_002_1103, w_002_1104, w_002_1105, w_002_1106, w_002_1107, w_002_1108, w_002_1109, w_002_1110, w_002_1111, w_002_1112, w_002_1113, w_002_1114, w_002_1115, w_002_1116, w_002_1117, w_002_1118, w_002_1119, w_002_1120, w_002_1121, w_002_1122, w_002_1123, w_002_1124, w_002_1125, w_002_1126, w_002_1127, w_002_1128, w_002_1129, w_002_1130, w_002_1131, w_002_1132, w_002_1133, w_002_1134, w_002_1135, w_002_1136, w_002_1137, w_002_1138, w_002_1139, w_002_1140, w_002_1141, w_002_1142, w_002_1143, w_002_1144, w_002_1145, w_002_1146, w_002_1147, w_002_1148, w_002_1149, w_002_1150, w_002_1151, w_002_1152, w_002_1153, w_002_1154, w_002_1155, w_002_1156, w_002_1157, w_002_1158, w_002_1159, w_002_1160, w_002_1161, w_002_1162, w_002_1163, w_002_1164, w_002_1165, w_002_1166, w_002_1167, w_002_1168, w_002_1169, w_002_1170, w_002_1171, w_002_1172, w_002_1173, w_002_1174, w_002_1175, w_002_1176, w_002_1177, w_002_1178, w_002_1179, w_002_1180, w_002_1181, w_002_1182, w_002_1183, w_002_1184, w_002_1185, w_002_1186, w_002_1187, w_002_1188, w_002_1189, w_002_1190, w_002_1191, w_002_1192, w_002_1193, w_002_1194, w_002_1195, w_002_1196, w_002_1197, w_002_1198, w_002_1199, w_002_1200, w_002_1201, w_002_1202, w_002_1203, w_002_1204, w_002_1205, w_002_1206, w_002_1207, w_002_1208, w_002_1209, w_002_1210, w_002_1211, w_002_1212, w_002_1213, w_002_1214, w_002_1215, w_002_1216, w_002_1217, w_002_1218, w_002_1219, w_002_1220, w_002_1221, w_002_1222, w_002_1223, w_002_1224, w_002_1225, w_002_1226, w_002_1227, w_002_1228, w_002_1229, w_002_1230, w_002_1231, w_002_1232, w_002_1233, w_002_1234, w_002_1235, w_002_1236, w_002_1237, w_002_1238, w_002_1239, w_002_1240, w_002_1241, w_002_1242, w_002_1243, w_002_1244, w_002_1245, w_002_1246, w_002_1247, w_002_1248, w_002_1249, w_002_1250, w_002_1251, w_002_1252, w_002_1253, w_002_1254, w_002_1255, w_002_1256, w_002_1257, w_002_1258, w_002_1259, w_002_1260, w_002_1261, w_002_1262, w_002_1263, w_002_1264, w_002_1265, w_002_1266, w_002_1267, w_002_1268, w_002_1269, w_002_1270, w_002_1271, w_002_1272, w_002_1273, w_002_1274, w_002_1275, w_002_1276, w_002_1277, w_002_1278, w_002_1279, w_002_1280, w_002_1281, w_002_1282, w_002_1283, w_002_1284, w_002_1285, w_002_1286, w_002_1287, w_002_1288, w_002_1289, w_002_1290, w_002_1291, w_002_1292, w_002_1293, w_002_1294, w_002_1295, w_002_1296, w_002_1297, w_002_1298, w_002_1299, w_002_1300, w_002_1301, w_002_1302, w_002_1303, w_002_1304, w_002_1305, w_002_1306, w_002_1307, w_002_1308, w_002_1309, w_002_1310, w_002_1311, w_002_1312, w_002_1313, w_002_1314, w_002_1315, w_002_1316, w_002_1317, w_002_1318, w_002_1319, w_002_1320, w_002_1321, w_002_1322, w_002_1323, w_002_1324, w_002_1325, w_002_1326, w_002_1327, w_002_1328, w_002_1329, w_002_1330, w_002_1331, w_002_1332, w_002_1333, w_002_1334, w_002_1335, w_002_1336, w_002_1337, w_002_1338, w_002_1339, w_002_1340, w_002_1341, w_002_1342, w_002_1343, w_002_1344, w_002_1345, w_002_1346, w_002_1347, w_002_1348, w_002_1349, w_002_1350, w_002_1351, w_002_1352, w_002_1353, w_002_1354, w_002_1355, w_002_1356, w_002_1357, w_002_1358, w_002_1359, w_002_1360, w_002_1361, w_002_1362, w_002_1363, w_002_1364, w_002_1365, w_002_1366, w_002_1367, w_002_1368, w_002_1369, w_002_1370, w_002_1371, w_002_1372, w_002_1373, w_002_1374, w_002_1375, w_002_1376, w_002_1377, w_002_1378, w_002_1379, w_002_1380, w_002_1381, w_002_1382, w_002_1383, w_002_1384, w_002_1385, w_002_1386, w_002_1387, w_002_1388, w_002_1389, w_002_1390, w_002_1391, w_002_1392, w_002_1393, w_002_1394, w_002_1395, w_002_1396, w_002_1397, w_002_1398, w_002_1399, w_002_1400, w_002_1401, w_002_1402, w_002_1403, w_002_1404, w_002_1405, w_002_1406, w_002_1407, w_002_1408, w_002_1409, w_002_1410, w_002_1411, w_002_1412, w_002_1413, w_002_1414, w_002_1415, w_002_1416, w_002_1417, w_002_1418, w_002_1419, w_002_1420, w_002_1421, w_002_1422, w_002_1423, w_002_1424, w_002_1425, w_002_1426, w_002_1427, w_002_1428, w_002_1429, w_002_1430, w_002_1431, w_002_1432, w_002_1433, w_002_1434, w_002_1435, w_002_1436, w_002_1437, w_002_1438, w_002_1439, w_002_1440, w_002_1441, w_002_1442, w_002_1443, w_002_1444, w_002_1445, w_002_1446, w_002_1447, w_002_1448, w_002_1449, w_002_1450, w_002_1451, w_002_1452, w_002_1453, w_002_1454, w_002_1455, w_002_1456, w_002_1457, w_002_1458, w_002_1459, w_002_1460, w_002_1461, w_002_1462, w_002_1463, w_002_1464, w_002_1465, w_002_1466, w_002_1467, w_002_1468, w_002_1469, w_002_1470, w_002_1471, w_002_1472, w_002_1473, w_002_1474, w_002_1475, w_002_1476, w_002_1477, w_002_1478, w_002_1479, w_002_1480, w_002_1481, w_002_1482, w_002_1483, w_002_1484, w_002_1485, w_002_1486, w_002_1487, w_002_1488, w_002_1489, w_002_1490, w_002_1491, w_002_1492, w_002_1493, w_002_1494, w_002_1495, w_002_1496, w_002_1497, w_002_1498, w_002_1499, w_002_1500, w_002_1501, w_002_1502, w_002_1503, w_002_1504, w_002_1505, w_002_1506, w_002_1507, w_002_1508, w_002_1509, w_002_1510, w_002_1511, w_002_1512, w_002_1513, w_002_1514, w_002_1515, w_002_1516, w_002_1517, w_002_1518, w_002_1519, w_002_1520, w_002_1521, w_002_1522, w_002_1523, w_002_1524, w_002_1525, w_002_1526, w_002_1527, w_002_1528, w_002_1529, w_002_1530, w_002_1531, w_002_1532, w_002_1533, w_002_1534, w_002_1535, w_002_1536, w_002_1537, w_002_1538, w_002_1539, w_002_1540, w_002_1541, w_002_1542, w_002_1543, w_002_1544, w_002_1545, w_002_1546, w_002_1547, w_002_1548, w_002_1549, w_002_1550, w_002_1551, w_002_1552, w_002_1553, w_002_1554, w_002_1555, w_002_1556, w_002_1557, w_002_1558, w_002_1559, w_002_1560, w_002_1561, w_002_1562, w_002_1563, w_002_1564, w_002_1565, w_002_1566, w_002_1567, w_002_1568, w_002_1569, w_002_1570, w_002_1571, w_002_1572, w_002_1573, w_002_1574, w_002_1575, w_002_1576, w_002_1577, w_002_1578, w_002_1579, w_002_1580, w_002_1581, w_002_1582, w_002_1583, w_002_1584, w_002_1585, w_002_1586, w_002_1587, w_002_1588, w_002_1589, w_002_1590, w_002_1591, w_002_1592, w_002_1593, w_002_1594, w_002_1595, w_002_1596, w_002_1597, w_002_1598, w_002_1599, w_002_1600, w_002_1601, w_002_1602, w_002_1603, w_002_1604, w_002_1605, w_002_1606, w_002_1607, w_002_1608, w_002_1609, w_002_1610, w_002_1611, w_002_1612, w_002_1613, w_002_1614, w_002_1615, w_002_1616, w_002_1617, w_002_1618, w_002_1619, w_002_1620, w_002_1621, w_002_1622, w_002_1623, w_002_1624, w_002_1625, w_002_1626, w_002_1627, w_002_1628, w_002_1629, w_002_1630, w_002_1631, w_002_1632, w_002_1633, w_002_1634, w_002_1635, w_002_1636, w_002_1637, w_002_1638, w_002_1639, w_002_1640, w_002_1641, w_002_1642, w_002_1643, w_002_1644, w_002_1645, w_002_1646, w_002_1647, w_002_1648, w_002_1649, w_002_1650, w_002_1651, w_002_1652, w_002_1653, w_002_1654, w_002_1655, w_002_1656, w_002_1657, w_002_1658, w_002_1659, w_002_1660, w_002_1661, w_002_1662, w_002_1663, w_002_1664, w_002_1665, w_002_1666, w_002_1667, w_002_1668, w_002_1669, w_002_1670, w_002_1671, w_002_1672, w_002_1673, w_002_1674, w_002_1675, w_002_1676, w_002_1677, w_002_1678, w_002_1679, w_002_1680, w_002_1681, w_002_1682, w_002_1683, w_002_1684, w_002_1685, w_002_1686, w_002_1687, w_002_1688, w_002_1689, w_002_1690, w_002_1691, w_002_1692, w_002_1693, w_002_1694, w_002_1695, w_002_1696, w_002_1697, w_002_1698, w_002_1699, w_002_1700, w_002_1701, w_002_1702, w_002_1703, w_002_1704, w_002_1705, w_002_1706, w_002_1707, w_002_1708, w_002_1709, w_002_1710, w_002_1711, w_002_1712, w_002_1713, w_002_1714, w_002_1715, w_002_1716, w_002_1717, w_002_1718, w_002_1719, w_002_1720, w_002_1721, w_002_1722, w_002_1723, w_002_1724, w_002_1725, w_002_1726, w_002_1727, w_002_1728, w_002_1729, w_002_1730, w_002_1731, w_002_1732, w_002_1733, w_002_1734, w_002_1735, w_002_1736, w_002_1737, w_002_1738, w_002_1739, w_002_1740, w_002_1741, w_002_1742, w_002_1743, w_002_1744, w_002_1745, w_002_1746, w_002_1747, w_002_1748, w_002_1749, w_002_1750, w_002_1751, w_002_1752, w_002_1753, w_002_1754, w_002_1755, w_002_1756, w_002_1757, w_002_1758, w_002_1759, w_002_1760, w_002_1761, w_002_1762, w_002_1763, w_002_1764, w_002_1765, w_002_1766, w_002_1767, w_002_1768, w_002_1769, w_002_1770, w_002_1771, w_002_1772, w_002_1773, w_002_1774, w_002_1775, w_002_1776, w_002_1777, w_002_1778, w_002_1779, w_002_1780, w_002_1781, w_002_1782, w_002_1783, w_002_1784, w_002_1785, w_002_1786, w_002_1787, w_002_1788, w_002_1789, w_002_1790, w_002_1791, w_002_1792, w_002_1793, w_002_1794, w_002_1795, w_002_1796, w_002_1797, w_002_1798, w_002_1799, w_002_1800, w_002_1801, w_002_1802, w_002_1803, w_002_1804, w_002_1805, w_002_1806, w_002_1807, w_002_1808, w_002_1809, w_002_1810, w_002_1811, w_002_1812, w_002_1813, w_002_1814, w_002_1815, w_002_1816, w_002_1817, w_002_1818, w_002_1819, w_002_1820, w_002_1821, w_002_1822, w_002_1823, w_002_1824, w_002_1825, w_002_1826, w_002_1827, w_002_1828, w_002_1829, w_002_1830, w_002_1831, w_002_1832, w_002_1833, w_002_1834, w_002_1835, w_002_1836, w_002_1837, w_002_1838, w_002_1839, w_002_1840, w_002_1841, w_002_1842, w_002_1843, w_002_1844, w_002_1845, w_002_1846, w_002_1847, w_002_1848, w_002_1849, w_002_1850, w_002_1851, w_002_1852, w_002_1853, w_002_1854, w_002_1855, w_002_1856, w_002_1857, w_002_1858, w_002_1859, w_002_1860, w_002_1861, w_002_1862, w_002_1863, w_002_1864, w_002_1865, w_002_1866, w_002_1867, w_002_1868, w_002_1869, w_002_1870, w_002_1871, w_002_1872, w_002_1873, w_002_1874, w_002_1875, w_002_1876, w_002_1877, w_002_1878, w_002_1879, w_002_1880, w_002_1881, w_002_1882, w_002_1883, w_002_1884, w_002_1885, w_002_1886, w_002_1887, w_002_1888, w_002_1889, w_002_1890, w_002_1891, w_002_1892, w_002_1893, w_002_1894, w_002_1895, w_002_1896, w_002_1897, w_002_1898, w_002_1899, w_002_1900, w_002_1901, w_002_1902, w_002_1903, w_002_1904, w_002_1905, w_002_1906, w_002_1907, w_002_1908, w_002_1909, w_002_1910, w_002_1911, w_002_1912, w_002_1913, w_002_1914, w_002_1915, w_002_1916, w_002_1917, w_002_1918, w_002_1919, w_002_1920, w_002_1921, w_002_1922, w_002_1923, w_002_1924, w_002_1925, w_002_1926, w_002_1927, w_002_1928, w_002_1929, w_002_1930, w_002_1931, w_002_1932, w_002_1933, w_002_1934, w_002_1935, w_002_1936, w_002_1937, w_002_1938, w_002_1939, w_002_1940, w_002_1941, w_002_1942, w_002_1943, w_002_1944, w_002_1945, w_002_1946, w_002_1947, w_002_1948, w_002_1949, w_002_1950, w_002_1951, w_002_1952, w_002_1953, w_002_1954, w_002_1955, w_002_1956, w_002_1957, w_002_1958, w_002_1959, w_002_1960, w_002_1961, w_002_1962, w_002_1963, w_002_1964, w_002_1965, w_002_1966, w_002_1967, w_002_1968, w_002_1969, w_002_1970, w_002_1971, w_002_1972, w_002_1973, w_002_1974, w_002_1975, w_002_1976, w_002_1977, w_002_1978, w_002_1979, w_002_1980, w_002_1981, w_002_1982, w_002_1983, w_002_1984, w_002_1985, w_002_1986, w_002_1987, w_002_1988, w_002_1989, w_002_1990, w_002_1991, w_002_1992, w_002_1993, w_002_1994, w_002_1995, w_002_1996, w_002_1997, w_002_1998, w_002_1999, w_002_2000, w_002_2001, w_002_2002, w_002_2003, w_002_2004, w_002_2005, w_002_2006, w_002_2007, w_002_2008, w_002_2009, w_002_2010, w_002_2011, w_002_2012, w_002_2013, w_002_2014, w_002_2015, w_002_2016, w_002_2017, w_002_2018, w_002_2019, w_002_2020, w_002_2021, w_002_2022, w_002_2023, w_002_2024, w_002_2025, w_002_2026, w_002_2027, w_002_2028, w_002_2029, w_002_2030, w_002_2031, w_002_2032, w_002_2033, w_002_2034, w_002_2035, w_002_2036, w_002_2037, w_002_2038, w_002_2039, w_002_2040, w_002_2041, w_002_2042, w_002_2043, w_002_2044, w_002_2045, w_002_2046, w_002_2047, w_002_2048, w_002_2049, w_002_2050, w_002_2051, w_002_2052, w_002_2053, w_002_2054, w_002_2055, w_002_2056, w_002_2057, w_002_2058, w_002_2059, w_002_2060, w_002_2061, w_002_2062, w_002_2063, w_002_2064, w_002_2065, w_002_2066, w_002_2067, w_002_2068, w_002_2069, w_002_2070, w_002_2071, w_002_2072, w_002_2073, w_002_2074, w_002_2075, w_002_2076, w_002_2077, w_002_2078, w_002_2079, w_002_2080, w_002_2081, w_002_2082, w_002_2083, w_002_2084, w_002_2085, w_002_2086, w_002_2087, w_002_2088, w_002_2089, w_002_2090, w_002_2091, w_002_2092, w_002_2093, w_002_2094, w_002_2095, w_002_2096, w_002_2097, w_002_2098, w_002_2099, w_002_2100, w_002_2101, w_002_2102, w_002_2103, w_002_2104, w_002_2105, w_002_2106, w_002_2107, w_002_2108, w_002_2109, w_002_2110, w_002_2111, w_002_2112, w_002_2113, w_002_2114, w_002_2115, w_002_2116, w_002_2117, w_002_2118, w_002_2119, w_002_2120, w_002_2121, w_002_2122, w_002_2123, w_002_2124, w_002_2125, w_002_2126, w_002_2127, w_002_2128, w_002_2129, w_002_2130, w_002_2131, w_002_2132, w_002_2133, w_002_2134, w_002_2135, w_002_2136, w_002_2137, w_002_2138, w_002_2139, w_002_2140, w_002_2141, w_002_2142, w_002_2143, w_002_2144, w_002_2145, w_002_2146, w_002_2147, w_002_2148, w_002_2149, w_002_2150, w_002_2151, w_002_2152, w_002_2153, w_002_2154, w_002_2155, w_002_2156, w_002_2157, w_002_2158, w_002_2159, w_002_2160, w_002_2161, w_002_2162, w_002_2163, w_002_2164, w_002_2165, w_002_2166, w_002_2167, w_002_2168, w_002_2169, w_002_2170, w_002_2171, w_002_2172, w_002_2173, w_002_2174, w_002_2175, w_002_2176, w_002_2177, w_002_2178, w_002_2179, w_002_2180, w_002_2181, w_002_2182, w_002_2183, w_002_2184, w_002_2185, w_002_2186, w_002_2187, w_002_2188, w_002_2189, w_002_2190, w_002_2191, w_002_2192, w_002_2193, w_002_2194, w_002_2195, w_002_2196, w_002_2197, w_002_2198, w_002_2199, w_002_2200, w_002_2201, w_002_2202, w_002_2203, w_002_2204, w_002_2205, w_002_2206, w_002_2207, w_002_2208, w_002_2209, w_002_2210, w_002_2211, w_002_2212, w_002_2213, w_002_2214, w_002_2215, w_002_2216, w_002_2217, w_002_2218, w_002_2219, w_002_2220, w_002_2221, w_002_2222, w_002_2223, w_002_2224, w_002_2225, w_002_2226, w_002_2227, w_002_2228, w_002_2229, w_002_2230, w_002_2231, w_002_2232, w_002_2233, w_002_2234, w_002_2235, w_002_2236, w_002_2237, w_002_2238, w_002_2239, w_002_2240, w_002_2241, w_002_2242, w_002_2243, w_002_2244, w_002_2245, w_002_2246, w_002_2247, w_002_2248, w_002_2249, w_002_2250, w_002_2251, w_002_2252, w_002_2253, w_002_2254, w_002_2255, w_002_2256, w_002_2257, w_002_2258, w_002_2259, w_002_2260, w_002_2261, w_002_2262, w_002_2263, w_002_2264, w_002_2265, w_002_2266, w_002_2267, w_002_2268, w_002_2269, w_002_2270, w_002_2271, w_002_2272, w_002_2273, w_002_2274, w_002_2275, w_002_2276, w_002_2277, w_002_2278, w_002_2279, w_002_2280, w_002_2281, w_002_2282, w_002_2283, w_002_2284, w_002_2285, w_002_2286, w_002_2287, w_002_2288, w_002_2289, w_002_2290, w_002_2291, w_002_2292, w_002_2293, w_002_2294, w_002_2295, w_002_2296, w_002_2297, w_002_2298, w_002_2299, w_002_2300, w_002_2301, w_002_2302, w_002_2303, w_002_2304, w_002_2305, w_002_2306, w_002_2307, w_002_2308, w_002_2309, w_002_2310, w_002_2311, w_002_2312, w_002_2313, w_002_2314, w_002_2315, w_002_2316, w_002_2317, w_002_2318, w_002_2319, w_002_2320, w_002_2321, w_002_2322, w_002_2323, w_002_2324, w_002_2325, w_002_2326, w_002_2327, w_002_2328, w_002_2329, w_002_2330, w_002_2331, w_002_2332, w_002_2333, w_002_2334, w_002_2335, w_002_2336, w_002_2337, w_002_2338, w_002_2339, w_002_2340, w_002_2341, w_002_2342, w_002_2343, w_002_2344, w_002_2345, w_002_2346, w_002_2347, w_002_2348, w_002_2349, w_002_2350, w_002_2351, w_002_2352, w_002_2353, w_002_2354, w_002_2355, w_002_2356, w_002_2357, w_002_2358, w_002_2359, w_002_2360, w_002_2361, w_002_2362, w_002_2363, w_002_2364, w_002_2365, w_002_2366, w_002_2367, w_002_2368, w_002_2369, w_002_2370, w_002_2371, w_002_2372, w_002_2373, w_002_2374, w_002_2375, w_002_2376, w_002_2377, w_002_2378, w_002_2379, w_002_2380, w_002_2381, w_002_2382, w_002_2383, w_002_2384, w_002_2385, w_002_2386, w_002_2387, w_002_2388, w_002_2389, w_002_2390, w_002_2391, w_002_2392, w_002_2393, w_002_2394, w_002_2395, w_002_2396, w_002_2397, w_002_2398, w_002_2399, w_002_2400, w_002_2401, w_002_2402, w_002_2403, w_002_2404, w_002_2405, w_002_2406, w_002_2407, w_002_2408, w_002_2409, w_002_2410, w_002_2411, w_002_2412, w_002_2413, w_002_2414, w_002_2415, w_002_2416, w_002_2417, w_002_2418, w_002_2419, w_002_2420, w_002_2421, w_002_2422, w_002_2423, w_002_2424, w_002_2425, w_002_2426, w_002_2427, w_002_2428, w_002_2429, w_002_2430, w_002_2431, w_002_2432, w_002_2433, w_002_2434, w_002_2435, w_002_2436, w_002_2437, w_002_2438, w_002_2439, w_002_2440, w_002_2441, w_002_2442, w_002_2443, w_002_2444, w_002_2445, w_002_2446, w_002_2447, w_002_2448, w_002_2449, w_002_2450, w_002_2451, w_002_2452, w_002_2453, w_002_2454, w_002_2455, w_002_2456, w_002_2457, w_002_2458, w_002_2459, w_002_2460, w_002_2461, w_002_2462, w_002_2463, w_002_2464, w_002_2465, w_002_2466, w_002_2467, w_002_2468, w_002_2469, w_002_2470, w_002_2471, w_002_2472, w_002_2473, w_002_2474, w_002_2475, w_002_2476, w_002_2477, w_002_2478, w_002_2479, w_002_2480, w_002_2481, w_002_2482, w_002_2483, w_002_2484, w_002_2485, w_002_2486, w_002_2487, w_002_2488, w_002_2489, w_002_2490, w_002_2491, w_002_2492, w_002_2493, w_002_2494, w_002_2495, w_002_2496, w_002_2497, w_002_2498, w_002_2499, w_002_2500, w_002_2501, w_002_2502, w_002_2503, w_002_2504, w_002_2505, w_002_2506, w_002_2507, w_002_2508, w_002_2509, w_002_2510, w_002_2511, w_002_2512, w_002_2513, w_002_2514, w_002_2515, w_002_2516, w_002_2517, w_002_2518, w_002_2519, w_002_2520, w_002_2521, w_002_2522, w_002_2523, w_002_2524, w_002_2525, w_002_2526, w_002_2527, w_002_2528, w_002_2529, w_002_2530, w_002_2531, w_002_2532, w_002_2533, w_002_2534, w_002_2535, w_002_2536, w_002_2537, w_002_2538, w_002_2539, w_002_2540, w_002_2541, w_002_2542, w_002_2543, w_002_2544, w_002_2545, w_002_2546, w_002_2547, w_002_2548, w_002_2549, w_002_2550, w_002_2551, w_002_2552, w_002_2553, w_002_2554, w_002_2555, w_002_2556, w_002_2557, w_002_2558, w_002_2559, w_002_2560, w_002_2561, w_002_2562, w_002_2563, w_002_2564, w_002_2565, w_002_2566, w_002_2567, w_002_2568, w_002_2569, w_002_2570, w_002_2571, w_002_2572, w_002_2573, w_002_2574, w_002_2575, w_002_2576, w_002_2577, w_002_2578, w_002_2579, w_002_2580, w_002_2581, w_002_2582, w_002_2583, w_002_2584, w_002_2585, w_002_2586, w_002_2587, w_002_2588, w_002_2589, w_002_2590, w_002_2591, w_002_2592, w_002_2593, w_002_2594, w_002_2595, w_002_2596, w_002_2597, w_002_2598, w_002_2599, w_002_2600, w_002_2601, w_002_2602, w_002_2603, w_002_2604, w_002_2605, w_002_2606, w_002_2607, w_002_2608, w_002_2609, w_002_2610, w_002_2611, w_002_2612, w_002_2613, w_002_2614, w_002_2615, w_002_2616, w_002_2617, w_002_2618, w_002_2619, w_002_2620, w_002_2621, w_002_2622, w_002_2623, w_002_2624, w_002_2625, w_002_2626, w_002_2627, w_002_2628, w_002_2629, w_002_2630, w_002_2631, w_002_2632, w_002_2633, w_002_2634, w_002_2635, w_002_2636, w_002_2637, w_002_2638, w_002_2639, w_002_2640, w_002_2641, w_002_2642, w_002_2643, w_002_2644, w_002_2645, w_002_2646, w_002_2647, w_002_2648, w_002_2649, w_002_2650, w_002_2651, w_002_2652, w_002_2653, w_002_2654, w_002_2655, w_002_2656, w_002_2657, w_002_2658, w_002_2659, w_002_2660, w_002_2661, w_002_2662, w_002_2663, w_002_2664, w_002_2665, w_002_2666, w_002_2667, w_002_2668, w_002_2669, w_002_2670, w_002_2671, w_002_2672, w_002_2673, w_002_2674, w_002_2675, w_002_2676, w_002_2677, w_002_2678, w_002_2679, w_002_2680, w_002_2681, w_002_2682, w_002_2683, w_002_2684, w_002_2685, w_002_2686, w_002_2687, w_002_2688, w_002_2689, w_002_2690, w_002_2691, w_002_2692, w_002_2693, w_002_2694, w_002_2695, w_002_2696, w_002_2697, w_002_2698, w_002_2699, w_002_2700, w_002_2701, w_002_2702, w_002_2703, w_002_2704, w_002_2705, w_002_2706, w_002_2707, w_002_2708, w_002_2709, w_002_2710, w_002_2711, w_002_2712, w_002_2713, w_002_2714, w_002_2715, w_002_2716, w_002_2717, w_002_2718, w_002_2719, w_002_2720, w_002_2721, w_002_2722, w_002_2723, w_002_2724, w_002_2725, w_002_2726, w_002_2727, w_002_2728, w_002_2729, w_002_2730, w_002_2731, w_002_2732, w_002_2733, w_002_2734, w_002_2735, w_002_2736, w_002_2737, w_002_2738, w_002_2739, w_002_2740, w_002_2741, w_002_2742, w_002_2743, w_002_2744, w_002_2745, w_002_2746, w_002_2747, w_002_2748, w_002_2749, w_002_2750, w_002_2751, w_002_2752, w_002_2753, w_002_2754, w_002_2755, w_002_2756, w_002_2757, w_002_2758, w_002_2759, w_002_2760, w_002_2761, w_002_2762, w_002_2763, w_002_2764, w_002_2765, w_002_2766, w_002_2767, w_002_2768, w_002_2769, w_002_2770, w_002_2771, w_002_2772, w_002_2773, w_002_2774, w_002_2775, w_002_2776, w_002_2777, w_002_2778, w_002_2779, w_002_2780, w_002_2781, w_002_2782, w_002_2783, w_002_2784, w_002_2785, w_002_2786, w_002_2787, w_002_2788, w_002_2789, w_002_2790, w_002_2791, w_002_2792, w_002_2793, w_002_2794, w_002_2795, w_002_2796, w_002_2797, w_002_2798, w_002_2799, w_002_2800, w_002_2801, w_002_2802, w_002_2803, w_002_2804, w_002_2805, w_002_2806, w_002_2807, w_002_2808, w_002_2809, w_002_2810, w_002_2811, w_002_2812, w_002_2813, w_002_2814, w_002_2815, w_002_2816, w_002_2817, w_002_2818, w_002_2819, w_002_2820, w_002_2821, w_002_2822, w_002_2823, w_002_2824, w_002_2825, w_002_2826, w_002_2827, w_002_2828, w_002_2829, w_002_2830, w_002_2831, w_002_2832, w_002_2833, w_002_2834, w_002_2835, w_002_2836, w_002_2837, w_002_2838, w_002_2839, w_002_2840, w_002_2841, w_002_2842, w_002_2843, w_002_2844, w_002_2845, w_002_2846, w_002_2847, w_002_2848, w_002_2849, w_002_2850, w_002_2851, w_002_2852, w_002_2853, w_002_2854, w_002_2855, w_002_2856, w_002_2857, w_002_2858, w_002_2859, w_002_2860, w_002_2861, w_002_2862, w_002_2863, w_002_2864, w_002_2865, w_002_2866, w_002_2867, w_002_2868, w_002_2869, w_002_2870, w_002_2871, w_002_2872, w_002_2873, w_002_2874, w_002_2875, w_002_2876, w_002_2877, w_002_2878, w_002_2879, w_002_2880, w_002_2881, w_002_2882, w_002_2883, w_002_2884, w_002_2885, w_002_2886, w_002_2887, w_002_2888, w_002_2889, w_002_2890, w_002_2891, w_002_2892, w_002_2893, w_002_2894, w_002_2895, w_002_2896, w_002_2897, w_002_2898, w_002_2899, w_002_2900, w_002_2901, w_002_2902, w_002_2903, w_002_2904, w_002_2905, w_002_2906, w_002_2907, w_002_2908, w_002_2909, w_002_2910, w_002_2911, w_002_2912, w_002_2913, w_002_2914, w_002_2915, w_002_2916, w_002_2917, w_002_2918, w_002_2919, w_002_2920, w_002_2921, w_002_2922, w_002_2923, w_002_2924, w_002_2925, w_002_2926, w_002_2927, w_002_2928, w_002_2929, w_002_2930, w_002_2931, w_002_2932, w_002_2933, w_002_2934, w_002_2935, w_002_2936, w_002_2937, w_002_2938, w_002_2939, w_002_2940, w_002_2941, w_002_2942, w_002_2943, w_002_2944, w_002_2945, w_002_2946, w_002_2947, w_002_2948, w_002_2949, w_002_2950, w_002_2951, w_002_2952, w_002_2953, w_002_2954, w_002_2955, w_002_2956, w_002_2957, w_002_2958, w_002_2959, w_002_2960, w_002_2961, w_002_2962, w_002_2963, w_002_2964, w_002_2965, w_002_2966, w_002_2967, w_002_2968, w_002_2969, w_002_2970, w_002_2971, w_002_2972, w_002_2973, w_002_2974, w_002_2975, w_002_2976, w_002_2977, w_002_2979, w_002_2980, w_002_2981, w_002_2982, w_002_2983, w_002_2984, w_002_2985, w_002_2986, w_002_2987, w_002_2988, w_002_2989, w_002_2990, w_002_2991, w_002_2992, w_002_2993, w_002_2994, w_002_2995, w_002_2996, w_002_2997, w_002_2998, w_002_2999, w_002_3000, w_002_3001, w_002_3002, w_002_3003, w_002_3004, w_002_3005, w_002_3006, w_002_3007, w_002_3008, w_002_3009, w_002_3010, w_002_3011, w_002_3012, w_002_3013, w_002_3014, w_002_3015, w_002_3016, w_002_3017, w_002_3018, w_002_3019, w_002_3020, w_002_3021, w_002_3022, w_002_3023, w_002_3024, w_002_3025, w_002_3026, w_002_3027, w_002_3028, w_002_3029, w_002_3030, w_002_3031, w_002_3032, w_002_3033, w_002_3034, w_002_3035, w_002_3036, w_002_3037, w_002_3038, w_002_3039, w_002_3040, w_002_3041, w_002_3042, w_002_3043, w_002_3044, w_002_3045, w_002_3046, w_002_3047, w_002_3048, w_002_3049, w_002_3050, w_002_3051, w_002_3052, w_002_3053, w_002_3054, w_002_3055, w_002_3056, w_002_3057, w_002_3058, w_002_3059, w_002_3060, w_002_3061, w_002_3062, w_002_3063, w_002_3064, w_002_3065, w_002_3066, w_002_3067, w_002_3068, w_002_3069, w_002_3070, w_002_3071, w_002_3072, w_002_3073, w_002_3074, w_002_3075, w_002_3076, w_002_3077, w_002_3078, w_002_3079, w_002_3080, w_002_3081, w_002_3082, w_002_3083, w_002_3084, w_002_3085, w_002_3086, w_002_3087, w_002_3088, w_002_3089, w_002_3090, w_002_3091, w_002_3092, w_002_3093, w_002_3094, w_002_3095, w_002_3096, w_002_3097, w_002_3098, w_002_3099, w_002_3100, w_002_3101, w_002_3102, w_002_3103, w_002_3104, w_002_3105, w_002_3106, w_002_3107, w_002_3108, w_002_3109, w_002_3110, w_002_3111, w_002_3112, w_002_3113, w_002_3114, w_002_3115, w_002_3116, w_002_3117, w_002_3118, w_002_3119, w_002_3120, w_002_3121, w_002_3122, w_002_3123, w_002_3124, w_002_3125, w_002_3126, w_002_3127, w_002_3128, w_002_3129, w_002_3130, w_002_3131, w_002_3132, w_002_3133, w_002_3134, w_002_3135, w_002_3136, w_002_3137, w_002_3138, w_002_3139, w_002_3140, w_002_3141, w_002_3142, w_002_3143, w_002_3144, w_002_3145, w_002_3146, w_002_3147, w_002_3148, w_002_3149, w_002_3150, w_002_3151, w_002_3152, w_002_3153, w_002_3154, w_002_3155, w_002_3156, w_002_3157, w_002_3158, w_002_3159, w_002_3160, w_002_3161, w_002_3162, w_002_3163, w_002_3164, w_002_3165, w_002_3166, w_002_3167, w_002_3168, w_002_3169, w_002_3170, w_002_3171, w_002_3172, w_002_3173, w_002_3174, w_002_3175, w_002_3176, w_002_3177, w_002_3178, w_002_3179, w_002_3180, w_002_3181, w_002_3182, w_002_3183, w_002_3184, w_002_3185, w_002_3186, w_002_3187, w_002_3188, w_002_3189, w_002_3190, w_002_3191, w_002_3192, w_002_3193, w_002_3194, w_002_3195, w_002_3196, w_002_3197, w_002_3198, w_002_3199, w_002_3200, w_002_3201, w_002_3202, w_002_3203, w_002_3204, w_002_3205, w_002_3206, w_002_3207, w_002_3208, w_002_3209, w_002_3210, w_002_3211, w_002_3212, w_002_3213, w_002_3214, w_002_3215, w_002_3216, w_002_3217, w_002_3218, w_002_3219, w_002_3220, w_002_3221, w_002_3222, w_002_3223, w_002_3224, w_002_3225, w_002_3226, w_002_3227, w_002_3228, w_002_3229, w_002_3230, w_002_3231, w_002_3232, w_002_3233, w_002_3234, w_002_3235, w_002_3236, w_002_3237, w_002_3238, w_002_3239, w_002_3240, w_002_3241, w_002_3242, w_002_3243, w_002_3244, w_002_3245, w_002_3246, w_002_3247, w_002_3248, w_002_3249, w_002_3250, w_002_3251, w_002_3252, w_002_3253, w_002_3254, w_002_3255, w_002_3256, w_002_3257, w_002_3258, w_002_3259, w_002_3260, w_002_3261, w_002_3262, w_002_3263, w_002_3264, w_002_3265, w_002_3266, w_002_3267, w_002_3268, w_002_3269, w_002_3270, w_002_3271, w_002_3272, w_002_3273, w_002_3274, w_002_3275, w_002_3276, w_002_3277, w_002_3278, w_002_3279, w_002_3280, w_002_3282, w_002_3283, w_002_3284, w_002_3285, w_002_3286, w_002_3287, w_002_3288, w_002_3289, w_002_3290, w_002_3291, w_002_3292, w_002_3293, w_002_3294, w_002_3295, w_002_3296, w_002_3297, w_002_3298, w_002_3299, w_002_3300, w_002_3301, w_002_3302, w_002_3303, w_002_3304, w_002_3305, w_002_3306, w_002_3307, w_002_3308, w_002_3309, w_002_3310, w_002_3311, w_002_3312, w_002_3313, w_002_3314, w_002_3315, w_002_3316, w_002_3317, w_002_3318, w_002_3319, w_002_3320, w_002_3321, w_002_3322, w_002_3323, w_002_3324, w_002_3325, w_002_3326, w_002_3327, w_002_3328, w_002_3329, w_002_3330, w_002_3331, w_002_3332, w_002_3333, w_002_3334, w_002_3335, w_002_3336, w_002_3337, w_002_3338, w_002_3339, w_002_3340, w_002_3341, w_002_3342, w_002_3343, w_002_3344, w_002_3345, w_002_3346, w_002_3347, w_002_3348, w_002_3349, w_002_3350, w_002_3351, w_002_3352, w_002_3353, w_002_3354, w_002_3355, w_002_3356, w_002_3357, w_002_3358, w_002_3359, w_002_3360, w_002_3361, w_002_3362, w_002_3363, w_002_3364, w_002_3365, w_002_3366, w_002_3367, w_002_3368, w_002_3369, w_002_3370, w_002_3371, w_002_3372, w_002_3373, w_002_3374, w_002_3375, w_002_3376, w_002_3377, w_002_3378, w_002_3379, w_002_3380, w_002_3381, w_002_3382, w_002_3383, w_002_3384, w_002_3385, w_002_3386, w_002_3387, w_002_3388, w_002_3389, w_002_3390, w_002_3391, w_002_3392, w_002_3393, w_002_3394, w_002_3395, w_002_3396, w_002_3397, w_002_3398, w_002_3399, w_002_3400, w_002_3401, w_002_3402, w_002_3403, w_002_3404, w_002_3405, w_002_3406, w_002_3407, w_002_3408, w_002_3409, w_002_3410, w_002_3411, w_002_3412, w_002_3413, w_002_3414, w_002_3415, w_002_3416, w_002_3417, w_002_3418, w_002_3419, w_002_3420, w_002_3421, w_002_3422;
  wire w_003_000, w_003_001, w_003_002, w_003_003, w_003_004, w_003_005, w_003_006, w_003_007, w_003_008, w_003_009, w_003_010, w_003_011, w_003_012, w_003_013, w_003_014, w_003_015, w_003_016, w_003_017, w_003_018, w_003_019, w_003_020, w_003_021, w_003_022, w_003_023, w_003_024, w_003_025, w_003_026, w_003_027, w_003_028, w_003_029, w_003_030, w_003_031, w_003_032, w_003_033, w_003_034, w_003_035, w_003_036, w_003_037, w_003_038, w_003_039, w_003_040, w_003_041, w_003_042, w_003_043, w_003_044, w_003_045, w_003_046, w_003_047, w_003_048, w_003_049, w_003_050, w_003_051, w_003_052, w_003_053, w_003_054, w_003_055, w_003_056, w_003_057, w_003_058, w_003_059, w_003_060, w_003_061, w_003_062, w_003_063, w_003_064, w_003_065, w_003_066, w_003_067, w_003_068, w_003_069, w_003_070, w_003_071, w_003_072, w_003_073, w_003_074, w_003_075, w_003_076, w_003_077, w_003_078, w_003_079, w_003_080, w_003_081, w_003_082, w_003_083, w_003_084, w_003_085, w_003_086, w_003_087, w_003_088, w_003_089, w_003_090, w_003_091, w_003_092, w_003_093, w_003_094, w_003_095, w_003_096, w_003_097, w_003_098, w_003_099, w_003_100, w_003_101, w_003_102, w_003_103, w_003_104, w_003_105, w_003_106, w_003_107, w_003_108, w_003_109, w_003_110, w_003_111, w_003_112, w_003_113, w_003_114, w_003_115, w_003_116, w_003_117, w_003_118, w_003_119, w_003_120, w_003_121, w_003_122, w_003_123, w_003_124, w_003_125, w_003_126, w_003_127, w_003_128, w_003_129, w_003_130, w_003_131, w_003_132, w_003_133, w_003_134, w_003_135, w_003_136, w_003_137, w_003_138, w_003_139, w_003_140, w_003_141, w_003_142, w_003_143, w_003_145, w_003_146, w_003_147, w_003_148, w_003_149, w_003_150, w_003_151, w_003_152, w_003_153, w_003_154, w_003_155, w_003_156, w_003_157, w_003_158, w_003_159, w_003_160, w_003_161, w_003_162, w_003_163, w_003_164, w_003_165, w_003_166, w_003_167, w_003_168, w_003_169, w_003_170, w_003_171, w_003_172, w_003_173, w_003_174, w_003_175, w_003_176, w_003_177, w_003_178, w_003_179, w_003_180, w_003_181, w_003_182, w_003_183, w_003_184, w_003_185, w_003_186, w_003_187, w_003_188, w_003_189, w_003_190, w_003_191, w_003_192, w_003_193, w_003_194, w_003_195, w_003_196, w_003_197, w_003_198, w_003_199, w_003_200, w_003_201, w_003_202, w_003_203, w_003_204, w_003_205, w_003_206, w_003_207, w_003_208, w_003_209, w_003_210, w_003_211, w_003_212, w_003_213, w_003_214, w_003_215, w_003_216, w_003_217, w_003_218, w_003_219, w_003_220, w_003_221, w_003_222, w_003_223, w_003_224, w_003_225, w_003_226, w_003_227, w_003_228, w_003_229, w_003_230, w_003_231, w_003_232, w_003_233, w_003_234, w_003_235, w_003_236, w_003_237, w_003_238, w_003_239, w_003_240, w_003_241, w_003_242, w_003_243, w_003_244, w_003_245, w_003_246, w_003_247, w_003_248, w_003_249, w_003_250, w_003_251, w_003_252, w_003_253, w_003_254, w_003_255, w_003_256, w_003_257, w_003_258, w_003_259, w_003_260, w_003_261, w_003_262, w_003_263, w_003_264, w_003_265, w_003_266, w_003_267, w_003_268, w_003_269, w_003_270, w_003_271, w_003_272, w_003_273, w_003_274, w_003_275, w_003_276, w_003_277, w_003_278, w_003_279, w_003_280, w_003_281, w_003_282, w_003_283, w_003_284, w_003_285, w_003_286, w_003_287, w_003_288, w_003_289, w_003_290, w_003_291, w_003_292, w_003_293, w_003_294, w_003_295, w_003_296, w_003_297, w_003_298, w_003_299, w_003_300, w_003_301, w_003_302, w_003_303, w_003_304, w_003_305, w_003_306, w_003_307, w_003_308, w_003_309, w_003_310, w_003_311, w_003_312, w_003_313, w_003_314, w_003_315, w_003_316, w_003_317, w_003_318, w_003_319, w_003_320, w_003_321, w_003_322, w_003_323, w_003_324, w_003_325, w_003_326, w_003_327, w_003_328, w_003_329, w_003_330, w_003_331, w_003_332, w_003_333, w_003_334, w_003_335, w_003_336, w_003_337, w_003_338, w_003_339, w_003_340, w_003_341, w_003_342, w_003_343, w_003_344, w_003_345, w_003_346, w_003_347, w_003_348, w_003_349, w_003_350, w_003_351, w_003_352, w_003_353, w_003_354, w_003_355, w_003_356, w_003_357, w_003_358, w_003_359, w_003_360, w_003_361, w_003_362, w_003_363, w_003_364, w_003_365, w_003_366, w_003_367, w_003_368, w_003_369, w_003_370, w_003_371, w_003_372, w_003_373, w_003_374, w_003_375, w_003_376, w_003_377, w_003_378, w_003_379, w_003_380, w_003_381, w_003_382, w_003_383, w_003_384, w_003_386, w_003_387, w_003_388, w_003_389, w_003_390, w_003_391, w_003_392, w_003_393, w_003_394, w_003_395, w_003_396, w_003_397, w_003_398, w_003_399, w_003_400, w_003_401, w_003_402, w_003_403, w_003_404, w_003_405, w_003_406, w_003_407, w_003_408, w_003_409, w_003_410, w_003_411, w_003_412, w_003_413, w_003_414, w_003_415, w_003_416, w_003_417, w_003_418, w_003_419, w_003_420, w_003_421, w_003_422, w_003_423, w_003_424, w_003_425, w_003_426, w_003_427, w_003_428, w_003_429, w_003_430, w_003_431, w_003_432, w_003_433, w_003_434, w_003_435, w_003_436, w_003_437, w_003_438, w_003_439, w_003_440, w_003_441, w_003_442, w_003_443, w_003_444, w_003_445, w_003_446, w_003_447, w_003_448, w_003_449, w_003_450, w_003_451, w_003_452, w_003_453, w_003_454, w_003_455, w_003_456, w_003_457, w_003_458, w_003_459, w_003_460, w_003_461, w_003_462, w_003_463, w_003_464, w_003_465, w_003_466, w_003_467, w_003_468, w_003_469, w_003_470, w_003_471, w_003_472, w_003_473, w_003_474, w_003_475, w_003_476, w_003_477, w_003_478, w_003_479, w_003_480, w_003_481, w_003_482, w_003_483, w_003_484, w_003_485, w_003_486, w_003_487, w_003_488, w_003_489, w_003_490, w_003_491, w_003_492, w_003_493, w_003_494, w_003_495, w_003_496, w_003_497, w_003_498, w_003_499, w_003_500, w_003_501, w_003_502, w_003_503, w_003_504, w_003_505, w_003_506, w_003_507, w_003_508, w_003_509, w_003_510, w_003_511, w_003_512, w_003_513, w_003_514, w_003_515, w_003_516, w_003_517, w_003_518, w_003_519, w_003_520, w_003_521, w_003_522, w_003_523, w_003_524, w_003_525, w_003_526, w_003_527, w_003_528, w_003_529, w_003_530, w_003_531, w_003_532, w_003_533, w_003_534, w_003_535, w_003_536, w_003_537, w_003_538, w_003_539, w_003_540, w_003_541, w_003_542, w_003_543, w_003_544, w_003_545, w_003_546, w_003_547, w_003_548, w_003_549, w_003_551, w_003_552, w_003_554, w_003_555, w_003_556, w_003_557, w_003_558, w_003_559, w_003_560, w_003_561, w_003_562, w_003_563, w_003_564, w_003_565, w_003_566, w_003_567, w_003_568, w_003_569, w_003_570, w_003_571, w_003_572, w_003_573, w_003_574, w_003_575, w_003_576, w_003_577, w_003_578, w_003_579, w_003_580, w_003_581, w_003_582, w_003_583, w_003_584, w_003_585, w_003_586, w_003_587, w_003_588, w_003_589, w_003_590, w_003_591, w_003_592, w_003_593, w_003_594, w_003_595, w_003_596, w_003_598, w_003_599, w_003_600, w_003_601, w_003_602, w_003_603, w_003_604, w_003_605, w_003_606, w_003_607, w_003_608, w_003_609, w_003_610, w_003_611, w_003_612, w_003_613, w_003_614, w_003_615, w_003_616, w_003_617, w_003_618, w_003_619, w_003_620, w_003_621, w_003_622, w_003_623, w_003_624, w_003_625, w_003_626, w_003_627, w_003_628, w_003_629, w_003_630, w_003_632, w_003_633, w_003_634, w_003_635, w_003_636, w_003_637, w_003_638, w_003_639, w_003_640, w_003_641, w_003_642, w_003_643, w_003_644, w_003_645, w_003_646, w_003_647, w_003_648, w_003_649, w_003_650, w_003_651, w_003_652, w_003_653, w_003_654, w_003_655, w_003_656, w_003_657, w_003_658, w_003_660, w_003_661, w_003_662, w_003_663, w_003_664, w_003_665, w_003_667, w_003_668, w_003_669, w_003_670, w_003_671, w_003_672, w_003_673, w_003_674, w_003_675, w_003_676, w_003_677, w_003_678, w_003_679, w_003_680, w_003_681, w_003_682, w_003_683, w_003_684, w_003_685, w_003_686, w_003_687, w_003_688, w_003_689, w_003_690, w_003_691, w_003_692, w_003_693, w_003_694, w_003_695, w_003_696, w_003_697, w_003_698, w_003_699, w_003_700, w_003_701, w_003_702, w_003_703, w_003_704, w_003_705, w_003_706, w_003_707, w_003_708, w_003_709, w_003_710, w_003_711, w_003_712, w_003_713, w_003_714, w_003_715, w_003_716, w_003_717, w_003_718, w_003_719, w_003_720, w_003_721, w_003_722, w_003_723, w_003_724, w_003_725, w_003_726, w_003_727, w_003_728, w_003_729, w_003_730, w_003_731, w_003_732, w_003_733, w_003_734, w_003_735, w_003_736, w_003_737, w_003_738, w_003_739, w_003_740, w_003_741, w_003_742, w_003_743, w_003_744, w_003_745, w_003_746, w_003_747, w_003_748, w_003_749, w_003_750, w_003_751, w_003_752, w_003_753, w_003_754, w_003_755, w_003_756, w_003_757, w_003_758, w_003_759, w_003_760, w_003_761, w_003_762, w_003_763, w_003_764, w_003_765, w_003_766, w_003_767, w_003_768, w_003_769, w_003_770, w_003_771, w_003_772, w_003_773, w_003_774, w_003_775, w_003_776, w_003_777, w_003_778, w_003_779, w_003_780, w_003_781, w_003_782, w_003_783, w_003_784, w_003_785, w_003_786, w_003_787, w_003_788, w_003_789, w_003_790, w_003_791, w_003_792, w_003_794, w_003_795, w_003_796, w_003_797, w_003_798, w_003_799, w_003_800, w_003_801, w_003_802, w_003_803, w_003_804, w_003_805, w_003_806, w_003_807, w_003_808, w_003_809, w_003_810, w_003_811, w_003_812, w_003_813, w_003_814, w_003_815, w_003_816, w_003_817, w_003_819, w_003_820, w_003_821, w_003_822, w_003_823, w_003_824, w_003_825, w_003_826, w_003_827, w_003_828, w_003_829, w_003_830, w_003_832, w_003_833, w_003_834, w_003_835, w_003_836, w_003_837, w_003_838, w_003_839, w_003_840, w_003_841, w_003_842, w_003_843, w_003_844, w_003_845, w_003_846, w_003_847, w_003_848, w_003_849, w_003_850, w_003_851, w_003_852, w_003_853, w_003_854, w_003_855, w_003_856, w_003_857, w_003_858, w_003_859, w_003_860, w_003_861, w_003_862, w_003_863, w_003_864, w_003_865, w_003_866, w_003_867, w_003_868, w_003_869, w_003_870, w_003_871, w_003_872, w_003_873, w_003_874, w_003_875, w_003_876, w_003_877, w_003_879, w_003_880, w_003_881, w_003_882, w_003_883, w_003_884, w_003_885, w_003_886, w_003_887, w_003_888, w_003_889, w_003_890, w_003_891, w_003_892, w_003_893, w_003_894, w_003_895, w_003_896, w_003_897, w_003_898, w_003_899, w_003_900, w_003_901, w_003_902, w_003_903, w_003_904, w_003_905, w_003_906, w_003_907, w_003_908, w_003_909, w_003_910, w_003_911, w_003_912, w_003_913, w_003_914, w_003_915, w_003_916, w_003_917, w_003_918, w_003_919, w_003_920, w_003_921, w_003_922, w_003_923, w_003_924, w_003_925, w_003_926, w_003_927, w_003_928, w_003_929, w_003_930, w_003_931, w_003_932, w_003_933, w_003_934, w_003_935, w_003_936, w_003_937, w_003_938, w_003_939, w_003_940, w_003_941, w_003_942, w_003_943, w_003_944, w_003_945, w_003_946, w_003_947, w_003_948, w_003_949, w_003_950, w_003_951, w_003_952, w_003_953, w_003_954, w_003_955, w_003_956, w_003_957, w_003_958, w_003_959, w_003_960, w_003_961, w_003_962, w_003_963, w_003_964, w_003_965, w_003_966, w_003_967, w_003_968, w_003_969, w_003_970, w_003_971, w_003_972, w_003_973, w_003_974, w_003_975, w_003_976, w_003_977, w_003_978, w_003_979, w_003_980, w_003_981, w_003_982, w_003_983, w_003_984, w_003_985, w_003_986, w_003_987, w_003_988, w_003_989, w_003_990, w_003_991, w_003_992, w_003_993, w_003_994, w_003_995, w_003_996, w_003_998, w_003_999, w_003_1000, w_003_1002, w_003_1003, w_003_1004, w_003_1005, w_003_1006, w_003_1007, w_003_1008, w_003_1009, w_003_1010, w_003_1011, w_003_1012, w_003_1013, w_003_1014, w_003_1015, w_003_1016, w_003_1018, w_003_1019, w_003_1020, w_003_1021, w_003_1022, w_003_1023, w_003_1024, w_003_1025, w_003_1026, w_003_1027, w_003_1028, w_003_1029, w_003_1030, w_003_1031, w_003_1032, w_003_1033, w_003_1034, w_003_1035, w_003_1036, w_003_1037, w_003_1038, w_003_1039, w_003_1040, w_003_1041, w_003_1042, w_003_1043, w_003_1044, w_003_1045, w_003_1046, w_003_1047, w_003_1048, w_003_1049, w_003_1050, w_003_1051, w_003_1052, w_003_1053, w_003_1054, w_003_1055, w_003_1056, w_003_1057, w_003_1058, w_003_1059, w_003_1060, w_003_1061, w_003_1062, w_003_1063, w_003_1064, w_003_1065, w_003_1066, w_003_1067, w_003_1068, w_003_1069, w_003_1070, w_003_1071, w_003_1072, w_003_1073, w_003_1074, w_003_1075, w_003_1076, w_003_1077, w_003_1078, w_003_1079, w_003_1080, w_003_1081, w_003_1082, w_003_1083, w_003_1084, w_003_1085, w_003_1086, w_003_1087, w_003_1088, w_003_1089, w_003_1090, w_003_1091, w_003_1092, w_003_1093, w_003_1094, w_003_1095, w_003_1096, w_003_1097, w_003_1098, w_003_1099, w_003_1100, w_003_1101, w_003_1102, w_003_1103, w_003_1104, w_003_1105, w_003_1106, w_003_1107, w_003_1108, w_003_1109, w_003_1110, w_003_1111, w_003_1112, w_003_1113, w_003_1114, w_003_1115, w_003_1116, w_003_1117, w_003_1118, w_003_1119, w_003_1120, w_003_1121, w_003_1122, w_003_1123, w_003_1124, w_003_1125, w_003_1126, w_003_1127, w_003_1128, w_003_1129, w_003_1131, w_003_1132, w_003_1133, w_003_1134, w_003_1136, w_003_1137, w_003_1138, w_003_1139, w_003_1140, w_003_1141, w_003_1142, w_003_1143, w_003_1144, w_003_1145, w_003_1147, w_003_1148, w_003_1149, w_003_1150, w_003_1151, w_003_1152, w_003_1153, w_003_1154, w_003_1155, w_003_1156, w_003_1157, w_003_1158, w_003_1159, w_003_1160, w_003_1161, w_003_1162, w_003_1163, w_003_1164, w_003_1165, w_003_1166, w_003_1167, w_003_1168, w_003_1169, w_003_1170, w_003_1171, w_003_1172, w_003_1173, w_003_1174, w_003_1175, w_003_1176, w_003_1177, w_003_1178, w_003_1179, w_003_1180, w_003_1181, w_003_1182, w_003_1183, w_003_1184, w_003_1185, w_003_1186, w_003_1187, w_003_1188, w_003_1189, w_003_1190, w_003_1191, w_003_1192, w_003_1193, w_003_1194, w_003_1195, w_003_1196, w_003_1197, w_003_1198, w_003_1199, w_003_1200, w_003_1201, w_003_1202, w_003_1203, w_003_1204, w_003_1205, w_003_1206, w_003_1207, w_003_1208, w_003_1209, w_003_1210, w_003_1211, w_003_1212, w_003_1213, w_003_1214, w_003_1215, w_003_1216, w_003_1217, w_003_1218, w_003_1219, w_003_1220, w_003_1221, w_003_1222, w_003_1223, w_003_1224, w_003_1225, w_003_1226, w_003_1227, w_003_1228, w_003_1229, w_003_1230, w_003_1231, w_003_1232, w_003_1233, w_003_1234, w_003_1235, w_003_1236, w_003_1237, w_003_1238, w_003_1239, w_003_1240, w_003_1241, w_003_1242, w_003_1243, w_003_1244, w_003_1245, w_003_1246, w_003_1247, w_003_1248, w_003_1249, w_003_1250, w_003_1251, w_003_1252, w_003_1253, w_003_1254, w_003_1255, w_003_1256, w_003_1257, w_003_1258, w_003_1259, w_003_1261, w_003_1262, w_003_1263, w_003_1264, w_003_1265, w_003_1266, w_003_1267, w_003_1268, w_003_1269, w_003_1270, w_003_1271, w_003_1272, w_003_1273, w_003_1274, w_003_1275, w_003_1276, w_003_1277, w_003_1278, w_003_1279, w_003_1280, w_003_1281, w_003_1282, w_003_1283, w_003_1284, w_003_1285, w_003_1286, w_003_1287, w_003_1288, w_003_1289, w_003_1290, w_003_1291, w_003_1292, w_003_1293, w_003_1294, w_003_1295, w_003_1296, w_003_1297, w_003_1298, w_003_1299, w_003_1300, w_003_1301, w_003_1302, w_003_1303, w_003_1304, w_003_1305, w_003_1306, w_003_1307, w_003_1308, w_003_1309, w_003_1310, w_003_1311, w_003_1312, w_003_1313, w_003_1314, w_003_1315, w_003_1316, w_003_1317, w_003_1318, w_003_1319, w_003_1320, w_003_1321, w_003_1322, w_003_1323, w_003_1324, w_003_1325, w_003_1326, w_003_1327, w_003_1328, w_003_1329, w_003_1330, w_003_1331, w_003_1332, w_003_1333, w_003_1334, w_003_1335, w_003_1336, w_003_1337, w_003_1338, w_003_1339, w_003_1340, w_003_1341, w_003_1343, w_003_1344, w_003_1345, w_003_1346, w_003_1347, w_003_1348, w_003_1349, w_003_1350, w_003_1351, w_003_1352, w_003_1353, w_003_1354, w_003_1355, w_003_1356, w_003_1357, w_003_1358, w_003_1359, w_003_1360, w_003_1361, w_003_1362, w_003_1363, w_003_1364, w_003_1365, w_003_1366, w_003_1367, w_003_1368, w_003_1369, w_003_1370, w_003_1371, w_003_1372, w_003_1373, w_003_1374, w_003_1375, w_003_1376, w_003_1377, w_003_1378, w_003_1379, w_003_1380, w_003_1382, w_003_1383, w_003_1384, w_003_1385, w_003_1386, w_003_1387, w_003_1388, w_003_1389, w_003_1390, w_003_1391, w_003_1392, w_003_1393, w_003_1394, w_003_1395, w_003_1396, w_003_1397, w_003_1398, w_003_1399, w_003_1400, w_003_1401, w_003_1402, w_003_1403, w_003_1404, w_003_1405, w_003_1406, w_003_1407, w_003_1408, w_003_1409, w_003_1410, w_003_1411, w_003_1412, w_003_1413, w_003_1414, w_003_1415, w_003_1416, w_003_1417, w_003_1418, w_003_1419, w_003_1420, w_003_1421, w_003_1423, w_003_1424, w_003_1425, w_003_1426, w_003_1427, w_003_1428, w_003_1429, w_003_1430, w_003_1431, w_003_1432, w_003_1433, w_003_1434, w_003_1435, w_003_1436, w_003_1437, w_003_1438, w_003_1439, w_003_1440, w_003_1441, w_003_1442, w_003_1443, w_003_1444, w_003_1445, w_003_1446, w_003_1447, w_003_1448, w_003_1449, w_003_1450, w_003_1451, w_003_1452, w_003_1453, w_003_1454, w_003_1455, w_003_1456, w_003_1457, w_003_1458, w_003_1459, w_003_1460, w_003_1461, w_003_1462, w_003_1463, w_003_1464, w_003_1465, w_003_1466, w_003_1467, w_003_1468, w_003_1469, w_003_1470, w_003_1471, w_003_1472, w_003_1473, w_003_1474, w_003_1475, w_003_1476, w_003_1477, w_003_1478, w_003_1479, w_003_1480, w_003_1481, w_003_1482, w_003_1483, w_003_1484, w_003_1485, w_003_1486, w_003_1487, w_003_1488, w_003_1489, w_003_1490, w_003_1491, w_003_1492, w_003_1493, w_003_1494, w_003_1495, w_003_1496, w_003_1497, w_003_1498, w_003_1499, w_003_1500, w_003_1501, w_003_1502, w_003_1503, w_003_1504, w_003_1505, w_003_1506, w_003_1507, w_003_1508, w_003_1509, w_003_1510, w_003_1511, w_003_1512, w_003_1513, w_003_1514, w_003_1515, w_003_1516, w_003_1517, w_003_1518, w_003_1519, w_003_1520, w_003_1521, w_003_1522, w_003_1523, w_003_1524, w_003_1525, w_003_1526, w_003_1527, w_003_1528, w_003_1529, w_003_1530, w_003_1531, w_003_1532, w_003_1533, w_003_1534, w_003_1535, w_003_1536, w_003_1537, w_003_1538, w_003_1539, w_003_1541, w_003_1542, w_003_1543, w_003_1544, w_003_1545, w_003_1546, w_003_1547, w_003_1548, w_003_1549, w_003_1550, w_003_1551, w_003_1552, w_003_1553, w_003_1554, w_003_1555, w_003_1556, w_003_1557, w_003_1558, w_003_1559, w_003_1560, w_003_1561, w_003_1562, w_003_1563, w_003_1564, w_003_1565, w_003_1566, w_003_1567, w_003_1568, w_003_1569, w_003_1570, w_003_1571, w_003_1572, w_003_1573, w_003_1574, w_003_1575, w_003_1576, w_003_1577, w_003_1578, w_003_1579, w_003_1580, w_003_1581, w_003_1582, w_003_1583, w_003_1584, w_003_1585, w_003_1586, w_003_1587, w_003_1588, w_003_1589, w_003_1590, w_003_1591, w_003_1592, w_003_1593, w_003_1594, w_003_1595, w_003_1596, w_003_1597, w_003_1598, w_003_1599, w_003_1600, w_003_1601, w_003_1602, w_003_1603, w_003_1604, w_003_1605, w_003_1606, w_003_1607, w_003_1608, w_003_1609, w_003_1610, w_003_1611, w_003_1612, w_003_1613, w_003_1614, w_003_1615, w_003_1616, w_003_1617, w_003_1618, w_003_1619, w_003_1620, w_003_1621, w_003_1622, w_003_1623, w_003_1624, w_003_1625, w_003_1626, w_003_1627, w_003_1628, w_003_1629, w_003_1630, w_003_1631, w_003_1632, w_003_1633, w_003_1634, w_003_1635, w_003_1636, w_003_1637, w_003_1638, w_003_1639, w_003_1640, w_003_1641, w_003_1642, w_003_1643, w_003_1644, w_003_1645, w_003_1646, w_003_1647, w_003_1648, w_003_1649, w_003_1650, w_003_1651, w_003_1652, w_003_1653, w_003_1654, w_003_1655, w_003_1656, w_003_1657, w_003_1658, w_003_1659, w_003_1661, w_003_1662, w_003_1663, w_003_1664, w_003_1665, w_003_1666, w_003_1667, w_003_1668, w_003_1669, w_003_1670, w_003_1671, w_003_1672, w_003_1673, w_003_1674, w_003_1675, w_003_1676, w_003_1677, w_003_1678, w_003_1679, w_003_1680, w_003_1681, w_003_1682, w_003_1683, w_003_1684, w_003_1685, w_003_1686, w_003_1687, w_003_1688, w_003_1689, w_003_1690, w_003_1691, w_003_1692, w_003_1693, w_003_1694, w_003_1695, w_003_1696, w_003_1697, w_003_1698, w_003_1699, w_003_1700, w_003_1701, w_003_1702, w_003_1703, w_003_1704, w_003_1705, w_003_1706, w_003_1707, w_003_1708, w_003_1709, w_003_1710, w_003_1711, w_003_1712, w_003_1713, w_003_1714, w_003_1715, w_003_1716, w_003_1717, w_003_1718, w_003_1719, w_003_1720, w_003_1721, w_003_1722, w_003_1723, w_003_1724, w_003_1725, w_003_1726, w_003_1727, w_003_1728, w_003_1729, w_003_1730, w_003_1731, w_003_1732, w_003_1733, w_003_1734, w_003_1735, w_003_1736, w_003_1737, w_003_1738, w_003_1739, w_003_1740, w_003_1741, w_003_1742, w_003_1743, w_003_1744, w_003_1745, w_003_1746, w_003_1747, w_003_1748, w_003_1749, w_003_1750, w_003_1751, w_003_1752, w_003_1753, w_003_1754, w_003_1756, w_003_1757, w_003_1758, w_003_1759, w_003_1760, w_003_1761, w_003_1762, w_003_1763, w_003_1764, w_003_1765, w_003_1766, w_003_1767, w_003_1768, w_003_1769, w_003_1770, w_003_1771, w_003_1772, w_003_1773, w_003_1774, w_003_1775, w_003_1776, w_003_1777, w_003_1778, w_003_1779, w_003_1780, w_003_1781, w_003_1782, w_003_1783, w_003_1784, w_003_1785, w_003_1786, w_003_1787, w_003_1788, w_003_1789, w_003_1790, w_003_1791, w_003_1792, w_003_1793, w_003_1794, w_003_1795, w_003_1796, w_003_1797, w_003_1798, w_003_1799, w_003_1800, w_003_1801, w_003_1802, w_003_1803, w_003_1804, w_003_1806, w_003_1807, w_003_1808, w_003_1809, w_003_1810, w_003_1811, w_003_1812, w_003_1813, w_003_1814, w_003_1815, w_003_1816, w_003_1817, w_003_1818, w_003_1819, w_003_1820, w_003_1821, w_003_1822, w_003_1823, w_003_1824, w_003_1825, w_003_1826, w_003_1827, w_003_1828, w_003_1829, w_003_1830, w_003_1831, w_003_1832, w_003_1833, w_003_1834, w_003_1835, w_003_1836, w_003_1837, w_003_1838, w_003_1839, w_003_1840, w_003_1841, w_003_1842, w_003_1843, w_003_1844, w_003_1845, w_003_1846, w_003_1847, w_003_1848, w_003_1849, w_003_1850, w_003_1851, w_003_1852, w_003_1853, w_003_1854, w_003_1855, w_003_1856, w_003_1857, w_003_1858, w_003_1859, w_003_1860, w_003_1861, w_003_1862, w_003_1864, w_003_1865, w_003_1866, w_003_1867, w_003_1868, w_003_1869, w_003_1870, w_003_1871, w_003_1872, w_003_1873, w_003_1874, w_003_1875, w_003_1876, w_003_1877, w_003_1878, w_003_1879, w_003_1880, w_003_1881, w_003_1882, w_003_1883, w_003_1884, w_003_1885, w_003_1886, w_003_1887, w_003_1888, w_003_1889, w_003_1890, w_003_1891, w_003_1892, w_003_1893, w_003_1894, w_003_1895, w_003_1896, w_003_1897, w_003_1898, w_003_1899, w_003_1900, w_003_1901, w_003_1902, w_003_1903, w_003_1904, w_003_1905, w_003_1906, w_003_1907, w_003_1908, w_003_1909, w_003_1910, w_003_1911, w_003_1912, w_003_1913, w_003_1914, w_003_1915, w_003_1916, w_003_1917, w_003_1918, w_003_1919, w_003_1920, w_003_1921, w_003_1922, w_003_1923, w_003_1924, w_003_1925, w_003_1926, w_003_1927, w_003_1928, w_003_1929, w_003_1930, w_003_1931, w_003_1932, w_003_1933, w_003_1934, w_003_1935, w_003_1936, w_003_1937, w_003_1938, w_003_1939, w_003_1940, w_003_1941, w_003_1942, w_003_1943, w_003_1944, w_003_1945, w_003_1946, w_003_1947, w_003_1948, w_003_1949, w_003_1950, w_003_1951, w_003_1952, w_003_1953, w_003_1954, w_003_1955, w_003_1956, w_003_1957, w_003_1958, w_003_1959, w_003_1960, w_003_1961, w_003_1962, w_003_1963, w_003_1964, w_003_1965, w_003_1966, w_003_1967, w_003_1968, w_003_1969, w_003_1970, w_003_1971, w_003_1972, w_003_1973, w_003_1974, w_003_1975, w_003_1976, w_003_1977, w_003_1978, w_003_1979, w_003_1980, w_003_1981, w_003_1982, w_003_1983, w_003_1984, w_003_1986, w_003_1987, w_003_1988, w_003_1989, w_003_1990, w_003_1991, w_003_1992, w_003_1993, w_003_1994, w_003_1995, w_003_1996, w_003_1997, w_003_1998, w_003_1999, w_003_2000, w_003_2001, w_003_2002, w_003_2003, w_003_2004, w_003_2005, w_003_2006, w_003_2007, w_003_2008, w_003_2009, w_003_2010, w_003_2011, w_003_2012, w_003_2013, w_003_2014, w_003_2015, w_003_2016, w_003_2017, w_003_2018, w_003_2019, w_003_2020, w_003_2021, w_003_2022, w_003_2023, w_003_2024, w_003_2025, w_003_2026, w_003_2027, w_003_2028, w_003_2029, w_003_2030, w_003_2031, w_003_2032, w_003_2033, w_003_2034, w_003_2035, w_003_2037, w_003_2038, w_003_2039, w_003_2040, w_003_2041, w_003_2042, w_003_2043, w_003_2044, w_003_2045, w_003_2046, w_003_2047, w_003_2048, w_003_2049, w_003_2050, w_003_2051, w_003_2052, w_003_2053, w_003_2054, w_003_2055, w_003_2056, w_003_2057, w_003_2058, w_003_2059, w_003_2060, w_003_2061, w_003_2062, w_003_2063, w_003_2065, w_003_2067, w_003_2068, w_003_2069, w_003_2070, w_003_2071, w_003_2072, w_003_2074, w_003_2076, w_003_2077, w_003_2080, w_003_2081, w_003_2082, w_003_2083, w_003_2084, w_003_2086, w_003_2087, w_003_2089, w_003_2090, w_003_2091, w_003_2092, w_003_2093, w_003_2094, w_003_2095, w_003_2096, w_003_2097, w_003_2098, w_003_2100, w_003_2101, w_003_2102, w_003_2104, w_003_2105, w_003_2106, w_003_2108, w_003_2109, w_003_2110, w_003_2111, w_003_2112, w_003_2114, w_003_2115, w_003_2116, w_003_2117, w_003_2118, w_003_2119, w_003_2120, w_003_2121, w_003_2122, w_003_2123, w_003_2124, w_003_2126, w_003_2128, w_003_2129, w_003_2130, w_003_2131, w_003_2132, w_003_2134, w_003_2135, w_003_2136, w_003_2137, w_003_2138, w_003_2140, w_003_2141, w_003_2142, w_003_2143, w_003_2144, w_003_2145, w_003_2146, w_003_2147, w_003_2149, w_003_2150, w_003_2151, w_003_2153, w_003_2154, w_003_2155, w_003_2156, w_003_2157, w_003_2158, w_003_2159, w_003_2162, w_003_2164, w_003_2165, w_003_2166, w_003_2167, w_003_2168, w_003_2170, w_003_2171, w_003_2172, w_003_2173, w_003_2174, w_003_2175, w_003_2176, w_003_2178, w_003_2179, w_003_2180, w_003_2181, w_003_2182, w_003_2183, w_003_2184, w_003_2185, w_003_2186, w_003_2187, w_003_2189, w_003_2190, w_003_2191, w_003_2192, w_003_2193, w_003_2194, w_003_2195, w_003_2196, w_003_2197, w_003_2198, w_003_2199, w_003_2200, w_003_2201, w_003_2202, w_003_2203, w_003_2204, w_003_2205, w_003_2206, w_003_2207, w_003_2208, w_003_2209, w_003_2210, w_003_2211, w_003_2212, w_003_2213, w_003_2214, w_003_2215, w_003_2217, w_003_2218, w_003_2219, w_003_2220, w_003_2221, w_003_2222, w_003_2224, w_003_2226, w_003_2227, w_003_2229, w_003_2231, w_003_2232, w_003_2233, w_003_2234, w_003_2235, w_003_2236, w_003_2237, w_003_2239, w_003_2240, w_003_2241, w_003_2242, w_003_2243, w_003_2244, w_003_2245, w_003_2246, w_003_2247, w_003_2248, w_003_2249, w_003_2250, w_003_2251, w_003_2252, w_003_2253, w_003_2255, w_003_2256, w_003_2258, w_003_2259, w_003_2260, w_003_2261, w_003_2262, w_003_2263, w_003_2264, w_003_2265, w_003_2266, w_003_2267, w_003_2268, w_003_2269, w_003_2271, w_003_2272, w_003_2273, w_003_2274, w_003_2275, w_003_2276, w_003_2277, w_003_2278, w_003_2279, w_003_2280, w_003_2282, w_003_2283, w_003_2284, w_003_2285, w_003_2286, w_003_2288, w_003_2289, w_003_2290, w_003_2291, w_003_2292, w_003_2293, w_003_2294, w_003_2295, w_003_2296, w_003_2297, w_003_2298, w_003_2299, w_003_2300, w_003_2302, w_003_2303, w_003_2304, w_003_2305, w_003_2306, w_003_2307, w_003_2308, w_003_2309, w_003_2310, w_003_2311, w_003_2312, w_003_2313, w_003_2314, w_003_2316, w_003_2318, w_003_2319, w_003_2320, w_003_2321, w_003_2322, w_003_2323, w_003_2324, w_003_2325, w_003_2326, w_003_2327, w_003_2328, w_003_2330, w_003_2331, w_003_2332, w_003_2333, w_003_2334, w_003_2335, w_003_2336, w_003_2337, w_003_2338, w_003_2339, w_003_2340, w_003_2342, w_003_2343, w_003_2344, w_003_2345, w_003_2346, w_003_2347, w_003_2350, w_003_2351, w_003_2352, w_003_2353, w_003_2354, w_003_2355, w_003_2356, w_003_2357, w_003_2358, w_003_2359, w_003_2360, w_003_2361, w_003_2362, w_003_2363, w_003_2364, w_003_2365, w_003_2366, w_003_2367, w_003_2368, w_003_2369, w_003_2370, w_003_2371, w_003_2372, w_003_2373, w_003_2374, w_003_2375, w_003_2378, w_003_2380, w_003_2382, w_003_2383, w_003_2384, w_003_2385, w_003_2386, w_003_2387, w_003_2388, w_003_2389, w_003_2390, w_003_2392, w_003_2393, w_003_2394, w_003_2395, w_003_2396, w_003_2397, w_003_2398, w_003_2400, w_003_2401, w_003_2402, w_003_2403, w_003_2404, w_003_2405, w_003_2406, w_003_2407, w_003_2408, w_003_2409, w_003_2410, w_003_2412, w_003_2413, w_003_2414, w_003_2415, w_003_2416, w_003_2417, w_003_2418, w_003_2419, w_003_2420, w_003_2421, w_003_2422, w_003_2423, w_003_2424, w_003_2425, w_003_2426, w_003_2427, w_003_2428, w_003_2429, w_003_2430, w_003_2431, w_003_2432, w_003_2433, w_003_2434, w_003_2435, w_003_2436, w_003_2437, w_003_2438, w_003_2439, w_003_2440, w_003_2441, w_003_2443, w_003_2444, w_003_2445, w_003_2446, w_003_2447, w_003_2448, w_003_2449, w_003_2451, w_003_2452, w_003_2453, w_003_2454, w_003_2455, w_003_2456, w_003_2458, w_003_2459, w_003_2460, w_003_2461, w_003_2463, w_003_2464, w_003_2467, w_003_2468, w_003_2469, w_003_2470, w_003_2471, w_003_2473, w_003_2474, w_003_2475, w_003_2477, w_003_2478, w_003_2479, w_003_2480, w_003_2481, w_003_2482, w_003_2483, w_003_2484, w_003_2485, w_003_2486, w_003_2487, w_003_2488, w_003_2489, w_003_2492, w_003_2493, w_003_2494, w_003_2495, w_003_2498, w_003_2499, w_003_2501, w_003_2502, w_003_2503, w_003_2506, w_003_2507, w_003_2508, w_003_2509, w_003_2510, w_003_2511, w_003_2512, w_003_2513, w_003_2515, w_003_2516, w_003_2518, w_003_2519, w_003_2520, w_003_2521, w_003_2522, w_003_2523, w_003_2524, w_003_2525, w_003_2526, w_003_2528, w_003_2529, w_003_2531, w_003_2533, w_003_2535, w_003_2536, w_003_2537, w_003_2538, w_003_2539, w_003_2540, w_003_2541, w_003_2542, w_003_2544, w_003_2545, w_003_2546, w_003_2547, w_003_2548, w_003_2549, w_003_2550, w_003_2551, w_003_2552, w_003_2554, w_003_2555, w_003_2556, w_003_2557, w_003_2558, w_003_2559, w_003_2561, w_003_2562, w_003_2563, w_003_2564, w_003_2565, w_003_2566, w_003_2567, w_003_2568, w_003_2569, w_003_2570, w_003_2571, w_003_2572, w_003_2573, w_003_2574, w_003_2576, w_003_2577, w_003_2578, w_003_2579, w_003_2581, w_003_2582, w_003_2583, w_003_2584, w_003_2585, w_003_2586, w_003_2588, w_003_2589, w_003_2590, w_003_2591, w_003_2592, w_003_2593, w_003_2594, w_003_2596, w_003_2598, w_003_2599, w_003_2600, w_003_2601, w_003_2602, w_003_2603, w_003_2604, w_003_2605, w_003_2606, w_003_2607, w_003_2608, w_003_2609, w_003_2612, w_003_2613, w_003_2614, w_003_2615, w_003_2616, w_003_2617, w_003_2618, w_003_2619, w_003_2620, w_003_2621, w_003_2622, w_003_2624, w_003_2625, w_003_2626, w_003_2627, w_003_2628, w_003_2629, w_003_2630, w_003_2631, w_003_2632, w_003_2633, w_003_2634, w_003_2635, w_003_2636, w_003_2637, w_003_2638, w_003_2639, w_003_2640, w_003_2641, w_003_2642, w_003_2643, w_003_2644, w_003_2645, w_003_2646, w_003_2647, w_003_2648, w_003_2649, w_003_2651, w_003_2652, w_003_2653, w_003_2654, w_003_2656, w_003_2657, w_003_2658, w_003_2659, w_003_2660, w_003_2661, w_003_2662, w_003_2663, w_003_2664, w_003_2665, w_003_2666, w_003_2668, w_003_2669, w_003_2670, w_003_2671, w_003_2672, w_003_2673, w_003_2674, w_003_2676, w_003_2677, w_003_2678, w_003_2679, w_003_2681, w_003_2682, w_003_2684, w_003_2685, w_003_2686, w_003_2687, w_003_2688, w_003_2689, w_003_2690, w_003_2691, w_003_2692, w_003_2693, w_003_2694, w_003_2695, w_003_2696, w_003_2697, w_003_2698, w_003_2699, w_003_2700, w_003_2701, w_003_2702, w_003_2703, w_003_2705, w_003_2706, w_003_2707, w_003_2708, w_003_2709, w_003_2710, w_003_2711, w_003_2712, w_003_2713, w_003_2714, w_003_2715, w_003_2716, w_003_2717, w_003_2718, w_003_2719, w_003_2720, w_003_2721, w_003_2722, w_003_2723, w_003_2724, w_003_2725, w_003_2726, w_003_2728, w_003_2730, w_003_2731, w_003_2732, w_003_2733, w_003_2735, w_003_2736, w_003_2737, w_003_2738, w_003_2739, w_003_2740, w_003_2741, w_003_2742, w_003_2743, w_003_2744, w_003_2745, w_003_2746, w_003_2747, w_003_2748, w_003_2749, w_003_2751, w_003_2752, w_003_2753, w_003_2754, w_003_2755, w_003_2756, w_003_2757, w_003_2758, w_003_2759, w_003_2760, w_003_2762, w_003_2763, w_003_2764, w_003_2765, w_003_2766, w_003_2767, w_003_2768, w_003_2770, w_003_2771, w_003_2772, w_003_2773, w_003_2774, w_003_2776, w_003_2777, w_003_2778, w_003_2779, w_003_2780, w_003_2781, w_003_2782, w_003_2783, w_003_2784, w_003_2785, w_003_2787, w_003_2788, w_003_2790, w_003_2791, w_003_2792, w_003_2793, w_003_2794, w_003_2796, w_003_2798, w_003_2799, w_003_2800, w_003_2801, w_003_2803, w_003_2804, w_003_2805, w_003_2806, w_003_2807, w_003_2808, w_003_2809, w_003_2810, w_003_2811, w_003_2812, w_003_2813, w_003_2814, w_003_2815, w_003_2816, w_003_2817, w_003_2819, w_003_2820, w_003_2821, w_003_2822, w_003_2823, w_003_2824, w_003_2826, w_003_2827, w_003_2829, w_003_2831, w_003_2832, w_003_2833, w_003_2834, w_003_2835, w_003_2836, w_003_2837, w_003_2838, w_003_2839, w_003_2841, w_003_2842, w_003_2843, w_003_2845, w_003_2846, w_003_2847, w_003_2849, w_003_2850, w_003_2851, w_003_2852, w_003_2853, w_003_2854, w_003_2855, w_003_2856, w_003_2857, w_003_2858, w_003_2859, w_003_2861, w_003_2862, w_003_2863, w_003_2864, w_003_2866, w_003_2867, w_003_2868, w_003_2869, w_003_2870, w_003_2871, w_003_2873, w_003_2874, w_003_2875, w_003_2877, w_003_2878, w_003_2879, w_003_2880, w_003_2881, w_003_2882, w_003_2884, w_003_2885, w_003_2886, w_003_2887, w_003_2888, w_003_2890, w_003_2892, w_003_2893, w_003_2894, w_003_2895, w_003_2896, w_003_2897, w_003_2898, w_003_2900, w_003_2901, w_003_2902, w_003_2903, w_003_2904, w_003_2906, w_003_2907, w_003_2908, w_003_2909, w_003_2910, w_003_2913, w_003_2914, w_003_2915, w_003_2916, w_003_2917, w_003_2918, w_003_2919, w_003_2920, w_003_2921, w_003_2922, w_003_2923, w_003_2924, w_003_2925, w_003_2926, w_003_2927, w_003_2928, w_003_2929, w_003_2930, w_003_2932, w_003_2933, w_003_2934, w_003_2935, w_003_2936, w_003_2938, w_003_2940, w_003_2941, w_003_2942, w_003_2943, w_003_2944, w_003_2945, w_003_2946, w_003_2948, w_003_2949, w_003_2950, w_003_2952, w_003_2953, w_003_2955, w_003_2956, w_003_2957, w_003_2958, w_003_2959, w_003_2960, w_003_2961, w_003_2962, w_003_2963, w_003_2964, w_003_2965, w_003_2966, w_003_2967, w_003_2968, w_003_2969, w_003_2970, w_003_2971, w_003_2972, w_003_2973, w_003_2974, w_003_2975, w_003_2976, w_003_2977, w_003_2978, w_003_2979, w_003_2980, w_003_2981, w_003_2982, w_003_2983, w_003_2984, w_003_2986, w_003_2987, w_003_2988, w_003_2989, w_003_2990, w_003_2991, w_003_2992, w_003_2993, w_003_2994, w_003_2995, w_003_2996, w_003_2997, w_003_2998, w_003_2999, w_003_3000, w_003_3001, w_003_3002, w_003_3003, w_003_3004, w_003_3006, w_003_3007, w_003_3008, w_003_3009, w_003_3010, w_003_3011, w_003_3012, w_003_3013, w_003_3014, w_003_3017, w_003_3018, w_003_3021, w_003_3022, w_003_3023, w_003_3024, w_003_3025, w_003_3026, w_003_3027, w_003_3028, w_003_3029, w_003_3030, w_003_3031, w_003_3032, w_003_3034, w_003_3035, w_003_3036, w_003_3037, w_003_3038, w_003_3039, w_003_3040, w_003_3041, w_003_3042, w_003_3043, w_003_3044, w_003_3045, w_003_3046, w_003_3047, w_003_3048, w_003_3049, w_003_3050, w_003_3051, w_003_3053, w_003_3054, w_003_3055, w_003_3056, w_003_3057, w_003_3058, w_003_3059, w_003_3060, w_003_3061, w_003_3062, w_003_3063, w_003_3064, w_003_3066, w_003_3067, w_003_3068, w_003_3070, w_003_3071, w_003_3072, w_003_3073, w_003_3074, w_003_3075, w_003_3076, w_003_3077, w_003_3079, w_003_3081, w_003_3082, w_003_3083, w_003_3084, w_003_3085, w_003_3086, w_003_3087, w_003_3088, w_003_3089, w_003_3090, w_003_3091, w_003_3092, w_003_3093, w_003_3094, w_003_3095, w_003_3096, w_003_3098, w_003_3099, w_003_3100, w_003_3101, w_003_3102, w_003_3103, w_003_3104, w_003_3105, w_003_3106, w_003_3107, w_003_3108, w_003_3109, w_003_3110, w_003_3111, w_003_3112, w_003_3113, w_003_3114, w_003_3115, w_003_3116, w_003_3117, w_003_3118, w_003_3119, w_003_3120, w_003_3121, w_003_3122, w_003_3123, w_003_3124, w_003_3125, w_003_3126, w_003_3127, w_003_3129, w_003_3130, w_003_3131, w_003_3132, w_003_3133, w_003_3134, w_003_3135, w_003_3136, w_003_3137, w_003_3138, w_003_3139, w_003_3140, w_003_3141, w_003_3142, w_003_3143, w_003_3145, w_003_3146, w_003_3147, w_003_3151, w_003_3152, w_003_3153, w_003_3154, w_003_3155, w_003_3156, w_003_3157, w_003_3158, w_003_3159, w_003_3160, w_003_3161, w_003_3163, w_003_3164, w_003_3165, w_003_3166, w_003_3167, w_003_3168, w_003_3169, w_003_3170, w_003_3171, w_003_3172, w_003_3173, w_003_3176, w_003_3177, w_003_3179, w_003_3180, w_003_3181, w_003_3182, w_003_3183, w_003_3184, w_003_3185, w_003_3186, w_003_3187, w_003_3188, w_003_3190, w_003_3191, w_003_3192, w_003_3193, w_003_3194, w_003_3195, w_003_3196, w_003_3198, w_003_3199, w_003_3200, w_003_3202, w_003_3203, w_003_3204, w_003_3205, w_003_3206, w_003_3207, w_003_3209, w_003_3210, w_003_3211, w_003_3212, w_003_3213, w_003_3214, w_003_3215, w_003_3216, w_003_3217, w_003_3219, w_003_3220, w_003_3221, w_003_3222, w_003_3223, w_003_3224, w_003_3225, w_003_3226, w_003_3227, w_003_3228, w_003_3231, w_003_3232, w_003_3234, w_003_3235, w_003_3236, w_003_3237, w_003_3238, w_003_3239, w_003_3240, w_003_3241, w_003_3242, w_003_3243, w_003_3244, w_003_3245, w_003_3249, w_003_3252, w_003_3253, w_003_3254, w_003_3255, w_003_3256, w_003_3258, w_003_3259, w_003_3260, w_003_3261, w_003_3262, w_003_3264, w_003_3265, w_003_3266, w_003_3267, w_003_3268, w_003_3269, w_003_3270, w_003_3271, w_003_3272, w_003_3273, w_003_3275, w_003_3276, w_003_3277, w_003_3278, w_003_3279, w_003_3280, w_003_3281, w_003_3282, w_003_3283, w_003_3285, w_003_3286, w_003_3287, w_003_3288, w_003_3289, w_003_3290, w_003_3291, w_003_3292, w_003_3293, w_003_3294, w_003_3295, w_003_3297, w_003_3299, w_003_3300, w_003_3301, w_003_3302, w_003_3303, w_003_3304, w_003_3305, w_003_3306, w_003_3307, w_003_3308, w_003_3310, w_003_3311, w_003_3315, w_003_3317, w_003_3318, w_003_3319, w_003_3320, w_003_3321, w_003_3322, w_003_3323, w_003_3324, w_003_3325, w_003_3326, w_003_3327, w_003_3328, w_003_3329, w_003_3330, w_003_3331, w_003_3332, w_003_3333, w_003_3334, w_003_3335, w_003_3336, w_003_3337, w_003_3338, w_003_3340, w_003_3341, w_003_3342, w_003_3343, w_003_3344, w_003_3345, w_003_3346, w_003_3347, w_003_3348, w_003_3350, w_003_3351, w_003_3352, w_003_3355, w_003_3357, w_003_3358, w_003_3360, w_003_3362, w_003_3363, w_003_3364, w_003_3365, w_003_3366, w_003_3367, w_003_3368, w_003_3369, w_003_3370, w_003_3371, w_003_3372, w_003_3373, w_003_3374, w_003_3375, w_003_3376, w_003_3377, w_003_3378, w_003_3379, w_003_3381, w_003_3383, w_003_3384, w_003_3386, w_003_3387, w_003_3388, w_003_3389, w_003_3390, w_003_3391, w_003_3392, w_003_3393, w_003_3394, w_003_3395, w_003_3397, w_003_3398, w_003_3399, w_003_3400, w_003_3402, w_003_3403, w_003_3404, w_003_3405, w_003_3406, w_003_3407, w_003_3408, w_003_3409, w_003_3410, w_003_3412, w_003_3414, w_003_3415, w_003_3417, w_003_3418, w_003_3420, w_003_3422, w_003_3423, w_003_3424, w_003_3425, w_003_3426, w_003_3427, w_003_3428, w_003_3429, w_003_3430, w_003_3431, w_003_3432, w_003_3433, w_003_3434, w_003_3435, w_003_3437, w_003_3438, w_003_3439, w_003_3440, w_003_3441, w_003_3442, w_003_3443, w_003_3444, w_003_3445, w_003_3446, w_003_3447, w_003_3448, w_003_3451, w_003_3452, w_003_3453, w_003_3454, w_003_3455, w_003_3456, w_003_3457, w_003_3458, w_003_3459, w_003_3460, w_003_3461, w_003_3462, w_003_3464, w_003_3466, w_003_3468, w_003_3469, w_003_3470, w_003_3471, w_003_3472, w_003_3474, w_003_3475, w_003_3478, w_003_3479, w_003_3480, w_003_3481, w_003_3482, w_003_3483, w_003_3484, w_003_3486, w_003_3488, w_003_3489, w_003_3490, w_003_3491, w_003_3493, w_003_3494, w_003_3495, w_003_3496, w_003_3497, w_003_3498, w_003_3499, w_003_3500, w_003_3501, w_003_3502, w_003_3504, w_003_3506, w_003_3507, w_003_3508, w_003_3509, w_003_3510, w_003_3511, w_003_3512, w_003_3513, w_003_3515, w_003_3516, w_003_3517, w_003_3519, w_003_3520, w_003_3521, w_003_3522, w_003_3523, w_003_3525, w_003_3526, w_003_3527, w_003_3528, w_003_3529, w_003_3530, w_003_3531, w_003_3532, w_003_3533, w_003_3537, w_003_3539, w_003_3540, w_003_3541, w_003_3542, w_003_3543, w_003_3544, w_003_3545, w_003_3546, w_003_3548, w_003_3549, w_003_3550, w_003_3551, w_003_3552, w_003_3553, w_003_3554, w_003_3555, w_003_3556, w_003_3557, w_003_3558, w_003_3559, w_003_3561, w_003_3562, w_003_3563, w_003_3564, w_003_3565, w_003_3567, w_003_3568, w_003_3569, w_003_3570, w_003_3571, w_003_3572, w_003_3573, w_003_3574, w_003_3576, w_003_3577, w_003_3578, w_003_3580, w_003_3581, w_003_3582, w_003_3583, w_003_3584, w_003_3585, w_003_3586, w_003_3587, w_003_3588, w_003_3589, w_003_3590, w_003_3591, w_003_3592, w_003_3593, w_003_3594, w_003_3595, w_003_3596, w_003_3597, w_003_3600, w_003_3601, w_003_3602, w_003_3603, w_003_3604, w_003_3605, w_003_3606, w_003_3607, w_003_3609, w_003_3610, w_003_3611, w_003_3612, w_003_3613, w_003_3614, w_003_3615, w_003_3616, w_003_3619, w_003_3620, w_003_3621, w_003_3622, w_003_3624, w_003_3626, w_003_3627, w_003_3628, w_003_3629, w_003_3630, w_003_3632, w_003_3633, w_003_3634, w_003_3635, w_003_3636, w_003_3637, w_003_3638, w_003_3639, w_003_3640, w_003_3641, w_003_3642, w_003_3644, w_003_3646, w_003_3648, w_003_3649, w_003_3651, w_003_3652, w_003_3654, w_003_3655, w_003_3656, w_003_3657, w_003_3658, w_003_3659, w_003_3662, w_003_3663, w_003_3664, w_003_3665, w_003_3666, w_003_3668, w_003_3669, w_003_3670, w_003_3671, w_003_3672, w_003_3673, w_003_3674, w_003_3675, w_003_3676, w_003_3678, w_003_3679, w_003_3680, w_003_3681, w_003_3682, w_003_3683, w_003_3684, w_003_3685, w_003_3686, w_003_3687, w_003_3688, w_003_3689, w_003_3690, w_003_3691, w_003_3692, w_003_3693, w_003_3696, w_003_3697, w_003_3698, w_003_3699, w_003_3701, w_003_3703, w_003_3704, w_003_3705, w_003_3706, w_003_3708, w_003_3709, w_003_3710, w_003_3711, w_003_3713, w_003_3714, w_003_3715, w_003_3716, w_003_3717, w_003_3718, w_003_3719, w_003_3721, w_003_3722, w_003_3724, w_003_3725, w_003_3726, w_003_3727, w_003_3728, w_003_3729, w_003_3730, w_003_3731, w_003_3732, w_003_3733, w_003_3734, w_003_3735, w_003_3737, w_003_3738, w_003_3739, w_003_3740, w_003_3741, w_003_3742, w_003_3743, w_003_3744, w_003_3747, w_003_3748, w_003_3749, w_003_3750, w_003_3751, w_003_3752, w_003_3753, w_003_3754, w_003_3755, w_003_3756, w_003_3757, w_003_3758, w_003_3759, w_003_3760, w_003_3761, w_003_3762, w_003_3763, w_003_3764, w_003_3765, w_003_3766, w_003_3767, w_003_3768, w_003_3769, w_003_3770, w_003_3771, w_003_3772, w_003_3774, w_003_3775, w_003_3776, w_003_3777, w_003_3778, w_003_3779, w_003_3780, w_003_3782, w_003_3783, w_003_3784, w_003_3785, w_003_3786, w_003_3787, w_003_3788, w_003_3789, w_003_3792, w_003_3793, w_003_3794, w_003_3795, w_003_3796, w_003_3797, w_003_3798, w_003_3799, w_003_3800, w_003_3802, w_003_3803, w_003_3804, w_003_3805, w_003_3806, w_003_3807, w_003_3808, w_003_3809, w_003_3811, w_003_3812, w_003_3813, w_003_3814, w_003_3815, w_003_3816, w_003_3817, w_003_3818, w_003_3820, w_003_3821, w_003_3822, w_003_3824, w_003_3825, w_003_3826, w_003_3827, w_003_3829, w_003_3831, w_003_3832, w_003_3834, w_003_3835, w_003_3836, w_003_3838, w_003_3839, w_003_3840, w_003_3841, w_003_3842, w_003_3843, w_003_3844, w_003_3845, w_003_3846, w_003_3847, w_003_3848, w_003_3849, w_003_3851, w_003_3852, w_003_3854, w_003_3855, w_003_3856, w_003_3857, w_003_3858, w_003_3860, w_003_3861, w_003_3862, w_003_3863, w_003_3864, w_003_3865, w_003_3866, w_003_3867, w_003_3869, w_003_3870, w_003_3872, w_003_3873, w_003_3874, w_003_3875, w_003_3876, w_003_3877, w_003_3878, w_003_3879, w_003_3880, w_003_3881, w_003_3883, w_003_3884, w_003_3886, w_003_3887, w_003_3888, w_003_3889, w_003_3890, w_003_3891, w_003_3892, w_003_3893, w_003_3894, w_003_3895, w_003_3896, w_003_3897, w_003_3898, w_003_3899, w_003_3900, w_003_3901, w_003_3902, w_003_3903, w_003_3905, w_003_3906, w_003_3907, w_003_3908, w_003_3909, w_003_3910, w_003_3911, w_003_3912, w_003_3913, w_003_3914, w_003_3915, w_003_3916, w_003_3917, w_003_3919, w_003_3921, w_003_3922, w_003_3923, w_003_3924, w_003_3925, w_003_3926, w_003_3927, w_003_3928, w_003_3929, w_003_3930, w_003_3931, w_003_3932, w_003_3933, w_003_3936, w_003_3937, w_003_3938, w_003_3939, w_003_3940, w_003_3941, w_003_3943, w_003_3944, w_003_3945, w_003_3946, w_003_3948, w_003_3949, w_003_3951, w_003_3952, w_003_3954, w_003_3955, w_003_3956, w_003_3957, w_003_3958, w_003_3959, w_003_3960, w_003_3961, w_003_3962, w_003_3963, w_003_3964, w_003_3965, w_003_3966, w_003_3967, w_003_3968, w_003_3969, w_003_3970, w_003_3971, w_003_3972, w_003_3974, w_003_3975, w_003_3976, w_003_3978, w_003_3979, w_003_3980, w_003_3981, w_003_3982, w_003_3984, w_003_3985, w_003_3986, w_003_3987, w_003_3988, w_003_3989, w_003_3990, w_003_3991, w_003_3992, w_003_3993, w_003_3994, w_003_3995, w_003_3996, w_003_3997, w_003_3998, w_003_3999, w_003_4000, w_003_4001, w_003_4002, w_003_4003, w_003_4005, w_003_4006, w_003_4007, w_003_4008, w_003_4009, w_003_4010, w_003_4011, w_003_4014, w_003_4015, w_003_4016, w_003_4017, w_003_4018, w_003_4019, w_003_4020, w_003_4021, w_003_4022, w_003_4023, w_003_4026, w_003_4027, w_003_4028, w_003_4029, w_003_4030, w_003_4031, w_003_4032, w_003_4033, w_003_4035, w_003_4036, w_003_4038, w_003_4039, w_003_4040, w_003_4041, w_003_4042, w_003_4043, w_003_4044, w_003_4045, w_003_4046, w_003_4047, w_003_4048, w_003_4049, w_003_4050, w_003_4051, w_003_4052, w_003_4053, w_003_4054, w_003_4055, w_003_4056, w_003_4057, w_003_4058, w_003_4059, w_003_4060, w_003_4061, w_003_4062, w_003_4063, w_003_4064, w_003_4065, w_003_4066, w_003_4067, w_003_4068, w_003_4069, w_003_4070, w_003_4071, w_003_4072, w_003_4073, w_003_4074, w_003_4075, w_003_4077, w_003_4078, w_003_4080, w_003_4081, w_003_4082, w_003_4083, w_003_4085, w_003_4086, w_003_4087, w_003_4088, w_003_4089, w_003_4090, w_003_4092, w_003_4093, w_003_4094, w_003_4095, w_003_4096, w_003_4097, w_003_4098, w_003_4099, w_003_4100, w_003_4101, w_003_4104, w_003_4105, w_003_4106, w_003_4107, w_003_4108, w_003_4109, w_003_4110, w_003_4111, w_003_4112, w_003_4113, w_003_4114, w_003_4115, w_003_4116, w_003_4117, w_003_4118, w_003_4119, w_003_4120, w_003_4121, w_003_4122, w_003_4123, w_003_4124, w_003_4125, w_003_4126, w_003_4127, w_003_4128, w_003_4129, w_003_4130, w_003_4131, w_003_4132, w_003_4133, w_003_4135, w_003_4136, w_003_4137, w_003_4138, w_003_4139, w_003_4140, w_003_4141, w_003_4142, w_003_4144, w_003_4145, w_003_4146, w_003_4147, w_003_4148, w_003_4149, w_003_4151, w_003_4153, w_003_4154, w_003_4155, w_003_4156, w_003_4157, w_003_4158, w_003_4159, w_003_4160, w_003_4161, w_003_4162, w_003_4165, w_003_4167, w_003_4168, w_003_4171, w_003_4172, w_003_4173, w_003_4174, w_003_4175, w_003_4176, w_003_4177, w_003_4178, w_003_4179, w_003_4180, w_003_4181, w_003_4182, w_003_4183, w_003_4185, w_003_4186, w_003_4187, w_003_4188, w_003_4189, w_003_4190, w_003_4191, w_003_4192, w_003_4193, w_003_4194, w_003_4195, w_003_4196, w_003_4197, w_003_4199, w_003_4200, w_003_4201, w_003_4202, w_003_4203, w_003_4204, w_003_4205, w_003_4206, w_003_4207, w_003_4208, w_003_4209, w_003_4210, w_003_4211, w_003_4212, w_003_4213, w_003_4214, w_003_4216, w_003_4217, w_003_4218, w_003_4219, w_003_4220, w_003_4221, w_003_4222, w_003_4223, w_003_4224, w_003_4225, w_003_4226, w_003_4227, w_003_4229, w_003_4230, w_003_4231, w_003_4232, w_003_4234, w_003_4235, w_003_4237, w_003_4239, w_003_4240, w_003_4242, w_003_4243, w_003_4244, w_003_4245, w_003_4246, w_003_4247, w_003_4248, w_003_4249, w_003_4250, w_003_4251, w_003_4252, w_003_4253, w_003_4254, w_003_4255, w_003_4256, w_003_4257, w_003_4258, w_003_4259, w_003_4260, w_003_4261, w_003_4262, w_003_4263, w_003_4264, w_003_4265, w_003_4266, w_003_4268, w_003_4270, w_003_4271, w_003_4273, w_003_4275, w_003_4277, w_003_4278, w_003_4279, w_003_4280, w_003_4281, w_003_4282, w_003_4283, w_003_4284, w_003_4285, w_003_4287, w_003_4288, w_003_4289, w_003_4290, w_003_4291, w_003_4293, w_003_4295, w_003_4296, w_003_4297, w_003_4299, w_003_4300, w_003_4301, w_003_4303, w_003_4304, w_003_4305, w_003_4307, w_003_4308, w_003_4309, w_003_4310, w_003_4311, w_003_4312, w_003_4313, w_003_4314, w_003_4315, w_003_4316, w_003_4317, w_003_4318, w_003_4319, w_003_4320, w_003_4321, w_003_4322, w_003_4323, w_003_4324, w_003_4325, w_003_4326, w_003_4327, w_003_4328, w_003_4329, w_003_4330, w_003_4331, w_003_4332, w_003_4333, w_003_4334, w_003_4336, w_003_4337, w_003_4338, w_003_4339, w_003_4340, w_003_4341, w_003_4342, w_003_4343, w_003_4344, w_003_4346, w_003_4347, w_003_4348, w_003_4349, w_003_4350, w_003_4352, w_003_4354, w_003_4355, w_003_4356, w_003_4357, w_003_4358, w_003_4359, w_003_4360, w_003_4361, w_003_4362, w_003_4363, w_003_4364, w_003_4365, w_003_4366, w_003_4368, w_003_4370, w_003_4371, w_003_4372, w_003_4373, w_003_4374, w_003_4375, w_003_4377, w_003_4378, w_003_4379, w_003_4380, w_003_4382, w_003_4383, w_003_4384, w_003_4385, w_003_4386, w_003_4387, w_003_4388, w_003_4389, w_003_4390, w_003_4391, w_003_4393, w_003_4394, w_003_4395, w_003_4396, w_003_4397, w_003_4398, w_003_4399, w_003_4400, w_003_4401, w_003_4402, w_003_4403, w_003_4404, w_003_4405, w_003_4406, w_003_4407, w_003_4408, w_003_4409, w_003_4410, w_003_4412, w_003_4413, w_003_4414, w_003_4415, w_003_4416, w_003_4417, w_003_4418, w_003_4419, w_003_4420, w_003_4421, w_003_4422, w_003_4424, w_003_4425, w_003_4426, w_003_4427, w_003_4428, w_003_4429, w_003_4430, w_003_4431, w_003_4433, w_003_4434, w_003_4435, w_003_4436, w_003_4437, w_003_4438, w_003_4440, w_003_4441, w_003_4442, w_003_4443, w_003_4444, w_003_4445, w_003_4446, w_003_4447, w_003_4448, w_003_4451, w_003_4452, w_003_4453, w_003_4455, w_003_4456, w_003_4457, w_003_4458, w_003_4459, w_003_4460, w_003_4461, w_003_4462, w_003_4463, w_003_4464, w_003_4465, w_003_4466, w_003_4467, w_003_4468, w_003_4469, w_003_4470, w_003_4471, w_003_4472, w_003_4473, w_003_4474, w_003_4475, w_003_4476, w_003_4477, w_003_4478, w_003_4479, w_003_4480, w_003_4481, w_003_4483, w_003_4484, w_003_4485, w_003_4486, w_003_4487, w_003_4488, w_003_4489, w_003_4490, w_003_4491, w_003_4492, w_003_4493, w_003_4494, w_003_4495, w_003_4496, w_003_4497, w_003_4498, w_003_4499, w_003_4500, w_003_4501, w_003_4502, w_003_4503, w_003_4504, w_003_4505, w_003_4506, w_003_4507, w_003_4508, w_003_4510, w_003_4511, w_003_4512, w_003_4513, w_003_4514, w_003_4516, w_003_4517, w_003_4518, w_003_4520, w_003_4523, w_003_4524, w_003_4525, w_003_4526, w_003_4527, w_003_4528, w_003_4529, w_003_4531, w_003_4532, w_003_4533, w_003_4535, w_003_4536, w_003_4537, w_003_4538, w_003_4539, w_003_4540, w_003_4541, w_003_4542, w_003_4543, w_003_4544, w_003_4545, w_003_4546, w_003_4547, w_003_4548, w_003_4550, w_003_4551, w_003_4552, w_003_4553, w_003_4554, w_003_4555, w_003_4556, w_003_4557, w_003_4559, w_003_4561, w_003_4562, w_003_4564, w_003_4565, w_003_4566, w_003_4567, w_003_4568, w_003_4569, w_003_4570, w_003_4571, w_003_4572, w_003_4573, w_003_4574, w_003_4575, w_003_4576, w_003_4577, w_003_4578, w_003_4579, w_003_4580, w_003_4581, w_003_4583, w_003_4585, w_003_4587, w_003_4588, w_003_4590, w_003_4591, w_003_4592, w_003_4593, w_003_4594, w_003_4595, w_003_4598, w_003_4599, w_003_4600, w_003_4601, w_003_4602, w_003_4603, w_003_4604, w_003_4605, w_003_4606, w_003_4607, w_003_4608, w_003_4609, w_003_4610, w_003_4612, w_003_4613, w_003_4616, w_003_4617, w_003_4619, w_003_4620, w_003_4621, w_003_4622, w_003_4623, w_003_4624, w_003_4625, w_003_4627, w_003_4628, w_003_4629, w_003_4631, w_003_4632, w_003_4633, w_003_4635, w_003_4636, w_003_4637, w_003_4638, w_003_4639, w_003_4640, w_003_4641, w_003_4642, w_003_4643, w_003_4644, w_003_4645, w_003_4646, w_003_4647, w_003_4648, w_003_4649, w_003_4650, w_003_4652, w_003_4653, w_003_4655, w_003_4656, w_003_4657, w_003_4658, w_003_4659, w_003_4660, w_003_4661, w_003_4662, w_003_4663, w_003_4664, w_003_4665, w_003_4666, w_003_4667, w_003_4668, w_003_4669, w_003_4670, w_003_4671, w_003_4672, w_003_4673, w_003_4674, w_003_4675, w_003_4677, w_003_4678, w_003_4679, w_003_4680, w_003_4681, w_003_4682, w_003_4683, w_003_4684, w_003_4685, w_003_4686, w_003_4687, w_003_4688, w_003_4689, w_003_4690, w_003_4691, w_003_4692, w_003_4693, w_003_4694, w_003_4695, w_003_4696, w_003_4697, w_003_4698, w_003_4700, w_003_4701, w_003_4703, w_003_4704, w_003_4706, w_003_4708, w_003_4709, w_003_4710, w_003_4712, w_003_4713, w_003_4714, w_003_4715, w_003_4716, w_003_4717, w_003_4718, w_003_4719, w_003_4720, w_003_4721, w_003_4722, w_003_4723, w_003_4724, w_003_4725, w_003_4726, w_003_4727, w_003_4728, w_003_4729, w_003_4730, w_003_4731, w_003_4732, w_003_4734, w_003_4735, w_003_4736, w_003_4738, w_003_4739, w_003_4740, w_003_4741, w_003_4742, w_003_4743, w_003_4744, w_003_4745, w_003_4746, w_003_4748, w_003_4750, w_003_4752, w_003_4754, w_003_4756, w_003_4757, w_003_4758, w_003_4759, w_003_4761, w_003_4762, w_003_4765, w_003_4766, w_003_4767, w_003_4768, w_003_4769, w_003_4770, w_003_4771, w_003_4772, w_003_4774, w_003_4776, w_003_4778, w_003_4779, w_003_4780, w_003_4781, w_003_4782, w_003_4783, w_003_4784, w_003_4786, w_003_4788, w_003_4789, w_003_4790, w_003_4791, w_003_4792, w_003_4793, w_003_4794, w_003_4795, w_003_4796, w_003_4797, w_003_4798, w_003_4799, w_003_4800, w_003_4801, w_003_4802, w_003_4803, w_003_4804, w_003_4806, w_003_4807, w_003_4809, w_003_4810, w_003_4812, w_003_4813, w_003_4814, w_003_4815, w_003_4816, w_003_4817, w_003_4818, w_003_4819, w_003_4820, w_003_4821, w_003_4823, w_003_4824, w_003_4825, w_003_4827, w_003_4828, w_003_4829, w_003_4830, w_003_4831, w_003_4832, w_003_4833, w_003_4834, w_003_4835, w_003_4836, w_003_4837, w_003_4839, w_003_4840, w_003_4841, w_003_4842, w_003_4844, w_003_4845, w_003_4846, w_003_4847, w_003_4848, w_003_4849, w_003_4850, w_003_4851, w_003_4852, w_003_4853, w_003_4854, w_003_4856, w_003_4857, w_003_4858, w_003_4859, w_003_4860, w_003_4861, w_003_4862, w_003_4863, w_003_4864, w_003_4866, w_003_4868, w_003_4869, w_003_4870, w_003_4871, w_003_4872, w_003_4873, w_003_4874, w_003_4875, w_003_4877, w_003_4878, w_003_4879, w_003_4880, w_003_4881, w_003_4882, w_003_4883, w_003_4884, w_003_4886, w_003_4888, w_003_4889, w_003_4890, w_003_4892, w_003_4894, w_003_4895, w_003_4896, w_003_4897, w_003_4898, w_003_4899, w_003_4900, w_003_4901, w_003_4903, w_003_4904, w_003_4905, w_003_4906, w_003_4907, w_003_4908, w_003_4910, w_003_4911, w_003_4914, w_003_4915, w_003_4916, w_003_4917, w_003_4918, w_003_4919, w_003_4920, w_003_4922, w_003_4923, w_003_4924, w_003_4925, w_003_4926, w_003_4927, w_003_4928, w_003_4929, w_003_4930, w_003_4931, w_003_4933, w_003_4934, w_003_4935, w_003_4936, w_003_4937, w_003_4938, w_003_4939, w_003_4940, w_003_4941, w_003_4942, w_003_4943, w_003_4944, w_003_4945, w_003_4946, w_003_4947, w_003_4948, w_003_4949, w_003_4950, w_003_4951, w_003_4952, w_003_4953, w_003_4954, w_003_4955, w_003_4956, w_003_4957, w_003_4958, w_003_4960, w_003_4961, w_003_4962, w_003_4963, w_003_4965, w_003_4966, w_003_4968, w_003_4969, w_003_4970, w_003_4971, w_003_4972, w_003_4973, w_003_4974, w_003_4975, w_003_4976, w_003_4977, w_003_4978, w_003_4979, w_003_4980, w_003_4984, w_003_4985, w_003_4986, w_003_4987, w_003_4988, w_003_4990, w_003_4991, w_003_4992, w_003_4993, w_003_4994, w_003_4995, w_003_4996, w_003_4997, w_003_4998, w_003_5000, w_003_5002, w_003_5003, w_003_5004, w_003_5006, w_003_5007, w_003_5008, w_003_5010, w_003_5011, w_003_5012, w_003_5013, w_003_5014, w_003_5015, w_003_5016, w_003_5018, w_003_5019, w_003_5020, w_003_5021, w_003_5022, w_003_5023, w_003_5024, w_003_5025, w_003_5026, w_003_5027, w_003_5028, w_003_5030, w_003_5031, w_003_5032, w_003_5033, w_003_5034, w_003_5036, w_003_5037, w_003_5038, w_003_5041, w_003_5042, w_003_5043, w_003_5045, w_003_5046, w_003_5047, w_003_5048, w_003_5051, w_003_5052, w_003_5053, w_003_5054, w_003_5057, w_003_5058, w_003_5059, w_003_5060, w_003_5061, w_003_5062, w_003_5063, w_003_5064, w_003_5065, w_003_5066, w_003_5067, w_003_5068, w_003_5069, w_003_5070, w_003_5071, w_003_5072, w_003_5073, w_003_5074, w_003_5075, w_003_5076, w_003_5077, w_003_5078, w_003_5079, w_003_5080, w_003_5081, w_003_5082, w_003_5083, w_003_5084, w_003_5085, w_003_5086, w_003_5087, w_003_5088, w_003_5089, w_003_5090, w_003_5091, w_003_5092, w_003_5093, w_003_5094, w_003_5095, w_003_5096, w_003_5097, w_003_5098, w_003_5099, w_003_5102, w_003_5103, w_003_5105, w_003_5106, w_003_5107, w_003_5108, w_003_5111, w_003_5112, w_003_5113, w_003_5114, w_003_5115, w_003_5116, w_003_5117, w_003_5118, w_003_5119, w_003_5120, w_003_5121, w_003_5122, w_003_5123, w_003_5125, w_003_5126, w_003_5129, w_003_5130, w_003_5131, w_003_5132, w_003_5133, w_003_5134, w_003_5135, w_003_5136, w_003_5137, w_003_5138, w_003_5139, w_003_5140, w_003_5141, w_003_5142, w_003_5143, w_003_5144, w_003_5145, w_003_5146, w_003_5147, w_003_5148, w_003_5149, w_003_5150, w_003_5152, w_003_5153, w_003_5154, w_003_5155, w_003_5158, w_003_5159, w_003_5160, w_003_5161, w_003_5162, w_003_5163, w_003_5165, w_003_5166, w_003_5167, w_003_5168, w_003_5170, w_003_5173, w_003_5174, w_003_5175, w_003_5176, w_003_5177, w_003_5178, w_003_5180, w_003_5183, w_003_5184, w_003_5185, w_003_5186, w_003_5187, w_003_5188, w_003_5190, w_003_5191, w_003_5192, w_003_5193, w_003_5194, w_003_5195, w_003_5196, w_003_5197, w_003_5198, w_003_5199, w_003_5200, w_003_5201, w_003_5203, w_003_5204, w_003_5205, w_003_5206, w_003_5207, w_003_5208, w_003_5209, w_003_5210, w_003_5211, w_003_5212, w_003_5213, w_003_5214, w_003_5215, w_003_5216, w_003_5217, w_003_5218, w_003_5219, w_003_5220, w_003_5221, w_003_5222, w_003_5223, w_003_5224, w_003_5225, w_003_5226, w_003_5227, w_003_5228, w_003_5229, w_003_5230, w_003_5231, w_003_5232, w_003_5235, w_003_5236, w_003_5237, w_003_5238, w_003_5239, w_003_5240, w_003_5241, w_003_5242, w_003_5243, w_003_5245, w_003_5246, w_003_5248, w_003_5249, w_003_5250, w_003_5253, w_003_5254, w_003_5255, w_003_5256, w_003_5257, w_003_5258, w_003_5260, w_003_5261, w_003_5262, w_003_5263, w_003_5266, w_003_5267, w_003_5268, w_003_5269, w_003_5270, w_003_5271, w_003_5273, w_003_5274, w_003_5275, w_003_5276, w_003_5278, w_003_5279, w_003_5280, w_003_5281, w_003_5282, w_003_5283, w_003_5284, w_003_5286, w_003_5287, w_003_5288, w_003_5289, w_003_5290, w_003_5291, w_003_5292, w_003_5293, w_003_5295, w_003_5296, w_003_5297, w_003_5299, w_003_5300, w_003_5301, w_003_5303, w_003_5305, w_003_5307, w_003_5308, w_003_5309, w_003_5310, w_003_5311, w_003_5312, w_003_5313, w_003_5314, w_003_5315, w_003_5317, w_003_5318, w_003_5319, w_003_5320, w_003_5321, w_003_5322, w_003_5324, w_003_5326, w_003_5327, w_003_5329, w_003_5330, w_003_5331, w_003_5332, w_003_5333, w_003_5334, w_003_5335, w_003_5337, w_003_5338, w_003_5339, w_003_5340, w_003_5341, w_003_5342, w_003_5343, w_003_5344, w_003_5345, w_003_5346, w_003_5347, w_003_5348, w_003_5350, w_003_5353, w_003_5355, w_003_5356, w_003_5357, w_003_5358, w_003_5359, w_003_5360, w_003_5361, w_003_5362, w_003_5364, w_003_5365, w_003_5366, w_003_5367, w_003_5370, w_003_5371, w_003_5373, w_003_5374, w_003_5375, w_003_5376, w_003_5377, w_003_5378, w_003_5379, w_003_5380, w_003_5381, w_003_5382, w_003_5383, w_003_5384, w_003_5385, w_003_5386, w_003_5388, w_003_5391, w_003_5392, w_003_5393, w_003_5395, w_003_5396, w_003_5398, w_003_5399, w_003_5401, w_003_5402, w_003_5403, w_003_5404, w_003_5405, w_003_5406, w_003_5407, w_003_5410, w_003_5411, w_003_5412, w_003_5413, w_003_5414, w_003_5415, w_003_5417, w_003_5418, w_003_5419, w_003_5420, w_003_5422, w_003_5424, w_003_5425, w_003_5426, w_003_5427, w_003_5428, w_003_5429, w_003_5430, w_003_5431, w_003_5432, w_003_5433, w_003_5434, w_003_5435, w_003_5436, w_003_5439, w_003_5440, w_003_5441, w_003_5442, w_003_5443, w_003_5444, w_003_5445, w_003_5448, w_003_5449, w_003_5450, w_003_5451, w_003_5452, w_003_5453, w_003_5454, w_003_5455, w_003_5456, w_003_5457, w_003_5458, w_003_5459, w_003_5460, w_003_5461, w_003_5462, w_003_5463, w_003_5464, w_003_5465, w_003_5466, w_003_5467, w_003_5468, w_003_5469, w_003_5470, w_003_5471, w_003_5473, w_003_5474, w_003_5475, w_003_5476, w_003_5480, w_003_5482, w_003_5483, w_003_5484, w_003_5485, w_003_5486, w_003_5487, w_003_5488, w_003_5489, w_003_5490, w_003_5491, w_003_5492, w_003_5495, w_003_5496, w_003_5497, w_003_5498, w_003_5499, w_003_5500, w_003_5501, w_003_5502, w_003_5504, w_003_5505, w_003_5506, w_003_5507, w_003_5508, w_003_5509, w_003_5510, w_003_5511, w_003_5512, w_003_5513, w_003_5514, w_003_5515, w_003_5516, w_003_5517, w_003_5518, w_003_5519, w_003_5520, w_003_5523, w_003_5524, w_003_5525, w_003_5527, w_003_5528, w_003_5529, w_003_5530, w_003_5531, w_003_5532, w_003_5534, w_003_5535, w_003_5536, w_003_5537, w_003_5538, w_003_5539, w_003_5540, w_003_5541, w_003_5542, w_003_5543, w_003_5544, w_003_5546, w_003_5547, w_003_5548, w_003_5549, w_003_5550, w_003_5551, w_003_5552, w_003_5553, w_003_5554, w_003_5555, w_003_5556, w_003_5557, w_003_5558, w_003_5559, w_003_5560, w_003_5561, w_003_5562, w_003_5563, w_003_5564, w_003_5565, w_003_5568, w_003_5569, w_003_5571, w_003_5572, w_003_5575, w_003_5576, w_003_5577, w_003_5578, w_003_5579, w_003_5581, w_003_5582, w_003_5583, w_003_5584, w_003_5585, w_003_5586, w_003_5587, w_003_5588, w_003_5589, w_003_5590, w_003_5591, w_003_5592, w_003_5593, w_003_5594, w_003_5595, w_003_5596, w_003_5597, w_003_5598, w_003_5599, w_003_5600, w_003_5601, w_003_5602, w_003_5603, w_003_5604, w_003_5605, w_003_5606, w_003_5607, w_003_5608, w_003_5609, w_003_5610, w_003_5611, w_003_5612, w_003_5614, w_003_5615, w_003_5617, w_003_5618, w_003_5619, w_003_5620, w_003_5621, w_003_5623, w_003_5624, w_003_5627, w_003_5628, w_003_5629, w_003_5630, w_003_5632, w_003_5633, w_003_5634, w_003_5636, w_003_5637, w_003_5638, w_003_5639, w_003_5640, w_003_5641, w_003_5642, w_003_5643, w_003_5644, w_003_5645, w_003_5646, w_003_5647, w_003_5648, w_003_5649, w_003_5650, w_003_5651, w_003_5652, w_003_5653, w_003_5654, w_003_5655, w_003_5656, w_003_5657, w_003_5658, w_003_5659, w_003_5660, w_003_5661, w_003_5662, w_003_5663, w_003_5664, w_003_5665, w_003_5666, w_003_5667, w_003_5668, w_003_5669, w_003_5670, w_003_5672, w_003_5673, w_003_5674, w_003_5675, w_003_5676, w_003_5678, w_003_5679, w_003_5680, w_003_5681, w_003_5682, w_003_5683, w_003_5684, w_003_5685, w_003_5686, w_003_5687, w_003_5688, w_003_5689, w_003_5690, w_003_5691, w_003_5693, w_003_5694, w_003_5695, w_003_5696, w_003_5697, w_003_5698, w_003_5699, w_003_5700, w_003_5701, w_003_5702, w_003_5703, w_003_5705, w_003_5706, w_003_5708, w_003_5709, w_003_5710, w_003_5711, w_003_5712, w_003_5713, w_003_5714, w_003_5716, w_003_5717, w_003_5718, w_003_5719, w_003_5720, w_003_5721, w_003_5722, w_003_5723, w_003_5724, w_003_5725, w_003_5726, w_003_5727, w_003_5728, w_003_5729, w_003_5730, w_003_5731, w_003_5732, w_003_5733, w_003_5734, w_003_5735, w_003_5736, w_003_5737, w_003_5739, w_003_5740, w_003_5741, w_003_5742, w_003_5743, w_003_5744, w_003_5745, w_003_5747, w_003_5749, w_003_5750, w_003_5752, w_003_5753, w_003_5754, w_003_5755, w_003_5756, w_003_5757, w_003_5759, w_003_5760, w_003_5761, w_003_5762, w_003_5763, w_003_5764, w_003_5765, w_003_5767, w_003_5768, w_003_5769, w_003_5770, w_003_5771, w_003_5772, w_003_5773, w_003_5774, w_003_5775, w_003_5776, w_003_5777, w_003_5779, w_003_5780, w_003_5781, w_003_5782, w_003_5783, w_003_5784, w_003_5785, w_003_5786, w_003_5787, w_003_5790, w_003_5791, w_003_5792, w_003_5793, w_003_5794, w_003_5797, w_003_5798, w_003_5799, w_003_5800, w_003_5801, w_003_5802, w_003_5803, w_003_5804, w_003_5805, w_003_5806, w_003_5807, w_003_5810, w_003_5812, w_003_5813, w_003_5814, w_003_5815, w_003_5816, w_003_5817, w_003_5818, w_003_5820, w_003_5821, w_003_5822, w_003_5823, w_003_5824, w_003_5826, w_003_5827, w_003_5828, w_003_5829, w_003_5830, w_003_5831, w_003_5832, w_003_5833, w_003_5834, w_003_5835, w_003_5836, w_003_5837, w_003_5839, w_003_5840, w_003_5841, w_003_5842, w_003_5843, w_003_5844, w_003_5845, w_003_5846, w_003_5847, w_003_5848, w_003_5849, w_003_5850, w_003_5851, w_003_5852, w_003_5854, w_003_5855, w_003_5856, w_003_5857, w_003_5860, w_003_5861, w_003_5862, w_003_5863, w_003_5864, w_003_5865, w_003_5866, w_003_5867, w_003_5868, w_003_5869, w_003_5870, w_003_5871, w_003_5872, w_003_5873, w_003_5874, w_003_5875, w_003_5876, w_003_5877, w_003_5878, w_003_5879, w_003_5880, w_003_5881, w_003_5882, w_003_5884, w_003_5885, w_003_5886, w_003_5887, w_003_5888, w_003_5889, w_003_5891, w_003_5892, w_003_5893, w_003_5894, w_003_5896, w_003_5897, w_003_5898, w_003_5899, w_003_5900, w_003_5901, w_003_5902, w_003_5903, w_003_5904, w_003_5905, w_003_5906, w_003_5907, w_003_5908, w_003_5909, w_003_5910, w_003_5911, w_003_5912, w_003_5913, w_003_5914, w_003_5915, w_003_5916, w_003_5918, w_003_5920, w_003_5921, w_003_5922, w_003_5923, w_003_5925, w_003_5926, w_003_5928, w_003_5930, w_003_5932, w_003_5933, w_003_5934, w_003_5935, w_003_5936, w_003_5937, w_003_5938, w_003_5939, w_003_5940, w_003_5941, w_003_5942, w_003_5943, w_003_5944, w_003_5945, w_003_5946, w_003_5948, w_003_5949, w_003_5950, w_003_5954, w_003_5955, w_003_5956, w_003_5957, w_003_5958, w_003_5959, w_003_5961, w_003_5964, w_003_5965, w_003_5966, w_003_5967, w_003_5968, w_003_5971, w_003_5972, w_003_5973, w_003_5974, w_003_5975, w_003_5977, w_003_5978, w_003_5979, w_003_5982, w_003_5983, w_003_5984, w_003_5985, w_003_5986, w_003_5987, w_003_5988, w_003_5989, w_003_5990, w_003_5991, w_003_5992, w_003_5993, w_003_5994, w_003_5995, w_003_5998, w_003_5999, w_003_6000, w_003_6001, w_003_6002, w_003_6003, w_003_6004, w_003_6006, w_003_6007, w_003_6008, w_003_6009, w_003_6010, w_003_6011, w_003_6012, w_003_6014, w_003_6015, w_003_6016, w_003_6017, w_003_6019, w_003_6021, w_003_6022, w_003_6023, w_003_6024, w_003_6025, w_003_6026, w_003_6027, w_003_6028, w_003_6029, w_003_6030, w_003_6031, w_003_6032, w_003_6033, w_003_6034, w_003_6035, w_003_6037, w_003_6038, w_003_6039, w_003_6040, w_003_6041, w_003_6042, w_003_6043, w_003_6044, w_003_6045, w_003_6046, w_003_6047, w_003_6048, w_003_6049, w_003_6051, w_003_6053, w_003_6054, w_003_6055, w_003_6056, w_003_6057, w_003_6058, w_003_6060, w_003_6061, w_003_6062, w_003_6063, w_003_6064, w_003_6065, w_003_6067, w_003_6068, w_003_6070, w_003_6071, w_003_6072, w_003_6073, w_003_6074, w_003_6075, w_003_6076, w_003_6077, w_003_6078, w_003_6079, w_003_6080, w_003_6081, w_003_6082, w_003_6083, w_003_6084, w_003_6085, w_003_6086, w_003_6087, w_003_6088, w_003_6089, w_003_6090, w_003_6091, w_003_6092, w_003_6093, w_003_6094, w_003_6095, w_003_6096, w_003_6097, w_003_6098, w_003_6100, w_003_6101, w_003_6102, w_003_6103, w_003_6104, w_003_6105, w_003_6106, w_003_6107, w_003_6108, w_003_6109, w_003_6110, w_003_6111, w_003_6112, w_003_6113, w_003_6114, w_003_6115, w_003_6116, w_003_6117, w_003_6118, w_003_6119, w_003_6120, w_003_6121, w_003_6122, w_003_6123, w_003_6127, w_003_6128, w_003_6129, w_003_6130, w_003_6131, w_003_6132, w_003_6133, w_003_6134, w_003_6135, w_003_6136, w_003_6137, w_003_6138, w_003_6139, w_003_6141, w_003_6142, w_003_6143, w_003_6145, w_003_6146, w_003_6147, w_003_6148, w_003_6149, w_003_6150, w_003_6151, w_003_6152, w_003_6153, w_003_6154, w_003_6155, w_003_6156, w_003_6157, w_003_6158, w_003_6159, w_003_6162, w_003_6164, w_003_6165, w_003_6166, w_003_6167, w_003_6168, w_003_6169, w_003_6170, w_003_6171, w_003_6172, w_003_6173, w_003_6174, w_003_6176, w_003_6177, w_003_6178, w_003_6179, w_003_6180, w_003_6181, w_003_6182, w_003_6184, w_003_6185, w_003_6186, w_003_6188, w_003_6189, w_003_6190, w_003_6191, w_003_6192, w_003_6193, w_003_6194, w_003_6196, w_003_6197, w_003_6198, w_003_6199, w_003_6200, w_003_6201, w_003_6202, w_003_6203, w_003_6204, w_003_6205, w_003_6206, w_003_6207, w_003_6208, w_003_6209, w_003_6210, w_003_6211, w_003_6212, w_003_6213, w_003_6214, w_003_6215, w_003_6217, w_003_6218, w_003_6219, w_003_6221, w_003_6222, w_003_6223, w_003_6225, w_003_6226, w_003_6227, w_003_6228, w_003_6229, w_003_6230, w_003_6231, w_003_6233, w_003_6234, w_003_6235, w_003_6236, w_003_6237, w_003_6238, w_003_6239, w_003_6241, w_003_6242, w_003_6243, w_003_6244, w_003_6246, w_003_6248, w_003_6249, w_003_6250, w_003_6251, w_003_6252, w_003_6253, w_003_6254, w_003_6256, w_003_6257, w_003_6258, w_003_6259, w_003_6260, w_003_6261, w_003_6262, w_003_6263, w_003_6264, w_003_6265, w_003_6266, w_003_6267, w_003_6268, w_003_6270, w_003_6271, w_003_6272, w_003_6273, w_003_6275, w_003_6276, w_003_6277, w_003_6278, w_003_6280, w_003_6281, w_003_6282, w_003_6283, w_003_6284, w_003_6285, w_003_6287, w_003_6288, w_003_6289, w_003_6290, w_003_6291, w_003_6293, w_003_6294, w_003_6295, w_003_6296, w_003_6297, w_003_6298, w_003_6299, w_003_6300, w_003_6301, w_003_6303, w_003_6304, w_003_6305, w_003_6306, w_003_6307, w_003_6308, w_003_6309, w_003_6310, w_003_6311, w_003_6312, w_003_6313, w_003_6314, w_003_6317, w_003_6318, w_003_6319, w_003_6320, w_003_6321, w_003_6322, w_003_6323, w_003_6324, w_003_6325, w_003_6326, w_003_6327, w_003_6328, w_003_6329, w_003_6331, w_003_6332, w_003_6333, w_003_6334, w_003_6335, w_003_6336, w_003_6337, w_003_6338, w_003_6339, w_003_6340, w_003_6341, w_003_6342, w_003_6343, w_003_6345, w_003_6346, w_003_6347, w_003_6348, w_003_6350, w_003_6351, w_003_6352, w_003_6353, w_003_6354, w_003_6356, w_003_6357, w_003_6358, w_003_6359, w_003_6360, w_003_6361, w_003_6362, w_003_6363, w_003_6364, w_003_6365, w_003_6366, w_003_6367, w_003_6368, w_003_6370, w_003_6372, w_003_6373, w_003_6374, w_003_6375, w_003_6376, w_003_6378, w_003_6380, w_003_6381, w_003_6382, w_003_6383, w_003_6384, w_003_6385, w_003_6386, w_003_6387, w_003_6390, w_003_6391, w_003_6392, w_003_6393, w_003_6394, w_003_6395, w_003_6396, w_003_6397, w_003_6398, w_003_6400, w_003_6401, w_003_6402, w_003_6403, w_003_6404, w_003_6405, w_003_6407, w_003_6408, w_003_6409, w_003_6410, w_003_6411, w_003_6412, w_003_6413, w_003_6414, w_003_6415, w_003_6416, w_003_6417, w_003_6418, w_003_6421, w_003_6422, w_003_6423, w_003_6424, w_003_6425, w_003_6426, w_003_6427, w_003_6428, w_003_6429, w_003_6430, w_003_6431, w_003_6432, w_003_6433, w_003_6434, w_003_6435, w_003_6437, w_003_6438, w_003_6439, w_003_6440, w_003_6441, w_003_6442, w_003_6443, w_003_6444, w_003_6445, w_003_6446, w_003_6447, w_003_6448, w_003_6449, w_003_6450, w_003_6451, w_003_6452, w_003_6453, w_003_6454, w_003_6455, w_003_6456, w_003_6458, w_003_6459, w_003_6460, w_003_6461, w_003_6462, w_003_6463, w_003_6464, w_003_6465, w_003_6466, w_003_6467, w_003_6468, w_003_6470, w_003_6471, w_003_6472, w_003_6473, w_003_6474, w_003_6475, w_003_6477, w_003_6478, w_003_6479, w_003_6481, w_003_6482, w_003_6484, w_003_6485, w_003_6486, w_003_6487, w_003_6488, w_003_6489, w_003_6490, w_003_6491, w_003_6492, w_003_6493, w_003_6494, w_003_6495, w_003_6496, w_003_6499, w_003_6502, w_003_6503, w_003_6504, w_003_6505, w_003_6506, w_003_6507, w_003_6508, w_003_6509, w_003_6510, w_003_6511, w_003_6512, w_003_6513, w_003_6514, w_003_6515, w_003_6517, w_003_6519, w_003_6520, w_003_6521, w_003_6522, w_003_6523, w_003_6524, w_003_6525, w_003_6526, w_003_6527, w_003_6528, w_003_6529, w_003_6530, w_003_6531, w_003_6532, w_003_6533, w_003_6534, w_003_6535, w_003_6537, w_003_6538, w_003_6539, w_003_6540, w_003_6542, w_003_6543, w_003_6544, w_003_6547, w_003_6551, w_003_6553, w_003_6555, w_003_6557, w_003_6558, w_003_6559, w_003_6560, w_003_6561, w_003_6562, w_003_6564, w_003_6565, w_003_6566, w_003_6567, w_003_6569, w_003_6570, w_003_6571, w_003_6572, w_003_6573, w_003_6574, w_003_6575, w_003_6576, w_003_6577, w_003_6578, w_003_6579, w_003_6580, w_003_6581, w_003_6582, w_003_6583, w_003_6587, w_003_6588, w_003_6589, w_003_6590, w_003_6591, w_003_6592, w_003_6593, w_003_6594, w_003_6595, w_003_6596, w_003_6597, w_003_6599, w_003_6600, w_003_6601, w_003_6602, w_003_6603, w_003_6604, w_003_6605, w_003_6606, w_003_6607, w_003_6608, w_003_6609, w_003_6610, w_003_6611, w_003_6612, w_003_6613, w_003_6614, w_003_6615, w_003_6616, w_003_6617, w_003_6618, w_003_6619, w_003_6620, w_003_6622, w_003_6623, w_003_6624, w_003_6625, w_003_6626, w_003_6628, w_003_6630, w_003_6631, w_003_6632, w_003_6634, w_003_6635, w_003_6636, w_003_6637, w_003_6639, w_003_6640, w_003_6641, w_003_6642, w_003_6643, w_003_6644, w_003_6645, w_003_6646, w_003_6648, w_003_6649, w_003_6650, w_003_6651, w_003_6652, w_003_6653, w_003_6654, w_003_6655, w_003_6656, w_003_6657, w_003_6658, w_003_6660, w_003_6661, w_003_6662, w_003_6664, w_003_6665, w_003_6666, w_003_6668, w_003_6669, w_003_6672, w_003_6673, w_003_6674, w_003_6676, w_003_6677, w_003_6678, w_003_6679, w_003_6680, w_003_6681, w_003_6682, w_003_6683, w_003_6684, w_003_6685, w_003_6686, w_003_6687, w_003_6688, w_003_6689, w_003_6690, w_003_6691, w_003_6692, w_003_6693, w_003_6695, w_003_6696, w_003_6697, w_003_6698, w_003_6700, w_003_6701, w_003_6702, w_003_6703, w_003_6704, w_003_6705, w_003_6706, w_003_6707, w_003_6708, w_003_6709, w_003_6710, w_003_6711, w_003_6712, w_003_6713, w_003_6714, w_003_6715, w_003_6716, w_003_6718, w_003_6719, w_003_6720, w_003_6721, w_003_6722, w_003_6723, w_003_6724, w_003_6725, w_003_6726, w_003_6727, w_003_6728, w_003_6729, w_003_6730, w_003_6731, w_003_6732, w_003_6733, w_003_6734, w_003_6736, w_003_6737, w_003_6738, w_003_6739, w_003_6741, w_003_6742, w_003_6743, w_003_6744, w_003_6745, w_003_6746, w_003_6747, w_003_6748, w_003_6749, w_003_6750, w_003_6751, w_003_6753, w_003_6754, w_003_6755, w_003_6756, w_003_6757, w_003_6758, w_003_6759, w_003_6760, w_003_6761, w_003_6762, w_003_6765, w_003_6766, w_003_6767, w_003_6768, w_003_6769, w_003_6770, w_003_6771, w_003_6772, w_003_6773, w_003_6774, w_003_6775, w_003_6777, w_003_6778, w_003_6779, w_003_6781, w_003_6782, w_003_6783, w_003_6784, w_003_6785, w_003_6786, w_003_6787, w_003_6788, w_003_6789, w_003_6790, w_003_6791, w_003_6792, w_003_6793, w_003_6794, w_003_6795, w_003_6796, w_003_6798, w_003_6799, w_003_6800, w_003_6801, w_003_6802, w_003_6803, w_003_6804, w_003_6805, w_003_6806, w_003_6807, w_003_6808, w_003_6809, w_003_6811, w_003_6812, w_003_6813, w_003_6815, w_003_6816, w_003_6817, w_003_6818, w_003_6819, w_003_6820, w_003_6821, w_003_6822, w_003_6823, w_003_6825, w_003_6826, w_003_6827, w_003_6828, w_003_6829, w_003_6830, w_003_6832, w_003_6833, w_003_6834, w_003_6835, w_003_6836, w_003_6837, w_003_6838, w_003_6839, w_003_6840, w_003_6841, w_003_6842, w_003_6843, w_003_6844, w_003_6845, w_003_6846, w_003_6847, w_003_6848, w_003_6849, w_003_6851, w_003_6852, w_003_6853, w_003_6854, w_003_6855, w_003_6856, w_003_6857, w_003_6858, w_003_6859, w_003_6860, w_003_6861, w_003_6862, w_003_6863, w_003_6864, w_003_6865, w_003_6866, w_003_6867, w_003_6868, w_003_6869, w_003_6870, w_003_6871, w_003_6872, w_003_6873, w_003_6874, w_003_6876, w_003_6877, w_003_6878, w_003_6879, w_003_6882, w_003_6883, w_003_6884, w_003_6885, w_003_6886, w_003_6887, w_003_6888, w_003_6889, w_003_6891, w_003_6892, w_003_6893, w_003_6894, w_003_6895, w_003_6896, w_003_6897, w_003_6898, w_003_6899, w_003_6900, w_003_6901, w_003_6902, w_003_6903, w_003_6904, w_003_6905, w_003_6906, w_003_6907, w_003_6908, w_003_6909, w_003_6910, w_003_6911, w_003_6912, w_003_6913, w_003_6914, w_003_6915, w_003_6916, w_003_6917, w_003_6918, w_003_6919, w_003_6920, w_003_6921, w_003_6922, w_003_6923, w_003_6924, w_003_6925, w_003_6926, w_003_6927, w_003_6928, w_003_6929, w_003_6930, w_003_6931, w_003_6932, w_003_6933, w_003_6934, w_003_6935, w_003_6936, w_003_6937, w_003_6940, w_003_6941, w_003_6942, w_003_6943, w_003_6944, w_003_6945, w_003_6946, w_003_6947, w_003_6949, w_003_6950, w_003_6951, w_003_6952, w_003_6953, w_003_6954, w_003_6956, w_003_6957, w_003_6958, w_003_6959, w_003_6961, w_003_6963, w_003_6964, w_003_6965, w_003_6967, w_003_6968, w_003_6971, w_003_6972, w_003_6973, w_003_6974, w_003_6975, w_003_6976, w_003_6978, w_003_6979, w_003_6981, w_003_6982, w_003_6983, w_003_6984, w_003_6985, w_003_6986, w_003_6987, w_003_6989, w_003_6990, w_003_6991, w_003_6992, w_003_6994, w_003_6995, w_003_6997, w_003_6998, w_003_6999, w_003_7000, w_003_7001, w_003_7003, w_003_7004, w_003_7005, w_003_7006, w_003_7007, w_003_7008, w_003_7009, w_003_7010, w_003_7011, w_003_7012, w_003_7013, w_003_7014, w_003_7015, w_003_7016, w_003_7017, w_003_7018, w_003_7019, w_003_7021, w_003_7022, w_003_7023, w_003_7024, w_003_7026, w_003_7027, w_003_7028, w_003_7029, w_003_7030, w_003_7031, w_003_7032, w_003_7033, w_003_7034, w_003_7035, w_003_7036, w_003_7037, w_003_7038, w_003_7039, w_003_7040, w_003_7041, w_003_7044, w_003_7045, w_003_7046, w_003_7047, w_003_7048, w_003_7049, w_003_7050, w_003_7051, w_003_7052, w_003_7053, w_003_7054, w_003_7055, w_003_7057, w_003_7058, w_003_7059, w_003_7060, w_003_7062, w_003_7063, w_003_7064, w_003_7066, w_003_7067, w_003_7068, w_003_7069, w_003_7070, w_003_7071, w_003_7072, w_003_7073, w_003_7074, w_003_7075, w_003_7076, w_003_7077, w_003_7078, w_003_7079, w_003_7080, w_003_7081, w_003_7082, w_003_7083, w_003_7084, w_003_7086, w_003_7087, w_003_7088, w_003_7089, w_003_7090, w_003_7091, w_003_7093, w_003_7094, w_003_7095, w_003_7096, w_003_7097, w_003_7099, w_003_7101, w_003_7103, w_003_7104, w_003_7105, w_003_7106, w_003_7107, w_003_7108, w_003_7109, w_003_7110, w_003_7112, w_003_7113, w_003_7114, w_003_7115, w_003_7116, w_003_7118, w_003_7119, w_003_7120, w_003_7121, w_003_7122, w_003_7123, w_003_7125, w_003_7126, w_003_7129, w_003_7130, w_003_7133, w_003_7134, w_003_7135, w_003_7136, w_003_7137, w_003_7138, w_003_7139, w_003_7140, w_003_7141, w_003_7142, w_003_7143, w_003_7144, w_003_7145, w_003_7146, w_003_7147, w_003_7148, w_003_7149, w_003_7150, w_003_7151, w_003_7152, w_003_7153, w_003_7154, w_003_7155, w_003_7156, w_003_7157, w_003_7158, w_003_7159, w_003_7161, w_003_7162, w_003_7163, w_003_7164, w_003_7165, w_003_7166, w_003_7167, w_003_7168, w_003_7169, w_003_7170, w_003_7172, w_003_7174, w_003_7175, w_003_7176, w_003_7177, w_003_7178, w_003_7179, w_003_7180, w_003_7181, w_003_7182, w_003_7183, w_003_7184, w_003_7185, w_003_7186, w_003_7187, w_003_7190, w_003_7191, w_003_7193, w_003_7194, w_003_7195, w_003_7196, w_003_7198, w_003_7199, w_003_7200, w_003_7201, w_003_7202, w_003_7203, w_003_7205, w_003_7206, w_003_7207, w_003_7208, w_003_7209, w_003_7210, w_003_7211, w_003_7212, w_003_7213, w_003_7214, w_003_7215, w_003_7216, w_003_7217, w_003_7218, w_003_7219, w_003_7220, w_003_7221, w_003_7222, w_003_7223, w_003_7224, w_003_7226, w_003_7227, w_003_7228, w_003_7229, w_003_7230, w_003_7231, w_003_7232, w_003_7233, w_003_7235, w_003_7236, w_003_7237, w_003_7238, w_003_7239, w_003_7240, w_003_7242, w_003_7243, w_003_7244, w_003_7246, w_003_7247, w_003_7248, w_003_7249, w_003_7250, w_003_7251, w_003_7252, w_003_7253, w_003_7254, w_003_7255, w_003_7256, w_003_7257, w_003_7258, w_003_7260, w_003_7261, w_003_7262, w_003_7263, w_003_7264, w_003_7265, w_003_7266, w_003_7267, w_003_7269, w_003_7270, w_003_7271, w_003_7273, w_003_7274, w_003_7275, w_003_7276, w_003_7277, w_003_7278, w_003_7279, w_003_7281, w_003_7282, w_003_7283, w_003_7284, w_003_7285, w_003_7286, w_003_7287, w_003_7288, w_003_7289, w_003_7290, w_003_7291, w_003_7292, w_003_7293, w_003_7295, w_003_7296, w_003_7297, w_003_7299, w_003_7301, w_003_7303, w_003_7304, w_003_7305, w_003_7307, w_003_7309, w_003_7311, w_003_7312, w_003_7313, w_003_7314, w_003_7316, w_003_7317, w_003_7318, w_003_7319, w_003_7320, w_003_7321, w_003_7322, w_003_7323, w_003_7324, w_003_7325, w_003_7326, w_003_7327, w_003_7328, w_003_7329, w_003_7330, w_003_7331, w_003_7332, w_003_7333, w_003_7334, w_003_7337, w_003_7339, w_003_7340, w_003_7341, w_003_7342, w_003_7343, w_003_7344, w_003_7346, w_003_7347, w_003_7348, w_003_7349, w_003_7350, w_003_7351, w_003_7352, w_003_7353, w_003_7354, w_003_7355, w_003_7356, w_003_7357, w_003_7358, w_003_7359, w_003_7360, w_003_7361, w_003_7362, w_003_7363, w_003_7364, w_003_7366, w_003_7368, w_003_7369, w_003_7371, w_003_7372, w_003_7373, w_003_7374, w_003_7375, w_003_7376, w_003_7377, w_003_7378, w_003_7379, w_003_7380, w_003_7381, w_003_7382, w_003_7383, w_003_7384, w_003_7385, w_003_7386, w_003_7387, w_003_7388, w_003_7389, w_003_7390, w_003_7391, w_003_7393, w_003_7394, w_003_7395, w_003_7396, w_003_7397, w_003_7398, w_003_7399, w_003_7400, w_003_7401, w_003_7402, w_003_7403, w_003_7405, w_003_7407, w_003_7408, w_003_7410, w_003_7411, w_003_7412, w_003_7413, w_003_7414, w_003_7415, w_003_7416, w_003_7417, w_003_7418, w_003_7419, w_003_7420, w_003_7421, w_003_7422, w_003_7423, w_003_7424, w_003_7427, w_003_7428, w_003_7429, w_003_7430, w_003_7431, w_003_7432, w_003_7433, w_003_7435, w_003_7436, w_003_7437, w_003_7438, w_003_7439, w_003_7440, w_003_7441, w_003_7442, w_003_7444, w_003_7445, w_003_7446, w_003_7447, w_003_7448, w_003_7450, w_003_7451, w_003_7452, w_003_7453, w_003_7454, w_003_7455, w_003_7456, w_003_7457, w_003_7458, w_003_7459, w_003_7460, w_003_7462, w_003_7463, w_003_7464, w_003_7466, w_003_7467, w_003_7468, w_003_7470, w_003_7471, w_003_7472, w_003_7473, w_003_7474, w_003_7475, w_003_7476, w_003_7477, w_003_7478, w_003_7480, w_003_7481, w_003_7482, w_003_7483, w_003_7484, w_003_7485, w_003_7486, w_003_7487, w_003_7488, w_003_7489, w_003_7490, w_003_7491, w_003_7492, w_003_7493, w_003_7494, w_003_7495, w_003_7496, w_003_7497, w_003_7498, w_003_7499, w_003_7500, w_003_7502, w_003_7503, w_003_7504, w_003_7505, w_003_7506, w_003_7507, w_003_7508, w_003_7509, w_003_7510, w_003_7512, w_003_7513, w_003_7514, w_003_7516, w_003_7517, w_003_7519, w_003_7520, w_003_7521, w_003_7522, w_003_7523, w_003_7524, w_003_7525, w_003_7526, w_003_7529, w_003_7530, w_003_7531, w_003_7532, w_003_7533, w_003_7535, w_003_7536, w_003_7537, w_003_7538, w_003_7539, w_003_7540, w_003_7541, w_003_7542, w_003_7543, w_003_7545, w_003_7546, w_003_7547, w_003_7548, w_003_7551, w_003_7552, w_003_7553, w_003_7554, w_003_7555, w_003_7556, w_003_7557, w_003_7559, w_003_7560, w_003_7561, w_003_7562, w_003_7563, w_003_7566, w_003_7567, w_003_7568, w_003_7570, w_003_7571, w_003_7572, w_003_7574, w_003_7575, w_003_7576, w_003_7577, w_003_7578, w_003_7579, w_003_7580, w_003_7581, w_003_7583, w_003_7584, w_003_7586, w_003_7587, w_003_7588, w_003_7589, w_003_7590, w_003_7591, w_003_7592, w_003_7593, w_003_7594, w_003_7596, w_003_7597, w_003_7598, w_003_7600, w_003_7601, w_003_7602, w_003_7603, w_003_7604, w_003_7605, w_003_7606, w_003_7607, w_003_7608, w_003_7610, w_003_7611, w_003_7613, w_003_7614, w_003_7615, w_003_7616, w_003_7617, w_003_7618, w_003_7619, w_003_7620, w_003_7621, w_003_7622, w_003_7623, w_003_7624, w_003_7625, w_003_7627, w_003_7628, w_003_7629, w_003_7630, w_003_7631, w_003_7632, w_003_7637, w_003_7638, w_003_7639, w_003_7640, w_003_7641, w_003_7642, w_003_7643, w_003_7644, w_003_7645, w_003_7646, w_003_7647, w_003_7648, w_003_7649, w_003_7650, w_003_7651, w_003_7652, w_003_7653, w_003_7654, w_003_7655, w_003_7656, w_003_7658, w_003_7659, w_003_7660, w_003_7661, w_003_7662, w_003_7663, w_003_7664, w_003_7665, w_003_7666, w_003_7667, w_003_7668, w_003_7669, w_003_7670, w_003_7672, w_003_7673, w_003_7674, w_003_7675, w_003_7676, w_003_7677, w_003_7678, w_003_7680, w_003_7681, w_003_7682, w_003_7683, w_003_7684, w_003_7685, w_003_7686, w_003_7687, w_003_7688, w_003_7689, w_003_7690, w_003_7692, w_003_7693, w_003_7694, w_003_7695, w_003_7697, w_003_7698, w_003_7699, w_003_7700, w_003_7701, w_003_7702, w_003_7703, w_003_7705, w_003_7706, w_003_7707, w_003_7708, w_003_7709, w_003_7710, w_003_7711, w_003_7712, w_003_7713, w_003_7714, w_003_7715, w_003_7716, w_003_7717, w_003_7719, w_003_7720, w_003_7721, w_003_7722, w_003_7724, w_003_7725, w_003_7726, w_003_7727, w_003_7728, w_003_7730, w_003_7731, w_003_7732, w_003_7733, w_003_7734, w_003_7735, w_003_7737, w_003_7738, w_003_7739, w_003_7740, w_003_7742, w_003_7743, w_003_7744, w_003_7746, w_003_7747, w_003_7748, w_003_7749, w_003_7750, w_003_7751, w_003_7752, w_003_7753, w_003_7754, w_003_7756, w_003_7757, w_003_7758, w_003_7759, w_003_7761, w_003_7762, w_003_7763, w_003_7764, w_003_7765, w_003_7766, w_003_7767, w_003_7768, w_003_7769, w_003_7770, w_003_7771, w_003_7772, w_003_7773, w_003_7774, w_003_7776, w_003_7779, w_003_7781, w_003_7783, w_003_7784, w_003_7786, w_003_7787, w_003_7788, w_003_7789, w_003_7791, w_003_7792, w_003_7793, w_003_7794, w_003_7795, w_003_7796, w_003_7797, w_003_7798, w_003_7799, w_003_7800, w_003_7801, w_003_7802, w_003_7803, w_003_7804, w_003_7805, w_003_7806, w_003_7808, w_003_7809, w_003_7810, w_003_7811, w_003_7812, w_003_7813, w_003_7814, w_003_7815, w_003_7817, w_003_7818, w_003_7819, w_003_7820, w_003_7821, w_003_7822, w_003_7823, w_003_7824, w_003_7825, w_003_7827, w_003_7828, w_003_7829, w_003_7830, w_003_7831, w_003_7832, w_003_7833, w_003_7834, w_003_7835, w_003_7836, w_003_7837, w_003_7839, w_003_7840, w_003_7841, w_003_7842, w_003_7843, w_003_7844, w_003_7845, w_003_7846, w_003_7847, w_003_7848, w_003_7849, w_003_7850, w_003_7851, w_003_7852, w_003_7853, w_003_7854, w_003_7855, w_003_7856, w_003_7857, w_003_7858, w_003_7860, w_003_7861, w_003_7862, w_003_7863, w_003_7864, w_003_7865, w_003_7866, w_003_7867, w_003_7868, w_003_7871, w_003_7872, w_003_7873, w_003_7874, w_003_7875, w_003_7876, w_003_7878, w_003_7879, w_003_7880, w_003_7881, w_003_7882, w_003_7883, w_003_7884, w_003_7885, w_003_7886, w_003_7887, w_003_7889, w_003_7890, w_003_7891, w_003_7892, w_003_7893, w_003_7894, w_003_7895, w_003_7896, w_003_7897, w_003_7898, w_003_7899, w_003_7901, w_003_7902, w_003_7903, w_003_7904, w_003_7905, w_003_7906, w_003_7907, w_003_7908, w_003_7909, w_003_7910, w_003_7913, w_003_7914, w_003_7915, w_003_7916, w_003_7917, w_003_7918, w_003_7919, w_003_7920, w_003_7922, w_003_7923, w_003_7925, w_003_7926, w_003_7927, w_003_7928, w_003_7929, w_003_7931, w_003_7932, w_003_7933, w_003_7934, w_003_7935, w_003_7936, w_003_7938, w_003_7939, w_003_7940, w_003_7941, w_003_7942;
  wire w_004_000, w_004_001, w_004_002, w_004_003, w_004_004, w_004_005, w_004_006, w_004_007, w_004_008, w_004_009, w_004_010, w_004_011, w_004_012, w_004_013, w_004_014, w_004_015, w_004_016, w_004_017, w_004_018, w_004_019, w_004_020, w_004_021, w_004_022, w_004_023, w_004_024, w_004_025, w_004_026, w_004_027, w_004_028, w_004_029, w_004_030, w_004_031, w_004_032, w_004_033, w_004_034, w_004_035, w_004_036, w_004_037, w_004_038, w_004_039, w_004_040, w_004_041, w_004_042, w_004_043, w_004_044, w_004_045, w_004_046, w_004_047, w_004_048, w_004_049, w_004_050, w_004_051, w_004_052, w_004_053, w_004_054, w_004_055, w_004_056, w_004_057, w_004_058, w_004_059, w_004_060, w_004_061, w_004_062, w_004_063, w_004_064, w_004_065, w_004_066, w_004_067, w_004_068, w_004_069, w_004_070, w_004_071, w_004_072, w_004_073, w_004_074, w_004_075, w_004_076, w_004_077, w_004_078, w_004_079, w_004_080, w_004_081, w_004_082, w_004_083, w_004_084, w_004_085, w_004_086, w_004_087, w_004_088, w_004_089, w_004_090, w_004_091, w_004_092, w_004_093, w_004_094, w_004_095, w_004_096, w_004_097, w_004_098, w_004_099, w_004_100, w_004_101, w_004_102, w_004_103, w_004_104, w_004_105, w_004_106, w_004_107, w_004_108, w_004_109, w_004_110, w_004_111, w_004_112, w_004_113, w_004_114, w_004_115, w_004_116, w_004_117, w_004_118, w_004_119, w_004_120, w_004_121, w_004_122, w_004_123, w_004_124, w_004_125, w_004_126, w_004_127, w_004_128, w_004_129, w_004_130, w_004_131, w_004_132, w_004_133, w_004_134, w_004_135, w_004_136, w_004_137, w_004_138, w_004_139, w_004_140, w_004_141, w_004_142, w_004_143, w_004_144, w_004_145, w_004_146, w_004_147, w_004_148, w_004_149, w_004_150, w_004_151, w_004_152, w_004_153, w_004_154, w_004_155, w_004_156, w_004_157, w_004_158, w_004_159, w_004_160, w_004_161, w_004_162, w_004_163, w_004_164, w_004_165, w_004_166, w_004_167, w_004_168, w_004_169, w_004_170, w_004_171, w_004_172, w_004_173, w_004_174, w_004_175, w_004_176, w_004_177, w_004_178, w_004_179, w_004_180, w_004_181, w_004_182, w_004_183, w_004_184, w_004_185, w_004_186, w_004_187, w_004_188, w_004_189, w_004_190, w_004_191, w_004_192, w_004_193, w_004_194, w_004_195, w_004_196, w_004_197, w_004_198, w_004_199, w_004_200, w_004_201, w_004_202, w_004_203, w_004_204, w_004_205, w_004_206, w_004_207, w_004_208, w_004_209, w_004_210, w_004_211, w_004_212, w_004_213, w_004_214, w_004_215, w_004_216, w_004_217, w_004_218, w_004_219, w_004_220, w_004_221, w_004_222, w_004_223, w_004_224, w_004_225, w_004_226, w_004_227, w_004_228, w_004_229, w_004_230, w_004_231, w_004_232, w_004_233, w_004_234, w_004_235, w_004_236, w_004_237, w_004_238, w_004_239, w_004_240, w_004_241, w_004_242, w_004_243, w_004_244, w_004_245, w_004_246, w_004_247, w_004_248, w_004_249, w_004_250, w_004_251, w_004_252, w_004_253, w_004_254, w_004_255, w_004_256, w_004_257, w_004_258, w_004_259, w_004_260, w_004_261, w_004_262, w_004_263, w_004_264, w_004_265, w_004_266, w_004_267, w_004_268, w_004_269, w_004_270, w_004_271, w_004_272, w_004_273, w_004_274, w_004_275, w_004_276, w_004_277, w_004_278, w_004_279, w_004_280, w_004_281, w_004_282, w_004_283, w_004_284, w_004_285, w_004_286, w_004_287, w_004_288, w_004_289, w_004_290, w_004_291, w_004_292, w_004_293, w_004_294, w_004_295, w_004_296, w_004_297, w_004_298, w_004_299, w_004_300, w_004_301, w_004_302, w_004_303, w_004_304, w_004_305, w_004_306, w_004_307, w_004_308, w_004_309, w_004_310, w_004_311, w_004_312, w_004_313, w_004_314, w_004_315, w_004_316, w_004_317, w_004_318, w_004_319, w_004_320, w_004_321, w_004_322, w_004_323, w_004_324, w_004_325, w_004_326, w_004_327, w_004_328, w_004_329, w_004_330, w_004_331, w_004_332, w_004_333, w_004_334, w_004_335, w_004_336, w_004_337, w_004_338, w_004_339, w_004_340, w_004_341, w_004_342, w_004_343, w_004_344, w_004_345, w_004_346, w_004_347, w_004_348, w_004_349, w_004_350, w_004_351, w_004_352, w_004_353, w_004_354, w_004_355, w_004_356, w_004_357, w_004_358, w_004_359, w_004_360, w_004_361, w_004_362, w_004_363, w_004_364, w_004_365, w_004_366, w_004_367, w_004_368, w_004_369, w_004_370, w_004_371, w_004_372, w_004_373, w_004_374, w_004_375, w_004_376, w_004_377, w_004_378, w_004_379, w_004_380, w_004_381, w_004_382, w_004_383, w_004_384, w_004_385, w_004_386, w_004_387, w_004_388, w_004_389, w_004_390, w_004_391, w_004_392, w_004_393, w_004_394, w_004_395, w_004_396, w_004_397, w_004_398, w_004_399, w_004_400, w_004_401, w_004_402, w_004_403, w_004_404, w_004_405, w_004_406, w_004_407, w_004_408, w_004_409, w_004_410, w_004_411, w_004_412, w_004_413, w_004_414, w_004_415, w_004_416, w_004_417, w_004_418, w_004_419, w_004_420, w_004_421, w_004_422, w_004_423, w_004_424, w_004_425, w_004_426, w_004_427, w_004_428, w_004_429, w_004_430, w_004_431, w_004_432, w_004_433, w_004_434, w_004_435, w_004_436, w_004_437, w_004_438, w_004_439, w_004_440, w_004_441, w_004_442, w_004_443, w_004_444, w_004_445, w_004_446, w_004_447, w_004_448, w_004_449, w_004_450, w_004_451, w_004_452, w_004_453, w_004_454, w_004_455, w_004_456, w_004_457, w_004_458, w_004_459, w_004_460, w_004_461, w_004_462, w_004_463, w_004_464, w_004_465, w_004_466, w_004_467, w_004_468, w_004_469, w_004_470, w_004_471, w_004_472, w_004_473, w_004_474, w_004_475, w_004_476, w_004_477, w_004_478, w_004_479, w_004_480, w_004_481, w_004_482, w_004_483, w_004_484, w_004_485, w_004_486, w_004_487, w_004_488, w_004_489, w_004_490, w_004_491, w_004_492, w_004_493, w_004_494, w_004_495, w_004_496, w_004_497, w_004_498, w_004_499, w_004_500, w_004_501, w_004_502, w_004_503, w_004_504, w_004_505, w_004_506, w_004_507, w_004_508, w_004_509, w_004_510, w_004_511, w_004_512, w_004_513, w_004_514, w_004_515, w_004_516, w_004_517, w_004_518, w_004_519, w_004_520, w_004_521, w_004_522, w_004_523, w_004_524, w_004_525, w_004_526, w_004_527, w_004_528, w_004_529, w_004_530, w_004_531, w_004_532, w_004_533, w_004_534, w_004_535, w_004_536, w_004_537, w_004_538, w_004_539, w_004_540, w_004_541, w_004_542, w_004_543, w_004_544, w_004_545, w_004_546, w_004_547, w_004_548, w_004_549, w_004_550, w_004_551, w_004_552, w_004_553, w_004_554, w_004_555, w_004_556, w_004_557, w_004_558, w_004_559, w_004_560, w_004_561, w_004_562, w_004_563, w_004_564, w_004_565, w_004_566, w_004_567, w_004_568, w_004_569, w_004_570, w_004_571, w_004_572, w_004_573, w_004_574, w_004_575, w_004_576, w_004_577, w_004_578, w_004_579, w_004_580, w_004_581, w_004_582, w_004_583, w_004_584, w_004_585, w_004_586, w_004_587, w_004_588, w_004_589, w_004_590, w_004_591, w_004_592, w_004_593, w_004_594, w_004_595, w_004_596, w_004_597, w_004_598, w_004_599, w_004_600, w_004_601, w_004_602, w_004_603, w_004_604, w_004_605, w_004_606, w_004_607, w_004_608, w_004_609, w_004_610, w_004_611, w_004_612, w_004_613, w_004_614, w_004_615, w_004_616, w_004_617, w_004_618, w_004_619, w_004_620, w_004_621, w_004_622, w_004_623, w_004_624, w_004_625, w_004_626, w_004_627, w_004_628, w_004_629, w_004_630, w_004_631, w_004_632, w_004_633, w_004_634, w_004_635, w_004_636, w_004_637, w_004_638, w_004_639, w_004_640, w_004_641, w_004_642, w_004_643, w_004_644, w_004_645, w_004_646, w_004_647, w_004_648, w_004_649, w_004_650, w_004_651, w_004_652, w_004_653, w_004_654, w_004_655, w_004_656, w_004_657, w_004_658, w_004_659, w_004_660, w_004_661, w_004_662, w_004_663, w_004_664, w_004_665, w_004_666, w_004_667, w_004_668, w_004_669, w_004_670, w_004_671, w_004_672, w_004_673, w_004_674, w_004_675, w_004_676, w_004_677, w_004_678, w_004_679, w_004_680, w_004_681, w_004_682, w_004_683, w_004_684, w_004_685, w_004_686, w_004_687, w_004_688, w_004_689, w_004_690, w_004_691, w_004_692, w_004_693, w_004_694, w_004_695, w_004_696, w_004_697, w_004_698, w_004_699, w_004_700, w_004_701, w_004_702, w_004_703, w_004_704, w_004_705, w_004_706, w_004_707, w_004_708, w_004_709, w_004_710, w_004_711, w_004_712, w_004_713, w_004_714, w_004_715, w_004_716, w_004_717, w_004_718, w_004_719, w_004_720, w_004_721, w_004_722, w_004_723, w_004_724, w_004_725, w_004_726, w_004_727, w_004_728, w_004_729, w_004_730, w_004_731, w_004_732, w_004_733, w_004_734, w_004_735, w_004_736, w_004_737, w_004_738, w_004_739, w_004_740, w_004_741, w_004_742, w_004_743, w_004_744, w_004_745, w_004_746, w_004_747, w_004_748, w_004_749, w_004_750, w_004_751, w_004_752, w_004_753, w_004_754, w_004_755, w_004_756, w_004_757, w_004_758, w_004_759, w_004_760, w_004_761, w_004_762, w_004_763, w_004_764, w_004_765, w_004_766, w_004_767, w_004_768, w_004_769, w_004_770, w_004_771, w_004_772, w_004_773, w_004_774, w_004_775, w_004_776, w_004_777, w_004_778, w_004_779, w_004_780, w_004_781, w_004_782, w_004_783, w_004_784, w_004_785, w_004_786, w_004_787, w_004_788, w_004_789, w_004_790, w_004_791, w_004_792, w_004_793, w_004_794, w_004_795, w_004_796, w_004_797, w_004_798, w_004_799, w_004_800, w_004_801, w_004_802, w_004_803, w_004_804, w_004_805, w_004_806, w_004_807, w_004_808, w_004_809, w_004_810, w_004_811, w_004_812, w_004_813, w_004_814, w_004_815, w_004_816, w_004_817, w_004_818, w_004_819, w_004_820, w_004_821, w_004_822, w_004_823, w_004_824, w_004_825, w_004_826, w_004_827, w_004_828, w_004_829, w_004_830, w_004_831, w_004_832, w_004_833, w_004_834, w_004_835, w_004_836, w_004_837, w_004_838, w_004_839, w_004_840, w_004_841, w_004_842, w_004_843, w_004_844, w_004_845, w_004_846, w_004_847, w_004_848, w_004_849, w_004_850, w_004_851, w_004_852, w_004_853, w_004_854, w_004_855, w_004_856, w_004_857, w_004_858, w_004_859, w_004_860, w_004_861, w_004_862, w_004_863, w_004_864, w_004_865, w_004_866, w_004_867, w_004_868, w_004_869, w_004_870, w_004_871, w_004_872, w_004_873, w_004_874, w_004_875, w_004_876, w_004_877, w_004_878, w_004_879, w_004_880, w_004_881, w_004_882, w_004_883, w_004_884, w_004_885, w_004_886, w_004_887, w_004_888, w_004_889, w_004_890, w_004_891, w_004_892, w_004_893, w_004_894, w_004_895, w_004_896, w_004_897, w_004_898, w_004_899, w_004_900, w_004_901, w_004_902, w_004_903, w_004_904, w_004_905, w_004_906, w_004_907, w_004_908, w_004_909, w_004_910, w_004_911, w_004_912, w_004_913, w_004_914, w_004_915, w_004_916, w_004_917, w_004_918, w_004_919, w_004_920, w_004_921, w_004_922, w_004_923, w_004_924, w_004_925, w_004_926, w_004_927, w_004_928, w_004_929, w_004_930, w_004_931, w_004_932, w_004_933, w_004_934, w_004_935, w_004_936, w_004_937, w_004_938, w_004_939, w_004_940, w_004_941, w_004_942, w_004_943, w_004_944, w_004_945, w_004_946, w_004_947, w_004_948, w_004_949, w_004_950, w_004_951, w_004_952, w_004_953, w_004_954, w_004_955, w_004_956, w_004_957, w_004_958, w_004_959, w_004_960, w_004_961, w_004_962, w_004_963, w_004_964, w_004_965, w_004_966, w_004_967, w_004_968, w_004_969, w_004_970, w_004_971, w_004_972, w_004_973, w_004_974, w_004_975, w_004_976, w_004_977, w_004_978, w_004_979, w_004_980, w_004_981, w_004_982, w_004_983, w_004_984, w_004_985, w_004_986, w_004_987, w_004_988, w_004_989, w_004_990, w_004_991, w_004_992, w_004_993, w_004_994, w_004_995, w_004_996, w_004_997, w_004_998, w_004_999, w_004_1000, w_004_1001, w_004_1002, w_004_1003, w_004_1004, w_004_1005, w_004_1006, w_004_1007, w_004_1008, w_004_1009, w_004_1010, w_004_1011, w_004_1012, w_004_1013, w_004_1014, w_004_1015, w_004_1016, w_004_1017, w_004_1018, w_004_1019, w_004_1020, w_004_1021, w_004_1022, w_004_1023, w_004_1024, w_004_1025, w_004_1026, w_004_1027, w_004_1028, w_004_1029, w_004_1030, w_004_1031, w_004_1032, w_004_1033, w_004_1034, w_004_1035, w_004_1036, w_004_1037, w_004_1038, w_004_1039, w_004_1040, w_004_1041, w_004_1042, w_004_1043, w_004_1044, w_004_1045, w_004_1046, w_004_1047, w_004_1048, w_004_1049, w_004_1050, w_004_1051, w_004_1052, w_004_1053, w_004_1054, w_004_1055, w_004_1056, w_004_1057, w_004_1058, w_004_1059, w_004_1060, w_004_1061, w_004_1062, w_004_1063, w_004_1064, w_004_1065, w_004_1066, w_004_1067, w_004_1068, w_004_1069, w_004_1070, w_004_1071, w_004_1072, w_004_1073, w_004_1074, w_004_1075, w_004_1076, w_004_1077, w_004_1078, w_004_1079, w_004_1080, w_004_1081, w_004_1082, w_004_1083, w_004_1084, w_004_1085, w_004_1086, w_004_1087, w_004_1088, w_004_1089, w_004_1090, w_004_1091, w_004_1092, w_004_1093, w_004_1094, w_004_1095, w_004_1096, w_004_1097, w_004_1098, w_004_1099, w_004_1100, w_004_1101, w_004_1102, w_004_1103, w_004_1104, w_004_1105, w_004_1106, w_004_1107, w_004_1108, w_004_1109, w_004_1110, w_004_1111, w_004_1112, w_004_1113, w_004_1114, w_004_1115, w_004_1116, w_004_1117, w_004_1118, w_004_1119, w_004_1120, w_004_1121, w_004_1122, w_004_1123, w_004_1124, w_004_1125, w_004_1126, w_004_1127, w_004_1128, w_004_1129, w_004_1130, w_004_1131, w_004_1132, w_004_1133, w_004_1134, w_004_1135, w_004_1136, w_004_1137, w_004_1138, w_004_1139, w_004_1140, w_004_1141, w_004_1142, w_004_1143, w_004_1144, w_004_1145, w_004_1146, w_004_1147, w_004_1148, w_004_1149, w_004_1150, w_004_1151, w_004_1152, w_004_1153, w_004_1154, w_004_1155, w_004_1156, w_004_1157, w_004_1158, w_004_1159, w_004_1160, w_004_1161, w_004_1162, w_004_1163, w_004_1164, w_004_1165, w_004_1166, w_004_1167, w_004_1168, w_004_1169, w_004_1170, w_004_1171, w_004_1172, w_004_1173, w_004_1174, w_004_1175, w_004_1176, w_004_1177, w_004_1178, w_004_1179, w_004_1180, w_004_1181, w_004_1182, w_004_1183, w_004_1184, w_004_1185, w_004_1186, w_004_1187, w_004_1188, w_004_1189, w_004_1190, w_004_1191, w_004_1192, w_004_1193, w_004_1194, w_004_1195, w_004_1196, w_004_1197, w_004_1198, w_004_1199, w_004_1200, w_004_1201, w_004_1202, w_004_1203, w_004_1204, w_004_1205, w_004_1206, w_004_1207, w_004_1208, w_004_1209, w_004_1210, w_004_1211, w_004_1212, w_004_1213, w_004_1214, w_004_1215, w_004_1216, w_004_1217, w_004_1218, w_004_1219, w_004_1220, w_004_1221, w_004_1222, w_004_1224, w_004_1225, w_004_1226, w_004_1227, w_004_1228, w_004_1229, w_004_1230, w_004_1231, w_004_1232, w_004_1233, w_004_1234, w_004_1235, w_004_1236, w_004_1237, w_004_1238, w_004_1239, w_004_1240, w_004_1241, w_004_1242, w_004_1243, w_004_1244, w_004_1245, w_004_1246, w_004_1247, w_004_1248, w_004_1249, w_004_1250, w_004_1251, w_004_1252, w_004_1253, w_004_1254, w_004_1255, w_004_1256, w_004_1257, w_004_1258, w_004_1259, w_004_1260, w_004_1261, w_004_1262, w_004_1263, w_004_1264, w_004_1265, w_004_1266, w_004_1267, w_004_1268, w_004_1269, w_004_1270, w_004_1271, w_004_1272, w_004_1273, w_004_1274, w_004_1275, w_004_1276, w_004_1277, w_004_1278, w_004_1279, w_004_1280, w_004_1281, w_004_1282, w_004_1283, w_004_1284, w_004_1285, w_004_1286, w_004_1287, w_004_1288, w_004_1289, w_004_1290, w_004_1291, w_004_1292, w_004_1293, w_004_1294, w_004_1295, w_004_1296, w_004_1297, w_004_1298, w_004_1299, w_004_1300, w_004_1301, w_004_1302, w_004_1303, w_004_1304, w_004_1305, w_004_1306, w_004_1307, w_004_1308, w_004_1309, w_004_1310, w_004_1311, w_004_1312, w_004_1313, w_004_1314, w_004_1315, w_004_1316, w_004_1317, w_004_1318, w_004_1319, w_004_1320, w_004_1321, w_004_1322, w_004_1323, w_004_1324, w_004_1325, w_004_1326, w_004_1327, w_004_1328, w_004_1329, w_004_1330, w_004_1331, w_004_1332, w_004_1333, w_004_1334, w_004_1335, w_004_1336, w_004_1337, w_004_1338, w_004_1339, w_004_1340, w_004_1341, w_004_1342, w_004_1343, w_004_1344, w_004_1345, w_004_1346, w_004_1347, w_004_1348, w_004_1349, w_004_1350, w_004_1351, w_004_1352, w_004_1353, w_004_1354, w_004_1355, w_004_1356, w_004_1357, w_004_1358, w_004_1359, w_004_1360, w_004_1361, w_004_1362, w_004_1363, w_004_1364, w_004_1365, w_004_1366, w_004_1367, w_004_1368, w_004_1369, w_004_1370, w_004_1371, w_004_1372, w_004_1373, w_004_1374, w_004_1375, w_004_1376, w_004_1377, w_004_1378, w_004_1379, w_004_1380, w_004_1381, w_004_1382, w_004_1383, w_004_1384, w_004_1385, w_004_1386, w_004_1387, w_004_1388, w_004_1389, w_004_1390, w_004_1391, w_004_1392, w_004_1393, w_004_1394, w_004_1395, w_004_1396, w_004_1397, w_004_1398, w_004_1399, w_004_1400, w_004_1401, w_004_1402, w_004_1403, w_004_1404, w_004_1405, w_004_1406, w_004_1407, w_004_1408, w_004_1409, w_004_1410, w_004_1411, w_004_1412, w_004_1413, w_004_1414, w_004_1415, w_004_1416, w_004_1417, w_004_1418, w_004_1419, w_004_1420, w_004_1421, w_004_1422, w_004_1423, w_004_1424, w_004_1425, w_004_1426, w_004_1427, w_004_1428, w_004_1429, w_004_1430, w_004_1431, w_004_1432, w_004_1433, w_004_1434, w_004_1435, w_004_1436, w_004_1437, w_004_1438, w_004_1439, w_004_1440, w_004_1441, w_004_1442, w_004_1443, w_004_1444, w_004_1445, w_004_1446, w_004_1447, w_004_1448, w_004_1449, w_004_1450, w_004_1451, w_004_1452, w_004_1453, w_004_1454, w_004_1455, w_004_1456, w_004_1457, w_004_1458, w_004_1459, w_004_1460, w_004_1461, w_004_1462, w_004_1463, w_004_1464, w_004_1465, w_004_1466, w_004_1467, w_004_1468, w_004_1469, w_004_1470, w_004_1471, w_004_1472, w_004_1473, w_004_1474, w_004_1475, w_004_1476, w_004_1477, w_004_1478, w_004_1479, w_004_1480, w_004_1481, w_004_1482, w_004_1483, w_004_1484, w_004_1485, w_004_1486, w_004_1487, w_004_1488, w_004_1489, w_004_1490, w_004_1491, w_004_1492, w_004_1493, w_004_1494, w_004_1495, w_004_1496, w_004_1497, w_004_1498, w_004_1499, w_004_1500, w_004_1501, w_004_1502, w_004_1503, w_004_1504, w_004_1505, w_004_1506, w_004_1507, w_004_1508, w_004_1509, w_004_1510, w_004_1511, w_004_1512, w_004_1513, w_004_1514, w_004_1515, w_004_1516, w_004_1517, w_004_1518, w_004_1519, w_004_1520, w_004_1521, w_004_1522, w_004_1523, w_004_1524, w_004_1525, w_004_1526, w_004_1527, w_004_1528, w_004_1529, w_004_1530, w_004_1531, w_004_1532, w_004_1533, w_004_1534, w_004_1535, w_004_1536, w_004_1537, w_004_1538, w_004_1539, w_004_1540, w_004_1541, w_004_1542, w_004_1543, w_004_1544, w_004_1545, w_004_1546, w_004_1547, w_004_1548, w_004_1549, w_004_1550, w_004_1551, w_004_1552, w_004_1553, w_004_1554, w_004_1555, w_004_1556, w_004_1557, w_004_1558, w_004_1559, w_004_1560, w_004_1561, w_004_1562, w_004_1563, w_004_1564, w_004_1565, w_004_1566, w_004_1567, w_004_1568, w_004_1569, w_004_1570, w_004_1571, w_004_1572, w_004_1573, w_004_1574, w_004_1575, w_004_1576, w_004_1577, w_004_1578, w_004_1579, w_004_1580, w_004_1581, w_004_1582, w_004_1583, w_004_1584, w_004_1585, w_004_1586, w_004_1587, w_004_1588, w_004_1589, w_004_1590, w_004_1591, w_004_1592, w_004_1593, w_004_1594, w_004_1595, w_004_1596, w_004_1597, w_004_1598, w_004_1599, w_004_1600, w_004_1601, w_004_1602, w_004_1603, w_004_1604, w_004_1605, w_004_1606, w_004_1607, w_004_1608, w_004_1609, w_004_1610, w_004_1611, w_004_1612, w_004_1613, w_004_1614, w_004_1615, w_004_1616, w_004_1617, w_004_1618, w_004_1619, w_004_1620, w_004_1621, w_004_1622, w_004_1623, w_004_1624, w_004_1625, w_004_1626, w_004_1627, w_004_1628, w_004_1629, w_004_1630, w_004_1631, w_004_1632, w_004_1633, w_004_1634, w_004_1635, w_004_1636, w_004_1637, w_004_1638, w_004_1639, w_004_1640, w_004_1641, w_004_1642, w_004_1643, w_004_1644, w_004_1645, w_004_1646, w_004_1647, w_004_1648, w_004_1649, w_004_1650, w_004_1651, w_004_1652, w_004_1653, w_004_1654, w_004_1655, w_004_1656, w_004_1657, w_004_1658, w_004_1659, w_004_1660, w_004_1661, w_004_1662, w_004_1663, w_004_1664, w_004_1665, w_004_1666, w_004_1667, w_004_1668, w_004_1669, w_004_1670, w_004_1671, w_004_1672, w_004_1673, w_004_1674, w_004_1675, w_004_1676, w_004_1677, w_004_1678, w_004_1679, w_004_1680, w_004_1681, w_004_1682, w_004_1683, w_004_1684, w_004_1685, w_004_1686, w_004_1687, w_004_1688, w_004_1689, w_004_1690, w_004_1691, w_004_1692, w_004_1693, w_004_1694, w_004_1695, w_004_1696, w_004_1697, w_004_1698, w_004_1699, w_004_1700, w_004_1701, w_004_1702, w_004_1703, w_004_1704, w_004_1705, w_004_1706, w_004_1707, w_004_1708, w_004_1709, w_004_1710, w_004_1711, w_004_1712, w_004_1713, w_004_1714, w_004_1715, w_004_1716, w_004_1717, w_004_1718, w_004_1719, w_004_1720, w_004_1721, w_004_1722, w_004_1723, w_004_1724, w_004_1725, w_004_1726, w_004_1727, w_004_1728, w_004_1729, w_004_1730, w_004_1731, w_004_1732, w_004_1733, w_004_1734, w_004_1735, w_004_1736, w_004_1737, w_004_1738, w_004_1739, w_004_1740, w_004_1741, w_004_1742, w_004_1743, w_004_1744, w_004_1745, w_004_1746, w_004_1747, w_004_1748, w_004_1749, w_004_1750, w_004_1751, w_004_1752, w_004_1753, w_004_1754, w_004_1755, w_004_1756, w_004_1757, w_004_1758, w_004_1759, w_004_1760, w_004_1761, w_004_1762, w_004_1763, w_004_1764, w_004_1765, w_004_1766, w_004_1767, w_004_1768, w_004_1769, w_004_1770, w_004_1771, w_004_1772, w_004_1773, w_004_1774, w_004_1775, w_004_1776, w_004_1777, w_004_1779, w_004_1780, w_004_1781, w_004_1782, w_004_1783, w_004_1784, w_004_1785, w_004_1786, w_004_1787, w_004_1788, w_004_1789, w_004_1790, w_004_1791, w_004_1792, w_004_1793, w_004_1794, w_004_1795, w_004_1796, w_004_1797, w_004_1798, w_004_1799, w_004_1800, w_004_1801, w_004_1802, w_004_1803, w_004_1804, w_004_1805, w_004_1806, w_004_1807, w_004_1808, w_004_1809, w_004_1811, w_004_1812, w_004_1813, w_004_1814, w_004_1815, w_004_1816, w_004_1817, w_004_1818, w_004_1819, w_004_1820, w_004_1821, w_004_1822, w_004_1823, w_004_1824, w_004_1825, w_004_1826, w_004_1827, w_004_1828, w_004_1829, w_004_1830, w_004_1831, w_004_1832, w_004_1833, w_004_1834, w_004_1835, w_004_1836, w_004_1837, w_004_1838, w_004_1839, w_004_1840, w_004_1841, w_004_1842, w_004_1843, w_004_1844, w_004_1845, w_004_1846, w_004_1847, w_004_1848, w_004_1849, w_004_1850, w_004_1851, w_004_1852, w_004_1853, w_004_1854, w_004_1855, w_004_1856, w_004_1857, w_004_1858, w_004_1859, w_004_1860, w_004_1861, w_004_1862, w_004_1863, w_004_1864, w_004_1865, w_004_1866, w_004_1867, w_004_1868, w_004_1869, w_004_1870, w_004_1871, w_004_1872, w_004_1873, w_004_1874, w_004_1875, w_004_1876, w_004_1877, w_004_1878, w_004_1879, w_004_1880, w_004_1881, w_004_1882, w_004_1883, w_004_1884, w_004_1885, w_004_1886, w_004_1887, w_004_1888, w_004_1889, w_004_1890, w_004_1891, w_004_1892, w_004_1893, w_004_1894, w_004_1895, w_004_1896, w_004_1897, w_004_1898, w_004_1899, w_004_1900, w_004_1901, w_004_1902, w_004_1903, w_004_1904, w_004_1905, w_004_1906, w_004_1907, w_004_1908, w_004_1909, w_004_1910, w_004_1911, w_004_1912, w_004_1913, w_004_1914, w_004_1915, w_004_1916, w_004_1917, w_004_1918, w_004_1919, w_004_1920, w_004_1921, w_004_1922, w_004_1923, w_004_1924, w_004_1925, w_004_1926, w_004_1927, w_004_1928, w_004_1929, w_004_1930, w_004_1931, w_004_1932, w_004_1933, w_004_1934, w_004_1935, w_004_1936, w_004_1937, w_004_1938, w_004_1939, w_004_1940, w_004_1941, w_004_1942, w_004_1943, w_004_1944, w_004_1945, w_004_1946, w_004_1947, w_004_1948, w_004_1949, w_004_1950, w_004_1951, w_004_1952, w_004_1953, w_004_1954, w_004_1955, w_004_1956, w_004_1957, w_004_1958, w_004_1959, w_004_1960, w_004_1961, w_004_1962, w_004_1963, w_004_1964, w_004_1965, w_004_1966, w_004_1967, w_004_1968, w_004_1969, w_004_1970, w_004_1971, w_004_1972, w_004_1973, w_004_1974, w_004_1975, w_004_1976, w_004_1977, w_004_1978, w_004_1979, w_004_1980, w_004_1981, w_004_1982, w_004_1983, w_004_1984, w_004_1985, w_004_1986, w_004_1987, w_004_1988, w_004_1989, w_004_1990, w_004_1991, w_004_1992, w_004_1993, w_004_1994, w_004_1995, w_004_1996, w_004_1997, w_004_1998, w_004_1999, w_004_2000, w_004_2001, w_004_2002, w_004_2003, w_004_2004, w_004_2005, w_004_2006, w_004_2007, w_004_2008, w_004_2009, w_004_2010, w_004_2011, w_004_2012, w_004_2013, w_004_2014, w_004_2015, w_004_2016, w_004_2017, w_004_2018, w_004_2019, w_004_2020, w_004_2021, w_004_2022, w_004_2023, w_004_2024, w_004_2025, w_004_2026, w_004_2027, w_004_2028, w_004_2029, w_004_2030, w_004_2031, w_004_2032, w_004_2033, w_004_2034, w_004_2035, w_004_2036, w_004_2037, w_004_2038, w_004_2039, w_004_2040, w_004_2041, w_004_2042, w_004_2043, w_004_2044, w_004_2045, w_004_2046, w_004_2047, w_004_2048, w_004_2049, w_004_2050, w_004_2051, w_004_2053, w_004_2054, w_004_2055, w_004_2056, w_004_2057, w_004_2058, w_004_2059, w_004_2060, w_004_2061, w_004_2062, w_004_2063, w_004_2064, w_004_2065, w_004_2066, w_004_2067, w_004_2068, w_004_2069, w_004_2070, w_004_2071, w_004_2072, w_004_2073, w_004_2074, w_004_2075, w_004_2076, w_004_2077, w_004_2078, w_004_2079, w_004_2080, w_004_2081, w_004_2082, w_004_2083, w_004_2084, w_004_2085, w_004_2086, w_004_2087, w_004_2088, w_004_2089, w_004_2090, w_004_2091, w_004_2092, w_004_2093, w_004_2094, w_004_2095, w_004_2096, w_004_2097, w_004_2098, w_004_2099, w_004_2100, w_004_2101, w_004_2102, w_004_2103, w_004_2104, w_004_2105, w_004_2106, w_004_2107, w_004_2108, w_004_2109, w_004_2110, w_004_2111, w_004_2112, w_004_2113, w_004_2114, w_004_2115, w_004_2116, w_004_2117, w_004_2118, w_004_2119, w_004_2120, w_004_2121, w_004_2122, w_004_2123, w_004_2124, w_004_2125, w_004_2126, w_004_2127, w_004_2128, w_004_2129, w_004_2130, w_004_2131, w_004_2132, w_004_2133, w_004_2134, w_004_2135, w_004_2136, w_004_2137, w_004_2138, w_004_2139, w_004_2140, w_004_2141, w_004_2142, w_004_2143, w_004_2144, w_004_2145, w_004_2146, w_004_2147, w_004_2148, w_004_2149, w_004_2150, w_004_2151, w_004_2152, w_004_2153, w_004_2154, w_004_2155, w_004_2156, w_004_2157, w_004_2158, w_004_2159, w_004_2160, w_004_2161, w_004_2162, w_004_2163, w_004_2164, w_004_2165, w_004_2166, w_004_2167, w_004_2168, w_004_2169, w_004_2170, w_004_2171, w_004_2172, w_004_2173, w_004_2174, w_004_2175, w_004_2176, w_004_2177, w_004_2178, w_004_2179, w_004_2180, w_004_2181, w_004_2182, w_004_2183, w_004_2184, w_004_2185, w_004_2186, w_004_2187, w_004_2188, w_004_2189, w_004_2190, w_004_2191, w_004_2192, w_004_2193, w_004_2194, w_004_2195, w_004_2196, w_004_2197, w_004_2198, w_004_2199, w_004_2200, w_004_2201, w_004_2202, w_004_2203, w_004_2204, w_004_2205, w_004_2206, w_004_2207, w_004_2208, w_004_2209, w_004_2210, w_004_2211, w_004_2212, w_004_2213, w_004_2214, w_004_2215, w_004_2216, w_004_2217, w_004_2218, w_004_2219, w_004_2220, w_004_2221, w_004_2222, w_004_2223, w_004_2224, w_004_2225, w_004_2226, w_004_2227, w_004_2228, w_004_2229, w_004_2230, w_004_2231, w_004_2232, w_004_2233, w_004_2234, w_004_2235, w_004_2236, w_004_2237, w_004_2238, w_004_2239, w_004_2240, w_004_2241, w_004_2242, w_004_2243, w_004_2244, w_004_2245, w_004_2246, w_004_2247, w_004_2248, w_004_2249, w_004_2250, w_004_2251, w_004_2252, w_004_2253, w_004_2254, w_004_2255, w_004_2256, w_004_2257, w_004_2258, w_004_2259, w_004_2260, w_004_2261, w_004_2262, w_004_2263, w_004_2264, w_004_2265, w_004_2266, w_004_2267, w_004_2268, w_004_2269, w_004_2270, w_004_2271, w_004_2272, w_004_2273, w_004_2274, w_004_2275, w_004_2276, w_004_2277, w_004_2278, w_004_2279, w_004_2280, w_004_2281, w_004_2282, w_004_2283, w_004_2284, w_004_2285, w_004_2286, w_004_2287, w_004_2288, w_004_2289, w_004_2290, w_004_2291, w_004_2292, w_004_2293, w_004_2294, w_004_2295, w_004_2296, w_004_2297, w_004_2298, w_004_2299, w_004_2300, w_004_2301, w_004_2302, w_004_2303, w_004_2304, w_004_2305, w_004_2306, w_004_2307, w_004_2308, w_004_2309, w_004_2310, w_004_2311, w_004_2312, w_004_2313, w_004_2314, w_004_2315, w_004_2316, w_004_2317, w_004_2318, w_004_2319, w_004_2320, w_004_2321, w_004_2322, w_004_2323, w_004_2324, w_004_2325, w_004_2326, w_004_2327, w_004_2328, w_004_2329, w_004_2330, w_004_2331, w_004_2332, w_004_2333, w_004_2334, w_004_2335, w_004_2336, w_004_2337, w_004_2338, w_004_2339, w_004_2340, w_004_2341, w_004_2342, w_004_2343, w_004_2344, w_004_2345, w_004_2346, w_004_2347, w_004_2348, w_004_2349, w_004_2350, w_004_2351, w_004_2352, w_004_2353, w_004_2354, w_004_2355, w_004_2356, w_004_2357, w_004_2358, w_004_2359, w_004_2360, w_004_2361, w_004_2362, w_004_2363, w_004_2364, w_004_2365, w_004_2366, w_004_2367, w_004_2368, w_004_2369, w_004_2370, w_004_2371, w_004_2372, w_004_2373, w_004_2374, w_004_2375, w_004_2376, w_004_2377, w_004_2378, w_004_2379, w_004_2380, w_004_2381, w_004_2382, w_004_2383, w_004_2384, w_004_2385, w_004_2386, w_004_2387, w_004_2388, w_004_2389, w_004_2390, w_004_2391, w_004_2392, w_004_2393, w_004_2394, w_004_2395, w_004_2396, w_004_2397, w_004_2398, w_004_2399, w_004_2400, w_004_2401, w_004_2402, w_004_2403, w_004_2404, w_004_2405, w_004_2406, w_004_2407, w_004_2408, w_004_2409, w_004_2410, w_004_2411, w_004_2412, w_004_2413, w_004_2414, w_004_2415, w_004_2416, w_004_2417, w_004_2418, w_004_2419, w_004_2420, w_004_2421, w_004_2422, w_004_2423, w_004_2424, w_004_2425, w_004_2426, w_004_2427, w_004_2428, w_004_2429, w_004_2430, w_004_2431, w_004_2432, w_004_2433, w_004_2434, w_004_2435, w_004_2436, w_004_2438, w_004_2439, w_004_2440, w_004_2441, w_004_2442, w_004_2443, w_004_2444, w_004_2445, w_004_2446, w_004_2447, w_004_2448, w_004_2449, w_004_2450, w_004_2451, w_004_2452, w_004_2453, w_004_2454, w_004_2455, w_004_2456, w_004_2457, w_004_2458, w_004_2459, w_004_2460, w_004_2461, w_004_2462, w_004_2463, w_004_2464, w_004_2465, w_004_2466, w_004_2467, w_004_2468, w_004_2469, w_004_2470, w_004_2471, w_004_2472, w_004_2473, w_004_2474, w_004_2475, w_004_2476, w_004_2477, w_004_2478, w_004_2479, w_004_2480, w_004_2481, w_004_2482, w_004_2483, w_004_2484, w_004_2485, w_004_2486, w_004_2487, w_004_2488, w_004_2489, w_004_2490, w_004_2491, w_004_2492, w_004_2493, w_004_2494, w_004_2495, w_004_2496, w_004_2497, w_004_2498, w_004_2499, w_004_2500, w_004_2501, w_004_2502, w_004_2503, w_004_2504, w_004_2505, w_004_2506, w_004_2507, w_004_2508, w_004_2509, w_004_2510, w_004_2511, w_004_2512, w_004_2513, w_004_2514, w_004_2515, w_004_2516, w_004_2517, w_004_2518, w_004_2519, w_004_2520, w_004_2521, w_004_2522, w_004_2523, w_004_2524, w_004_2525, w_004_2526, w_004_2527, w_004_2528, w_004_2529, w_004_2530, w_004_2531, w_004_2532, w_004_2533, w_004_2534, w_004_2535, w_004_2536, w_004_2537, w_004_2538, w_004_2539, w_004_2540, w_004_2541, w_004_2542, w_004_2543, w_004_2544, w_004_2545, w_004_2546, w_004_2547, w_004_2548, w_004_2549, w_004_2550, w_004_2551, w_004_2552, w_004_2553, w_004_2554, w_004_2555, w_004_2556, w_004_2557, w_004_2558, w_004_2559, w_004_2560, w_004_2561, w_004_2562, w_004_2563, w_004_2564, w_004_2565, w_004_2566, w_004_2567, w_004_2568, w_004_2569, w_004_2570, w_004_2571, w_004_2572, w_004_2573, w_004_2574, w_004_2575, w_004_2576, w_004_2577, w_004_2578, w_004_2579, w_004_2580, w_004_2581, w_004_2582, w_004_2583, w_004_2584, w_004_2585, w_004_2586, w_004_2587, w_004_2588, w_004_2589, w_004_2590, w_004_2591, w_004_2592, w_004_2593, w_004_2594, w_004_2595, w_004_2596, w_004_2597, w_004_2598, w_004_2599, w_004_2600, w_004_2601, w_004_2602, w_004_2603, w_004_2604, w_004_2605, w_004_2606, w_004_2607, w_004_2608, w_004_2609, w_004_2610, w_004_2611, w_004_2612, w_004_2613, w_004_2614, w_004_2615, w_004_2616, w_004_2617, w_004_2618, w_004_2619, w_004_2620, w_004_2621, w_004_2622, w_004_2623, w_004_2624, w_004_2625, w_004_2626, w_004_2627, w_004_2628, w_004_2629, w_004_2630, w_004_2631, w_004_2632, w_004_2633, w_004_2634, w_004_2635, w_004_2636, w_004_2637, w_004_2638, w_004_2639, w_004_2640, w_004_2641, w_004_2642, w_004_2643, w_004_2644, w_004_2645, w_004_2646, w_004_2647, w_004_2648, w_004_2649, w_004_2650, w_004_2651, w_004_2652, w_004_2653, w_004_2654, w_004_2655, w_004_2656, w_004_2657, w_004_2658, w_004_2659, w_004_2660, w_004_2661, w_004_2662, w_004_2663, w_004_2664, w_004_2665, w_004_2666, w_004_2667, w_004_2668, w_004_2669, w_004_2670, w_004_2671, w_004_2672, w_004_2673, w_004_2674, w_004_2675, w_004_2676, w_004_2677, w_004_2678, w_004_2679, w_004_2680, w_004_2681, w_004_2682, w_004_2683, w_004_2684, w_004_2685, w_004_2686, w_004_2687, w_004_2688, w_004_2689, w_004_2690, w_004_2691, w_004_2692, w_004_2693, w_004_2694, w_004_2695, w_004_2696, w_004_2697, w_004_2698, w_004_2699, w_004_2700, w_004_2701, w_004_2702, w_004_2703, w_004_2704, w_004_2705, w_004_2706, w_004_2707, w_004_2708, w_004_2709, w_004_2710, w_004_2711, w_004_2712, w_004_2713, w_004_2714, w_004_2715, w_004_2716, w_004_2717, w_004_2718, w_004_2719, w_004_2720, w_004_2721, w_004_2722, w_004_2723, w_004_2724, w_004_2725, w_004_2726, w_004_2727, w_004_2728, w_004_2729, w_004_2730, w_004_2731, w_004_2732, w_004_2733, w_004_2734, w_004_2735, w_004_2736, w_004_2737, w_004_2738, w_004_2739, w_004_2740, w_004_2741, w_004_2742, w_004_2743, w_004_2744, w_004_2745, w_004_2746, w_004_2747, w_004_2748, w_004_2749, w_004_2750, w_004_2751, w_004_2752, w_004_2753, w_004_2754, w_004_2755, w_004_2756, w_004_2757, w_004_2758, w_004_2759, w_004_2760, w_004_2761, w_004_2762, w_004_2763, w_004_2764, w_004_2765, w_004_2766, w_004_2767, w_004_2768, w_004_2769, w_004_2770, w_004_2771, w_004_2772, w_004_2773, w_004_2774, w_004_2775, w_004_2776, w_004_2777, w_004_2778, w_004_2779, w_004_2780, w_004_2781, w_004_2782, w_004_2783, w_004_2784, w_004_2785, w_004_2786, w_004_2787, w_004_2788, w_004_2789, w_004_2790, w_004_2791, w_004_2792, w_004_2793, w_004_2794, w_004_2795, w_004_2796, w_004_2797, w_004_2798, w_004_2799, w_004_2800, w_004_2801, w_004_2802, w_004_2803, w_004_2804, w_004_2805, w_004_2806, w_004_2807, w_004_2808, w_004_2809, w_004_2810, w_004_2811, w_004_2812, w_004_2813, w_004_2814, w_004_2815, w_004_2816, w_004_2817, w_004_2818, w_004_2819, w_004_2820, w_004_2821, w_004_2822, w_004_2823, w_004_2824, w_004_2825, w_004_2826, w_004_2827, w_004_2828, w_004_2829, w_004_2830, w_004_2831, w_004_2832;
  wire w_005_000, w_005_001, w_005_002, w_005_003, w_005_004, w_005_005, w_005_006, w_005_007, w_005_008, w_005_009, w_005_010, w_005_011, w_005_012, w_005_013, w_005_014, w_005_015, w_005_016, w_005_017, w_005_018, w_005_019, w_005_020, w_005_021, w_005_022, w_005_023, w_005_024, w_005_025, w_005_026, w_005_027, w_005_028, w_005_029, w_005_030, w_005_031, w_005_032, w_005_033, w_005_034, w_005_035, w_005_036, w_005_037, w_005_038, w_005_039, w_005_040, w_005_041, w_005_042, w_005_043, w_005_044, w_005_045, w_005_046, w_005_047, w_005_048, w_005_049, w_005_050, w_005_051, w_005_052, w_005_053, w_005_054, w_005_055, w_005_056, w_005_057, w_005_058, w_005_059, w_005_060, w_005_061, w_005_062, w_005_063, w_005_064, w_005_065, w_005_066, w_005_067, w_005_068, w_005_069, w_005_070, w_005_071, w_005_072, w_005_073, w_005_074, w_005_075, w_005_076, w_005_077, w_005_078, w_005_079, w_005_080, w_005_081, w_005_082, w_005_083, w_005_084, w_005_085, w_005_086, w_005_087, w_005_088, w_005_089, w_005_090, w_005_091, w_005_092, w_005_093, w_005_094, w_005_095, w_005_096, w_005_097, w_005_098, w_005_099, w_005_100, w_005_101, w_005_102, w_005_103, w_005_104, w_005_105, w_005_106, w_005_107, w_005_108, w_005_109, w_005_110, w_005_111, w_005_112, w_005_113, w_005_114, w_005_115, w_005_116, w_005_117, w_005_118, w_005_119, w_005_120, w_005_121, w_005_122, w_005_123, w_005_124, w_005_125, w_005_126, w_005_127, w_005_128, w_005_129, w_005_130, w_005_131, w_005_132, w_005_133, w_005_134, w_005_135, w_005_136, w_005_137, w_005_138, w_005_139, w_005_140, w_005_141, w_005_142, w_005_143, w_005_144, w_005_145, w_005_146, w_005_147, w_005_148, w_005_149, w_005_150, w_005_151, w_005_152, w_005_153, w_005_154, w_005_155, w_005_156, w_005_157, w_005_158, w_005_159, w_005_160, w_005_161, w_005_162, w_005_163, w_005_164, w_005_165, w_005_166, w_005_167, w_005_168, w_005_169, w_005_170, w_005_171, w_005_172, w_005_173, w_005_174, w_005_175, w_005_176, w_005_177, w_005_178, w_005_179, w_005_180, w_005_181, w_005_182, w_005_183, w_005_184, w_005_185, w_005_186, w_005_187, w_005_188, w_005_189, w_005_190, w_005_191, w_005_192, w_005_193, w_005_194, w_005_195, w_005_196, w_005_197, w_005_198, w_005_199, w_005_200, w_005_201, w_005_202, w_005_203, w_005_204, w_005_205, w_005_206, w_005_207, w_005_208, w_005_209, w_005_210, w_005_211, w_005_212, w_005_213, w_005_214, w_005_215, w_005_216, w_005_217, w_005_218, w_005_219, w_005_220, w_005_221, w_005_222, w_005_223, w_005_224, w_005_225, w_005_226, w_005_227, w_005_228, w_005_229, w_005_230, w_005_231, w_005_232, w_005_233, w_005_234, w_005_235, w_005_236, w_005_237, w_005_238, w_005_239, w_005_240, w_005_241, w_005_242, w_005_243, w_005_244, w_005_245, w_005_246, w_005_247, w_005_248, w_005_249, w_005_250, w_005_251, w_005_252, w_005_253, w_005_254, w_005_255, w_005_256, w_005_257, w_005_258, w_005_259, w_005_260, w_005_261, w_005_262, w_005_263, w_005_264, w_005_265, w_005_266, w_005_267, w_005_268, w_005_269, w_005_270, w_005_271, w_005_272, w_005_273, w_005_274, w_005_275, w_005_276, w_005_277, w_005_278, w_005_279, w_005_280, w_005_281, w_005_282, w_005_283, w_005_284, w_005_285, w_005_286, w_005_287, w_005_288, w_005_289, w_005_290, w_005_291, w_005_292, w_005_293, w_005_294, w_005_295, w_005_296, w_005_297, w_005_298, w_005_299, w_005_300, w_005_301, w_005_302, w_005_303, w_005_304, w_005_305, w_005_306, w_005_307, w_005_308, w_005_309, w_005_310, w_005_311, w_005_312, w_005_313, w_005_314, w_005_315, w_005_316, w_005_317, w_005_318, w_005_319, w_005_320, w_005_321, w_005_322, w_005_323, w_005_324, w_005_325, w_005_326, w_005_327, w_005_328, w_005_329, w_005_330, w_005_331, w_005_332, w_005_333, w_005_334, w_005_335, w_005_336, w_005_337, w_005_338, w_005_339, w_005_340, w_005_341, w_005_342, w_005_343, w_005_344, w_005_345, w_005_346, w_005_347, w_005_348, w_005_349, w_005_350, w_005_351, w_005_352, w_005_353, w_005_354, w_005_355, w_005_356, w_005_357, w_005_358, w_005_359, w_005_360, w_005_361, w_005_362, w_005_363, w_005_364, w_005_365, w_005_366, w_005_367, w_005_368, w_005_369, w_005_370, w_005_371, w_005_372, w_005_373, w_005_374, w_005_375, w_005_376, w_005_377, w_005_378, w_005_379, w_005_380, w_005_381, w_005_382, w_005_383, w_005_384, w_005_385, w_005_386, w_005_387, w_005_388, w_005_389, w_005_390, w_005_391, w_005_392, w_005_393, w_005_394, w_005_395, w_005_396, w_005_397, w_005_398, w_005_399, w_005_400, w_005_401, w_005_402, w_005_403, w_005_404, w_005_405, w_005_406, w_005_407, w_005_408, w_005_409, w_005_410, w_005_411, w_005_412, w_005_413, w_005_414, w_005_415, w_005_416, w_005_417, w_005_418, w_005_419, w_005_420, w_005_421, w_005_422, w_005_423, w_005_424, w_005_425, w_005_426, w_005_427, w_005_428, w_005_429, w_005_430, w_005_431, w_005_432, w_005_433, w_005_434, w_005_435, w_005_436, w_005_437, w_005_438, w_005_439, w_005_440, w_005_441, w_005_442, w_005_443, w_005_444, w_005_445, w_005_446, w_005_447, w_005_448, w_005_449, w_005_450, w_005_451, w_005_452, w_005_453, w_005_454, w_005_455, w_005_456, w_005_457, w_005_458, w_005_459, w_005_460, w_005_461, w_005_462, w_005_463, w_005_464, w_005_465, w_005_466, w_005_467, w_005_468, w_005_469, w_005_470, w_005_471, w_005_472, w_005_473, w_005_474, w_005_475, w_005_476, w_005_477, w_005_478, w_005_479, w_005_480, w_005_481, w_005_482, w_005_483, w_005_484, w_005_485, w_005_486, w_005_487, w_005_488, w_005_489, w_005_490, w_005_491, w_005_492, w_005_493, w_005_494, w_005_495, w_005_496, w_005_497, w_005_498, w_005_499, w_005_500, w_005_501, w_005_502, w_005_503, w_005_504, w_005_505, w_005_506, w_005_507, w_005_508, w_005_509, w_005_510, w_005_511, w_005_512, w_005_513, w_005_514, w_005_515, w_005_516, w_005_517, w_005_518, w_005_519, w_005_520, w_005_521, w_005_522, w_005_523, w_005_524, w_005_525, w_005_526, w_005_527, w_005_528, w_005_529, w_005_530, w_005_531, w_005_532, w_005_533, w_005_534, w_005_535, w_005_536, w_005_537, w_005_538, w_005_539, w_005_540, w_005_541, w_005_542, w_005_543, w_005_544, w_005_545, w_005_546, w_005_547, w_005_548, w_005_549, w_005_550, w_005_551, w_005_552, w_005_553, w_005_554, w_005_555, w_005_556, w_005_557, w_005_558, w_005_559, w_005_560, w_005_561, w_005_562, w_005_563, w_005_564, w_005_565, w_005_566, w_005_567, w_005_568, w_005_569, w_005_570, w_005_571, w_005_572, w_005_573, w_005_574, w_005_575, w_005_576, w_005_577, w_005_578, w_005_579, w_005_580, w_005_581, w_005_582, w_005_583, w_005_584, w_005_585, w_005_586, w_005_587, w_005_588, w_005_589, w_005_590, w_005_591, w_005_592, w_005_593, w_005_594, w_005_595, w_005_596, w_005_597, w_005_598, w_005_599, w_005_600, w_005_601, w_005_602, w_005_603, w_005_604, w_005_605, w_005_606, w_005_607, w_005_608, w_005_609, w_005_610, w_005_611, w_005_612, w_005_613, w_005_614, w_005_615, w_005_616, w_005_617, w_005_618, w_005_619, w_005_620, w_005_621, w_005_622, w_005_623, w_005_624, w_005_625, w_005_626, w_005_627, w_005_628, w_005_629, w_005_630, w_005_631, w_005_632, w_005_633, w_005_634, w_005_635, w_005_636, w_005_637, w_005_638, w_005_639, w_005_640, w_005_641, w_005_642, w_005_643, w_005_644, w_005_645, w_005_646, w_005_647, w_005_648, w_005_649, w_005_650, w_005_651, w_005_652, w_005_653, w_005_654, w_005_655, w_005_656, w_005_657, w_005_658, w_005_659, w_005_660, w_005_661, w_005_662, w_005_663, w_005_664, w_005_665, w_005_666, w_005_667, w_005_668, w_005_669, w_005_670, w_005_671, w_005_672, w_005_673, w_005_674, w_005_675, w_005_676, w_005_677, w_005_678, w_005_679, w_005_680, w_005_681, w_005_682, w_005_683, w_005_684, w_005_685, w_005_686, w_005_687, w_005_688, w_005_689, w_005_690, w_005_691, w_005_692, w_005_693, w_005_694, w_005_695, w_005_696, w_005_697, w_005_698, w_005_699, w_005_700, w_005_701, w_005_702, w_005_703, w_005_704, w_005_705, w_005_706, w_005_707, w_005_708, w_005_709, w_005_710, w_005_711, w_005_712, w_005_713, w_005_714, w_005_715, w_005_716, w_005_717, w_005_718, w_005_719, w_005_720, w_005_721, w_005_722, w_005_723, w_005_724, w_005_725, w_005_726, w_005_727, w_005_728, w_005_729, w_005_730, w_005_731, w_005_732, w_005_733, w_005_734, w_005_735, w_005_736, w_005_737, w_005_738, w_005_739, w_005_740, w_005_741, w_005_742, w_005_743, w_005_744, w_005_745, w_005_746, w_005_747, w_005_748, w_005_749, w_005_750, w_005_751, w_005_752, w_005_753, w_005_754, w_005_755, w_005_756, w_005_757, w_005_758, w_005_759, w_005_760, w_005_761, w_005_762, w_005_763, w_005_764, w_005_765, w_005_766, w_005_767, w_005_768, w_005_769, w_005_770, w_005_771, w_005_772, w_005_773, w_005_774, w_005_775, w_005_776, w_005_777, w_005_778, w_005_779, w_005_780, w_005_781, w_005_782, w_005_783, w_005_784, w_005_785, w_005_786, w_005_787, w_005_788, w_005_789, w_005_790, w_005_791, w_005_792, w_005_793, w_005_794, w_005_795, w_005_796, w_005_797, w_005_798, w_005_799, w_005_800, w_005_801, w_005_802, w_005_803, w_005_804, w_005_805, w_005_806, w_005_807, w_005_808, w_005_809, w_005_810, w_005_811, w_005_812, w_005_813, w_005_814, w_005_815, w_005_816, w_005_817, w_005_818, w_005_819, w_005_820, w_005_821, w_005_822, w_005_823, w_005_824, w_005_825, w_005_826, w_005_827, w_005_828, w_005_829, w_005_830, w_005_831, w_005_832, w_005_833, w_005_834, w_005_835, w_005_836, w_005_837, w_005_838, w_005_839, w_005_840, w_005_841, w_005_842, w_005_843, w_005_844, w_005_845, w_005_846, w_005_847, w_005_848, w_005_849, w_005_850, w_005_851, w_005_852, w_005_853, w_005_854, w_005_855, w_005_856, w_005_857, w_005_858, w_005_859, w_005_860, w_005_861, w_005_862, w_005_863, w_005_864, w_005_865, w_005_866, w_005_867, w_005_868, w_005_869, w_005_870, w_005_871, w_005_872, w_005_873, w_005_874, w_005_875, w_005_876, w_005_877, w_005_878, w_005_879, w_005_880, w_005_881, w_005_882, w_005_883, w_005_884, w_005_885, w_005_886, w_005_887, w_005_888, w_005_889, w_005_890, w_005_891, w_005_892, w_005_893, w_005_894, w_005_895, w_005_896, w_005_897, w_005_898, w_005_899, w_005_900, w_005_901, w_005_902, w_005_903, w_005_904, w_005_905, w_005_906, w_005_907, w_005_908, w_005_909, w_005_910, w_005_911, w_005_912, w_005_913, w_005_914, w_005_915, w_005_916, w_005_917, w_005_918, w_005_919, w_005_920, w_005_921, w_005_922, w_005_923, w_005_924, w_005_925, w_005_926, w_005_927, w_005_928, w_005_929, w_005_930, w_005_931, w_005_932, w_005_933, w_005_934, w_005_935, w_005_936, w_005_937, w_005_938, w_005_939, w_005_940, w_005_941, w_005_942, w_005_943, w_005_944, w_005_945, w_005_946, w_005_947, w_005_948, w_005_949, w_005_950, w_005_951, w_005_952, w_005_953, w_005_954, w_005_955, w_005_956, w_005_957, w_005_958, w_005_959, w_005_960, w_005_961, w_005_962, w_005_963, w_005_964, w_005_965, w_005_966, w_005_967, w_005_968, w_005_969, w_005_970, w_005_971, w_005_972, w_005_973, w_005_974, w_005_975, w_005_976, w_005_977, w_005_978, w_005_979, w_005_980, w_005_981, w_005_982, w_005_983, w_005_984, w_005_985, w_005_986, w_005_987, w_005_988, w_005_989, w_005_990, w_005_991, w_005_992, w_005_993, w_005_994, w_005_995, w_005_996, w_005_997, w_005_998, w_005_999, w_005_1000, w_005_1001, w_005_1002, w_005_1003, w_005_1004, w_005_1005, w_005_1006, w_005_1007, w_005_1008, w_005_1009, w_005_1010, w_005_1011, w_005_1012, w_005_1013, w_005_1014, w_005_1015, w_005_1016, w_005_1017, w_005_1018, w_005_1019, w_005_1020, w_005_1021, w_005_1022, w_005_1023, w_005_1024, w_005_1025, w_005_1026, w_005_1027, w_005_1028, w_005_1029, w_005_1030, w_005_1031, w_005_1032, w_005_1033, w_005_1034, w_005_1035, w_005_1036, w_005_1037, w_005_1038, w_005_1039, w_005_1040, w_005_1041, w_005_1042, w_005_1043, w_005_1044, w_005_1045, w_005_1046, w_005_1047, w_005_1048, w_005_1049, w_005_1050, w_005_1051, w_005_1052, w_005_1053, w_005_1054, w_005_1055, w_005_1056, w_005_1057, w_005_1058, w_005_1059, w_005_1060, w_005_1061, w_005_1062, w_005_1063, w_005_1064, w_005_1065, w_005_1066, w_005_1067, w_005_1068, w_005_1069, w_005_1070, w_005_1071, w_005_1072, w_005_1073, w_005_1074, w_005_1075, w_005_1076, w_005_1077, w_005_1078, w_005_1079, w_005_1080, w_005_1081, w_005_1082, w_005_1083, w_005_1084, w_005_1085, w_005_1086, w_005_1087, w_005_1088, w_005_1089, w_005_1090, w_005_1091, w_005_1092, w_005_1093, w_005_1094, w_005_1095, w_005_1096, w_005_1097, w_005_1098, w_005_1099, w_005_1100, w_005_1101, w_005_1102, w_005_1103, w_005_1104, w_005_1105, w_005_1106, w_005_1107, w_005_1108, w_005_1109, w_005_1110, w_005_1111, w_005_1112, w_005_1113, w_005_1114, w_005_1115, w_005_1116, w_005_1117, w_005_1118, w_005_1119, w_005_1120, w_005_1121, w_005_1122, w_005_1123, w_005_1124, w_005_1125, w_005_1126, w_005_1127, w_005_1128, w_005_1129, w_005_1130, w_005_1131, w_005_1132, w_005_1133, w_005_1134, w_005_1135, w_005_1136, w_005_1137, w_005_1138, w_005_1139, w_005_1140, w_005_1141, w_005_1142, w_005_1143, w_005_1144, w_005_1145, w_005_1146, w_005_1147, w_005_1148, w_005_1149, w_005_1150, w_005_1151, w_005_1152, w_005_1153, w_005_1154, w_005_1155, w_005_1156, w_005_1157, w_005_1158, w_005_1159, w_005_1160, w_005_1161, w_005_1162, w_005_1163, w_005_1164, w_005_1165, w_005_1166, w_005_1167, w_005_1168, w_005_1169, w_005_1170, w_005_1171, w_005_1172, w_005_1173, w_005_1174, w_005_1175, w_005_1176, w_005_1177, w_005_1178, w_005_1179, w_005_1180, w_005_1181, w_005_1182, w_005_1183, w_005_1184, w_005_1185, w_005_1186, w_005_1187, w_005_1188, w_005_1189, w_005_1190, w_005_1191, w_005_1192, w_005_1193, w_005_1194, w_005_1195, w_005_1196, w_005_1197, w_005_1198, w_005_1199, w_005_1200, w_005_1201, w_005_1202, w_005_1203, w_005_1204, w_005_1205, w_005_1206, w_005_1207, w_005_1208, w_005_1209, w_005_1210, w_005_1211, w_005_1212, w_005_1213, w_005_1214, w_005_1215, w_005_1216, w_005_1217, w_005_1218, w_005_1219, w_005_1220, w_005_1221, w_005_1222, w_005_1223, w_005_1224, w_005_1225, w_005_1226, w_005_1227, w_005_1228, w_005_1229, w_005_1230, w_005_1231, w_005_1232, w_005_1233, w_005_1234, w_005_1235, w_005_1236, w_005_1237, w_005_1238, w_005_1239, w_005_1240, w_005_1241, w_005_1242, w_005_1243, w_005_1244, w_005_1245, w_005_1246, w_005_1247, w_005_1248, w_005_1249, w_005_1250, w_005_1251, w_005_1252, w_005_1253, w_005_1254, w_005_1255, w_005_1256, w_005_1257, w_005_1258, w_005_1259, w_005_1260, w_005_1261, w_005_1262, w_005_1263, w_005_1264, w_005_1265, w_005_1266, w_005_1267, w_005_1268, w_005_1269, w_005_1270, w_005_1271, w_005_1272, w_005_1273, w_005_1274, w_005_1275, w_005_1276, w_005_1277, w_005_1278, w_005_1279, w_005_1280, w_005_1281, w_005_1282, w_005_1283, w_005_1284, w_005_1285, w_005_1286, w_005_1287, w_005_1288, w_005_1289, w_005_1290, w_005_1291, w_005_1292, w_005_1293, w_005_1294, w_005_1295, w_005_1296, w_005_1297, w_005_1298, w_005_1299, w_005_1300, w_005_1301, w_005_1302, w_005_1303, w_005_1304, w_005_1305, w_005_1306, w_005_1307, w_005_1308, w_005_1309, w_005_1310, w_005_1311, w_005_1312, w_005_1313, w_005_1314, w_005_1315, w_005_1316, w_005_1317, w_005_1318, w_005_1319, w_005_1320, w_005_1321, w_005_1322, w_005_1323, w_005_1324, w_005_1325, w_005_1326, w_005_1327, w_005_1328, w_005_1329, w_005_1330, w_005_1331, w_005_1332, w_005_1333, w_005_1334, w_005_1335, w_005_1336, w_005_1337, w_005_1338, w_005_1339, w_005_1340, w_005_1341, w_005_1342, w_005_1343, w_005_1344, w_005_1345, w_005_1346, w_005_1347, w_005_1348, w_005_1349, w_005_1350, w_005_1351, w_005_1352, w_005_1353, w_005_1354, w_005_1355, w_005_1356, w_005_1357, w_005_1358, w_005_1359, w_005_1360, w_005_1361, w_005_1362, w_005_1363, w_005_1364, w_005_1365, w_005_1366, w_005_1367, w_005_1368, w_005_1369, w_005_1370, w_005_1371, w_005_1372, w_005_1373, w_005_1374, w_005_1375, w_005_1376, w_005_1377, w_005_1378, w_005_1379, w_005_1380, w_005_1381, w_005_1382, w_005_1383, w_005_1384, w_005_1385, w_005_1386, w_005_1387, w_005_1388, w_005_1389, w_005_1390, w_005_1391, w_005_1392, w_005_1393, w_005_1394, w_005_1395, w_005_1396, w_005_1397, w_005_1398, w_005_1399, w_005_1400, w_005_1401, w_005_1402, w_005_1403, w_005_1404, w_005_1405, w_005_1406, w_005_1407, w_005_1408, w_005_1409, w_005_1410, w_005_1411, w_005_1412, w_005_1413, w_005_1414, w_005_1415, w_005_1416, w_005_1417, w_005_1418, w_005_1419, w_005_1420, w_005_1421, w_005_1422, w_005_1423, w_005_1424, w_005_1425, w_005_1426, w_005_1427, w_005_1428, w_005_1429, w_005_1430, w_005_1431, w_005_1432, w_005_1433, w_005_1434, w_005_1435, w_005_1436, w_005_1437, w_005_1438, w_005_1439, w_005_1440, w_005_1441, w_005_1442, w_005_1443, w_005_1444, w_005_1445, w_005_1446, w_005_1447, w_005_1448, w_005_1449, w_005_1450, w_005_1451, w_005_1452, w_005_1453, w_005_1454, w_005_1455, w_005_1456, w_005_1457, w_005_1458, w_005_1459, w_005_1460, w_005_1461, w_005_1462, w_005_1463, w_005_1464, w_005_1465, w_005_1466, w_005_1467, w_005_1468, w_005_1469, w_005_1470, w_005_1471, w_005_1472, w_005_1473, w_005_1474, w_005_1475, w_005_1476, w_005_1477, w_005_1478, w_005_1479, w_005_1480, w_005_1481, w_005_1482, w_005_1483, w_005_1484, w_005_1485, w_005_1486, w_005_1487, w_005_1488, w_005_1489, w_005_1490, w_005_1491, w_005_1492, w_005_1493, w_005_1494, w_005_1495, w_005_1496, w_005_1497, w_005_1498, w_005_1499, w_005_1500, w_005_1501, w_005_1502, w_005_1503, w_005_1504, w_005_1505, w_005_1506, w_005_1507, w_005_1508, w_005_1509, w_005_1510, w_005_1511, w_005_1512, w_005_1513, w_005_1514, w_005_1515, w_005_1516, w_005_1517, w_005_1518, w_005_1519, w_005_1520, w_005_1521, w_005_1522, w_005_1523, w_005_1524, w_005_1525, w_005_1526, w_005_1527, w_005_1528, w_005_1529, w_005_1530, w_005_1531, w_005_1532, w_005_1533, w_005_1534, w_005_1535, w_005_1536, w_005_1537, w_005_1538, w_005_1539, w_005_1540, w_005_1541, w_005_1542, w_005_1543, w_005_1544, w_005_1545, w_005_1546, w_005_1547, w_005_1548, w_005_1549, w_005_1550, w_005_1551, w_005_1552, w_005_1553, w_005_1554, w_005_1555, w_005_1556, w_005_1557, w_005_1558, w_005_1559, w_005_1560, w_005_1561, w_005_1562, w_005_1563, w_005_1564, w_005_1565, w_005_1566, w_005_1567, w_005_1568, w_005_1569, w_005_1570, w_005_1571, w_005_1572, w_005_1573, w_005_1574, w_005_1575, w_005_1576, w_005_1577, w_005_1578, w_005_1579, w_005_1580, w_005_1581, w_005_1582, w_005_1583, w_005_1584, w_005_1585, w_005_1586, w_005_1587;
  wire w_006_000, w_006_001, w_006_002, w_006_003, w_006_004, w_006_005, w_006_006, w_006_007, w_006_008, w_006_009, w_006_010, w_006_011, w_006_012, w_006_013, w_006_014, w_006_015, w_006_016, w_006_017, w_006_018, w_006_019, w_006_020, w_006_021, w_006_022, w_006_023, w_006_024, w_006_025, w_006_026, w_006_027, w_006_028, w_006_029, w_006_030, w_006_031, w_006_032, w_006_033, w_006_034, w_006_035, w_006_036, w_006_037, w_006_038, w_006_039, w_006_040, w_006_041, w_006_042, w_006_043, w_006_044, w_006_045, w_006_046, w_006_047, w_006_048, w_006_049, w_006_050, w_006_051, w_006_052, w_006_053, w_006_054, w_006_055, w_006_056, w_006_057, w_006_058, w_006_059, w_006_060, w_006_061, w_006_062, w_006_063, w_006_064, w_006_065, w_006_066, w_006_067, w_006_068, w_006_069, w_006_070, w_006_071, w_006_072, w_006_073, w_006_074, w_006_075, w_006_076, w_006_077, w_006_078, w_006_079, w_006_080, w_006_081, w_006_082, w_006_083, w_006_084, w_006_085, w_006_086, w_006_087, w_006_088, w_006_089, w_006_090, w_006_091, w_006_092, w_006_093, w_006_094, w_006_095, w_006_096, w_006_097, w_006_098, w_006_099, w_006_100, w_006_101, w_006_102, w_006_103, w_006_104, w_006_105, w_006_106, w_006_107, w_006_108, w_006_109, w_006_110, w_006_111, w_006_112, w_006_113, w_006_114, w_006_115, w_006_116, w_006_117, w_006_118, w_006_119, w_006_120, w_006_121, w_006_122, w_006_123, w_006_124, w_006_125, w_006_126, w_006_127, w_006_128, w_006_129, w_006_130, w_006_131, w_006_132, w_006_133, w_006_134, w_006_135, w_006_136, w_006_137, w_006_138, w_006_139, w_006_140, w_006_141, w_006_142, w_006_143, w_006_144, w_006_145, w_006_146, w_006_147, w_006_148, w_006_149, w_006_150, w_006_151, w_006_152, w_006_153, w_006_154, w_006_155, w_006_156, w_006_157, w_006_158, w_006_159, w_006_160, w_006_161, w_006_162, w_006_163, w_006_164, w_006_165, w_006_166, w_006_167, w_006_168, w_006_169, w_006_170, w_006_171, w_006_172, w_006_173, w_006_174, w_006_175, w_006_176, w_006_177, w_006_178, w_006_179, w_006_180, w_006_181, w_006_182, w_006_183, w_006_184, w_006_185, w_006_186, w_006_187, w_006_188, w_006_189, w_006_190, w_006_191, w_006_192, w_006_193, w_006_194, w_006_195, w_006_196, w_006_197, w_006_198, w_006_199, w_006_200, w_006_201, w_006_202, w_006_203, w_006_204, w_006_205, w_006_206, w_006_207, w_006_208, w_006_209, w_006_210, w_006_211, w_006_212, w_006_213, w_006_214, w_006_215, w_006_216, w_006_217, w_006_218, w_006_219, w_006_220, w_006_221, w_006_222, w_006_223, w_006_224, w_006_225, w_006_226, w_006_227, w_006_228, w_006_229, w_006_230, w_006_231, w_006_232, w_006_233, w_006_234, w_006_235, w_006_236, w_006_237, w_006_238, w_006_239, w_006_240, w_006_241, w_006_242, w_006_243, w_006_244, w_006_245, w_006_246, w_006_247, w_006_248, w_006_249, w_006_250, w_006_251, w_006_252, w_006_253, w_006_254, w_006_255, w_006_256, w_006_257, w_006_258, w_006_259, w_006_260, w_006_261, w_006_262, w_006_263, w_006_264, w_006_265, w_006_266, w_006_267, w_006_268, w_006_269, w_006_270, w_006_271, w_006_272, w_006_273, w_006_274, w_006_275, w_006_276, w_006_277, w_006_278, w_006_279, w_006_280, w_006_281, w_006_282, w_006_283, w_006_284, w_006_285, w_006_286, w_006_287, w_006_288, w_006_289, w_006_290, w_006_291, w_006_292, w_006_293, w_006_294, w_006_295, w_006_296, w_006_297, w_006_298, w_006_299, w_006_300, w_006_301, w_006_302, w_006_303, w_006_304, w_006_305, w_006_306, w_006_307, w_006_308, w_006_309, w_006_310, w_006_312, w_006_313, w_006_314, w_006_315, w_006_316, w_006_317, w_006_318, w_006_319, w_006_320, w_006_321, w_006_322, w_006_323, w_006_324, w_006_325, w_006_326, w_006_327, w_006_328, w_006_329, w_006_330, w_006_331, w_006_332, w_006_333, w_006_334, w_006_335, w_006_336, w_006_337, w_006_338, w_006_339, w_006_340, w_006_341, w_006_342, w_006_343, w_006_344, w_006_345, w_006_346, w_006_347, w_006_348, w_006_349, w_006_350, w_006_351, w_006_352, w_006_353, w_006_354, w_006_355, w_006_356, w_006_357, w_006_358, w_006_359, w_006_360, w_006_361, w_006_362, w_006_363, w_006_364, w_006_365, w_006_366, w_006_367, w_006_368, w_006_369, w_006_370, w_006_371, w_006_372, w_006_373, w_006_374, w_006_375, w_006_376, w_006_377, w_006_378, w_006_379, w_006_380, w_006_381, w_006_382, w_006_383, w_006_384, w_006_385, w_006_386, w_006_387, w_006_388, w_006_389, w_006_390, w_006_391, w_006_392, w_006_393, w_006_394, w_006_395, w_006_396, w_006_397, w_006_398, w_006_399, w_006_400, w_006_401, w_006_402, w_006_403, w_006_404, w_006_405, w_006_406, w_006_407, w_006_408, w_006_409, w_006_410, w_006_411, w_006_412, w_006_413, w_006_414, w_006_415, w_006_416, w_006_417, w_006_418, w_006_419, w_006_420, w_006_421, w_006_422, w_006_423, w_006_424, w_006_425, w_006_426, w_006_427, w_006_428, w_006_429, w_006_430, w_006_431, w_006_432, w_006_433, w_006_434, w_006_435, w_006_436, w_006_437, w_006_438, w_006_439, w_006_440, w_006_441, w_006_442, w_006_443, w_006_444, w_006_445, w_006_446, w_006_447, w_006_448, w_006_449, w_006_450, w_006_451, w_006_452, w_006_453, w_006_454, w_006_455, w_006_456, w_006_457, w_006_458, w_006_459, w_006_460, w_006_461, w_006_462, w_006_463, w_006_464, w_006_465, w_006_466, w_006_467, w_006_468, w_006_469, w_006_470, w_006_471, w_006_472, w_006_473, w_006_474, w_006_475, w_006_476, w_006_477, w_006_478, w_006_480, w_006_481, w_006_482, w_006_483, w_006_484, w_006_485, w_006_486, w_006_487, w_006_488, w_006_489, w_006_490, w_006_491, w_006_492, w_006_493, w_006_494, w_006_495, w_006_496, w_006_497, w_006_498, w_006_499, w_006_500, w_006_501, w_006_502, w_006_503, w_006_504, w_006_505, w_006_506, w_006_507, w_006_508, w_006_509, w_006_510, w_006_511, w_006_512, w_006_513, w_006_514, w_006_515, w_006_516, w_006_517, w_006_518, w_006_519, w_006_520, w_006_521, w_006_522, w_006_523, w_006_524, w_006_525, w_006_526, w_006_527, w_006_528, w_006_529, w_006_530, w_006_531, w_006_532, w_006_533, w_006_534, w_006_535, w_006_536, w_006_537, w_006_538, w_006_539, w_006_540, w_006_541, w_006_542, w_006_543, w_006_544, w_006_545, w_006_546, w_006_547, w_006_548, w_006_549, w_006_550, w_006_551, w_006_552, w_006_553, w_006_554, w_006_555, w_006_556, w_006_557, w_006_558, w_006_559, w_006_560, w_006_561, w_006_562, w_006_563, w_006_564, w_006_565, w_006_566, w_006_567, w_006_568, w_006_569, w_006_570, w_006_571, w_006_572, w_006_573, w_006_574, w_006_575, w_006_576, w_006_577, w_006_578, w_006_579, w_006_580, w_006_581, w_006_582, w_006_583, w_006_584, w_006_585, w_006_586, w_006_587, w_006_588, w_006_589, w_006_590, w_006_591, w_006_592, w_006_593, w_006_594, w_006_595, w_006_596, w_006_597, w_006_598, w_006_599, w_006_600, w_006_601, w_006_602, w_006_603, w_006_604, w_006_605, w_006_606, w_006_607, w_006_608, w_006_609, w_006_610, w_006_611, w_006_612, w_006_613, w_006_614, w_006_615, w_006_616, w_006_617, w_006_618, w_006_619, w_006_620, w_006_621, w_006_622, w_006_623, w_006_624, w_006_625, w_006_626, w_006_627, w_006_628, w_006_629, w_006_630, w_006_631, w_006_632, w_006_633, w_006_634, w_006_635, w_006_636, w_006_637, w_006_638, w_006_639, w_006_640, w_006_641, w_006_642, w_006_643, w_006_644, w_006_645, w_006_646, w_006_647, w_006_648, w_006_649, w_006_650, w_006_651, w_006_652, w_006_653, w_006_654, w_006_655, w_006_656, w_006_657, w_006_658, w_006_659, w_006_660, w_006_661, w_006_662, w_006_663, w_006_664, w_006_665, w_006_666, w_006_667, w_006_668, w_006_669, w_006_670, w_006_671, w_006_672, w_006_673, w_006_674, w_006_675, w_006_676, w_006_677, w_006_678, w_006_679, w_006_680, w_006_681, w_006_682, w_006_683, w_006_684, w_006_685, w_006_686, w_006_687, w_006_688, w_006_689, w_006_690, w_006_691, w_006_692, w_006_693, w_006_694, w_006_695, w_006_696, w_006_697, w_006_698, w_006_699, w_006_700, w_006_701, w_006_702, w_006_703, w_006_704, w_006_705, w_006_706, w_006_707, w_006_708, w_006_709, w_006_710, w_006_711, w_006_712, w_006_713, w_006_714, w_006_715, w_006_716, w_006_717, w_006_718, w_006_719, w_006_720, w_006_721, w_006_722, w_006_723, w_006_724, w_006_725, w_006_726, w_006_727, w_006_728, w_006_729, w_006_730, w_006_731, w_006_732, w_006_733, w_006_734, w_006_735, w_006_736, w_006_737, w_006_738, w_006_739, w_006_740, w_006_741, w_006_742, w_006_743, w_006_744, w_006_745, w_006_746, w_006_747, w_006_748, w_006_749, w_006_750, w_006_751, w_006_752, w_006_753, w_006_754, w_006_755, w_006_756, w_006_757, w_006_758, w_006_759, w_006_760, w_006_761, w_006_762, w_006_763, w_006_764, w_006_765, w_006_766, w_006_767, w_006_768, w_006_769, w_006_770, w_006_771, w_006_772, w_006_773, w_006_774, w_006_775, w_006_776, w_006_777, w_006_778, w_006_779, w_006_780, w_006_781, w_006_782, w_006_783, w_006_784, w_006_785, w_006_786, w_006_787, w_006_788, w_006_789, w_006_790, w_006_791, w_006_792, w_006_793, w_006_794, w_006_795, w_006_796, w_006_797, w_006_798, w_006_799, w_006_800, w_006_801, w_006_802, w_006_803, w_006_804, w_006_805, w_006_806, w_006_807, w_006_808, w_006_809, w_006_810, w_006_811, w_006_812, w_006_813, w_006_814, w_006_815, w_006_816, w_006_817, w_006_818, w_006_819, w_006_820, w_006_821, w_006_822, w_006_823, w_006_824, w_006_825, w_006_826, w_006_827, w_006_828, w_006_829, w_006_830, w_006_831, w_006_832, w_006_833, w_006_834, w_006_835, w_006_836, w_006_837, w_006_838, w_006_839, w_006_840, w_006_841, w_006_842, w_006_843, w_006_844, w_006_845, w_006_846, w_006_847, w_006_848, w_006_849, w_006_850, w_006_851, w_006_852, w_006_853, w_006_854, w_006_855, w_006_856, w_006_857, w_006_858, w_006_859, w_006_860, w_006_861, w_006_862, w_006_863, w_006_864, w_006_865, w_006_866, w_006_867, w_006_868, w_006_869, w_006_870, w_006_871, w_006_872, w_006_873, w_006_874, w_006_875, w_006_876, w_006_877, w_006_878, w_006_879, w_006_880, w_006_881, w_006_882, w_006_883, w_006_884, w_006_885, w_006_886, w_006_888, w_006_889, w_006_890, w_006_891, w_006_892, w_006_893, w_006_894, w_006_895, w_006_896, w_006_897, w_006_898, w_006_899, w_006_900, w_006_901, w_006_902, w_006_903, w_006_904, w_006_905, w_006_906, w_006_907, w_006_908, w_006_909, w_006_910, w_006_911, w_006_912, w_006_913, w_006_914, w_006_915, w_006_916, w_006_917, w_006_918, w_006_919, w_006_920, w_006_921, w_006_922, w_006_923, w_006_924, w_006_925, w_006_926, w_006_927, w_006_928, w_006_929, w_006_930, w_006_931, w_006_932, w_006_934, w_006_935, w_006_936, w_006_937, w_006_938, w_006_939, w_006_940, w_006_941, w_006_942, w_006_943, w_006_944, w_006_945, w_006_946, w_006_947, w_006_948, w_006_949, w_006_950, w_006_951, w_006_952, w_006_953, w_006_954, w_006_955, w_006_956, w_006_957, w_006_958, w_006_959, w_006_960, w_006_961, w_006_962, w_006_963, w_006_964, w_006_965, w_006_966, w_006_967, w_006_968, w_006_969, w_006_970, w_006_971, w_006_972, w_006_973, w_006_974, w_006_975, w_006_976, w_006_977, w_006_978, w_006_979, w_006_980, w_006_981, w_006_982, w_006_983, w_006_984, w_006_985, w_006_986, w_006_987, w_006_988, w_006_989, w_006_990, w_006_991, w_006_992, w_006_993, w_006_994, w_006_995, w_006_996, w_006_997, w_006_998, w_006_999, w_006_1000, w_006_1001, w_006_1002, w_006_1003, w_006_1004, w_006_1005, w_006_1006, w_006_1007, w_006_1008, w_006_1009, w_006_1010, w_006_1011, w_006_1012, w_006_1013, w_006_1014, w_006_1015, w_006_1016, w_006_1017, w_006_1018, w_006_1019, w_006_1020, w_006_1021, w_006_1022, w_006_1023, w_006_1024, w_006_1025, w_006_1026, w_006_1027, w_006_1028, w_006_1029, w_006_1030, w_006_1031, w_006_1032, w_006_1033, w_006_1034, w_006_1035, w_006_1036, w_006_1037, w_006_1038, w_006_1039, w_006_1040, w_006_1041, w_006_1042, w_006_1043, w_006_1044, w_006_1045, w_006_1046, w_006_1047, w_006_1048, w_006_1049, w_006_1050, w_006_1051, w_006_1052, w_006_1053, w_006_1054, w_006_1055, w_006_1056, w_006_1057, w_006_1058, w_006_1059, w_006_1060, w_006_1061, w_006_1062, w_006_1063, w_006_1064, w_006_1065, w_006_1066, w_006_1067, w_006_1068, w_006_1069, w_006_1070, w_006_1071, w_006_1072, w_006_1073, w_006_1074, w_006_1075, w_006_1076, w_006_1077, w_006_1078, w_006_1079, w_006_1080, w_006_1081, w_006_1082, w_006_1083, w_006_1084, w_006_1085, w_006_1086, w_006_1087, w_006_1088, w_006_1089, w_006_1090, w_006_1091, w_006_1092, w_006_1093, w_006_1094, w_006_1095, w_006_1096, w_006_1097, w_006_1098, w_006_1099, w_006_1100, w_006_1101, w_006_1102, w_006_1103, w_006_1104, w_006_1105, w_006_1106, w_006_1107, w_006_1108, w_006_1109, w_006_1110, w_006_1111, w_006_1112, w_006_1113, w_006_1114, w_006_1115, w_006_1116, w_006_1117, w_006_1118, w_006_1119, w_006_1120, w_006_1121, w_006_1122, w_006_1123, w_006_1124, w_006_1125, w_006_1126, w_006_1127, w_006_1128, w_006_1129, w_006_1130, w_006_1131, w_006_1132, w_006_1133, w_006_1134, w_006_1135, w_006_1136, w_006_1137, w_006_1138, w_006_1139, w_006_1140, w_006_1141, w_006_1142, w_006_1143, w_006_1144, w_006_1145, w_006_1146, w_006_1147, w_006_1148, w_006_1149, w_006_1150, w_006_1151, w_006_1152, w_006_1153, w_006_1154, w_006_1155, w_006_1156, w_006_1157, w_006_1158, w_006_1159, w_006_1160, w_006_1161, w_006_1162, w_006_1163, w_006_1164, w_006_1165, w_006_1166, w_006_1167, w_006_1168, w_006_1169, w_006_1170, w_006_1171, w_006_1172, w_006_1173, w_006_1174, w_006_1175, w_006_1176, w_006_1177, w_006_1178, w_006_1179, w_006_1180, w_006_1181, w_006_1182, w_006_1183, w_006_1184, w_006_1185, w_006_1186, w_006_1187, w_006_1188, w_006_1189, w_006_1190, w_006_1191, w_006_1192, w_006_1193, w_006_1194, w_006_1195, w_006_1196, w_006_1197, w_006_1198, w_006_1199, w_006_1200, w_006_1201, w_006_1202, w_006_1203, w_006_1204, w_006_1205, w_006_1206, w_006_1207, w_006_1208, w_006_1209, w_006_1210, w_006_1211, w_006_1212, w_006_1213, w_006_1214, w_006_1215, w_006_1216, w_006_1217, w_006_1218, w_006_1219, w_006_1221, w_006_1222, w_006_1223, w_006_1224, w_006_1225, w_006_1226, w_006_1227, w_006_1228, w_006_1229, w_006_1230, w_006_1231, w_006_1232, w_006_1233, w_006_1234, w_006_1235, w_006_1236, w_006_1237, w_006_1238, w_006_1239, w_006_1240, w_006_1241, w_006_1242, w_006_1243, w_006_1244, w_006_1245, w_006_1246, w_006_1247, w_006_1248, w_006_1249, w_006_1250, w_006_1251, w_006_1252, w_006_1253, w_006_1254, w_006_1255, w_006_1256, w_006_1257, w_006_1258, w_006_1259, w_006_1260, w_006_1261, w_006_1262, w_006_1263, w_006_1264, w_006_1265, w_006_1266, w_006_1267, w_006_1268, w_006_1269, w_006_1270, w_006_1271, w_006_1272, w_006_1273, w_006_1274, w_006_1275, w_006_1276, w_006_1277, w_006_1278, w_006_1279, w_006_1280, w_006_1281, w_006_1282, w_006_1283, w_006_1284, w_006_1285, w_006_1286, w_006_1287, w_006_1288, w_006_1289, w_006_1290, w_006_1291, w_006_1292, w_006_1293, w_006_1294, w_006_1295, w_006_1296, w_006_1297, w_006_1298, w_006_1299, w_006_1300, w_006_1301, w_006_1302, w_006_1303, w_006_1304, w_006_1305, w_006_1306, w_006_1307, w_006_1308, w_006_1309, w_006_1310, w_006_1311, w_006_1312, w_006_1313, w_006_1314, w_006_1315, w_006_1316, w_006_1317, w_006_1318, w_006_1319, w_006_1320, w_006_1321, w_006_1322, w_006_1323, w_006_1324, w_006_1325, w_006_1326, w_006_1327, w_006_1328, w_006_1329, w_006_1330, w_006_1331, w_006_1332, w_006_1333, w_006_1334, w_006_1335, w_006_1336, w_006_1337, w_006_1338, w_006_1339, w_006_1340, w_006_1341, w_006_1342, w_006_1343, w_006_1344, w_006_1345, w_006_1346, w_006_1347, w_006_1348, w_006_1349, w_006_1350, w_006_1351, w_006_1352, w_006_1353, w_006_1354, w_006_1355, w_006_1356, w_006_1357, w_006_1358, w_006_1359, w_006_1360, w_006_1361, w_006_1362, w_006_1363, w_006_1364, w_006_1365, w_006_1366, w_006_1367, w_006_1368, w_006_1369, w_006_1370, w_006_1371, w_006_1372, w_006_1373, w_006_1374, w_006_1375, w_006_1376, w_006_1377, w_006_1378, w_006_1379, w_006_1380, w_006_1382, w_006_1383, w_006_1384, w_006_1385, w_006_1386, w_006_1387, w_006_1388, w_006_1389, w_006_1390, w_006_1391, w_006_1392, w_006_1393, w_006_1394, w_006_1395, w_006_1396, w_006_1397, w_006_1398, w_006_1399, w_006_1400, w_006_1401, w_006_1402, w_006_1403, w_006_1404, w_006_1405, w_006_1406, w_006_1407, w_006_1408, w_006_1409, w_006_1410, w_006_1411, w_006_1412, w_006_1413, w_006_1414, w_006_1415, w_006_1416, w_006_1417, w_006_1418, w_006_1419, w_006_1420, w_006_1421, w_006_1422, w_006_1423, w_006_1424, w_006_1425, w_006_1426, w_006_1427, w_006_1428, w_006_1429, w_006_1430, w_006_1431, w_006_1432, w_006_1433, w_006_1434, w_006_1435, w_006_1436, w_006_1437, w_006_1438, w_006_1439, w_006_1440, w_006_1441, w_006_1442, w_006_1443, w_006_1444, w_006_1445, w_006_1446, w_006_1447, w_006_1448, w_006_1449, w_006_1450, w_006_1451, w_006_1452, w_006_1453, w_006_1454, w_006_1455, w_006_1456, w_006_1457, w_006_1458, w_006_1459, w_006_1460, w_006_1461, w_006_1462, w_006_1463, w_006_1464, w_006_1465, w_006_1466, w_006_1467, w_006_1468, w_006_1469, w_006_1470, w_006_1471, w_006_1472, w_006_1473, w_006_1474, w_006_1475, w_006_1476, w_006_1477, w_006_1478, w_006_1479, w_006_1480, w_006_1481, w_006_1482, w_006_1483, w_006_1484, w_006_1485, w_006_1486, w_006_1487, w_006_1488, w_006_1489, w_006_1490, w_006_1491, w_006_1492, w_006_1493, w_006_1494, w_006_1495, w_006_1496, w_006_1497, w_006_1498, w_006_1499, w_006_1500, w_006_1501, w_006_1502, w_006_1503, w_006_1504, w_006_1505, w_006_1506, w_006_1507, w_006_1508, w_006_1509, w_006_1510, w_006_1511, w_006_1512, w_006_1513, w_006_1514, w_006_1515, w_006_1516, w_006_1517, w_006_1519, w_006_1520, w_006_1521, w_006_1522, w_006_1523, w_006_1524, w_006_1525, w_006_1526, w_006_1527, w_006_1528, w_006_1529, w_006_1530, w_006_1531, w_006_1532, w_006_1533, w_006_1534, w_006_1535, w_006_1536, w_006_1537, w_006_1538, w_006_1539, w_006_1540, w_006_1541, w_006_1542, w_006_1543, w_006_1544, w_006_1545, w_006_1546, w_006_1547, w_006_1548, w_006_1549, w_006_1550, w_006_1551, w_006_1552, w_006_1553, w_006_1554, w_006_1555, w_006_1556, w_006_1557, w_006_1558, w_006_1559, w_006_1560, w_006_1561, w_006_1562, w_006_1563, w_006_1564, w_006_1565, w_006_1566, w_006_1567, w_006_1569, w_006_1570, w_006_1571, w_006_1572, w_006_1573, w_006_1574, w_006_1575, w_006_1576, w_006_1577, w_006_1578, w_006_1579, w_006_1580, w_006_1581, w_006_1582, w_006_1583, w_006_1584, w_006_1585, w_006_1586, w_006_1587, w_006_1588, w_006_1589, w_006_1590, w_006_1591, w_006_1592, w_006_1593, w_006_1594, w_006_1595, w_006_1596, w_006_1597, w_006_1598, w_006_1599, w_006_1600, w_006_1601, w_006_1602, w_006_1603, w_006_1604, w_006_1605, w_006_1606, w_006_1607, w_006_1608, w_006_1609, w_006_1610, w_006_1611, w_006_1612, w_006_1613, w_006_1614, w_006_1615, w_006_1616, w_006_1617, w_006_1618, w_006_1619, w_006_1620, w_006_1621, w_006_1622, w_006_1623, w_006_1624, w_006_1625, w_006_1626, w_006_1627, w_006_1629, w_006_1630, w_006_1631, w_006_1632, w_006_1633, w_006_1634, w_006_1635, w_006_1636, w_006_1637, w_006_1639, w_006_1640, w_006_1641, w_006_1642, w_006_1643, w_006_1644, w_006_1645, w_006_1646, w_006_1647, w_006_1648, w_006_1649, w_006_1650, w_006_1651, w_006_1652, w_006_1653, w_006_1654, w_006_1655, w_006_1656, w_006_1657, w_006_1658, w_006_1659, w_006_1660, w_006_1661, w_006_1662, w_006_1663, w_006_1664, w_006_1665, w_006_1666, w_006_1667, w_006_1668, w_006_1669, w_006_1670, w_006_1671, w_006_1672, w_006_1673, w_006_1674, w_006_1675, w_006_1676, w_006_1677, w_006_1678, w_006_1679, w_006_1680, w_006_1681, w_006_1682, w_006_1683, w_006_1684, w_006_1685, w_006_1686, w_006_1687, w_006_1688, w_006_1689, w_006_1690, w_006_1691, w_006_1692, w_006_1693, w_006_1694, w_006_1695, w_006_1696, w_006_1697, w_006_1698, w_006_1699, w_006_1700, w_006_1701, w_006_1702, w_006_1703, w_006_1704, w_006_1705, w_006_1706, w_006_1707, w_006_1708, w_006_1709, w_006_1710, w_006_1711, w_006_1712, w_006_1713, w_006_1714, w_006_1715, w_006_1716, w_006_1717, w_006_1718, w_006_1719, w_006_1720, w_006_1721, w_006_1722, w_006_1723, w_006_1724, w_006_1725, w_006_1726, w_006_1727, w_006_1728, w_006_1729, w_006_1730, w_006_1731, w_006_1732, w_006_1733, w_006_1734, w_006_1735, w_006_1736, w_006_1737, w_006_1738, w_006_1739, w_006_1740, w_006_1741, w_006_1742, w_006_1743, w_006_1744, w_006_1745, w_006_1746, w_006_1747, w_006_1748, w_006_1749, w_006_1750, w_006_1751, w_006_1752, w_006_1753, w_006_1754, w_006_1755, w_006_1756, w_006_1757, w_006_1758, w_006_1759, w_006_1760, w_006_1761, w_006_1762, w_006_1763, w_006_1764, w_006_1765, w_006_1766, w_006_1767, w_006_1768, w_006_1769, w_006_1770, w_006_1771, w_006_1772, w_006_1773, w_006_1774, w_006_1775, w_006_1776, w_006_1777, w_006_1778, w_006_1779, w_006_1780, w_006_1781, w_006_1782, w_006_1783, w_006_1784, w_006_1785, w_006_1786, w_006_1787, w_006_1788, w_006_1789, w_006_1790, w_006_1791, w_006_1792, w_006_1793, w_006_1794, w_006_1795, w_006_1796, w_006_1797, w_006_1798, w_006_1799, w_006_1800, w_006_1801, w_006_1802, w_006_1803, w_006_1804, w_006_1805, w_006_1806, w_006_1807, w_006_1808, w_006_1809, w_006_1810, w_006_1811, w_006_1812, w_006_1813, w_006_1814, w_006_1815, w_006_1816, w_006_1817, w_006_1818, w_006_1819, w_006_1820, w_006_1821, w_006_1822, w_006_1823, w_006_1824, w_006_1825, w_006_1826, w_006_1827, w_006_1828, w_006_1829, w_006_1830, w_006_1831, w_006_1832, w_006_1833, w_006_1834, w_006_1835, w_006_1836, w_006_1837, w_006_1838, w_006_1839, w_006_1840, w_006_1841, w_006_1842, w_006_1843, w_006_1844, w_006_1845, w_006_1846, w_006_1847, w_006_1848, w_006_1849, w_006_1850, w_006_1851, w_006_1852, w_006_1853, w_006_1854, w_006_1855, w_006_1856, w_006_1857, w_006_1858, w_006_1859, w_006_1860, w_006_1861, w_006_1862, w_006_1863, w_006_1864, w_006_1865, w_006_1866, w_006_1867, w_006_1868, w_006_1869, w_006_1870, w_006_1871, w_006_1872, w_006_1873, w_006_1874, w_006_1875, w_006_1876, w_006_1877, w_006_1878, w_006_1879, w_006_1880, w_006_1881, w_006_1882, w_006_1883, w_006_1884, w_006_1885, w_006_1886, w_006_1887, w_006_1888, w_006_1889, w_006_1890, w_006_1891, w_006_1892, w_006_1893, w_006_1894, w_006_1895, w_006_1896, w_006_1897, w_006_1898, w_006_1899, w_006_1900, w_006_1901, w_006_1902, w_006_1903, w_006_1904, w_006_1905, w_006_1906, w_006_1907, w_006_1908, w_006_1909, w_006_1910, w_006_1911, w_006_1912, w_006_1913, w_006_1914, w_006_1915, w_006_1916, w_006_1917, w_006_1918, w_006_1919, w_006_1920, w_006_1921, w_006_1922, w_006_1923, w_006_1924, w_006_1925, w_006_1927, w_006_1928, w_006_1929, w_006_1930, w_006_1931, w_006_1932, w_006_1933, w_006_1934, w_006_1935, w_006_1936, w_006_1937, w_006_1938, w_006_1939, w_006_1940, w_006_1941, w_006_1942, w_006_1943, w_006_1944, w_006_1945, w_006_1946, w_006_1947, w_006_1948, w_006_1949, w_006_1950, w_006_1951, w_006_1952, w_006_1953, w_006_1954, w_006_1955, w_006_1956, w_006_1957, w_006_1958, w_006_1959, w_006_1960, w_006_1961, w_006_1962, w_006_1963, w_006_1964, w_006_1965, w_006_1966, w_006_1967, w_006_1968, w_006_1969, w_006_1970, w_006_1971, w_006_1972, w_006_1973, w_006_1974, w_006_1975, w_006_1976, w_006_1977, w_006_1978, w_006_1979, w_006_1980, w_006_1981, w_006_1982, w_006_1983, w_006_1984, w_006_1985, w_006_1986, w_006_1987, w_006_1988, w_006_1989, w_006_1990, w_006_1991, w_006_1992, w_006_1993, w_006_1994, w_006_1995, w_006_1996, w_006_1997, w_006_1998, w_006_1999, w_006_2000, w_006_2001, w_006_2002, w_006_2003, w_006_2004, w_006_2005, w_006_2006, w_006_2007, w_006_2008, w_006_2009, w_006_2010, w_006_2011, w_006_2012, w_006_2013, w_006_2014, w_006_2015, w_006_2016, w_006_2017, w_006_2018, w_006_2019, w_006_2020, w_006_2021, w_006_2022, w_006_2023, w_006_2024, w_006_2025, w_006_2026, w_006_2027, w_006_2028, w_006_2029, w_006_2030, w_006_2031, w_006_2032, w_006_2033, w_006_2034, w_006_2035, w_006_2036, w_006_2037, w_006_2038, w_006_2039, w_006_2040, w_006_2041, w_006_2042, w_006_2043, w_006_2044, w_006_2045, w_006_2046, w_006_2047, w_006_2048, w_006_2049, w_006_2050, w_006_2051, w_006_2052, w_006_2053, w_006_2054, w_006_2055, w_006_2056, w_006_2057, w_006_2058, w_006_2059, w_006_2060, w_006_2061, w_006_2062, w_006_2063, w_006_2065, w_006_2066, w_006_2067, w_006_2068, w_006_2069, w_006_2070, w_006_2071, w_006_2072, w_006_2073, w_006_2074, w_006_2075, w_006_2076, w_006_2077, w_006_2078, w_006_2079, w_006_2080, w_006_2081, w_006_2082, w_006_2083, w_006_2084, w_006_2085, w_006_2086, w_006_2087, w_006_2088, w_006_2089, w_006_2090, w_006_2091, w_006_2092, w_006_2093, w_006_2094, w_006_2095, w_006_2096, w_006_2097, w_006_2098, w_006_2099, w_006_2100, w_006_2101, w_006_2102, w_006_2103, w_006_2104, w_006_2105, w_006_2106, w_006_2107, w_006_2108, w_006_2109, w_006_2110, w_006_2111, w_006_2112, w_006_2113, w_006_2114, w_006_2115, w_006_2116, w_006_2117, w_006_2118, w_006_2119, w_006_2120, w_006_2121, w_006_2122, w_006_2123, w_006_2124, w_006_2125, w_006_2126, w_006_2127, w_006_2128, w_006_2129, w_006_2130, w_006_2131, w_006_2132, w_006_2133, w_006_2134, w_006_2135, w_006_2136, w_006_2137, w_006_2138, w_006_2139, w_006_2140, w_006_2141, w_006_2142, w_006_2143, w_006_2144, w_006_2145, w_006_2146, w_006_2147, w_006_2148, w_006_2149, w_006_2150, w_006_2151, w_006_2152, w_006_2153, w_006_2154, w_006_2155, w_006_2156, w_006_2157, w_006_2158, w_006_2159, w_006_2160, w_006_2161, w_006_2162, w_006_2163, w_006_2164, w_006_2165, w_006_2166, w_006_2167, w_006_2168, w_006_2169, w_006_2170, w_006_2171, w_006_2172, w_006_2173, w_006_2174, w_006_2175, w_006_2176, w_006_2177, w_006_2178, w_006_2179, w_006_2180, w_006_2181, w_006_2182, w_006_2183, w_006_2184, w_006_2185, w_006_2186, w_006_2187, w_006_2188, w_006_2189, w_006_2190, w_006_2191, w_006_2192, w_006_2193, w_006_2194, w_006_2195, w_006_2196, w_006_2197, w_006_2198, w_006_2199, w_006_2200, w_006_2201, w_006_2202, w_006_2203, w_006_2204, w_006_2205, w_006_2206, w_006_2207, w_006_2208, w_006_2209, w_006_2210, w_006_2211, w_006_2212, w_006_2213, w_006_2215, w_006_2216, w_006_2217, w_006_2218, w_006_2219, w_006_2220, w_006_2221, w_006_2222, w_006_2223, w_006_2224, w_006_2225, w_006_2226, w_006_2227, w_006_2228, w_006_2229, w_006_2230, w_006_2231, w_006_2232, w_006_2233, w_006_2234, w_006_2235, w_006_2236, w_006_2237, w_006_2238, w_006_2239, w_006_2240, w_006_2241, w_006_2242, w_006_2243, w_006_2244, w_006_2245, w_006_2246, w_006_2247, w_006_2248, w_006_2249, w_006_2250, w_006_2251, w_006_2252, w_006_2253, w_006_2254, w_006_2255, w_006_2256, w_006_2257, w_006_2258, w_006_2259, w_006_2260, w_006_2261, w_006_2262, w_006_2263, w_006_2264, w_006_2265, w_006_2266, w_006_2267, w_006_2268, w_006_2269, w_006_2270, w_006_2271, w_006_2272, w_006_2273, w_006_2274, w_006_2275, w_006_2276, w_006_2277, w_006_2278, w_006_2279, w_006_2280, w_006_2281, w_006_2282, w_006_2283, w_006_2284, w_006_2285, w_006_2286, w_006_2287, w_006_2288, w_006_2289, w_006_2290, w_006_2291, w_006_2292, w_006_2293, w_006_2294, w_006_2295, w_006_2296, w_006_2297, w_006_2298, w_006_2299, w_006_2300, w_006_2301, w_006_2302, w_006_2303, w_006_2304, w_006_2305, w_006_2306, w_006_2307, w_006_2308, w_006_2309, w_006_2310, w_006_2311, w_006_2312, w_006_2313, w_006_2314, w_006_2315, w_006_2316, w_006_2317, w_006_2318, w_006_2319, w_006_2320, w_006_2321, w_006_2322, w_006_2323, w_006_2324, w_006_2325, w_006_2326, w_006_2327, w_006_2328, w_006_2329, w_006_2330, w_006_2331, w_006_2332, w_006_2333, w_006_2334, w_006_2335, w_006_2336, w_006_2337, w_006_2338, w_006_2339, w_006_2340, w_006_2341, w_006_2342, w_006_2343, w_006_2344, w_006_2345, w_006_2346, w_006_2347, w_006_2348, w_006_2349, w_006_2350, w_006_2351, w_006_2352, w_006_2353, w_006_2354, w_006_2355, w_006_2356, w_006_2357, w_006_2358, w_006_2359, w_006_2360, w_006_2361, w_006_2362, w_006_2363, w_006_2364, w_006_2365, w_006_2366, w_006_2367, w_006_2368, w_006_2369, w_006_2370, w_006_2371, w_006_2372, w_006_2373, w_006_2374, w_006_2375, w_006_2376, w_006_2377, w_006_2378, w_006_2379, w_006_2380, w_006_2381, w_006_2382, w_006_2383, w_006_2384, w_006_2385, w_006_2386, w_006_2387, w_006_2388, w_006_2389, w_006_2390, w_006_2391, w_006_2392, w_006_2393, w_006_2394, w_006_2395, w_006_2396, w_006_2397, w_006_2398, w_006_2399, w_006_2400, w_006_2401, w_006_2402, w_006_2403, w_006_2404, w_006_2405, w_006_2406, w_006_2407, w_006_2408, w_006_2409, w_006_2410, w_006_2411, w_006_2412, w_006_2413, w_006_2414, w_006_2415, w_006_2416, w_006_2417, w_006_2418, w_006_2419, w_006_2420, w_006_2421, w_006_2422, w_006_2423, w_006_2424, w_006_2425, w_006_2426, w_006_2427, w_006_2428, w_006_2429, w_006_2430, w_006_2431, w_006_2432, w_006_2433, w_006_2434, w_006_2435, w_006_2436, w_006_2437, w_006_2438, w_006_2439, w_006_2440, w_006_2441, w_006_2442, w_006_2443, w_006_2444, w_006_2445, w_006_2446, w_006_2447, w_006_2448, w_006_2449, w_006_2450, w_006_2451, w_006_2452, w_006_2453, w_006_2454, w_006_2455, w_006_2456, w_006_2457, w_006_2458, w_006_2459, w_006_2460, w_006_2461, w_006_2462, w_006_2463, w_006_2464, w_006_2465, w_006_2466, w_006_2467, w_006_2468, w_006_2469, w_006_2470, w_006_2471, w_006_2472, w_006_2473, w_006_2474, w_006_2475, w_006_2476, w_006_2477, w_006_2478, w_006_2479, w_006_2480, w_006_2481, w_006_2482, w_006_2483, w_006_2484, w_006_2485, w_006_2486, w_006_2487, w_006_2488, w_006_2489, w_006_2490, w_006_2491, w_006_2492, w_006_2493, w_006_2494, w_006_2495, w_006_2496, w_006_2497, w_006_2498, w_006_2499, w_006_2500, w_006_2501, w_006_2502, w_006_2503, w_006_2504, w_006_2505, w_006_2506, w_006_2507, w_006_2508, w_006_2509, w_006_2510, w_006_2511, w_006_2512, w_006_2513, w_006_2514, w_006_2515, w_006_2516, w_006_2517, w_006_2518, w_006_2519, w_006_2520, w_006_2521, w_006_2522, w_006_2523, w_006_2524, w_006_2525, w_006_2526, w_006_2527, w_006_2528, w_006_2529, w_006_2530, w_006_2531, w_006_2532, w_006_2533, w_006_2534, w_006_2535, w_006_2536, w_006_2537, w_006_2538, w_006_2539, w_006_2540, w_006_2541, w_006_2542, w_006_2543, w_006_2544, w_006_2545, w_006_2546, w_006_2547, w_006_2548, w_006_2549, w_006_2550, w_006_2551, w_006_2552, w_006_2553, w_006_2554, w_006_2555, w_006_2556, w_006_2557, w_006_2558, w_006_2559, w_006_2560, w_006_2561, w_006_2562, w_006_2563, w_006_2564, w_006_2565, w_006_2566, w_006_2567, w_006_2568, w_006_2569, w_006_2570, w_006_2571, w_006_2572, w_006_2573, w_006_2574, w_006_2575, w_006_2576, w_006_2577, w_006_2578, w_006_2579, w_006_2580, w_006_2581, w_006_2582, w_006_2583, w_006_2584, w_006_2585, w_006_2586, w_006_2587, w_006_2588, w_006_2589, w_006_2590, w_006_2591, w_006_2592, w_006_2593, w_006_2594, w_006_2595, w_006_2596, w_006_2597, w_006_2598, w_006_2599, w_006_2600, w_006_2601, w_006_2602, w_006_2603, w_006_2604, w_006_2605, w_006_2606, w_006_2607, w_006_2608, w_006_2609, w_006_2610, w_006_2611, w_006_2612, w_006_2613, w_006_2614, w_006_2615, w_006_2616, w_006_2617, w_006_2618, w_006_2619, w_006_2620, w_006_2621, w_006_2622, w_006_2623, w_006_2624, w_006_2625, w_006_2626, w_006_2627, w_006_2628, w_006_2629, w_006_2630, w_006_2631, w_006_2632, w_006_2633, w_006_2634, w_006_2635, w_006_2636, w_006_2637, w_006_2638, w_006_2639, w_006_2640, w_006_2641, w_006_2642, w_006_2643, w_006_2644, w_006_2645, w_006_2646, w_006_2647, w_006_2648, w_006_2649, w_006_2650, w_006_2651, w_006_2652, w_006_2653, w_006_2654, w_006_2655, w_006_2656, w_006_2657, w_006_2658, w_006_2659, w_006_2660, w_006_2661, w_006_2662, w_006_2663, w_006_2664, w_006_2665, w_006_2666, w_006_2667, w_006_2668, w_006_2669, w_006_2670, w_006_2671, w_006_2672, w_006_2673, w_006_2674, w_006_2675, w_006_2676, w_006_2677, w_006_2678, w_006_2679, w_006_2680, w_006_2681, w_006_2682, w_006_2683, w_006_2684, w_006_2685, w_006_2686, w_006_2687, w_006_2688, w_006_2689, w_006_2690, w_006_2691, w_006_2692, w_006_2693, w_006_2694, w_006_2695, w_006_2696, w_006_2697, w_006_2698, w_006_2699, w_006_2700, w_006_2701, w_006_2702, w_006_2703, w_006_2704, w_006_2705, w_006_2706, w_006_2707, w_006_2708, w_006_2709, w_006_2710, w_006_2711, w_006_2712, w_006_2713, w_006_2714, w_006_2715, w_006_2716, w_006_2717, w_006_2718, w_006_2719, w_006_2720, w_006_2721, w_006_2722, w_006_2723, w_006_2724, w_006_2725, w_006_2726, w_006_2727, w_006_2728, w_006_2729, w_006_2730, w_006_2731, w_006_2732, w_006_2733, w_006_2734, w_006_2735, w_006_2736, w_006_2737, w_006_2738, w_006_2739, w_006_2740, w_006_2741, w_006_2742, w_006_2743, w_006_2744, w_006_2745, w_006_2746, w_006_2747, w_006_2748, w_006_2749, w_006_2750, w_006_2751, w_006_2752, w_006_2753, w_006_2754, w_006_2755, w_006_2756, w_006_2757, w_006_2758, w_006_2759, w_006_2760, w_006_2761, w_006_2762, w_006_2763, w_006_2764, w_006_2765, w_006_2766, w_006_2767, w_006_2768, w_006_2769, w_006_2770, w_006_2771, w_006_2772, w_006_2773, w_006_2774, w_006_2775, w_006_2776, w_006_2777, w_006_2778, w_006_2779, w_006_2780, w_006_2781, w_006_2782, w_006_2783, w_006_2784, w_006_2785, w_006_2786, w_006_2787, w_006_2788, w_006_2789, w_006_2790, w_006_2791, w_006_2792, w_006_2793, w_006_2794, w_006_2795, w_006_2796, w_006_2797, w_006_2798, w_006_2799, w_006_2800, w_006_2801, w_006_2802, w_006_2803, w_006_2804, w_006_2805, w_006_2806, w_006_2807, w_006_2808, w_006_2809, w_006_2810, w_006_2811, w_006_2812, w_006_2813, w_006_2814, w_006_2815, w_006_2816, w_006_2817, w_006_2818, w_006_2819, w_006_2820, w_006_2821, w_006_2822, w_006_2823, w_006_2824, w_006_2825, w_006_2826, w_006_2827, w_006_2828, w_006_2829, w_006_2830, w_006_2831, w_006_2832, w_006_2833, w_006_2834, w_006_2835, w_006_2836, w_006_2837, w_006_2838, w_006_2839, w_006_2840, w_006_2841, w_006_2842, w_006_2843, w_006_2844, w_006_2845, w_006_2846, w_006_2847, w_006_2848, w_006_2849, w_006_2850, w_006_2851, w_006_2852, w_006_2853, w_006_2854, w_006_2855, w_006_2856, w_006_2857, w_006_2858, w_006_2859, w_006_2860, w_006_2861, w_006_2862, w_006_2863, w_006_2864, w_006_2865, w_006_2866, w_006_2867, w_006_2868, w_006_2869, w_006_2870, w_006_2871, w_006_2872, w_006_2873, w_006_2874, w_006_2875, w_006_2876, w_006_2877, w_006_2878, w_006_2879, w_006_2880, w_006_2881, w_006_2882, w_006_2883, w_006_2884, w_006_2885, w_006_2886, w_006_2887, w_006_2888, w_006_2889, w_006_2890, w_006_2891, w_006_2892, w_006_2893, w_006_2894, w_006_2895, w_006_2896, w_006_2897, w_006_2898, w_006_2899, w_006_2900, w_006_2901, w_006_2902, w_006_2903, w_006_2904, w_006_2905, w_006_2906, w_006_2907, w_006_2908, w_006_2909, w_006_2910, w_006_2911, w_006_2912, w_006_2913, w_006_2914, w_006_2915, w_006_2916, w_006_2917, w_006_2918, w_006_2919, w_006_2920, w_006_2921, w_006_2922, w_006_2923, w_006_2925, w_006_2926, w_006_2927, w_006_2928, w_006_2929, w_006_2930, w_006_2931, w_006_2932, w_006_2933, w_006_2934, w_006_2935, w_006_2936, w_006_2937, w_006_2938, w_006_2939, w_006_2940, w_006_2941, w_006_2942, w_006_2943, w_006_2944, w_006_2945, w_006_2946, w_006_2947, w_006_2948, w_006_2949, w_006_2950, w_006_2951, w_006_2952, w_006_2953, w_006_2954, w_006_2955, w_006_2956, w_006_2957, w_006_2958, w_006_2959, w_006_2960, w_006_2961, w_006_2962, w_006_2963, w_006_2964, w_006_2965, w_006_2966, w_006_2967, w_006_2968, w_006_2969, w_006_2970, w_006_2971, w_006_2972, w_006_2973, w_006_2974, w_006_2975, w_006_2976, w_006_2977, w_006_2978, w_006_2979, w_006_2980, w_006_2981, w_006_2982, w_006_2983, w_006_2984, w_006_2985, w_006_2986, w_006_2987, w_006_2988, w_006_2989, w_006_2990, w_006_2991, w_006_2992, w_006_2993, w_006_2994, w_006_2995, w_006_2996, w_006_2997, w_006_2998, w_006_2999, w_006_3000, w_006_3001, w_006_3002, w_006_3003, w_006_3004, w_006_3005, w_006_3006, w_006_3007, w_006_3008, w_006_3009, w_006_3010, w_006_3011, w_006_3012, w_006_3013, w_006_3014, w_006_3015, w_006_3016, w_006_3017, w_006_3018, w_006_3019, w_006_3020, w_006_3021, w_006_3022, w_006_3023, w_006_3024, w_006_3025, w_006_3026, w_006_3027, w_006_3028, w_006_3029, w_006_3030, w_006_3031, w_006_3032, w_006_3033, w_006_3034, w_006_3035, w_006_3036, w_006_3037, w_006_3038, w_006_3039, w_006_3040, w_006_3041, w_006_3042, w_006_3043, w_006_3044, w_006_3045, w_006_3046, w_006_3047, w_006_3048, w_006_3049, w_006_3050, w_006_3051, w_006_3052, w_006_3053, w_006_3054, w_006_3055, w_006_3056, w_006_3057, w_006_3058, w_006_3059, w_006_3060, w_006_3061, w_006_3062, w_006_3063, w_006_3064, w_006_3065, w_006_3066, w_006_3067, w_006_3068, w_006_3069, w_006_3070, w_006_3071, w_006_3072, w_006_3073, w_006_3074, w_006_3075, w_006_3076, w_006_3077, w_006_3078, w_006_3079, w_006_3080, w_006_3081, w_006_3082, w_006_3083, w_006_3084, w_006_3085, w_006_3086, w_006_3087, w_006_3088, w_006_3089, w_006_3090, w_006_3091, w_006_3092, w_006_3093, w_006_3094, w_006_3095, w_006_3096, w_006_3097, w_006_3098, w_006_3099, w_006_3100, w_006_3101, w_006_3102, w_006_3103, w_006_3104, w_006_3105, w_006_3106, w_006_3107, w_006_3108, w_006_3109, w_006_3110, w_006_3111, w_006_3112, w_006_3113, w_006_3114, w_006_3115, w_006_3116, w_006_3117, w_006_3118, w_006_3119, w_006_3120, w_006_3121, w_006_3122, w_006_3123, w_006_3124, w_006_3125, w_006_3126, w_006_3127, w_006_3128, w_006_3129, w_006_3130, w_006_3131, w_006_3132, w_006_3133, w_006_3134, w_006_3135, w_006_3136, w_006_3137, w_006_3138, w_006_3139, w_006_3140, w_006_3141, w_006_3142, w_006_3143, w_006_3144, w_006_3145, w_006_3146, w_006_3147, w_006_3148, w_006_3149, w_006_3150, w_006_3151, w_006_3152, w_006_3153, w_006_3154, w_006_3155, w_006_3156, w_006_3157, w_006_3158, w_006_3159, w_006_3160, w_006_3161, w_006_3162, w_006_3163, w_006_3164, w_006_3165, w_006_3166, w_006_3167, w_006_3168, w_006_3169, w_006_3170, w_006_3171, w_006_3172, w_006_3173, w_006_3174, w_006_3175, w_006_3176, w_006_3177, w_006_3178, w_006_3179, w_006_3180, w_006_3181, w_006_3182, w_006_3183, w_006_3184, w_006_3185, w_006_3186, w_006_3187, w_006_3188, w_006_3189, w_006_3190, w_006_3191, w_006_3192, w_006_3193, w_006_3194, w_006_3195, w_006_3196, w_006_3197, w_006_3198, w_006_3199, w_006_3200, w_006_3201, w_006_3202, w_006_3203, w_006_3204, w_006_3205, w_006_3206, w_006_3207, w_006_3208, w_006_3210, w_006_3211, w_006_3212, w_006_3213, w_006_3214, w_006_3215, w_006_3216, w_006_3217, w_006_3218, w_006_3219, w_006_3220, w_006_3221, w_006_3222, w_006_3223, w_006_3224, w_006_3225, w_006_3226, w_006_3227, w_006_3228, w_006_3229, w_006_3230, w_006_3231, w_006_3232, w_006_3233, w_006_3234, w_006_3235, w_006_3236, w_006_3237, w_006_3238, w_006_3239, w_006_3240, w_006_3241, w_006_3242, w_006_3243, w_006_3244;
  wire w_007_000, w_007_001, w_007_002, w_007_003, w_007_004, w_007_005, w_007_006, w_007_007, w_007_008, w_007_009, w_007_010, w_007_011, w_007_012, w_007_013, w_007_014, w_007_015, w_007_016, w_007_017, w_007_018, w_007_019, w_007_020, w_007_021, w_007_022, w_007_023, w_007_024, w_007_025, w_007_026, w_007_027, w_007_028, w_007_029, w_007_030, w_007_031, w_007_032, w_007_033, w_007_034, w_007_035, w_007_036, w_007_037, w_007_038, w_007_039, w_007_040, w_007_041, w_007_042, w_007_043, w_007_044, w_007_045, w_007_046, w_007_047, w_007_048, w_007_049, w_007_050, w_007_051, w_007_052, w_007_053, w_007_054, w_007_055, w_007_056, w_007_057, w_007_058, w_007_059, w_007_060, w_007_061, w_007_062, w_007_063, w_007_064, w_007_065, w_007_066, w_007_067, w_007_068, w_007_069, w_007_070, w_007_071, w_007_072, w_007_073, w_007_074, w_007_075, w_007_076, w_007_077, w_007_078, w_007_079, w_007_080, w_007_081, w_007_082, w_007_083, w_007_084, w_007_085, w_007_086, w_007_087, w_007_088, w_007_089, w_007_090, w_007_091, w_007_092, w_007_093, w_007_094, w_007_095, w_007_096, w_007_097, w_007_098, w_007_099, w_007_100, w_007_101, w_007_102, w_007_103, w_007_104, w_007_105, w_007_106, w_007_107, w_007_108, w_007_109, w_007_110, w_007_111, w_007_112, w_007_113, w_007_114, w_007_115, w_007_116, w_007_117, w_007_118, w_007_119, w_007_120, w_007_121, w_007_122, w_007_123, w_007_124, w_007_125, w_007_126, w_007_127, w_007_128, w_007_129, w_007_130, w_007_131, w_007_132, w_007_133, w_007_134, w_007_135, w_007_136, w_007_137, w_007_138, w_007_139, w_007_140, w_007_141, w_007_142, w_007_143, w_007_144, w_007_145, w_007_146, w_007_147, w_007_148, w_007_149, w_007_150, w_007_151, w_007_152, w_007_153, w_007_154, w_007_155, w_007_156, w_007_157, w_007_158, w_007_159, w_007_160, w_007_161, w_007_162, w_007_163, w_007_164, w_007_165, w_007_166, w_007_167, w_007_168, w_007_169, w_007_170, w_007_171, w_007_172, w_007_173, w_007_174, w_007_175, w_007_176, w_007_177, w_007_178, w_007_179, w_007_180, w_007_181, w_007_182, w_007_183, w_007_184, w_007_185, w_007_186, w_007_187, w_007_188, w_007_189, w_007_190, w_007_191, w_007_192, w_007_193, w_007_194, w_007_195, w_007_196, w_007_197, w_007_198, w_007_199, w_007_200, w_007_201, w_007_202, w_007_203, w_007_204, w_007_205, w_007_206, w_007_207, w_007_208, w_007_209, w_007_210, w_007_211, w_007_212, w_007_213, w_007_214, w_007_215, w_007_216, w_007_217, w_007_218, w_007_219, w_007_220, w_007_221, w_007_222, w_007_223, w_007_224, w_007_225, w_007_226, w_007_227, w_007_228, w_007_229, w_007_230, w_007_231, w_007_232, w_007_233, w_007_234, w_007_235, w_007_236, w_007_237, w_007_238, w_007_239, w_007_240, w_007_241, w_007_242, w_007_243, w_007_244, w_007_245, w_007_246, w_007_247, w_007_248, w_007_249, w_007_250, w_007_251, w_007_252, w_007_253, w_007_254, w_007_255, w_007_256, w_007_257, w_007_258, w_007_259, w_007_260, w_007_261, w_007_262, w_007_263, w_007_264, w_007_265, w_007_266, w_007_267, w_007_268, w_007_269, w_007_270, w_007_271, w_007_272, w_007_273, w_007_274, w_007_275, w_007_276, w_007_277, w_007_278, w_007_279, w_007_280, w_007_281, w_007_282, w_007_283, w_007_284, w_007_285, w_007_286, w_007_287, w_007_288, w_007_289, w_007_290, w_007_291, w_007_292, w_007_293, w_007_294, w_007_295, w_007_296, w_007_297, w_007_298, w_007_299, w_007_300, w_007_301, w_007_302, w_007_303, w_007_304, w_007_305, w_007_306, w_007_307, w_007_308, w_007_309, w_007_310, w_007_311, w_007_312, w_007_313, w_007_314, w_007_315, w_007_316, w_007_317, w_007_318, w_007_319, w_007_320, w_007_321, w_007_322, w_007_323, w_007_324, w_007_325, w_007_326, w_007_327, w_007_328, w_007_329, w_007_330, w_007_331, w_007_332, w_007_333, w_007_334, w_007_335, w_007_336, w_007_337, w_007_338, w_007_339, w_007_340, w_007_341, w_007_342, w_007_343, w_007_344, w_007_345, w_007_346, w_007_347, w_007_348, w_007_349, w_007_350, w_007_351, w_007_352, w_007_353, w_007_354, w_007_355, w_007_356, w_007_357, w_007_358, w_007_359, w_007_360, w_007_361, w_007_362, w_007_363, w_007_364, w_007_365, w_007_366, w_007_367, w_007_368, w_007_369, w_007_370, w_007_371, w_007_372, w_007_373, w_007_374, w_007_375, w_007_376, w_007_377, w_007_378, w_007_379, w_007_380, w_007_381, w_007_382, w_007_383, w_007_384, w_007_385, w_007_386, w_007_387, w_007_388, w_007_389, w_007_390, w_007_391, w_007_392, w_007_393, w_007_394, w_007_395, w_007_396, w_007_397, w_007_398, w_007_399, w_007_400, w_007_401, w_007_402, w_007_403, w_007_404, w_007_405, w_007_406, w_007_407, w_007_408, w_007_409, w_007_410, w_007_411, w_007_412, w_007_413, w_007_414, w_007_415, w_007_416, w_007_417, w_007_418, w_007_419, w_007_420, w_007_421, w_007_422, w_007_423, w_007_424, w_007_425, w_007_426, w_007_427, w_007_428, w_007_429, w_007_430, w_007_431, w_007_432, w_007_433, w_007_434, w_007_435, w_007_436, w_007_437, w_007_438, w_007_439, w_007_440, w_007_441, w_007_442, w_007_443, w_007_444, w_007_445, w_007_446, w_007_447, w_007_448, w_007_449, w_007_450, w_007_451, w_007_452, w_007_453, w_007_454, w_007_455, w_007_456, w_007_457, w_007_458, w_007_459, w_007_460, w_007_461, w_007_462, w_007_463, w_007_464, w_007_465, w_007_466, w_007_467, w_007_468, w_007_469, w_007_470, w_007_471, w_007_472, w_007_473, w_007_474, w_007_475, w_007_476, w_007_477, w_007_478, w_007_479, w_007_480, w_007_481, w_007_482, w_007_483, w_007_484, w_007_485, w_007_486, w_007_487, w_007_488, w_007_489, w_007_490, w_007_491, w_007_492, w_007_493, w_007_494, w_007_495, w_007_496, w_007_497, w_007_498, w_007_499, w_007_500, w_007_501, w_007_502, w_007_503, w_007_504, w_007_505, w_007_506, w_007_507, w_007_508, w_007_509, w_007_510, w_007_511, w_007_512, w_007_513, w_007_514, w_007_515, w_007_516, w_007_517, w_007_518, w_007_519, w_007_520, w_007_521, w_007_522, w_007_523, w_007_524, w_007_525, w_007_526, w_007_527, w_007_528, w_007_529, w_007_530, w_007_531, w_007_532, w_007_533, w_007_534, w_007_535, w_007_536, w_007_537, w_007_538, w_007_539, w_007_540, w_007_541, w_007_542, w_007_543, w_007_544, w_007_545, w_007_546, w_007_547, w_007_548, w_007_549, w_007_550, w_007_551, w_007_552, w_007_553, w_007_554, w_007_555, w_007_556, w_007_557, w_007_558, w_007_559, w_007_560, w_007_561, w_007_562, w_007_563, w_007_564, w_007_565, w_007_566, w_007_567, w_007_568, w_007_569, w_007_570, w_007_571, w_007_572, w_007_573, w_007_574, w_007_575, w_007_576, w_007_577, w_007_578, w_007_579, w_007_580, w_007_581, w_007_582, w_007_583, w_007_584, w_007_585, w_007_586, w_007_587, w_007_588, w_007_589, w_007_590, w_007_591, w_007_592, w_007_593, w_007_594, w_007_595, w_007_596, w_007_597, w_007_598, w_007_599, w_007_600, w_007_601, w_007_602, w_007_603, w_007_604, w_007_605, w_007_606, w_007_607, w_007_608, w_007_609, w_007_610, w_007_611, w_007_612, w_007_613, w_007_614, w_007_615, w_007_616, w_007_617, w_007_618, w_007_619, w_007_620, w_007_621, w_007_622, w_007_623, w_007_624, w_007_625, w_007_626, w_007_627, w_007_628, w_007_629, w_007_630, w_007_631, w_007_632, w_007_633, w_007_634, w_007_635, w_007_636, w_007_637, w_007_638, w_007_639, w_007_640, w_007_641, w_007_642, w_007_643, w_007_644, w_007_645, w_007_646, w_007_647, w_007_648, w_007_649, w_007_650, w_007_651, w_007_652, w_007_653, w_007_654, w_007_655, w_007_656, w_007_657, w_007_658, w_007_659, w_007_660, w_007_661, w_007_662, w_007_663, w_007_664, w_007_665, w_007_666, w_007_667, w_007_668, w_007_669, w_007_670, w_007_671, w_007_672, w_007_673, w_007_674, w_007_675, w_007_676, w_007_677, w_007_678, w_007_679, w_007_680, w_007_681, w_007_682, w_007_683, w_007_684, w_007_685, w_007_686, w_007_687, w_007_688, w_007_689, w_007_690, w_007_691, w_007_692, w_007_693, w_007_694, w_007_695, w_007_696, w_007_697, w_007_698, w_007_699, w_007_700, w_007_701, w_007_702, w_007_703, w_007_704, w_007_705, w_007_706, w_007_707, w_007_708, w_007_709, w_007_710, w_007_711, w_007_712, w_007_713, w_007_714, w_007_715, w_007_716, w_007_717, w_007_718, w_007_719, w_007_720, w_007_721, w_007_722, w_007_723, w_007_724, w_007_725, w_007_726, w_007_727, w_007_728, w_007_729, w_007_730, w_007_731, w_007_732, w_007_733, w_007_734, w_007_735, w_007_736, w_007_737, w_007_738, w_007_739, w_007_740, w_007_741, w_007_742, w_007_743, w_007_744, w_007_745, w_007_746, w_007_747, w_007_748, w_007_749, w_007_750, w_007_751, w_007_752, w_007_753, w_007_754, w_007_755, w_007_756, w_007_757, w_007_758, w_007_759, w_007_760, w_007_761, w_007_762, w_007_763, w_007_764, w_007_765, w_007_766, w_007_767, w_007_768, w_007_769, w_007_770, w_007_771, w_007_772, w_007_773, w_007_774, w_007_775, w_007_776, w_007_777, w_007_778, w_007_779, w_007_780, w_007_781, w_007_782, w_007_783, w_007_784, w_007_785, w_007_786, w_007_787, w_007_788, w_007_789, w_007_790, w_007_791, w_007_792, w_007_793, w_007_794, w_007_795, w_007_796, w_007_797, w_007_798, w_007_799, w_007_800, w_007_801, w_007_802, w_007_803, w_007_804, w_007_805, w_007_806, w_007_807, w_007_808, w_007_809, w_007_810, w_007_811, w_007_812, w_007_813, w_007_814, w_007_815, w_007_816, w_007_817, w_007_818, w_007_819, w_007_820, w_007_821, w_007_822, w_007_823, w_007_824, w_007_825, w_007_826, w_007_827, w_007_828, w_007_829, w_007_830, w_007_831, w_007_832, w_007_833, w_007_834, w_007_835, w_007_836, w_007_837, w_007_838, w_007_839, w_007_840, w_007_841, w_007_842, w_007_843, w_007_844, w_007_845, w_007_846, w_007_847, w_007_848, w_007_849, w_007_850, w_007_851, w_007_852, w_007_853, w_007_854, w_007_855, w_007_856, w_007_857, w_007_858, w_007_859, w_007_860, w_007_861, w_007_862, w_007_863, w_007_864, w_007_865, w_007_866, w_007_867, w_007_868, w_007_869, w_007_870, w_007_871, w_007_872, w_007_873, w_007_874, w_007_875, w_007_876, w_007_877, w_007_878, w_007_879, w_007_880, w_007_881, w_007_882, w_007_883, w_007_884, w_007_885, w_007_886, w_007_887, w_007_888, w_007_889, w_007_890, w_007_891, w_007_892, w_007_893, w_007_894, w_007_895, w_007_896, w_007_897, w_007_898, w_007_899, w_007_900, w_007_901, w_007_902, w_007_903, w_007_904, w_007_905, w_007_906, w_007_907, w_007_908, w_007_909, w_007_910, w_007_911, w_007_912, w_007_913, w_007_914, w_007_915, w_007_916, w_007_917, w_007_918, w_007_919, w_007_920, w_007_921, w_007_922, w_007_923, w_007_924, w_007_925, w_007_926, w_007_927, w_007_928, w_007_929, w_007_930, w_007_931, w_007_932, w_007_933, w_007_934, w_007_935, w_007_936, w_007_937, w_007_938, w_007_939, w_007_940, w_007_941, w_007_942, w_007_943, w_007_944, w_007_945, w_007_946, w_007_947, w_007_948, w_007_949, w_007_950, w_007_951, w_007_952, w_007_953, w_007_954, w_007_955, w_007_956, w_007_957, w_007_958, w_007_959, w_007_960, w_007_961, w_007_962, w_007_963, w_007_964, w_007_965, w_007_966, w_007_967, w_007_968, w_007_969, w_007_970, w_007_971, w_007_972, w_007_973, w_007_974, w_007_975, w_007_976, w_007_977, w_007_978, w_007_979, w_007_980, w_007_981, w_007_982, w_007_983, w_007_984, w_007_985, w_007_986, w_007_987, w_007_988, w_007_989, w_007_990, w_007_991, w_007_992, w_007_993, w_007_994, w_007_995, w_007_996, w_007_997, w_007_998, w_007_999, w_007_1000, w_007_1001, w_007_1002, w_007_1003, w_007_1004, w_007_1005, w_007_1006, w_007_1007, w_007_1008, w_007_1009, w_007_1010, w_007_1011, w_007_1012, w_007_1013, w_007_1014, w_007_1015, w_007_1016, w_007_1017, w_007_1018, w_007_1019, w_007_1020, w_007_1021, w_007_1022, w_007_1023, w_007_1024, w_007_1025, w_007_1026, w_007_1027, w_007_1028, w_007_1029, w_007_1030, w_007_1031, w_007_1032, w_007_1033, w_007_1034, w_007_1035, w_007_1036, w_007_1037, w_007_1038, w_007_1039, w_007_1040, w_007_1041, w_007_1042, w_007_1043, w_007_1044, w_007_1045, w_007_1046, w_007_1047, w_007_1048, w_007_1049, w_007_1050, w_007_1051, w_007_1052, w_007_1053, w_007_1054, w_007_1055, w_007_1056, w_007_1057, w_007_1058, w_007_1059, w_007_1060, w_007_1061, w_007_1062, w_007_1063, w_007_1064, w_007_1065, w_007_1066, w_007_1067, w_007_1068, w_007_1069, w_007_1070, w_007_1071, w_007_1072, w_007_1073, w_007_1074, w_007_1075, w_007_1076, w_007_1077, w_007_1078, w_007_1079, w_007_1080, w_007_1081, w_007_1082, w_007_1083, w_007_1084, w_007_1085, w_007_1086, w_007_1087, w_007_1088, w_007_1089, w_007_1090, w_007_1091, w_007_1092, w_007_1093, w_007_1094, w_007_1095, w_007_1096, w_007_1097, w_007_1098, w_007_1099, w_007_1100, w_007_1101, w_007_1102, w_007_1103, w_007_1104, w_007_1105, w_007_1106, w_007_1107, w_007_1108, w_007_1109, w_007_1110, w_007_1111, w_007_1112, w_007_1113, w_007_1114, w_007_1115, w_007_1116, w_007_1117, w_007_1118, w_007_1119, w_007_1120, w_007_1121, w_007_1122, w_007_1123, w_007_1124, w_007_1125, w_007_1126, w_007_1127, w_007_1128, w_007_1129, w_007_1130, w_007_1131, w_007_1132, w_007_1133, w_007_1134, w_007_1135, w_007_1136, w_007_1137, w_007_1138, w_007_1139, w_007_1140, w_007_1141, w_007_1142, w_007_1143, w_007_1144, w_007_1145, w_007_1146, w_007_1147, w_007_1148, w_007_1149, w_007_1150, w_007_1151, w_007_1152, w_007_1153, w_007_1154, w_007_1155, w_007_1156, w_007_1157, w_007_1158, w_007_1159, w_007_1160, w_007_1161, w_007_1162, w_007_1163, w_007_1164, w_007_1165, w_007_1166, w_007_1167, w_007_1168, w_007_1169, w_007_1170, w_007_1171, w_007_1172, w_007_1173, w_007_1174, w_007_1175, w_007_1176, w_007_1177, w_007_1178, w_007_1179, w_007_1180, w_007_1181, w_007_1182, w_007_1183, w_007_1184, w_007_1185, w_007_1186, w_007_1187, w_007_1188, w_007_1189, w_007_1190, w_007_1191, w_007_1192, w_007_1193, w_007_1194, w_007_1195, w_007_1196, w_007_1197, w_007_1198, w_007_1199, w_007_1200, w_007_1201, w_007_1202, w_007_1203, w_007_1204, w_007_1205, w_007_1206, w_007_1207, w_007_1208, w_007_1209, w_007_1210, w_007_1211, w_007_1212, w_007_1213, w_007_1214, w_007_1215, w_007_1216, w_007_1217, w_007_1218, w_007_1219, w_007_1220, w_007_1221, w_007_1222, w_007_1223, w_007_1224, w_007_1225, w_007_1226, w_007_1227, w_007_1228, w_007_1229, w_007_1230, w_007_1231, w_007_1232, w_007_1233, w_007_1234, w_007_1235, w_007_1236, w_007_1237, w_007_1238, w_007_1239, w_007_1240, w_007_1241, w_007_1242, w_007_1243, w_007_1244, w_007_1245, w_007_1246, w_007_1247, w_007_1248, w_007_1249, w_007_1250, w_007_1251, w_007_1252, w_007_1253, w_007_1254, w_007_1255, w_007_1256, w_007_1257, w_007_1258, w_007_1259, w_007_1260, w_007_1261, w_007_1262, w_007_1263, w_007_1264, w_007_1265, w_007_1266, w_007_1267, w_007_1268, w_007_1269, w_007_1270, w_007_1271, w_007_1272, w_007_1273, w_007_1274, w_007_1275, w_007_1276, w_007_1277, w_007_1278, w_007_1279, w_007_1280, w_007_1281, w_007_1282, w_007_1283, w_007_1284, w_007_1285, w_007_1286, w_007_1287, w_007_1288, w_007_1289, w_007_1290, w_007_1291, w_007_1292, w_007_1293, w_007_1294, w_007_1295, w_007_1296, w_007_1297, w_007_1298, w_007_1299, w_007_1300, w_007_1301, w_007_1302, w_007_1303, w_007_1304, w_007_1305, w_007_1306, w_007_1307, w_007_1308, w_007_1309, w_007_1310, w_007_1311, w_007_1312, w_007_1313, w_007_1314, w_007_1315, w_007_1316, w_007_1317, w_007_1318, w_007_1319, w_007_1320, w_007_1321, w_007_1322, w_007_1323, w_007_1324, w_007_1325, w_007_1326, w_007_1327, w_007_1328, w_007_1329, w_007_1330, w_007_1331, w_007_1332, w_007_1333, w_007_1334, w_007_1335, w_007_1336, w_007_1337, w_007_1338, w_007_1339, w_007_1340, w_007_1341, w_007_1342, w_007_1343, w_007_1344, w_007_1345, w_007_1346, w_007_1347, w_007_1348, w_007_1349, w_007_1350, w_007_1351, w_007_1352, w_007_1353, w_007_1354, w_007_1355, w_007_1356, w_007_1357, w_007_1358, w_007_1359, w_007_1360, w_007_1361, w_007_1362, w_007_1363, w_007_1364, w_007_1365, w_007_1366, w_007_1367, w_007_1368, w_007_1369, w_007_1370, w_007_1371, w_007_1372, w_007_1373, w_007_1374, w_007_1375, w_007_1376, w_007_1377, w_007_1378, w_007_1379, w_007_1380, w_007_1381, w_007_1382, w_007_1383, w_007_1384, w_007_1385, w_007_1386, w_007_1387, w_007_1388, w_007_1389, w_007_1390, w_007_1391, w_007_1392, w_007_1393, w_007_1394, w_007_1395, w_007_1396, w_007_1397, w_007_1398, w_007_1399, w_007_1400, w_007_1401, w_007_1402, w_007_1403, w_007_1404, w_007_1405, w_007_1406, w_007_1407, w_007_1408, w_007_1409, w_007_1410, w_007_1411, w_007_1412, w_007_1413, w_007_1414, w_007_1415, w_007_1416, w_007_1417, w_007_1418, w_007_1419, w_007_1420, w_007_1421, w_007_1422, w_007_1423, w_007_1424, w_007_1425, w_007_1426, w_007_1427, w_007_1428, w_007_1429, w_007_1430, w_007_1431, w_007_1432, w_007_1433, w_007_1434, w_007_1435, w_007_1436, w_007_1437, w_007_1438, w_007_1439, w_007_1440, w_007_1441, w_007_1442, w_007_1443, w_007_1444, w_007_1445, w_007_1446, w_007_1447, w_007_1448, w_007_1449, w_007_1450, w_007_1451, w_007_1452, w_007_1453, w_007_1454, w_007_1455, w_007_1456, w_007_1457, w_007_1458, w_007_1459, w_007_1460, w_007_1461, w_007_1462, w_007_1463, w_007_1464, w_007_1465, w_007_1466, w_007_1467, w_007_1468, w_007_1469, w_007_1470, w_007_1471, w_007_1472, w_007_1473, w_007_1474, w_007_1475, w_007_1476, w_007_1477, w_007_1478, w_007_1479, w_007_1480, w_007_1481, w_007_1482, w_007_1483, w_007_1484, w_007_1485, w_007_1486, w_007_1487, w_007_1488, w_007_1489, w_007_1490, w_007_1491, w_007_1492, w_007_1493, w_007_1494, w_007_1495, w_007_1496, w_007_1497, w_007_1498, w_007_1499, w_007_1500, w_007_1501, w_007_1502, w_007_1503, w_007_1504, w_007_1505, w_007_1506, w_007_1507, w_007_1508, w_007_1509, w_007_1510, w_007_1511, w_007_1512, w_007_1513, w_007_1514, w_007_1515, w_007_1516, w_007_1517, w_007_1518, w_007_1519, w_007_1520, w_007_1521, w_007_1522, w_007_1523, w_007_1524, w_007_1525, w_007_1526, w_007_1527, w_007_1528, w_007_1529, w_007_1530, w_007_1531, w_007_1532, w_007_1533, w_007_1534, w_007_1535, w_007_1536, w_007_1537, w_007_1538, w_007_1539, w_007_1540, w_007_1541, w_007_1542, w_007_1543, w_007_1544, w_007_1545, w_007_1546, w_007_1547, w_007_1548, w_007_1549, w_007_1550, w_007_1551, w_007_1552, w_007_1553, w_007_1554, w_007_1555, w_007_1556, w_007_1557, w_007_1558, w_007_1559, w_007_1560, w_007_1561, w_007_1562, w_007_1563, w_007_1564, w_007_1565, w_007_1566, w_007_1567, w_007_1568, w_007_1569, w_007_1570, w_007_1571, w_007_1572, w_007_1573, w_007_1574, w_007_1575, w_007_1576, w_007_1577, w_007_1578, w_007_1579, w_007_1580, w_007_1581, w_007_1582, w_007_1583, w_007_1584, w_007_1585, w_007_1586, w_007_1587, w_007_1588, w_007_1589, w_007_1590, w_007_1591, w_007_1592, w_007_1593, w_007_1594, w_007_1595, w_007_1596, w_007_1597, w_007_1598, w_007_1599, w_007_1600, w_007_1601, w_007_1602, w_007_1603, w_007_1604, w_007_1605, w_007_1606, w_007_1607, w_007_1608, w_007_1609, w_007_1610, w_007_1611, w_007_1612, w_007_1613, w_007_1614, w_007_1615, w_007_1616, w_007_1617, w_007_1618, w_007_1619, w_007_1620, w_007_1621, w_007_1622, w_007_1623, w_007_1624, w_007_1625, w_007_1626, w_007_1627, w_007_1628, w_007_1629, w_007_1630, w_007_1631, w_007_1632, w_007_1633, w_007_1634, w_007_1635, w_007_1636, w_007_1637, w_007_1638, w_007_1639, w_007_1640, w_007_1641, w_007_1642, w_007_1643, w_007_1644, w_007_1645, w_007_1646, w_007_1647, w_007_1648, w_007_1649, w_007_1650, w_007_1651, w_007_1652, w_007_1653, w_007_1654, w_007_1655, w_007_1656, w_007_1657, w_007_1658, w_007_1659, w_007_1660, w_007_1661, w_007_1662, w_007_1663, w_007_1664, w_007_1665, w_007_1666, w_007_1667, w_007_1668, w_007_1669, w_007_1670, w_007_1671, w_007_1672, w_007_1673, w_007_1674, w_007_1675, w_007_1676, w_007_1677, w_007_1678, w_007_1679, w_007_1680, w_007_1681, w_007_1682, w_007_1683, w_007_1684, w_007_1685, w_007_1686, w_007_1687, w_007_1688, w_007_1689, w_007_1690, w_007_1691, w_007_1692, w_007_1693, w_007_1694, w_007_1695, w_007_1696, w_007_1697, w_007_1698, w_007_1699, w_007_1700, w_007_1701, w_007_1702, w_007_1703, w_007_1704, w_007_1705, w_007_1706, w_007_1707, w_007_1708, w_007_1709, w_007_1710, w_007_1711, w_007_1712, w_007_1713, w_007_1714, w_007_1715, w_007_1716, w_007_1717, w_007_1718, w_007_1719, w_007_1720, w_007_1721, w_007_1722, w_007_1723, w_007_1724, w_007_1725, w_007_1726, w_007_1727, w_007_1728, w_007_1729, w_007_1730, w_007_1731, w_007_1732, w_007_1733, w_007_1734, w_007_1735, w_007_1736, w_007_1737, w_007_1738, w_007_1739, w_007_1740, w_007_1741, w_007_1742, w_007_1743, w_007_1744, w_007_1745, w_007_1746, w_007_1747, w_007_1748, w_007_1749, w_007_1750, w_007_1751, w_007_1752, w_007_1753, w_007_1754, w_007_1755, w_007_1756, w_007_1757, w_007_1758, w_007_1759, w_007_1760, w_007_1761, w_007_1762, w_007_1763, w_007_1764, w_007_1765, w_007_1766, w_007_1767, w_007_1768, w_007_1769, w_007_1770, w_007_1771, w_007_1772, w_007_1773, w_007_1774, w_007_1775, w_007_1776, w_007_1777, w_007_1778, w_007_1779, w_007_1780, w_007_1781, w_007_1782, w_007_1783, w_007_1784, w_007_1785, w_007_1786, w_007_1787, w_007_1788, w_007_1789, w_007_1790, w_007_1791, w_007_1792, w_007_1793, w_007_1794, w_007_1795, w_007_1796, w_007_1797, w_007_1798, w_007_1799, w_007_1800, w_007_1801, w_007_1802, w_007_1803, w_007_1804, w_007_1805, w_007_1806, w_007_1807, w_007_1808, w_007_1809, w_007_1810, w_007_1811, w_007_1812, w_007_1813, w_007_1814, w_007_1815, w_007_1816, w_007_1817, w_007_1818, w_007_1819, w_007_1820, w_007_1821, w_007_1822, w_007_1823, w_007_1824, w_007_1825, w_007_1826, w_007_1827, w_007_1828, w_007_1829, w_007_1830, w_007_1831, w_007_1832, w_007_1833, w_007_1834, w_007_1835, w_007_1836, w_007_1837, w_007_1838, w_007_1839, w_007_1840, w_007_1841, w_007_1842, w_007_1843, w_007_1844, w_007_1845, w_007_1846, w_007_1847, w_007_1848, w_007_1849, w_007_1850, w_007_1851, w_007_1852;
  wire w_008_000, w_008_001, w_008_002, w_008_004, w_008_005, w_008_006, w_008_007, w_008_008, w_008_009, w_008_010, w_008_011, w_008_012, w_008_013, w_008_014, w_008_015, w_008_016, w_008_017, w_008_018, w_008_019, w_008_020, w_008_021, w_008_022, w_008_023, w_008_024, w_008_025, w_008_026, w_008_027, w_008_028, w_008_029, w_008_030, w_008_031, w_008_032, w_008_033, w_008_034, w_008_035, w_008_036, w_008_037, w_008_038, w_008_039, w_008_040, w_008_041, w_008_042, w_008_043, w_008_044, w_008_045, w_008_046, w_008_047, w_008_048, w_008_049, w_008_050, w_008_052, w_008_053, w_008_054, w_008_055, w_008_056, w_008_057, w_008_058, w_008_059, w_008_060, w_008_061, w_008_062, w_008_063, w_008_064, w_008_066, w_008_067, w_008_068, w_008_069, w_008_070, w_008_071, w_008_072, w_008_073, w_008_074, w_008_075, w_008_076, w_008_077, w_008_078, w_008_080, w_008_081, w_008_082, w_008_083, w_008_084, w_008_085, w_008_086, w_008_087, w_008_088, w_008_089, w_008_090, w_008_091, w_008_092, w_008_093, w_008_094, w_008_095, w_008_096, w_008_097, w_008_098, w_008_099, w_008_100, w_008_102, w_008_103, w_008_104, w_008_105, w_008_106, w_008_107, w_008_108, w_008_109, w_008_110, w_008_111, w_008_112, w_008_113, w_008_114, w_008_115, w_008_116, w_008_117, w_008_118, w_008_119, w_008_120, w_008_121, w_008_122, w_008_123, w_008_124, w_008_125, w_008_126, w_008_127, w_008_128, w_008_129, w_008_130, w_008_131, w_008_132, w_008_133, w_008_134, w_008_135, w_008_136, w_008_137, w_008_138, w_008_139, w_008_140, w_008_141, w_008_142, w_008_143, w_008_144, w_008_145, w_008_146, w_008_147, w_008_148, w_008_149, w_008_150, w_008_151, w_008_152, w_008_153, w_008_154, w_008_155, w_008_156, w_008_157, w_008_158, w_008_159, w_008_160, w_008_161, w_008_162, w_008_163, w_008_164, w_008_165, w_008_166, w_008_167, w_008_170, w_008_171, w_008_172, w_008_173, w_008_174, w_008_175, w_008_176, w_008_177, w_008_178, w_008_179, w_008_180, w_008_181, w_008_182, w_008_183, w_008_184, w_008_185, w_008_186, w_008_187, w_008_188, w_008_189, w_008_190, w_008_191, w_008_193, w_008_194, w_008_195, w_008_196, w_008_197, w_008_198, w_008_199, w_008_200, w_008_201, w_008_202, w_008_203, w_008_204, w_008_205, w_008_206, w_008_208, w_008_209, w_008_210, w_008_211, w_008_212, w_008_213, w_008_214, w_008_215, w_008_216, w_008_217, w_008_218, w_008_219, w_008_220, w_008_221, w_008_222, w_008_223, w_008_224, w_008_225, w_008_226, w_008_227, w_008_228, w_008_229, w_008_230, w_008_231, w_008_232, w_008_233, w_008_234, w_008_235, w_008_236, w_008_237, w_008_238, w_008_239, w_008_240, w_008_241, w_008_242, w_008_243, w_008_244, w_008_245, w_008_246, w_008_247, w_008_248, w_008_249, w_008_250, w_008_251, w_008_252, w_008_253, w_008_254, w_008_255, w_008_256, w_008_257, w_008_258, w_008_259, w_008_260, w_008_261, w_008_262, w_008_263, w_008_264, w_008_265, w_008_266, w_008_267, w_008_268, w_008_269, w_008_270, w_008_271, w_008_272, w_008_273, w_008_274, w_008_275, w_008_276, w_008_277, w_008_278, w_008_279, w_008_280, w_008_281, w_008_282, w_008_283, w_008_284, w_008_285, w_008_286, w_008_287, w_008_288, w_008_289, w_008_290, w_008_291, w_008_292, w_008_293, w_008_294, w_008_295, w_008_296, w_008_297, w_008_298, w_008_299, w_008_300, w_008_301, w_008_302, w_008_303, w_008_304, w_008_305, w_008_306, w_008_307, w_008_308, w_008_309, w_008_310, w_008_311, w_008_312, w_008_313, w_008_314, w_008_315, w_008_316, w_008_317, w_008_318, w_008_319, w_008_320, w_008_321, w_008_322, w_008_323, w_008_324, w_008_325, w_008_327, w_008_328, w_008_329, w_008_330, w_008_331, w_008_332, w_008_333, w_008_335, w_008_336, w_008_337, w_008_338, w_008_339, w_008_340, w_008_341, w_008_342, w_008_343, w_008_344, w_008_345, w_008_346, w_008_347, w_008_349, w_008_350, w_008_351, w_008_352, w_008_353, w_008_355, w_008_356, w_008_357, w_008_358, w_008_359, w_008_360, w_008_361, w_008_362, w_008_363, w_008_364, w_008_365, w_008_366, w_008_367, w_008_368, w_008_369, w_008_370, w_008_371, w_008_373, w_008_374, w_008_375, w_008_376, w_008_377, w_008_378, w_008_379, w_008_380, w_008_382, w_008_383, w_008_384, w_008_385, w_008_386, w_008_387, w_008_388, w_008_389, w_008_390, w_008_391, w_008_392, w_008_393, w_008_394, w_008_395, w_008_396, w_008_397, w_008_398, w_008_399, w_008_400, w_008_401, w_008_402, w_008_403, w_008_404, w_008_405, w_008_406, w_008_407, w_008_408, w_008_409, w_008_410, w_008_411, w_008_412, w_008_413, w_008_414, w_008_415, w_008_416, w_008_417, w_008_418, w_008_419, w_008_420, w_008_421, w_008_423, w_008_424, w_008_425, w_008_426, w_008_427, w_008_428, w_008_429, w_008_430, w_008_431, w_008_432, w_008_433, w_008_434, w_008_435, w_008_436, w_008_437, w_008_438, w_008_439, w_008_440, w_008_441, w_008_442, w_008_443, w_008_444, w_008_445, w_008_446, w_008_447, w_008_449, w_008_450, w_008_451, w_008_452, w_008_454, w_008_455, w_008_456, w_008_457, w_008_458, w_008_459, w_008_460, w_008_461, w_008_462, w_008_463, w_008_464, w_008_465, w_008_466, w_008_467, w_008_468, w_008_469, w_008_470, w_008_471, w_008_472, w_008_473, w_008_474, w_008_475, w_008_476, w_008_477, w_008_478, w_008_479, w_008_480, w_008_481, w_008_482, w_008_483, w_008_484, w_008_485, w_008_486, w_008_487, w_008_488, w_008_489, w_008_490, w_008_491, w_008_492, w_008_493, w_008_494, w_008_495, w_008_496, w_008_497, w_008_498, w_008_499, w_008_500, w_008_501, w_008_502, w_008_503, w_008_504, w_008_505, w_008_506, w_008_507, w_008_508, w_008_509, w_008_510, w_008_512, w_008_513, w_008_514, w_008_515, w_008_516, w_008_517, w_008_518, w_008_519, w_008_520, w_008_521, w_008_522, w_008_524, w_008_525, w_008_526, w_008_527, w_008_528, w_008_529, w_008_530, w_008_531, w_008_532, w_008_533, w_008_534, w_008_535, w_008_536, w_008_537, w_008_538, w_008_539, w_008_540, w_008_541, w_008_542, w_008_543, w_008_544, w_008_545, w_008_546, w_008_547, w_008_548, w_008_549, w_008_550, w_008_551, w_008_552, w_008_554, w_008_555, w_008_556, w_008_557, w_008_558, w_008_559, w_008_560, w_008_561, w_008_562, w_008_563, w_008_564, w_008_565, w_008_566, w_008_567, w_008_568, w_008_569, w_008_571, w_008_572, w_008_573, w_008_574, w_008_575, w_008_576, w_008_577, w_008_578, w_008_579, w_008_580, w_008_581, w_008_582, w_008_583, w_008_584, w_008_585, w_008_586, w_008_587, w_008_588, w_008_589, w_008_590, w_008_592, w_008_593, w_008_594, w_008_595, w_008_596, w_008_597, w_008_598, w_008_599, w_008_600, w_008_601, w_008_602, w_008_603, w_008_604, w_008_605, w_008_606, w_008_607, w_008_608, w_008_609, w_008_610, w_008_611, w_008_612, w_008_613, w_008_614, w_008_615, w_008_616, w_008_617, w_008_618, w_008_619, w_008_620, w_008_621, w_008_622, w_008_623, w_008_624, w_008_625, w_008_626, w_008_627, w_008_628, w_008_629, w_008_630, w_008_631, w_008_632, w_008_633, w_008_634, w_008_635, w_008_636, w_008_638, w_008_639, w_008_640, w_008_641, w_008_642, w_008_643, w_008_644, w_008_645, w_008_646, w_008_647, w_008_648, w_008_649, w_008_650, w_008_651, w_008_652, w_008_653, w_008_654, w_008_655, w_008_656, w_008_657, w_008_658, w_008_659, w_008_660, w_008_661, w_008_662, w_008_663, w_008_664, w_008_665, w_008_666, w_008_667, w_008_668, w_008_669, w_008_670, w_008_671, w_008_672, w_008_673, w_008_674, w_008_675, w_008_676, w_008_677, w_008_678, w_008_679, w_008_680, w_008_681, w_008_682, w_008_683, w_008_684, w_008_685, w_008_686, w_008_687, w_008_688, w_008_689, w_008_690, w_008_691, w_008_692, w_008_693, w_008_694, w_008_695, w_008_696, w_008_697, w_008_698, w_008_699, w_008_700, w_008_701, w_008_703, w_008_704, w_008_705, w_008_706, w_008_707, w_008_708, w_008_709, w_008_710, w_008_712, w_008_713, w_008_714, w_008_715, w_008_716, w_008_717, w_008_718, w_008_719, w_008_720, w_008_721, w_008_722, w_008_723, w_008_724, w_008_725, w_008_726, w_008_727, w_008_728, w_008_729, w_008_730, w_008_731, w_008_732, w_008_733, w_008_734, w_008_735, w_008_736, w_008_737, w_008_738, w_008_740, w_008_741, w_008_742, w_008_743, w_008_744, w_008_745, w_008_746, w_008_747, w_008_748, w_008_749, w_008_750, w_008_751, w_008_752, w_008_753, w_008_754, w_008_755, w_008_756, w_008_757, w_008_758, w_008_759, w_008_760, w_008_761, w_008_762, w_008_763, w_008_764, w_008_765, w_008_766, w_008_767, w_008_768, w_008_769, w_008_770, w_008_771, w_008_772, w_008_773, w_008_774, w_008_775, w_008_776, w_008_777, w_008_778, w_008_779, w_008_780, w_008_781, w_008_782, w_008_783, w_008_784, w_008_785, w_008_786, w_008_788, w_008_789, w_008_790, w_008_791, w_008_792, w_008_793, w_008_794, w_008_795, w_008_796, w_008_797, w_008_798, w_008_799, w_008_800, w_008_801, w_008_802, w_008_803, w_008_804, w_008_805, w_008_806, w_008_807, w_008_808, w_008_809, w_008_810, w_008_811, w_008_812, w_008_813, w_008_814, w_008_815, w_008_816, w_008_817, w_008_818, w_008_819, w_008_820, w_008_821, w_008_822, w_008_823, w_008_824, w_008_825, w_008_827, w_008_829, w_008_830, w_008_831, w_008_833, w_008_834, w_008_835, w_008_836, w_008_837, w_008_838, w_008_839, w_008_840, w_008_841, w_008_842, w_008_843, w_008_844, w_008_845, w_008_846, w_008_847, w_008_848, w_008_849, w_008_850, w_008_851, w_008_852, w_008_853, w_008_854, w_008_855, w_008_856, w_008_857, w_008_858, w_008_859, w_008_860, w_008_861, w_008_862, w_008_863, w_008_864, w_008_865, w_008_866, w_008_867, w_008_868, w_008_869, w_008_870, w_008_871, w_008_872, w_008_873, w_008_874, w_008_875, w_008_876, w_008_877, w_008_878, w_008_879, w_008_880, w_008_881, w_008_882, w_008_883, w_008_884, w_008_885, w_008_886, w_008_887, w_008_888, w_008_889, w_008_890, w_008_891, w_008_894, w_008_895, w_008_896, w_008_897, w_008_898, w_008_899, w_008_900, w_008_901, w_008_902, w_008_903, w_008_904, w_008_905, w_008_907, w_008_908, w_008_909, w_008_910, w_008_911, w_008_912, w_008_913, w_008_914, w_008_915, w_008_916, w_008_917, w_008_919, w_008_920, w_008_921, w_008_922, w_008_923, w_008_924, w_008_925, w_008_926, w_008_927, w_008_928, w_008_929, w_008_930, w_008_931, w_008_932, w_008_933, w_008_934, w_008_935, w_008_936, w_008_937, w_008_938, w_008_939, w_008_941, w_008_942, w_008_943, w_008_944, w_008_945, w_008_946, w_008_947, w_008_948, w_008_949, w_008_950, w_008_951, w_008_952, w_008_953, w_008_954, w_008_955, w_008_956, w_008_957, w_008_958, w_008_959, w_008_960, w_008_962, w_008_963, w_008_964, w_008_965, w_008_966, w_008_967, w_008_968, w_008_969, w_008_970, w_008_971, w_008_972, w_008_973, w_008_976, w_008_977, w_008_978, w_008_979, w_008_980, w_008_981, w_008_982, w_008_984, w_008_985, w_008_986, w_008_987, w_008_988, w_008_989, w_008_990, w_008_991, w_008_992, w_008_993, w_008_994, w_008_995, w_008_996, w_008_997, w_008_999, w_008_1000, w_008_1001, w_008_1002, w_008_1003, w_008_1004, w_008_1005, w_008_1006, w_008_1007, w_008_1008, w_008_1009, w_008_1010, w_008_1011, w_008_1013, w_008_1014, w_008_1015, w_008_1016, w_008_1017, w_008_1018, w_008_1019, w_008_1020, w_008_1021, w_008_1022, w_008_1024, w_008_1025, w_008_1026, w_008_1027, w_008_1028, w_008_1030, w_008_1031, w_008_1032, w_008_1033, w_008_1034, w_008_1035, w_008_1036, w_008_1037, w_008_1038, w_008_1039, w_008_1040, w_008_1041, w_008_1042, w_008_1043, w_008_1044, w_008_1045, w_008_1046, w_008_1047, w_008_1048, w_008_1049, w_008_1050, w_008_1051, w_008_1052, w_008_1053, w_008_1054, w_008_1055, w_008_1056, w_008_1057, w_008_1058, w_008_1059, w_008_1060, w_008_1061, w_008_1062, w_008_1063, w_008_1064, w_008_1065, w_008_1066, w_008_1067, w_008_1068, w_008_1069, w_008_1071, w_008_1072, w_008_1073, w_008_1074, w_008_1075, w_008_1076, w_008_1077, w_008_1078, w_008_1079, w_008_1080, w_008_1081, w_008_1082, w_008_1083, w_008_1084, w_008_1085, w_008_1086, w_008_1087, w_008_1088, w_008_1089, w_008_1090, w_008_1091, w_008_1092, w_008_1093, w_008_1094, w_008_1095, w_008_1096, w_008_1097, w_008_1098, w_008_1099, w_008_1100, w_008_1101, w_008_1102, w_008_1103, w_008_1104, w_008_1105, w_008_1106, w_008_1107, w_008_1108, w_008_1109, w_008_1110, w_008_1111, w_008_1112, w_008_1113, w_008_1114, w_008_1115, w_008_1116, w_008_1117, w_008_1118, w_008_1120, w_008_1121, w_008_1122, w_008_1123, w_008_1124, w_008_1125, w_008_1126, w_008_1127, w_008_1128, w_008_1129, w_008_1130, w_008_1131, w_008_1132, w_008_1133, w_008_1134, w_008_1135, w_008_1136, w_008_1137, w_008_1138, w_008_1139, w_008_1140, w_008_1141, w_008_1142, w_008_1143, w_008_1144, w_008_1145, w_008_1146, w_008_1147, w_008_1148, w_008_1149, w_008_1150, w_008_1151, w_008_1152, w_008_1153, w_008_1154, w_008_1155, w_008_1156, w_008_1157, w_008_1158, w_008_1159, w_008_1160, w_008_1161, w_008_1162, w_008_1163, w_008_1164, w_008_1166, w_008_1167, w_008_1168, w_008_1169, w_008_1170, w_008_1171, w_008_1172, w_008_1173, w_008_1174, w_008_1175, w_008_1176, w_008_1177, w_008_1178, w_008_1179, w_008_1180, w_008_1181, w_008_1182, w_008_1183, w_008_1184, w_008_1185, w_008_1186, w_008_1187, w_008_1188, w_008_1189, w_008_1190, w_008_1191, w_008_1192, w_008_1193, w_008_1194, w_008_1195, w_008_1196, w_008_1197, w_008_1198, w_008_1199, w_008_1200, w_008_1201, w_008_1202, w_008_1203, w_008_1204, w_008_1205, w_008_1206, w_008_1207, w_008_1208, w_008_1209, w_008_1210, w_008_1212, w_008_1213, w_008_1214, w_008_1215, w_008_1216, w_008_1217, w_008_1218, w_008_1219, w_008_1220, w_008_1221, w_008_1222, w_008_1223, w_008_1224, w_008_1225, w_008_1226, w_008_1227, w_008_1228, w_008_1229, w_008_1230, w_008_1231, w_008_1232, w_008_1233, w_008_1234, w_008_1235, w_008_1236, w_008_1237, w_008_1238, w_008_1239, w_008_1240, w_008_1241, w_008_1242, w_008_1243, w_008_1244, w_008_1245, w_008_1246, w_008_1247, w_008_1248, w_008_1249, w_008_1250, w_008_1251, w_008_1252, w_008_1253, w_008_1254, w_008_1255, w_008_1256, w_008_1257, w_008_1258, w_008_1259, w_008_1260, w_008_1261, w_008_1262, w_008_1263, w_008_1264, w_008_1265, w_008_1267, w_008_1268, w_008_1271, w_008_1272, w_008_1273, w_008_1274, w_008_1275, w_008_1276, w_008_1277, w_008_1278, w_008_1279, w_008_1280, w_008_1281, w_008_1282, w_008_1283, w_008_1284, w_008_1285, w_008_1286, w_008_1287, w_008_1288, w_008_1289, w_008_1290, w_008_1291, w_008_1292, w_008_1293, w_008_1294, w_008_1295, w_008_1296, w_008_1297, w_008_1298, w_008_1299, w_008_1300, w_008_1301, w_008_1302, w_008_1303, w_008_1304, w_008_1305, w_008_1307, w_008_1308, w_008_1309, w_008_1310, w_008_1312, w_008_1313, w_008_1314, w_008_1315, w_008_1316, w_008_1317, w_008_1318, w_008_1319, w_008_1320, w_008_1321, w_008_1322, w_008_1323, w_008_1324, w_008_1325, w_008_1326, w_008_1327, w_008_1328, w_008_1329, w_008_1330, w_008_1331, w_008_1332, w_008_1333, w_008_1334, w_008_1335, w_008_1336, w_008_1337, w_008_1338, w_008_1339, w_008_1340, w_008_1341, w_008_1342, w_008_1343, w_008_1344, w_008_1345, w_008_1346, w_008_1347, w_008_1348, w_008_1349, w_008_1350, w_008_1351, w_008_1352, w_008_1353, w_008_1354, w_008_1355, w_008_1356, w_008_1357, w_008_1358, w_008_1359, w_008_1360, w_008_1361, w_008_1362, w_008_1363, w_008_1364, w_008_1365, w_008_1366, w_008_1367, w_008_1368, w_008_1369, w_008_1370, w_008_1371, w_008_1372, w_008_1373, w_008_1374, w_008_1375, w_008_1376, w_008_1377, w_008_1378, w_008_1379, w_008_1380, w_008_1381, w_008_1382, w_008_1383, w_008_1384, w_008_1385, w_008_1386, w_008_1387, w_008_1388, w_008_1389, w_008_1390, w_008_1391, w_008_1392, w_008_1393, w_008_1394, w_008_1395, w_008_1396, w_008_1397, w_008_1398, w_008_1399, w_008_1400, w_008_1401, w_008_1402, w_008_1404, w_008_1405, w_008_1406, w_008_1407, w_008_1408, w_008_1409, w_008_1410, w_008_1411, w_008_1412, w_008_1413, w_008_1415, w_008_1416, w_008_1417, w_008_1418, w_008_1419, w_008_1420, w_008_1421, w_008_1422, w_008_1423, w_008_1424, w_008_1425, w_008_1426, w_008_1427, w_008_1428, w_008_1429, w_008_1430, w_008_1431, w_008_1432, w_008_1433, w_008_1434, w_008_1435, w_008_1436, w_008_1437, w_008_1438, w_008_1439, w_008_1440, w_008_1441, w_008_1442, w_008_1443, w_008_1444, w_008_1445, w_008_1446, w_008_1447, w_008_1448, w_008_1449, w_008_1450, w_008_1451, w_008_1452, w_008_1453, w_008_1454, w_008_1455, w_008_1456, w_008_1457, w_008_1458, w_008_1459, w_008_1460, w_008_1461, w_008_1462, w_008_1463, w_008_1464, w_008_1465, w_008_1466, w_008_1467, w_008_1468, w_008_1469, w_008_1470, w_008_1471, w_008_1472, w_008_1473, w_008_1474, w_008_1475, w_008_1476, w_008_1477, w_008_1478, w_008_1479, w_008_1480, w_008_1481, w_008_1482, w_008_1483, w_008_1484, w_008_1485, w_008_1486, w_008_1487, w_008_1488, w_008_1489, w_008_1490, w_008_1491, w_008_1492, w_008_1493, w_008_1494, w_008_1495, w_008_1496, w_008_1497, w_008_1498, w_008_1499, w_008_1500, w_008_1501, w_008_1503, w_008_1504, w_008_1505, w_008_1506, w_008_1507, w_008_1509, w_008_1510, w_008_1511, w_008_1512, w_008_1513, w_008_1514, w_008_1515, w_008_1516, w_008_1517, w_008_1518, w_008_1519, w_008_1520, w_008_1521, w_008_1523, w_008_1524, w_008_1525, w_008_1526, w_008_1527, w_008_1528, w_008_1529, w_008_1530, w_008_1532, w_008_1533, w_008_1534, w_008_1535, w_008_1536, w_008_1537, w_008_1538, w_008_1539, w_008_1540, w_008_1541, w_008_1542, w_008_1543, w_008_1544, w_008_1545, w_008_1546, w_008_1547, w_008_1548, w_008_1549, w_008_1550, w_008_1551, w_008_1552, w_008_1553, w_008_1554, w_008_1555, w_008_1556, w_008_1557, w_008_1558, w_008_1559, w_008_1560, w_008_1561, w_008_1562, w_008_1563, w_008_1564, w_008_1565, w_008_1566, w_008_1567, w_008_1568, w_008_1569, w_008_1570, w_008_1571, w_008_1572, w_008_1573, w_008_1574, w_008_1575, w_008_1576, w_008_1577, w_008_1578, w_008_1579, w_008_1580, w_008_1581, w_008_1582, w_008_1583, w_008_1584, w_008_1585, w_008_1586, w_008_1587, w_008_1588, w_008_1589, w_008_1590, w_008_1591, w_008_1592, w_008_1593, w_008_1594, w_008_1595, w_008_1596, w_008_1597, w_008_1598, w_008_1599, w_008_1600, w_008_1601, w_008_1602, w_008_1603, w_008_1604, w_008_1605, w_008_1606, w_008_1607, w_008_1608, w_008_1609, w_008_1610, w_008_1611, w_008_1612, w_008_1613, w_008_1614, w_008_1615, w_008_1616, w_008_1617, w_008_1618, w_008_1620, w_008_1621, w_008_1622, w_008_1623, w_008_1624, w_008_1625, w_008_1626, w_008_1627, w_008_1628, w_008_1629, w_008_1630, w_008_1631, w_008_1632, w_008_1633, w_008_1634, w_008_1635, w_008_1636, w_008_1637, w_008_1638, w_008_1639, w_008_1640, w_008_1641, w_008_1643, w_008_1644, w_008_1645, w_008_1646, w_008_1647, w_008_1648, w_008_1649, w_008_1650, w_008_1651, w_008_1652, w_008_1653, w_008_1654, w_008_1655, w_008_1656, w_008_1657, w_008_1658, w_008_1659, w_008_1660, w_008_1661, w_008_1662, w_008_1663, w_008_1664, w_008_1665, w_008_1666, w_008_1667, w_008_1668, w_008_1669, w_008_1670, w_008_1671, w_008_1672, w_008_1673, w_008_1674, w_008_1675, w_008_1676, w_008_1677, w_008_1678, w_008_1679, w_008_1680, w_008_1681, w_008_1682, w_008_1683, w_008_1685, w_008_1686, w_008_1687, w_008_1688, w_008_1689, w_008_1690, w_008_1691, w_008_1692, w_008_1693, w_008_1694, w_008_1695, w_008_1696, w_008_1697, w_008_1698, w_008_1699, w_008_1700, w_008_1701, w_008_1702, w_008_1703, w_008_1704, w_008_1705, w_008_1706, w_008_1707, w_008_1708, w_008_1709, w_008_1710, w_008_1711, w_008_1712, w_008_1713, w_008_1714, w_008_1715, w_008_1716, w_008_1717, w_008_1718, w_008_1719, w_008_1720, w_008_1721, w_008_1722, w_008_1723, w_008_1724, w_008_1725, w_008_1726, w_008_1727, w_008_1728, w_008_1729, w_008_1730, w_008_1731, w_008_1732, w_008_1733, w_008_1734, w_008_1735, w_008_1736, w_008_1738, w_008_1739, w_008_1740, w_008_1742, w_008_1743, w_008_1744, w_008_1745, w_008_1746, w_008_1747, w_008_1748, w_008_1749, w_008_1750, w_008_1751, w_008_1752, w_008_1753, w_008_1754, w_008_1755, w_008_1756, w_008_1757, w_008_1758, w_008_1759, w_008_1760, w_008_1761, w_008_1762, w_008_1763, w_008_1764, w_008_1765, w_008_1766, w_008_1767, w_008_1768, w_008_1769, w_008_1770, w_008_1771, w_008_1772, w_008_1773, w_008_1774, w_008_1775, w_008_1776, w_008_1777, w_008_1778, w_008_1779, w_008_1780, w_008_1781, w_008_1782, w_008_1783, w_008_1784, w_008_1785, w_008_1786, w_008_1787, w_008_1788, w_008_1789, w_008_1790, w_008_1791, w_008_1792, w_008_1793, w_008_1794, w_008_1795, w_008_1796, w_008_1797, w_008_1798, w_008_1799, w_008_1800, w_008_1801, w_008_1802, w_008_1803, w_008_1804, w_008_1805, w_008_1807, w_008_1808, w_008_1809, w_008_1810, w_008_1811, w_008_1812, w_008_1813, w_008_1815, w_008_1816, w_008_1817, w_008_1818, w_008_1819, w_008_1820, w_008_1821, w_008_1822, w_008_1823, w_008_1824, w_008_1825, w_008_1826, w_008_1827, w_008_1828, w_008_1829, w_008_1830, w_008_1831, w_008_1832, w_008_1833, w_008_1834, w_008_1835, w_008_1836, w_008_1837, w_008_1838, w_008_1839, w_008_1840, w_008_1841, w_008_1842, w_008_1843, w_008_1844, w_008_1845, w_008_1846, w_008_1847, w_008_1848, w_008_1849, w_008_1850, w_008_1851, w_008_1852, w_008_1853, w_008_1854, w_008_1855, w_008_1856, w_008_1857, w_008_1858, w_008_1859, w_008_1860, w_008_1861, w_008_1862, w_008_1863, w_008_1864, w_008_1865, w_008_1866, w_008_1867, w_008_1868, w_008_1869, w_008_1870, w_008_1871, w_008_1872, w_008_1873, w_008_1874, w_008_1875, w_008_1876, w_008_1877, w_008_1878, w_008_1879, w_008_1880, w_008_1881, w_008_1882, w_008_1883, w_008_1884, w_008_1885, w_008_1887, w_008_1888, w_008_1890, w_008_1891, w_008_1892, w_008_1893, w_008_1894, w_008_1895, w_008_1896, w_008_1897, w_008_1898, w_008_1900, w_008_1901, w_008_1903, w_008_1904, w_008_1906, w_008_1907, w_008_1908, w_008_1909, w_008_1910, w_008_1911, w_008_1913, w_008_1914, w_008_1915, w_008_1916, w_008_1917, w_008_1918, w_008_1919, w_008_1920, w_008_1921, w_008_1922, w_008_1923, w_008_1924, w_008_1925, w_008_1926, w_008_1927, w_008_1928, w_008_1929, w_008_1931, w_008_1932, w_008_1933, w_008_1934, w_008_1935, w_008_1936, w_008_1937, w_008_1938, w_008_1939, w_008_1940, w_008_1941, w_008_1942, w_008_1943, w_008_1944, w_008_1945, w_008_1946, w_008_1947, w_008_1948, w_008_1949, w_008_1950, w_008_1951, w_008_1952, w_008_1953, w_008_1954, w_008_1955, w_008_1956, w_008_1957, w_008_1959, w_008_1960, w_008_1961, w_008_1962, w_008_1963, w_008_1964, w_008_1965, w_008_1966, w_008_1967, w_008_1968, w_008_1969, w_008_1970, w_008_1971, w_008_1972, w_008_1973, w_008_1974, w_008_1975, w_008_1976, w_008_1977, w_008_1978, w_008_1979, w_008_1980, w_008_1981, w_008_1982, w_008_1983, w_008_1984, w_008_1985, w_008_1986, w_008_1987, w_008_1988, w_008_1989, w_008_1990, w_008_1991, w_008_1992, w_008_1993, w_008_1994, w_008_1995, w_008_1996, w_008_1997, w_008_1998, w_008_1999, w_008_2000, w_008_2001, w_008_2002, w_008_2003, w_008_2004, w_008_2005, w_008_2006, w_008_2007, w_008_2008, w_008_2009, w_008_2010, w_008_2011, w_008_2012, w_008_2013, w_008_2014, w_008_2015, w_008_2016, w_008_2017, w_008_2018, w_008_2019, w_008_2020, w_008_2021, w_008_2022, w_008_2023, w_008_2024, w_008_2025, w_008_2026, w_008_2027, w_008_2028, w_008_2029, w_008_2030, w_008_2031, w_008_2032, w_008_2033, w_008_2034, w_008_2035, w_008_2036, w_008_2037, w_008_2038, w_008_2039, w_008_2040, w_008_2041, w_008_2042, w_008_2044, w_008_2045, w_008_2046, w_008_2047, w_008_2048, w_008_2049, w_008_2050, w_008_2051, w_008_2052, w_008_2053, w_008_2054, w_008_2055, w_008_2056, w_008_2057, w_008_2058, w_008_2059, w_008_2060, w_008_2061, w_008_2062, w_008_2063, w_008_2065, w_008_2066, w_008_2067, w_008_2068, w_008_2069, w_008_2070, w_008_2071, w_008_2072, w_008_2073, w_008_2074, w_008_2075, w_008_2076, w_008_2077, w_008_2078, w_008_2079, w_008_2080, w_008_2081, w_008_2082, w_008_2083, w_008_2084, w_008_2085, w_008_2086, w_008_2087, w_008_2088, w_008_2089, w_008_2090, w_008_2091, w_008_2092, w_008_2093, w_008_2094, w_008_2095, w_008_2096, w_008_2097, w_008_2098, w_008_2099, w_008_2100, w_008_2101, w_008_2102, w_008_2103, w_008_2104, w_008_2105, w_008_2106, w_008_2107, w_008_2108, w_008_2109, w_008_2110, w_008_2111, w_008_2112, w_008_2113, w_008_2114, w_008_2115, w_008_2116, w_008_2118, w_008_2119, w_008_2120, w_008_2121, w_008_2122, w_008_2123, w_008_2124, w_008_2125, w_008_2126, w_008_2127, w_008_2128, w_008_2129, w_008_2130, w_008_2131, w_008_2132, w_008_2133, w_008_2134, w_008_2135, w_008_2136, w_008_2137, w_008_2138, w_008_2139, w_008_2140, w_008_2141, w_008_2142, w_008_2143, w_008_2144, w_008_2145, w_008_2146, w_008_2147, w_008_2148, w_008_2149, w_008_2150, w_008_2151, w_008_2152, w_008_2153, w_008_2154, w_008_2155, w_008_2156, w_008_2157, w_008_2158, w_008_2159, w_008_2160, w_008_2161, w_008_2162, w_008_2163, w_008_2164, w_008_2165, w_008_2166, w_008_2167, w_008_2169, w_008_2170, w_008_2171, w_008_2172, w_008_2173, w_008_2174, w_008_2175, w_008_2176, w_008_2177, w_008_2178, w_008_2179, w_008_2180, w_008_2181, w_008_2182, w_008_2183, w_008_2184, w_008_2185, w_008_2186, w_008_2187, w_008_2188, w_008_2189, w_008_2190, w_008_2191, w_008_2192, w_008_2193, w_008_2194, w_008_2195, w_008_2196, w_008_2197, w_008_2198, w_008_2199, w_008_2200, w_008_2201, w_008_2202, w_008_2203, w_008_2204, w_008_2205, w_008_2206, w_008_2207, w_008_2208, w_008_2209, w_008_2210, w_008_2211, w_008_2212, w_008_2214, w_008_2215, w_008_2216, w_008_2217, w_008_2218, w_008_2219, w_008_2222, w_008_2223, w_008_2224, w_008_2225, w_008_2226, w_008_2227, w_008_2228, w_008_2229, w_008_2230, w_008_2231, w_008_2232, w_008_2233, w_008_2234, w_008_2235, w_008_2236, w_008_2237, w_008_2238, w_008_2239, w_008_2240, w_008_2241, w_008_2242, w_008_2243, w_008_2244, w_008_2245, w_008_2246, w_008_2247, w_008_2248, w_008_2249, w_008_2250, w_008_2251, w_008_2252, w_008_2253, w_008_2254, w_008_2255, w_008_2256, w_008_2257, w_008_2258, w_008_2259, w_008_2260, w_008_2261, w_008_2262, w_008_2263, w_008_2264, w_008_2265, w_008_2266, w_008_2267, w_008_2268, w_008_2269, w_008_2270, w_008_2271, w_008_2272, w_008_2273, w_008_2274, w_008_2275, w_008_2276, w_008_2277, w_008_2278, w_008_2279, w_008_2280, w_008_2281, w_008_2282, w_008_2283, w_008_2284, w_008_2286, w_008_2287, w_008_2288, w_008_2289, w_008_2290, w_008_2291, w_008_2292, w_008_2293, w_008_2294, w_008_2295, w_008_2296, w_008_2297, w_008_2298, w_008_2299, w_008_2300, w_008_2301, w_008_2302, w_008_2303, w_008_2304, w_008_2305, w_008_2306, w_008_2307, w_008_2308, w_008_2310, w_008_2311, w_008_2312, w_008_2313, w_008_2315, w_008_2316, w_008_2317, w_008_2318, w_008_2319, w_008_2320, w_008_2321, w_008_2322, w_008_2323, w_008_2324, w_008_2325, w_008_2326, w_008_2327, w_008_2328, w_008_2329, w_008_2330, w_008_2331, w_008_2332, w_008_2333, w_008_2334, w_008_2335, w_008_2336, w_008_2337, w_008_2338, w_008_2339, w_008_2340, w_008_2341, w_008_2343, w_008_2344, w_008_2345, w_008_2346, w_008_2347, w_008_2348, w_008_2349, w_008_2350, w_008_2351, w_008_2352, w_008_2353, w_008_2354, w_008_2355, w_008_2357, w_008_2358, w_008_2359, w_008_2360, w_008_2361, w_008_2362, w_008_2363, w_008_2364, w_008_2365, w_008_2366, w_008_2367, w_008_2368, w_008_2369, w_008_2370, w_008_2371, w_008_2372, w_008_2373, w_008_2374, w_008_2375, w_008_2376, w_008_2377, w_008_2378, w_008_2379, w_008_2380, w_008_2382, w_008_2384, w_008_2385, w_008_2386, w_008_2387, w_008_2388, w_008_2389, w_008_2390, w_008_2392, w_008_2393, w_008_2394, w_008_2395, w_008_2396, w_008_2397, w_008_2398, w_008_2399, w_008_2400, w_008_2401, w_008_2402, w_008_2403, w_008_2404, w_008_2405, w_008_2406, w_008_2407, w_008_2409, w_008_2410, w_008_2411, w_008_2412, w_008_2413, w_008_2414, w_008_2415, w_008_2416, w_008_2417, w_008_2418, w_008_2419, w_008_2420, w_008_2421, w_008_2422, w_008_2423, w_008_2424, w_008_2425, w_008_2426, w_008_2427, w_008_2428, w_008_2429, w_008_2430, w_008_2432, w_008_2433, w_008_2434, w_008_2435, w_008_2436, w_008_2437, w_008_2438, w_008_2440, w_008_2441, w_008_2442, w_008_2443, w_008_2444, w_008_2446, w_008_2447, w_008_2448, w_008_2449, w_008_2450, w_008_2451, w_008_2452, w_008_2453, w_008_2454, w_008_2455, w_008_2456, w_008_2457, w_008_2458, w_008_2459, w_008_2460, w_008_2461, w_008_2462, w_008_2463, w_008_2464, w_008_2465, w_008_2466, w_008_2467, w_008_2468, w_008_2469, w_008_2470, w_008_2471, w_008_2472, w_008_2473, w_008_2474, w_008_2475, w_008_2476, w_008_2477, w_008_2478, w_008_2479, w_008_2480, w_008_2481, w_008_2482, w_008_2483, w_008_2484, w_008_2485, w_008_2486, w_008_2487, w_008_2488, w_008_2489, w_008_2490, w_008_2491, w_008_2492, w_008_2494, w_008_2495, w_008_2496, w_008_2497, w_008_2498, w_008_2499, w_008_2500, w_008_2501, w_008_2502, w_008_2503, w_008_2504, w_008_2505, w_008_2506, w_008_2507, w_008_2508, w_008_2509, w_008_2510, w_008_2511, w_008_2512, w_008_2513, w_008_2514, w_008_2516, w_008_2517, w_008_2518, w_008_2519, w_008_2520, w_008_2521, w_008_2522, w_008_2523, w_008_2524, w_008_2525, w_008_2526, w_008_2527, w_008_2528, w_008_2529, w_008_2530, w_008_2531, w_008_2532, w_008_2533, w_008_2534, w_008_2535, w_008_2536, w_008_2537, w_008_2538, w_008_2539, w_008_2540, w_008_2541, w_008_2542, w_008_2543, w_008_2544, w_008_2545, w_008_2546, w_008_2547, w_008_2548, w_008_2550, w_008_2552, w_008_2553, w_008_2554, w_008_2555, w_008_2556, w_008_2557, w_008_2558, w_008_2559, w_008_2560, w_008_2561, w_008_2562, w_008_2563, w_008_2564, w_008_2565, w_008_2567, w_008_2568, w_008_2569, w_008_2570, w_008_2571, w_008_2572, w_008_2573, w_008_2574, w_008_2575, w_008_2576, w_008_2577, w_008_2578, w_008_2579, w_008_2580, w_008_2581, w_008_2582, w_008_2583, w_008_2584, w_008_2585, w_008_2586, w_008_2587, w_008_2588, w_008_2589, w_008_2590, w_008_2591, w_008_2592, w_008_2593, w_008_2594, w_008_2595, w_008_2596, w_008_2598, w_008_2599, w_008_2600, w_008_2601, w_008_2602, w_008_2603, w_008_2604, w_008_2605, w_008_2606, w_008_2608, w_008_2609, w_008_2610, w_008_2611, w_008_2612, w_008_2613, w_008_2614, w_008_2615, w_008_2616, w_008_2618, w_008_2619, w_008_2620, w_008_2621, w_008_2622, w_008_2623, w_008_2624, w_008_2625, w_008_2626, w_008_2627, w_008_2629, w_008_2630, w_008_2631, w_008_2632, w_008_2633, w_008_2634, w_008_2635, w_008_2636, w_008_2637, w_008_2638, w_008_2640, w_008_2641, w_008_2642, w_008_2643, w_008_2644, w_008_2645, w_008_2646, w_008_2647, w_008_2648, w_008_2649, w_008_2650, w_008_2651, w_008_2653, w_008_2654, w_008_2655, w_008_2656, w_008_2657, w_008_2658, w_008_2659, w_008_2660, w_008_2661, w_008_2662, w_008_2663, w_008_2664, w_008_2665, w_008_2666, w_008_2667, w_008_2668, w_008_2669, w_008_2670, w_008_2671, w_008_2672, w_008_2673, w_008_2674, w_008_2675, w_008_2676, w_008_2677, w_008_2678, w_008_2679, w_008_2680, w_008_2681, w_008_2682, w_008_2683, w_008_2684, w_008_2685, w_008_2686, w_008_2687, w_008_2688, w_008_2689, w_008_2690, w_008_2691, w_008_2692, w_008_2693, w_008_2694, w_008_2695, w_008_2696, w_008_2697, w_008_2698, w_008_2699, w_008_2700, w_008_2701, w_008_2702, w_008_2703, w_008_2704, w_008_2705, w_008_2706, w_008_2707, w_008_2708, w_008_2709, w_008_2710, w_008_2711, w_008_2712, w_008_2713, w_008_2714, w_008_2715, w_008_2716, w_008_2717, w_008_2718, w_008_2719, w_008_2720, w_008_2721, w_008_2722, w_008_2723, w_008_2724, w_008_2725, w_008_2726, w_008_2727, w_008_2729, w_008_2730, w_008_2731, w_008_2732, w_008_2733, w_008_2734, w_008_2735, w_008_2736, w_008_2737, w_008_2738, w_008_2739, w_008_2740, w_008_2741, w_008_2742, w_008_2743, w_008_2744, w_008_2745, w_008_2746, w_008_2747, w_008_2748, w_008_2749, w_008_2750, w_008_2751, w_008_2752, w_008_2753, w_008_2754, w_008_2755, w_008_2756, w_008_2758, w_008_2759, w_008_2760, w_008_2761, w_008_2762, w_008_2763, w_008_2764, w_008_2766, w_008_2767, w_008_2768, w_008_2769, w_008_2770, w_008_2771, w_008_2772, w_008_2773, w_008_2774, w_008_2775, w_008_2776, w_008_2777, w_008_2779, w_008_2780, w_008_2781, w_008_2782, w_008_2784, w_008_2785, w_008_2786, w_008_2787, w_008_2788, w_008_2790, w_008_2791, w_008_2792, w_008_2793, w_008_2794, w_008_2795, w_008_2796, w_008_2797, w_008_2798, w_008_2799, w_008_2800, w_008_2801, w_008_2802, w_008_2803, w_008_2804, w_008_2805, w_008_2806, w_008_2807, w_008_2808, w_008_2809, w_008_2810, w_008_2811, w_008_2812, w_008_2813, w_008_2814, w_008_2815, w_008_2816, w_008_2817, w_008_2818, w_008_2819, w_008_2820, w_008_2822, w_008_2823, w_008_2824, w_008_2825, w_008_2827, w_008_2828, w_008_2829, w_008_2830, w_008_2832, w_008_2833, w_008_2834, w_008_2835, w_008_2836, w_008_2837, w_008_2838, w_008_2839, w_008_2840, w_008_2841, w_008_2842, w_008_2843, w_008_2844, w_008_2845, w_008_2846, w_008_2847, w_008_2848, w_008_2849, w_008_2850, w_008_2851, w_008_2852, w_008_2853, w_008_2854, w_008_2855, w_008_2857, w_008_2858, w_008_2859, w_008_2860, w_008_2861, w_008_2862, w_008_2863, w_008_2864, w_008_2865, w_008_2866, w_008_2867, w_008_2868, w_008_2869, w_008_2870, w_008_2871, w_008_2873, w_008_2874, w_008_2875, w_008_2876, w_008_2877, w_008_2878, w_008_2880, w_008_2881, w_008_2882, w_008_2883, w_008_2884, w_008_2885, w_008_2886, w_008_2887, w_008_2888, w_008_2889, w_008_2890, w_008_2891, w_008_2892, w_008_2893, w_008_2894, w_008_2895, w_008_2896, w_008_2897, w_008_2898, w_008_2899, w_008_2900, w_008_2901, w_008_2902, w_008_2903, w_008_2904, w_008_2905, w_008_2906, w_008_2907, w_008_2908, w_008_2909, w_008_2910, w_008_2911, w_008_2912, w_008_2913, w_008_2914, w_008_2915, w_008_2916, w_008_2917, w_008_2918, w_008_2919, w_008_2920, w_008_2921, w_008_2923, w_008_2924, w_008_2925, w_008_2926, w_008_2927, w_008_2928, w_008_2929, w_008_2932, w_008_2934, w_008_2935, w_008_2936, w_008_2937, w_008_2938, w_008_2939, w_008_2940, w_008_2941, w_008_2942, w_008_2944, w_008_2945, w_008_2946, w_008_2947, w_008_2948, w_008_2949, w_008_2950, w_008_2951, w_008_2952, w_008_2953, w_008_2954, w_008_2955, w_008_2956, w_008_2957, w_008_2958, w_008_2961, w_008_2962, w_008_2963, w_008_2964, w_008_2965, w_008_2966, w_008_2967, w_008_2968, w_008_2969, w_008_2970, w_008_2971, w_008_2972, w_008_2973, w_008_2974, w_008_2975, w_008_2976, w_008_2977, w_008_2978, w_008_2979, w_008_2980, w_008_2981, w_008_2982, w_008_2983, w_008_2984, w_008_2985, w_008_2986, w_008_2987, w_008_2988, w_008_2989, w_008_2990, w_008_2991, w_008_2992, w_008_2993, w_008_2994, w_008_2995, w_008_2996, w_008_2997, w_008_2998, w_008_2999, w_008_3000, w_008_3001, w_008_3002, w_008_3003, w_008_3004, w_008_3005, w_008_3006, w_008_3008, w_008_3009, w_008_3010, w_008_3011, w_008_3012, w_008_3013, w_008_3014, w_008_3015, w_008_3016, w_008_3017, w_008_3018, w_008_3019, w_008_3020, w_008_3021, w_008_3022, w_008_3023, w_008_3024, w_008_3025, w_008_3026, w_008_3027, w_008_3028, w_008_3029, w_008_3030, w_008_3031, w_008_3032, w_008_3033, w_008_3034, w_008_3035, w_008_3036, w_008_3037, w_008_3038, w_008_3039, w_008_3040, w_008_3041, w_008_3042, w_008_3043, w_008_3044, w_008_3045, w_008_3046, w_008_3047, w_008_3048, w_008_3049, w_008_3050, w_008_3051, w_008_3052, w_008_3053, w_008_3054, w_008_3055, w_008_3056, w_008_3057, w_008_3058, w_008_3059, w_008_3060, w_008_3062, w_008_3063, w_008_3064, w_008_3065, w_008_3066, w_008_3067, w_008_3068, w_008_3069, w_008_3070, w_008_3071, w_008_3073, w_008_3074, w_008_3075, w_008_3076, w_008_3077, w_008_3078, w_008_3079, w_008_3080, w_008_3081, w_008_3083, w_008_3084, w_008_3085, w_008_3086, w_008_3087, w_008_3088, w_008_3089, w_008_3090, w_008_3091, w_008_3092, w_008_3093, w_008_3094, w_008_3096, w_008_3097, w_008_3098, w_008_3099, w_008_3100, w_008_3101, w_008_3102, w_008_3103, w_008_3104, w_008_3105, w_008_3106, w_008_3107, w_008_3108, w_008_3109, w_008_3110, w_008_3111, w_008_3112, w_008_3113, w_008_3114, w_008_3115, w_008_3116, w_008_3117, w_008_3118, w_008_3121, w_008_3122, w_008_3123, w_008_3124, w_008_3125, w_008_3126, w_008_3127, w_008_3128, w_008_3129, w_008_3130, w_008_3131, w_008_3132, w_008_3133, w_008_3134, w_008_3136, w_008_3137, w_008_3138, w_008_3139, w_008_3141, w_008_3142, w_008_3143, w_008_3144, w_008_3145, w_008_3146, w_008_3147, w_008_3148, w_008_3149, w_008_3150, w_008_3151, w_008_3152, w_008_3153, w_008_3154, w_008_3155, w_008_3156, w_008_3157, w_008_3158, w_008_3159, w_008_3160, w_008_3161, w_008_3162, w_008_3163, w_008_3164, w_008_3165, w_008_3166, w_008_3167, w_008_3168, w_008_3169, w_008_3170, w_008_3171, w_008_3172, w_008_3174, w_008_3175, w_008_3176, w_008_3177, w_008_3178, w_008_3179, w_008_3180, w_008_3181, w_008_3182, w_008_3183, w_008_3184, w_008_3186, w_008_3187, w_008_3188, w_008_3190, w_008_3191, w_008_3192, w_008_3193, w_008_3194, w_008_3195, w_008_3196, w_008_3197, w_008_3198, w_008_3199, w_008_3200, w_008_3201, w_008_3202, w_008_3203, w_008_3204, w_008_3205, w_008_3206, w_008_3207, w_008_3208, w_008_3209, w_008_3210, w_008_3211, w_008_3212, w_008_3213, w_008_3214, w_008_3215, w_008_3216, w_008_3217, w_008_3219, w_008_3220, w_008_3221, w_008_3222, w_008_3223, w_008_3224, w_008_3225, w_008_3226, w_008_3227, w_008_3228, w_008_3229, w_008_3230, w_008_3231, w_008_3232, w_008_3233, w_008_3234, w_008_3235, w_008_3236, w_008_3237, w_008_3238, w_008_3239, w_008_3240, w_008_3241, w_008_3242, w_008_3243, w_008_3244, w_008_3245, w_008_3246, w_008_3247, w_008_3248, w_008_3249, w_008_3250, w_008_3251, w_008_3252, w_008_3253, w_008_3254, w_008_3255, w_008_3256, w_008_3257, w_008_3258, w_008_3259, w_008_3260, w_008_3261, w_008_3262, w_008_3263, w_008_3264, w_008_3265, w_008_3266, w_008_3267, w_008_3268, w_008_3269, w_008_3270, w_008_3271, w_008_3272, w_008_3273, w_008_3274, w_008_3275, w_008_3276, w_008_3277, w_008_3278, w_008_3279, w_008_3280, w_008_3281, w_008_3282, w_008_3283, w_008_3284, w_008_3285, w_008_3286, w_008_3287, w_008_3288, w_008_3289, w_008_3290, w_008_3291, w_008_3292, w_008_3293, w_008_3294, w_008_3295, w_008_3296, w_008_3297, w_008_3298, w_008_3299, w_008_3300, w_008_3301, w_008_3302, w_008_3303, w_008_3304, w_008_3305, w_008_3306, w_008_3307, w_008_3308, w_008_3310, w_008_3311, w_008_3312, w_008_3313, w_008_3314, w_008_3315, w_008_3316, w_008_3317, w_008_3318, w_008_3319, w_008_3320, w_008_3321, w_008_3322, w_008_3323, w_008_3324, w_008_3325, w_008_3326, w_008_3327, w_008_3329, w_008_3330, w_008_3331, w_008_3332, w_008_3333, w_008_3334, w_008_3335, w_008_3336, w_008_3337, w_008_3338, w_008_3339, w_008_3340, w_008_3341, w_008_3342, w_008_3343, w_008_3344, w_008_3345, w_008_3346, w_008_3347, w_008_3348, w_008_3349, w_008_3350, w_008_3351, w_008_3352, w_008_3353, w_008_3354, w_008_3355, w_008_3356, w_008_3357, w_008_3358, w_008_3360, w_008_3361, w_008_3362, w_008_3363, w_008_3364, w_008_3365, w_008_3366, w_008_3367, w_008_3368, w_008_3369, w_008_3370, w_008_3371, w_008_3372, w_008_3373, w_008_3374, w_008_3375, w_008_3376, w_008_3377, w_008_3378, w_008_3379, w_008_3380, w_008_3381, w_008_3382, w_008_3383, w_008_3384, w_008_3385, w_008_3386, w_008_3387, w_008_3389, w_008_3390, w_008_3391, w_008_3392, w_008_3393, w_008_3394, w_008_3395, w_008_3396, w_008_3397, w_008_3398, w_008_3399, w_008_3400, w_008_3401, w_008_3402, w_008_3403, w_008_3404, w_008_3405, w_008_3406, w_008_3407, w_008_3408, w_008_3409, w_008_3410, w_008_3411, w_008_3412, w_008_3413, w_008_3414, w_008_3415, w_008_3416, w_008_3417, w_008_3418, w_008_3419, w_008_3420, w_008_3421, w_008_3422, w_008_3423, w_008_3424, w_008_3425, w_008_3426, w_008_3427, w_008_3428, w_008_3429, w_008_3430, w_008_3431, w_008_3432, w_008_3433, w_008_3434, w_008_3435, w_008_3436, w_008_3437, w_008_3438, w_008_3439, w_008_3441, w_008_3443, w_008_3444, w_008_3445, w_008_3446, w_008_3447, w_008_3448, w_008_3449, w_008_3450, w_008_3451, w_008_3452, w_008_3453, w_008_3454, w_008_3455, w_008_3456, w_008_3457, w_008_3458, w_008_3459, w_008_3460, w_008_3461, w_008_3462, w_008_3463, w_008_3464, w_008_3465, w_008_3466, w_008_3467, w_008_3468, w_008_3469, w_008_3470, w_008_3471, w_008_3472, w_008_3473, w_008_3474, w_008_3475, w_008_3476, w_008_3477, w_008_3478, w_008_3479, w_008_3480, w_008_3481, w_008_3482, w_008_3483, w_008_3484, w_008_3485, w_008_3486, w_008_3488, w_008_3489, w_008_3490, w_008_3491, w_008_3492, w_008_3493, w_008_3494, w_008_3495, w_008_3496, w_008_3497, w_008_3498, w_008_3499, w_008_3500, w_008_3501, w_008_3502, w_008_3503, w_008_3504, w_008_3505, w_008_3506, w_008_3507, w_008_3508, w_008_3509, w_008_3510, w_008_3511, w_008_3512, w_008_3513, w_008_3514, w_008_3515, w_008_3516, w_008_3517, w_008_3518, w_008_3519, w_008_3520, w_008_3521, w_008_3522, w_008_3523, w_008_3524, w_008_3525, w_008_3526, w_008_3527, w_008_3528, w_008_3529, w_008_3530, w_008_3531, w_008_3532, w_008_3533, w_008_3534, w_008_3535, w_008_3536, w_008_3537, w_008_3538, w_008_3539, w_008_3540, w_008_3541, w_008_3542, w_008_3543, w_008_3544, w_008_3545, w_008_3546, w_008_3547, w_008_3548, w_008_3549, w_008_3550, w_008_3551, w_008_3552, w_008_3553, w_008_3554, w_008_3555, w_008_3556, w_008_3557, w_008_3558, w_008_3559, w_008_3560, w_008_3561, w_008_3562, w_008_3563, w_008_3564, w_008_3565, w_008_3566, w_008_3567, w_008_3568, w_008_3569, w_008_3570, w_008_3571, w_008_3572, w_008_3573, w_008_3574, w_008_3575, w_008_3576, w_008_3577, w_008_3578, w_008_3579, w_008_3581, w_008_3583, w_008_3584, w_008_3585, w_008_3586, w_008_3587, w_008_3588, w_008_3589, w_008_3590, w_008_3591, w_008_3592, w_008_3593, w_008_3594, w_008_3595, w_008_3596, w_008_3597, w_008_3598, w_008_3599, w_008_3600, w_008_3601, w_008_3602, w_008_3603, w_008_3604, w_008_3605, w_008_3606, w_008_3607, w_008_3608, w_008_3609, w_008_3610, w_008_3612, w_008_3613, w_008_3614, w_008_3615, w_008_3616, w_008_3617, w_008_3618, w_008_3619, w_008_3621, w_008_3623, w_008_3624, w_008_3625, w_008_3626, w_008_3627, w_008_3628, w_008_3629, w_008_3630, w_008_3631, w_008_3632, w_008_3633, w_008_3634, w_008_3635, w_008_3636, w_008_3637, w_008_3638, w_008_3639, w_008_3640, w_008_3641, w_008_3642, w_008_3645, w_008_3646, w_008_3647, w_008_3648, w_008_3649, w_008_3650, w_008_3651, w_008_3652, w_008_3653, w_008_3654, w_008_3655, w_008_3656, w_008_3657, w_008_3658, w_008_3659, w_008_3660, w_008_3661, w_008_3662, w_008_3663, w_008_3664, w_008_3665, w_008_3666, w_008_3668, w_008_3669, w_008_3670, w_008_3671, w_008_3672, w_008_3673, w_008_3674, w_008_3675, w_008_3676, w_008_3677, w_008_3678, w_008_3679, w_008_3680, w_008_3681, w_008_3682, w_008_3683, w_008_3684, w_008_3685, w_008_3686, w_008_3687, w_008_3688, w_008_3689, w_008_3690, w_008_3691, w_008_3692, w_008_3693, w_008_3694, w_008_3695, w_008_3696, w_008_3697, w_008_3698, w_008_3699, w_008_3700, w_008_3701, w_008_3702, w_008_3703, w_008_3704, w_008_3705, w_008_3706, w_008_3707, w_008_3708, w_008_3709, w_008_3710, w_008_3711, w_008_3712, w_008_3713, w_008_3714, w_008_3715, w_008_3716, w_008_3717, w_008_3718, w_008_3719, w_008_3720, w_008_3721, w_008_3722, w_008_3723, w_008_3724, w_008_3725, w_008_3726, w_008_3727, w_008_3728, w_008_3729, w_008_3730, w_008_3731, w_008_3732, w_008_3733, w_008_3734, w_008_3735, w_008_3736, w_008_3737, w_008_3738, w_008_3739, w_008_3741, w_008_3742, w_008_3743, w_008_3744, w_008_3745, w_008_3746, w_008_3747, w_008_3748, w_008_3749, w_008_3750, w_008_3751, w_008_3752, w_008_3753, w_008_3754, w_008_3755, w_008_3756, w_008_3757, w_008_3758, w_008_3759, w_008_3760, w_008_3761, w_008_3762, w_008_3764, w_008_3765, w_008_3766, w_008_3767, w_008_3768, w_008_3769, w_008_3770, w_008_3771, w_008_3772, w_008_3773, w_008_3774, w_008_3775, w_008_3776, w_008_3777, w_008_3779, w_008_3780, w_008_3781, w_008_3782, w_008_3784, w_008_3785, w_008_3786, w_008_3787, w_008_3788, w_008_3789, w_008_3790, w_008_3791, w_008_3792, w_008_3793, w_008_3794, w_008_3795, w_008_3796, w_008_3797, w_008_3798, w_008_3799, w_008_3800, w_008_3801, w_008_3802, w_008_3803, w_008_3804, w_008_3805, w_008_3806, w_008_3807, w_008_3808, w_008_3809, w_008_3810, w_008_3811, w_008_3812, w_008_3813, w_008_3814, w_008_3815, w_008_3816, w_008_3817, w_008_3818, w_008_3819, w_008_3820, w_008_3821, w_008_3822, w_008_3823, w_008_3824, w_008_3825, w_008_3826, w_008_3827, w_008_3828, w_008_3829, w_008_3830, w_008_3831, w_008_3832, w_008_3833, w_008_3834, w_008_3835, w_008_3836, w_008_3837, w_008_3838, w_008_3839, w_008_3840, w_008_3841, w_008_3842, w_008_3843, w_008_3844, w_008_3845, w_008_3846, w_008_3847, w_008_3848, w_008_3849, w_008_3850, w_008_3851, w_008_3852, w_008_3853, w_008_3854, w_008_3855, w_008_3856, w_008_3857, w_008_3858, w_008_3859, w_008_3860, w_008_3861, w_008_3862, w_008_3863, w_008_3864, w_008_3865, w_008_3866, w_008_3867, w_008_3868, w_008_3869, w_008_3870, w_008_3871, w_008_3872, w_008_3873, w_008_3874, w_008_3875, w_008_3876, w_008_3877, w_008_3878, w_008_3879, w_008_3880, w_008_3881, w_008_3882, w_008_3883, w_008_3884, w_008_3885, w_008_3886, w_008_3887, w_008_3888, w_008_3889, w_008_3891, w_008_3892, w_008_3893, w_008_3894, w_008_3895, w_008_3896, w_008_3897, w_008_3898, w_008_3899, w_008_3900, w_008_3901, w_008_3902, w_008_3903, w_008_3904, w_008_3905, w_008_3906, w_008_3907, w_008_3908, w_008_3909, w_008_3910, w_008_3911, w_008_3912, w_008_3913, w_008_3914, w_008_3915, w_008_3916, w_008_3917, w_008_3918, w_008_3919, w_008_3920, w_008_3921, w_008_3922, w_008_3923, w_008_3924, w_008_3925, w_008_3926, w_008_3927, w_008_3928, w_008_3929, w_008_3930, w_008_3931, w_008_3932, w_008_3933, w_008_3934, w_008_3935, w_008_3936, w_008_3937, w_008_3938, w_008_3940, w_008_3941, w_008_3942, w_008_3944, w_008_3945, w_008_3946, w_008_3947, w_008_3948, w_008_3949, w_008_3950, w_008_3951, w_008_3953, w_008_3954, w_008_3955, w_008_3956, w_008_3957, w_008_3958, w_008_3959, w_008_3960, w_008_3961, w_008_3962, w_008_3963, w_008_3964, w_008_3965, w_008_3966, w_008_3967, w_008_3968, w_008_3969, w_008_3970, w_008_3971, w_008_3972, w_008_3973, w_008_3974, w_008_3975, w_008_3976, w_008_3977, w_008_3978, w_008_3979, w_008_3980, w_008_3981, w_008_3982, w_008_3983, w_008_3984, w_008_3986, w_008_3987, w_008_3988, w_008_3989, w_008_3990, w_008_3991, w_008_3992, w_008_3993, w_008_3994, w_008_3995, w_008_3996, w_008_3997, w_008_3998, w_008_3999, w_008_4000, w_008_4001, w_008_4002, w_008_4003, w_008_4004, w_008_4005, w_008_4006, w_008_4007, w_008_4008, w_008_4009, w_008_4010, w_008_4011, w_008_4012, w_008_4013, w_008_4014, w_008_4015, w_008_4016, w_008_4017, w_008_4018, w_008_4019, w_008_4020, w_008_4021, w_008_4022, w_008_4023, w_008_4025, w_008_4026, w_008_4027, w_008_4028, w_008_4029, w_008_4030, w_008_4031, w_008_4032, w_008_4033, w_008_4034, w_008_4035, w_008_4036, w_008_4037, w_008_4038, w_008_4039, w_008_4040, w_008_4041, w_008_4042, w_008_4043, w_008_4044, w_008_4045, w_008_4048, w_008_4049, w_008_4050, w_008_4051, w_008_4052, w_008_4053, w_008_4054, w_008_4055, w_008_4056, w_008_4057, w_008_4058, w_008_4059, w_008_4061, w_008_4062, w_008_4063, w_008_4064, w_008_4065, w_008_4066, w_008_4067, w_008_4068, w_008_4069, w_008_4070, w_008_4071, w_008_4072, w_008_4073, w_008_4074, w_008_4075, w_008_4076, w_008_4077, w_008_4078, w_008_4079, w_008_4080, w_008_4081, w_008_4082, w_008_4083, w_008_4084, w_008_4085, w_008_4086, w_008_4087, w_008_4088, w_008_4089, w_008_4090, w_008_4091, w_008_4092, w_008_4093, w_008_4094, w_008_4095, w_008_4096, w_008_4097, w_008_4098, w_008_4099, w_008_4100, w_008_4101, w_008_4102, w_008_4103, w_008_4104, w_008_4105, w_008_4106, w_008_4107, w_008_4108, w_008_4109, w_008_4110, w_008_4111, w_008_4112, w_008_4113, w_008_4114, w_008_4115, w_008_4116, w_008_4117, w_008_4118, w_008_4119, w_008_4120, w_008_4121, w_008_4122, w_008_4123, w_008_4124, w_008_4125, w_008_4126, w_008_4127, w_008_4128, w_008_4129, w_008_4130, w_008_4131, w_008_4132, w_008_4134, w_008_4135, w_008_4136, w_008_4137, w_008_4138, w_008_4139, w_008_4140, w_008_4141, w_008_4142, w_008_4143, w_008_4144, w_008_4146, w_008_4147, w_008_4148, w_008_4149, w_008_4150, w_008_4151, w_008_4152, w_008_4153, w_008_4154, w_008_4155, w_008_4156, w_008_4157, w_008_4158, w_008_4159, w_008_4160, w_008_4161, w_008_4162, w_008_4163, w_008_4164, w_008_4165, w_008_4166, w_008_4167, w_008_4168, w_008_4169, w_008_4170, w_008_4171, w_008_4172, w_008_4174, w_008_4175, w_008_4177, w_008_4178, w_008_4179, w_008_4180, w_008_4181, w_008_4182, w_008_4183, w_008_4184, w_008_4185, w_008_4186, w_008_4187, w_008_4188, w_008_4189, w_008_4190, w_008_4191, w_008_4192, w_008_4194, w_008_4195, w_008_4197, w_008_4198, w_008_4200, w_008_4201, w_008_4203, w_008_4205, w_008_4206, w_008_4207, w_008_4208, w_008_4210, w_008_4213, w_008_4214, w_008_4215, w_008_4216, w_008_4218, w_008_4220, w_008_4221, w_008_4222, w_008_4223, w_008_4224, w_008_4225, w_008_4226, w_008_4227, w_008_4228, w_008_4229, w_008_4230, w_008_4231, w_008_4233, w_008_4234, w_008_4235, w_008_4236, w_008_4237, w_008_4239, w_008_4240, w_008_4242, w_008_4243, w_008_4244, w_008_4245, w_008_4246, w_008_4247, w_008_4249, w_008_4250, w_008_4251, w_008_4253, w_008_4254, w_008_4255, w_008_4256, w_008_4257, w_008_4258, w_008_4259, w_008_4260, w_008_4262, w_008_4263, w_008_4264, w_008_4265, w_008_4266, w_008_4267, w_008_4268, w_008_4269, w_008_4270, w_008_4272, w_008_4273, w_008_4274, w_008_4275, w_008_4276, w_008_4278, w_008_4280, w_008_4281, w_008_4283, w_008_4285, w_008_4286, w_008_4287, w_008_4289, w_008_4290, w_008_4291, w_008_4292, w_008_4293, w_008_4294, w_008_4295, w_008_4296, w_008_4297, w_008_4298, w_008_4299, w_008_4301, w_008_4302, w_008_4303, w_008_4304, w_008_4306, w_008_4307, w_008_4309, w_008_4310, w_008_4311, w_008_4313, w_008_4314, w_008_4317, w_008_4319, w_008_4323, w_008_4324, w_008_4325, w_008_4326, w_008_4327, w_008_4328, w_008_4331, w_008_4333, w_008_4334, w_008_4335, w_008_4336, w_008_4337, w_008_4338, w_008_4341, w_008_4342, w_008_4344, w_008_4345, w_008_4346, w_008_4347, w_008_4348, w_008_4349, w_008_4350, w_008_4353, w_008_4355, w_008_4356, w_008_4357, w_008_4358, w_008_4359, w_008_4361, w_008_4367, w_008_4368, w_008_4369, w_008_4370, w_008_4373, w_008_4374, w_008_4376, w_008_4377, w_008_4378, w_008_4379, w_008_4382, w_008_4383, w_008_4384, w_008_4385, w_008_4386, w_008_4387, w_008_4388, w_008_4389, w_008_4392, w_008_4393, w_008_4395, w_008_4396, w_008_4397, w_008_4398, w_008_4399, w_008_4400, w_008_4401, w_008_4402, w_008_4403, w_008_4404, w_008_4406, w_008_4408, w_008_4411, w_008_4412, w_008_4413, w_008_4416, w_008_4417, w_008_4419, w_008_4420, w_008_4421, w_008_4424, w_008_4426, w_008_4428, w_008_4430, w_008_4431, w_008_4432, w_008_4433, w_008_4434, w_008_4435, w_008_4436, w_008_4439, w_008_4440, w_008_4441, w_008_4442, w_008_4443, w_008_4444, w_008_4445, w_008_4446, w_008_4447, w_008_4448, w_008_4449, w_008_4450, w_008_4452, w_008_4453, w_008_4454, w_008_4457, w_008_4458, w_008_4459, w_008_4460, w_008_4463, w_008_4464, w_008_4465, w_008_4466, w_008_4467, w_008_4468, w_008_4469, w_008_4470, w_008_4472, w_008_4473, w_008_4474, w_008_4475, w_008_4476, w_008_4479, w_008_4480, w_008_4481, w_008_4483, w_008_4484, w_008_4485, w_008_4486, w_008_4487, w_008_4489, w_008_4490, w_008_4491, w_008_4492, w_008_4493, w_008_4495, w_008_4497, w_008_4498, w_008_4499, w_008_4500, w_008_4501, w_008_4502, w_008_4503, w_008_4504, w_008_4505, w_008_4506, w_008_4507, w_008_4508, w_008_4509, w_008_4510, w_008_4511, w_008_4512, w_008_4513, w_008_4514, w_008_4515, w_008_4516, w_008_4518, w_008_4519, w_008_4521, w_008_4522, w_008_4523, w_008_4524, w_008_4525, w_008_4526, w_008_4527, w_008_4528, w_008_4529, w_008_4530, w_008_4533, w_008_4535, w_008_4536, w_008_4539, w_008_4540, w_008_4541, w_008_4544, w_008_4545, w_008_4546, w_008_4547, w_008_4548, w_008_4550, w_008_4551, w_008_4552, w_008_4553, w_008_4554, w_008_4555, w_008_4557, w_008_4558, w_008_4559, w_008_4560, w_008_4561, w_008_4562, w_008_4563, w_008_4564, w_008_4565, w_008_4566, w_008_4567, w_008_4568, w_008_4570, w_008_4571, w_008_4573, w_008_4574, w_008_4575, w_008_4576, w_008_4578, w_008_4579, w_008_4580, w_008_4581, w_008_4583, w_008_4584, w_008_4586, w_008_4588, w_008_4590, w_008_4591, w_008_4592, w_008_4593, w_008_4594, w_008_4595, w_008_4596, w_008_4597, w_008_4598, w_008_4599, w_008_4600, w_008_4601, w_008_4602, w_008_4603, w_008_4604, w_008_4605, w_008_4608, w_008_4611, w_008_4612, w_008_4614, w_008_4615, w_008_4617, w_008_4618, w_008_4619, w_008_4620, w_008_4622, w_008_4624, w_008_4625, w_008_4626, w_008_4627, w_008_4629, w_008_4630, w_008_4634, w_008_4635, w_008_4636, w_008_4637, w_008_4638, w_008_4639, w_008_4640, w_008_4641, w_008_4643, w_008_4646, w_008_4647, w_008_4648, w_008_4649, w_008_4651, w_008_4653, w_008_4654, w_008_4655, w_008_4658, w_008_4659, w_008_4661, w_008_4662, w_008_4663, w_008_4664, w_008_4665, w_008_4666, w_008_4668, w_008_4669, w_008_4671, w_008_4672, w_008_4673, w_008_4674, w_008_4675, w_008_4676, w_008_4677, w_008_4678, w_008_4679, w_008_4680, w_008_4683, w_008_4684, w_008_4685, w_008_4686, w_008_4687, w_008_4688, w_008_4689, w_008_4690, w_008_4691, w_008_4693, w_008_4694, w_008_4695, w_008_4696, w_008_4697, w_008_4698, w_008_4699, w_008_4700, w_008_4702, w_008_4703, w_008_4704, w_008_4705, w_008_4706, w_008_4707, w_008_4709, w_008_4710, w_008_4711, w_008_4712, w_008_4713, w_008_4714, w_008_4716, w_008_4718, w_008_4719, w_008_4721, w_008_4722, w_008_4723, w_008_4724, w_008_4726, w_008_4727, w_008_4728, w_008_4729, w_008_4730, w_008_4732, w_008_4733, w_008_4734, w_008_4735, w_008_4736, w_008_4738, w_008_4739, w_008_4740, w_008_4742, w_008_4744, w_008_4745, w_008_4747, w_008_4748, w_008_4749, w_008_4750, w_008_4752, w_008_4753, w_008_4755, w_008_4756, w_008_4757, w_008_4758, w_008_4759, w_008_4760, w_008_4761, w_008_4762, w_008_4763, w_008_4765, w_008_4766, w_008_4768, w_008_4770, w_008_4771, w_008_4772, w_008_4773, w_008_4774, w_008_4776, w_008_4777, w_008_4778, w_008_4779, w_008_4780, w_008_4782, w_008_4783, w_008_4784, w_008_4785, w_008_4786, w_008_4788, w_008_4789, w_008_4790, w_008_4791, w_008_4793, w_008_4794, w_008_4795, w_008_4796, w_008_4797, w_008_4798, w_008_4799, w_008_4801, w_008_4803, w_008_4804, w_008_4805, w_008_4809, w_008_4811, w_008_4812, w_008_4813, w_008_4814, w_008_4815, w_008_4816, w_008_4817, w_008_4818, w_008_4820, w_008_4821, w_008_4822, w_008_4823, w_008_4824, w_008_4825, w_008_4826, w_008_4828, w_008_4831, w_008_4832, w_008_4835, w_008_4836, w_008_4838, w_008_4839, w_008_4840, w_008_4841, w_008_4842, w_008_4844, w_008_4846, w_008_4848, w_008_4850, w_008_4852, w_008_4853, w_008_4854, w_008_4855, w_008_4857, w_008_4858, w_008_4859, w_008_4861, w_008_4862, w_008_4863, w_008_4864, w_008_4865, w_008_4867, w_008_4870, w_008_4871, w_008_4872, w_008_4874, w_008_4875, w_008_4876, w_008_4877, w_008_4879, w_008_4880, w_008_4883, w_008_4886, w_008_4887, w_008_4888, w_008_4890, w_008_4891, w_008_4892, w_008_4893, w_008_4894, w_008_4895, w_008_4896, w_008_4897, w_008_4898, w_008_4899, w_008_4900, w_008_4901, w_008_4902, w_008_4903, w_008_4905, w_008_4906, w_008_4908, w_008_4909, w_008_4910, w_008_4911, w_008_4913, w_008_4914, w_008_4915, w_008_4916, w_008_4917, w_008_4918, w_008_4919, w_008_4920, w_008_4921, w_008_4923, w_008_4924, w_008_4926, w_008_4927, w_008_4928, w_008_4929, w_008_4930, w_008_4931, w_008_4932, w_008_4933, w_008_4934, w_008_4936, w_008_4937, w_008_4939, w_008_4941, w_008_4942, w_008_4943, w_008_4944, w_008_4945, w_008_4946, w_008_4947, w_008_4951, w_008_4953, w_008_4955, w_008_4956, w_008_4957, w_008_4959, w_008_4960, w_008_4961, w_008_4962, w_008_4963, w_008_4964, w_008_4965, w_008_4966, w_008_4968, w_008_4969, w_008_4970, w_008_4971, w_008_4972, w_008_4973, w_008_4974, w_008_4975, w_008_4976, w_008_4979, w_008_4980, w_008_4981, w_008_4982, w_008_4983, w_008_4987, w_008_4988, w_008_4989, w_008_4990, w_008_4991, w_008_4992, w_008_4993, w_008_4994, w_008_4995, w_008_4996, w_008_4997, w_008_4998, w_008_4999, w_008_5000, w_008_5001, w_008_5002, w_008_5003, w_008_5004, w_008_5005, w_008_5008, w_008_5009, w_008_5010, w_008_5011, w_008_5015, w_008_5016, w_008_5018, w_008_5019, w_008_5020, w_008_5021, w_008_5022, w_008_5023, w_008_5024, w_008_5025, w_008_5026, w_008_5029, w_008_5030, w_008_5031, w_008_5032, w_008_5033, w_008_5034, w_008_5036, w_008_5037, w_008_5038, w_008_5039, w_008_5040, w_008_5041, w_008_5043, w_008_5044, w_008_5047, w_008_5050, w_008_5051, w_008_5052, w_008_5053, w_008_5056, w_008_5057, w_008_5058, w_008_5059, w_008_5061, w_008_5062, w_008_5063, w_008_5065, w_008_5066, w_008_5069, w_008_5071, w_008_5072, w_008_5073, w_008_5075, w_008_5077, w_008_5078, w_008_5079, w_008_5080, w_008_5081, w_008_5082, w_008_5083, w_008_5084, w_008_5085, w_008_5086, w_008_5087, w_008_5089, w_008_5091, w_008_5093, w_008_5094, w_008_5095, w_008_5096, w_008_5097, w_008_5098, w_008_5099, w_008_5100, w_008_5101, w_008_5102, w_008_5105, w_008_5107, w_008_5108, w_008_5109, w_008_5110, w_008_5111, w_008_5112, w_008_5114, w_008_5116, w_008_5117, w_008_5118, w_008_5119, w_008_5120, w_008_5121, w_008_5122, w_008_5123, w_008_5124, w_008_5125, w_008_5126, w_008_5127, w_008_5128, w_008_5129, w_008_5130, w_008_5131, w_008_5132, w_008_5133, w_008_5134, w_008_5137, w_008_5138, w_008_5140, w_008_5141, w_008_5142, w_008_5143, w_008_5144, w_008_5145, w_008_5146, w_008_5147, w_008_5149, w_008_5150, w_008_5152, w_008_5153, w_008_5154, w_008_5155, w_008_5156, w_008_5157, w_008_5158, w_008_5159, w_008_5160, w_008_5161, w_008_5162, w_008_5163, w_008_5164, w_008_5165, w_008_5166, w_008_5167, w_008_5168, w_008_5169, w_008_5172, w_008_5174, w_008_5175, w_008_5176, w_008_5178, w_008_5180, w_008_5181, w_008_5182, w_008_5183, w_008_5184, w_008_5186, w_008_5187, w_008_5188, w_008_5189, w_008_5190, w_008_5192, w_008_5196, w_008_5199, w_008_5200, w_008_5201, w_008_5202, w_008_5204, w_008_5206, w_008_5207, w_008_5208, w_008_5209, w_008_5210, w_008_5211, w_008_5213, w_008_5214, w_008_5215, w_008_5217, w_008_5218, w_008_5220, w_008_5221, w_008_5224, w_008_5225, w_008_5226, w_008_5227, w_008_5228, w_008_5229, w_008_5230, w_008_5231, w_008_5232, w_008_5234, w_008_5236, w_008_5239, w_008_5240, w_008_5241, w_008_5242, w_008_5243, w_008_5244, w_008_5245, w_008_5246, w_008_5247, w_008_5248, w_008_5249, w_008_5250, w_008_5251, w_008_5252, w_008_5253, w_008_5255, w_008_5257, w_008_5258, w_008_5259, w_008_5260, w_008_5261, w_008_5262, w_008_5263, w_008_5264, w_008_5265, w_008_5266, w_008_5267, w_008_5268, w_008_5270, w_008_5271, w_008_5272, w_008_5274, w_008_5278, w_008_5279, w_008_5280, w_008_5282, w_008_5283, w_008_5284, w_008_5286, w_008_5287, w_008_5288, w_008_5289, w_008_5290, w_008_5291, w_008_5292, w_008_5293, w_008_5294, w_008_5295, w_008_5297, w_008_5298, w_008_5299, w_008_5301, w_008_5302, w_008_5303, w_008_5304, w_008_5305, w_008_5309, w_008_5310, w_008_5311, w_008_5312, w_008_5313, w_008_5314, w_008_5316, w_008_5319, w_008_5320, w_008_5321, w_008_5322, w_008_5323, w_008_5324, w_008_5325, w_008_5327, w_008_5329, w_008_5330, w_008_5331, w_008_5332, w_008_5333, w_008_5334, w_008_5335, w_008_5336, w_008_5337, w_008_5339, w_008_5340, w_008_5342, w_008_5343, w_008_5344, w_008_5345, w_008_5346, w_008_5347, w_008_5348, w_008_5349, w_008_5352, w_008_5353, w_008_5354, w_008_5355, w_008_5356, w_008_5357, w_008_5358, w_008_5359, w_008_5360, w_008_5362, w_008_5364, w_008_5366, w_008_5367, w_008_5368, w_008_5369, w_008_5372, w_008_5373, w_008_5374, w_008_5376, w_008_5377, w_008_5378, w_008_5379, w_008_5380, w_008_5382, w_008_5383, w_008_5384, w_008_5385, w_008_5386, w_008_5387, w_008_5388, w_008_5389, w_008_5391, w_008_5392, w_008_5393, w_008_5394, w_008_5395, w_008_5397, w_008_5398, w_008_5399, w_008_5400, w_008_5401, w_008_5402, w_008_5403, w_008_5404, w_008_5405, w_008_5406, w_008_5407, w_008_5409, w_008_5410, w_008_5411, w_008_5412, w_008_5414, w_008_5415, w_008_5416, w_008_5417, w_008_5419, w_008_5420, w_008_5421, w_008_5422, w_008_5423, w_008_5424, w_008_5425, w_008_5426, w_008_5427, w_008_5428, w_008_5429, w_008_5430, w_008_5431, w_008_5432, w_008_5433, w_008_5434, w_008_5435, w_008_5436, w_008_5437, w_008_5438, w_008_5439, w_008_5440, w_008_5441, w_008_5442, w_008_5443, w_008_5445, w_008_5446, w_008_5447, w_008_5448, w_008_5449, w_008_5450, w_008_5451, w_008_5453, w_008_5455, w_008_5456, w_008_5457, w_008_5458, w_008_5459, w_008_5460, w_008_5461, w_008_5463, w_008_5466, w_008_5467, w_008_5468, w_008_5470, w_008_5471, w_008_5472, w_008_5473, w_008_5474, w_008_5475, w_008_5476, w_008_5477, w_008_5478, w_008_5479, w_008_5482, w_008_5483, w_008_5484, w_008_5485, w_008_5486, w_008_5488, w_008_5489, w_008_5490, w_008_5492, w_008_5494, w_008_5495, w_008_5497, w_008_5498, w_008_5499, w_008_5500, w_008_5501, w_008_5502, w_008_5503, w_008_5504, w_008_5505, w_008_5506, w_008_5507, w_008_5510, w_008_5511, w_008_5512, w_008_5513, w_008_5514, w_008_5515, w_008_5516, w_008_5518, w_008_5519, w_008_5520, w_008_5521, w_008_5522, w_008_5524, w_008_5525, w_008_5526, w_008_5527, w_008_5528, w_008_5529, w_008_5530, w_008_5531, w_008_5532, w_008_5533, w_008_5534, w_008_5535, w_008_5536, w_008_5537, w_008_5539, w_008_5540, w_008_5541, w_008_5542, w_008_5543, w_008_5544, w_008_5545, w_008_5546, w_008_5547, w_008_5548, w_008_5550, w_008_5551, w_008_5552, w_008_5553, w_008_5555, w_008_5556, w_008_5557, w_008_5558, w_008_5559, w_008_5560, w_008_5561, w_008_5562, w_008_5563, w_008_5564, w_008_5565, w_008_5566, w_008_5568, w_008_5569, w_008_5570, w_008_5572, w_008_5573, w_008_5574, w_008_5575, w_008_5577, w_008_5578, w_008_5579, w_008_5580, w_008_5581, w_008_5583, w_008_5585, w_008_5587, w_008_5588, w_008_5589, w_008_5592, w_008_5593, w_008_5594, w_008_5596, w_008_5597, w_008_5598, w_008_5600, w_008_5602, w_008_5603, w_008_5604, w_008_5605, w_008_5606, w_008_5607, w_008_5609, w_008_5610, w_008_5611, w_008_5613, w_008_5614, w_008_5615, w_008_5616, w_008_5617, w_008_5618, w_008_5619, w_008_5620, w_008_5622, w_008_5623, w_008_5624, w_008_5625, w_008_5626, w_008_5627, w_008_5628, w_008_5629, w_008_5630, w_008_5631, w_008_5632, w_008_5633, w_008_5634, w_008_5636, w_008_5637, w_008_5638, w_008_5640, w_008_5641, w_008_5644, w_008_5647, w_008_5648, w_008_5650, w_008_5652, w_008_5653, w_008_5654, w_008_5655, w_008_5656, w_008_5657, w_008_5658, w_008_5660, w_008_5661, w_008_5662, w_008_5664, w_008_5665, w_008_5667, w_008_5668, w_008_5669, w_008_5670, w_008_5671, w_008_5672, w_008_5673, w_008_5677, w_008_5678, w_008_5680, w_008_5682, w_008_5683, w_008_5684, w_008_5685, w_008_5686, w_008_5687, w_008_5688, w_008_5691, w_008_5692, w_008_5693, w_008_5694, w_008_5695, w_008_5696, w_008_5698, w_008_5699, w_008_5700, w_008_5701, w_008_5702, w_008_5703, w_008_5705, w_008_5706, w_008_5707, w_008_5708, w_008_5709, w_008_5710, w_008_5711, w_008_5712, w_008_5713, w_008_5714, w_008_5715, w_008_5716, w_008_5717, w_008_5718, w_008_5719, w_008_5721, w_008_5722, w_008_5723, w_008_5724, w_008_5725, w_008_5726, w_008_5729, w_008_5730, w_008_5731, w_008_5732, w_008_5733, w_008_5734, w_008_5735, w_008_5736, w_008_5737, w_008_5738, w_008_5740, w_008_5741, w_008_5743, w_008_5744, w_008_5745, w_008_5747, w_008_5748, w_008_5749, w_008_5750, w_008_5751, w_008_5752, w_008_5754, w_008_5755, w_008_5756, w_008_5757, w_008_5758, w_008_5759, w_008_5760, w_008_5762, w_008_5763, w_008_5764, w_008_5765, w_008_5766, w_008_5767, w_008_5768, w_008_5770, w_008_5771, w_008_5772, w_008_5773, w_008_5774, w_008_5775, w_008_5776, w_008_5778, w_008_5779, w_008_5780, w_008_5782, w_008_5783, w_008_5784, w_008_5785, w_008_5786, w_008_5787, w_008_5788, w_008_5789, w_008_5790, w_008_5791, w_008_5794, w_008_5797, w_008_5798, w_008_5799, w_008_5800, w_008_5801, w_008_5802, w_008_5803, w_008_5804, w_008_5805, w_008_5806, w_008_5807, w_008_5808, w_008_5809, w_008_5811, w_008_5812, w_008_5815, w_008_5816;
  wire w_009_000, w_009_001, w_009_002, w_009_003, w_009_004, w_009_005, w_009_006, w_009_007, w_009_008, w_009_009, w_009_010, w_009_011, w_009_012, w_009_013, w_009_014, w_009_015, w_009_016, w_009_017, w_009_018, w_009_019, w_009_020, w_009_021, w_009_022, w_009_023, w_009_024, w_009_025, w_009_026, w_009_027, w_009_028, w_009_029, w_009_030, w_009_031, w_009_032, w_009_033, w_009_034, w_009_035, w_009_036, w_009_037, w_009_038, w_009_039, w_009_040, w_009_041, w_009_042, w_009_043, w_009_044, w_009_045, w_009_046, w_009_047, w_009_048, w_009_049, w_009_050, w_009_051, w_009_052, w_009_053, w_009_054, w_009_055, w_009_056, w_009_057, w_009_058, w_009_059, w_009_060, w_009_061, w_009_062, w_009_063, w_009_064, w_009_065, w_009_066, w_009_067, w_009_068, w_009_069, w_009_070, w_009_071, w_009_072, w_009_073, w_009_074, w_009_075, w_009_076, w_009_077, w_009_078, w_009_079, w_009_080, w_009_081, w_009_082, w_009_083, w_009_084, w_009_085, w_009_086, w_009_087, w_009_088, w_009_089, w_009_090, w_009_091, w_009_092, w_009_093, w_009_094, w_009_095, w_009_096, w_009_097, w_009_098, w_009_099, w_009_100, w_009_101, w_009_102, w_009_103, w_009_104, w_009_105, w_009_106, w_009_107, w_009_108, w_009_109, w_009_110, w_009_111, w_009_112, w_009_113, w_009_114, w_009_115, w_009_116, w_009_117, w_009_118, w_009_119, w_009_120, w_009_121, w_009_122, w_009_123, w_009_124, w_009_125, w_009_126, w_009_127, w_009_128, w_009_129, w_009_130, w_009_131, w_009_132, w_009_133, w_009_134, w_009_135, w_009_136, w_009_137, w_009_138, w_009_139, w_009_140, w_009_141, w_009_142, w_009_143, w_009_144, w_009_145, w_009_146, w_009_147, w_009_148, w_009_149, w_009_150, w_009_151, w_009_152, w_009_153, w_009_154, w_009_155, w_009_156, w_009_157, w_009_158, w_009_159, w_009_160, w_009_161, w_009_162, w_009_163, w_009_164, w_009_165, w_009_166, w_009_167, w_009_168, w_009_169, w_009_170, w_009_171, w_009_172, w_009_173, w_009_174, w_009_175, w_009_176, w_009_177, w_009_178, w_009_179, w_009_180, w_009_181, w_009_182, w_009_183, w_009_184, w_009_185, w_009_186, w_009_187, w_009_188, w_009_189, w_009_190, w_009_191, w_009_192, w_009_193, w_009_194, w_009_195, w_009_196, w_009_197, w_009_198, w_009_199, w_009_200, w_009_201, w_009_202, w_009_203, w_009_204, w_009_205, w_009_206, w_009_207, w_009_208, w_009_209, w_009_210, w_009_211, w_009_212, w_009_213, w_009_214, w_009_215, w_009_216, w_009_217, w_009_218, w_009_219, w_009_220, w_009_221, w_009_222, w_009_223, w_009_224, w_009_225, w_009_226, w_009_227, w_009_228, w_009_229, w_009_230, w_009_231, w_009_232, w_009_233, w_009_234, w_009_235, w_009_236, w_009_237, w_009_238, w_009_239, w_009_240, w_009_241, w_009_242, w_009_243, w_009_244, w_009_245, w_009_246, w_009_247, w_009_248, w_009_249, w_009_250, w_009_252, w_009_253, w_009_254, w_009_255, w_009_256, w_009_257, w_009_258, w_009_259, w_009_260, w_009_261, w_009_262, w_009_263, w_009_264, w_009_265, w_009_266, w_009_267, w_009_268, w_009_269, w_009_270, w_009_271, w_009_272, w_009_273, w_009_274, w_009_275, w_009_276, w_009_277, w_009_278, w_009_279, w_009_280, w_009_281, w_009_282, w_009_283, w_009_284, w_009_285, w_009_286, w_009_287, w_009_288, w_009_289, w_009_290, w_009_291, w_009_292, w_009_293, w_009_294, w_009_295, w_009_296, w_009_297, w_009_298, w_009_299, w_009_300, w_009_301, w_009_302, w_009_303, w_009_304, w_009_305, w_009_306, w_009_307, w_009_308, w_009_309, w_009_310, w_009_311, w_009_312, w_009_313, w_009_314, w_009_315, w_009_316, w_009_317, w_009_318, w_009_319, w_009_320, w_009_321, w_009_322, w_009_323, w_009_324, w_009_325, w_009_326, w_009_327, w_009_328, w_009_329, w_009_330, w_009_331, w_009_332, w_009_333, w_009_334, w_009_335, w_009_336, w_009_337, w_009_338, w_009_339, w_009_340, w_009_341, w_009_342, w_009_344, w_009_345, w_009_346, w_009_347, w_009_348, w_009_349, w_009_350, w_009_351, w_009_352, w_009_353, w_009_354, w_009_355, w_009_356, w_009_357, w_009_358, w_009_359, w_009_360, w_009_361, w_009_362, w_009_363, w_009_364, w_009_365, w_009_366, w_009_367, w_009_368, w_009_369, w_009_370, w_009_371, w_009_373, w_009_374, w_009_375, w_009_376, w_009_377, w_009_378, w_009_379, w_009_380, w_009_381, w_009_382, w_009_383, w_009_385, w_009_386, w_009_387, w_009_388, w_009_389, w_009_390, w_009_391, w_009_392, w_009_393, w_009_394, w_009_395, w_009_396, w_009_397, w_009_398, w_009_399, w_009_400, w_009_401, w_009_402, w_009_403, w_009_404, w_009_405, w_009_406, w_009_407, w_009_408, w_009_409, w_009_410, w_009_411, w_009_412, w_009_413, w_009_414, w_009_415, w_009_416, w_009_417, w_009_418, w_009_419, w_009_420, w_009_421, w_009_422, w_009_423, w_009_424, w_009_425, w_009_426, w_009_427, w_009_429, w_009_430, w_009_431, w_009_432, w_009_433, w_009_434, w_009_435, w_009_436, w_009_437, w_009_438, w_009_439, w_009_440, w_009_441, w_009_442, w_009_443, w_009_444, w_009_445, w_009_446, w_009_447, w_009_448, w_009_449, w_009_450, w_009_451, w_009_452, w_009_454, w_009_455, w_009_456, w_009_457, w_009_458, w_009_459, w_009_460, w_009_461, w_009_462, w_009_463, w_009_464, w_009_465, w_009_466, w_009_467, w_009_468, w_009_469, w_009_470, w_009_471, w_009_472, w_009_473, w_009_474, w_009_475, w_009_476, w_009_477, w_009_478, w_009_479, w_009_480, w_009_481, w_009_482, w_009_483, w_009_484, w_009_485, w_009_486, w_009_487, w_009_488, w_009_489, w_009_490, w_009_491, w_009_492, w_009_493, w_009_494, w_009_495, w_009_496, w_009_497, w_009_498, w_009_499, w_009_500, w_009_501, w_009_502, w_009_503, w_009_504, w_009_505, w_009_506, w_009_507, w_009_508, w_009_509, w_009_510, w_009_511, w_009_512, w_009_513, w_009_514, w_009_515, w_009_516, w_009_517, w_009_518, w_009_519, w_009_520, w_009_521, w_009_522, w_009_523, w_009_524, w_009_525, w_009_526, w_009_527, w_009_528, w_009_529, w_009_530, w_009_531, w_009_532, w_009_533, w_009_534, w_009_535, w_009_536, w_009_537, w_009_538, w_009_539, w_009_540, w_009_541, w_009_542, w_009_543, w_009_544, w_009_545, w_009_546, w_009_547, w_009_548, w_009_549, w_009_550, w_009_551, w_009_552, w_009_553, w_009_554, w_009_555, w_009_556, w_009_557, w_009_558, w_009_559, w_009_560, w_009_561, w_009_562, w_009_563, w_009_564, w_009_565, w_009_566, w_009_567, w_009_568, w_009_569, w_009_570, w_009_571, w_009_572, w_009_573, w_009_574, w_009_575, w_009_576, w_009_577, w_009_578, w_009_579, w_009_580, w_009_581, w_009_582, w_009_583, w_009_584, w_009_585, w_009_586, w_009_587, w_009_588, w_009_589, w_009_590, w_009_591, w_009_592, w_009_593, w_009_594, w_009_595, w_009_596, w_009_597, w_009_598, w_009_599, w_009_600, w_009_601, w_009_602, w_009_603, w_009_604, w_009_605, w_009_606, w_009_607, w_009_608, w_009_609, w_009_610, w_009_611, w_009_612, w_009_614, w_009_615, w_009_616, w_009_617, w_009_618, w_009_619, w_009_620, w_009_621, w_009_622, w_009_623, w_009_624, w_009_625, w_009_626, w_009_627, w_009_628, w_009_629, w_009_630, w_009_632, w_009_633, w_009_634, w_009_635, w_009_636, w_009_637, w_009_638, w_009_639, w_009_640, w_009_641, w_009_642, w_009_643, w_009_644, w_009_645, w_009_646, w_009_647, w_009_648, w_009_649, w_009_650, w_009_651, w_009_652, w_009_653, w_009_654, w_009_655, w_009_656, w_009_657, w_009_658, w_009_659, w_009_660, w_009_661, w_009_662, w_009_663, w_009_664, w_009_665, w_009_666, w_009_667, w_009_668, w_009_669, w_009_670, w_009_671, w_009_672, w_009_673, w_009_674, w_009_675, w_009_676, w_009_677, w_009_678, w_009_679, w_009_680, w_009_681, w_009_682, w_009_683, w_009_684, w_009_685, w_009_686, w_009_687, w_009_688, w_009_689, w_009_690, w_009_691, w_009_692, w_009_693, w_009_694, w_009_695, w_009_696, w_009_697, w_009_698, w_009_699, w_009_700, w_009_701, w_009_702, w_009_703, w_009_704, w_009_705, w_009_706, w_009_707, w_009_708, w_009_709, w_009_710, w_009_711, w_009_712, w_009_713, w_009_714, w_009_715, w_009_716, w_009_717, w_009_718, w_009_719, w_009_720, w_009_721, w_009_722, w_009_723, w_009_724, w_009_725, w_009_726, w_009_727, w_009_728, w_009_729, w_009_730, w_009_731, w_009_732, w_009_733, w_009_734, w_009_735, w_009_736, w_009_737, w_009_738, w_009_739, w_009_740, w_009_741, w_009_742, w_009_743, w_009_744, w_009_745, w_009_746, w_009_747, w_009_748, w_009_749, w_009_750, w_009_751, w_009_752, w_009_753, w_009_754, w_009_755, w_009_756, w_009_757, w_009_758, w_009_759, w_009_760, w_009_761, w_009_762, w_009_763, w_009_764, w_009_765, w_009_766, w_009_767, w_009_768, w_009_769, w_009_770, w_009_771, w_009_772, w_009_773, w_009_774, w_009_775, w_009_776, w_009_777, w_009_778, w_009_779, w_009_780, w_009_781, w_009_782, w_009_783, w_009_784, w_009_785, w_009_786, w_009_787, w_009_788, w_009_789, w_009_790, w_009_791, w_009_792, w_009_793, w_009_794, w_009_795, w_009_796, w_009_797, w_009_798, w_009_799, w_009_800, w_009_801, w_009_802, w_009_803, w_009_804, w_009_805, w_009_806, w_009_807, w_009_808, w_009_810, w_009_811, w_009_812, w_009_813, w_009_814, w_009_815, w_009_816, w_009_817, w_009_818, w_009_819, w_009_820, w_009_821, w_009_822, w_009_823, w_009_824, w_009_825, w_009_826, w_009_827, w_009_828, w_009_829, w_009_830, w_009_831, w_009_832, w_009_833, w_009_834, w_009_835, w_009_836, w_009_837, w_009_838, w_009_839, w_009_840, w_009_841, w_009_842, w_009_843, w_009_844, w_009_845, w_009_846, w_009_848, w_009_849, w_009_850, w_009_851, w_009_852, w_009_853, w_009_855, w_009_856, w_009_857, w_009_858, w_009_859, w_009_860, w_009_861, w_009_862, w_009_863, w_009_864, w_009_865, w_009_866, w_009_867, w_009_868, w_009_869, w_009_870, w_009_871, w_009_872, w_009_873, w_009_874, w_009_875, w_009_876, w_009_877, w_009_878, w_009_879, w_009_880, w_009_881, w_009_882, w_009_883, w_009_884, w_009_885, w_009_887, w_009_888, w_009_889, w_009_890, w_009_891, w_009_892, w_009_893, w_009_894, w_009_895, w_009_896, w_009_897, w_009_898, w_009_899, w_009_900, w_009_901, w_009_902, w_009_903, w_009_904, w_009_905, w_009_906, w_009_907, w_009_908, w_009_909, w_009_910, w_009_911, w_009_912, w_009_913, w_009_914, w_009_915, w_009_916, w_009_917, w_009_919, w_009_920, w_009_921, w_009_922, w_009_923, w_009_924, w_009_925, w_009_926, w_009_927, w_009_928, w_009_929, w_009_930, w_009_931, w_009_932, w_009_933, w_009_934, w_009_935, w_009_936, w_009_937, w_009_938, w_009_940, w_009_941, w_009_942, w_009_943, w_009_945, w_009_947, w_009_948, w_009_949, w_009_950, w_009_951, w_009_952, w_009_953, w_009_954, w_009_956, w_009_957, w_009_959, w_009_960, w_009_961, w_009_962, w_009_963, w_009_964, w_009_965, w_009_966, w_009_967, w_009_968, w_009_969, w_009_970, w_009_971, w_009_972, w_009_973, w_009_974, w_009_975, w_009_976, w_009_977, w_009_978, w_009_979, w_009_980, w_009_981, w_009_982, w_009_983, w_009_985, w_009_986, w_009_987, w_009_988, w_009_989, w_009_990, w_009_991, w_009_992, w_009_993, w_009_994, w_009_995, w_009_996, w_009_998, w_009_999, w_009_1000, w_009_1001, w_009_1002, w_009_1003, w_009_1004, w_009_1005, w_009_1006, w_009_1007, w_009_1008, w_009_1009, w_009_1010, w_009_1011, w_009_1012, w_009_1013, w_009_1014, w_009_1015, w_009_1016, w_009_1017, w_009_1018, w_009_1019, w_009_1020, w_009_1021, w_009_1022, w_009_1023, w_009_1024, w_009_1025, w_009_1026, w_009_1027, w_009_1028, w_009_1029, w_009_1030, w_009_1031, w_009_1032, w_009_1034, w_009_1035, w_009_1036, w_009_1037, w_009_1038, w_009_1039, w_009_1040, w_009_1041, w_009_1042, w_009_1043, w_009_1044, w_009_1045, w_009_1046, w_009_1047, w_009_1048, w_009_1049, w_009_1050, w_009_1051, w_009_1052, w_009_1053, w_009_1054, w_009_1055, w_009_1056, w_009_1057, w_009_1058, w_009_1059, w_009_1060, w_009_1061, w_009_1062, w_009_1063, w_009_1064, w_009_1065, w_009_1066, w_009_1067, w_009_1068, w_009_1069, w_009_1070, w_009_1071, w_009_1072, w_009_1073, w_009_1074, w_009_1075, w_009_1076, w_009_1077, w_009_1079, w_009_1080, w_009_1081, w_009_1082, w_009_1083, w_009_1084, w_009_1085, w_009_1086, w_009_1087, w_009_1088, w_009_1089, w_009_1090, w_009_1091, w_009_1092, w_009_1093, w_009_1094, w_009_1095, w_009_1096, w_009_1097, w_009_1098, w_009_1099, w_009_1100, w_009_1101, w_009_1102, w_009_1103, w_009_1105, w_009_1106, w_009_1107, w_009_1108, w_009_1109, w_009_1110, w_009_1111, w_009_1112, w_009_1113, w_009_1114, w_009_1115, w_009_1116, w_009_1117, w_009_1118, w_009_1119, w_009_1120, w_009_1121, w_009_1122, w_009_1123, w_009_1124, w_009_1125, w_009_1126, w_009_1127, w_009_1128, w_009_1129, w_009_1130, w_009_1131, w_009_1132, w_009_1133, w_009_1134, w_009_1135, w_009_1136, w_009_1137, w_009_1138, w_009_1139, w_009_1140, w_009_1141, w_009_1142, w_009_1143, w_009_1144, w_009_1145, w_009_1146, w_009_1147, w_009_1148, w_009_1149, w_009_1150, w_009_1151, w_009_1152, w_009_1153, w_009_1154, w_009_1155, w_009_1156, w_009_1157, w_009_1158, w_009_1159, w_009_1161, w_009_1162, w_009_1163, w_009_1164, w_009_1165, w_009_1166, w_009_1167, w_009_1168, w_009_1169, w_009_1170, w_009_1171, w_009_1172, w_009_1173, w_009_1174, w_009_1175, w_009_1177, w_009_1178, w_009_1179, w_009_1180, w_009_1181, w_009_1182, w_009_1183, w_009_1184, w_009_1185, w_009_1186, w_009_1187, w_009_1188, w_009_1189, w_009_1190, w_009_1191, w_009_1192, w_009_1193, w_009_1194, w_009_1195, w_009_1196, w_009_1197, w_009_1198, w_009_1199, w_009_1200, w_009_1201, w_009_1202, w_009_1203, w_009_1204, w_009_1205, w_009_1206, w_009_1207, w_009_1208, w_009_1209, w_009_1210, w_009_1211, w_009_1212, w_009_1213, w_009_1214, w_009_1215, w_009_1216, w_009_1217, w_009_1218, w_009_1219, w_009_1220, w_009_1221, w_009_1222, w_009_1223, w_009_1224, w_009_1225, w_009_1226, w_009_1227, w_009_1228, w_009_1229, w_009_1230, w_009_1232, w_009_1233, w_009_1234, w_009_1235, w_009_1236, w_009_1237, w_009_1238, w_009_1239, w_009_1240, w_009_1241, w_009_1242, w_009_1243, w_009_1244, w_009_1245, w_009_1246, w_009_1247, w_009_1248, w_009_1249, w_009_1250, w_009_1251, w_009_1252, w_009_1253, w_009_1254, w_009_1255, w_009_1256, w_009_1257, w_009_1258, w_009_1259, w_009_1260, w_009_1261, w_009_1263, w_009_1264, w_009_1265, w_009_1266, w_009_1267, w_009_1268, w_009_1269, w_009_1270, w_009_1271, w_009_1272, w_009_1273, w_009_1274, w_009_1275, w_009_1276, w_009_1277, w_009_1278, w_009_1279, w_009_1280, w_009_1281, w_009_1282, w_009_1283, w_009_1284, w_009_1285, w_009_1286, w_009_1287, w_009_1288, w_009_1289, w_009_1290, w_009_1291, w_009_1293, w_009_1294, w_009_1295, w_009_1296, w_009_1298, w_009_1299, w_009_1300, w_009_1301, w_009_1302, w_009_1303, w_009_1304, w_009_1305, w_009_1306, w_009_1307, w_009_1308, w_009_1309, w_009_1310, w_009_1311, w_009_1312, w_009_1313, w_009_1314, w_009_1315, w_009_1316, w_009_1317, w_009_1318, w_009_1320, w_009_1321, w_009_1322, w_009_1323, w_009_1324, w_009_1325, w_009_1326, w_009_1327, w_009_1328, w_009_1329, w_009_1330, w_009_1331, w_009_1332, w_009_1333, w_009_1334, w_009_1335, w_009_1336, w_009_1337, w_009_1338, w_009_1339, w_009_1340, w_009_1341, w_009_1342, w_009_1343, w_009_1344, w_009_1345, w_009_1346, w_009_1347, w_009_1348, w_009_1349, w_009_1350, w_009_1351, w_009_1352, w_009_1353, w_009_1354, w_009_1355, w_009_1356, w_009_1357, w_009_1358, w_009_1359, w_009_1360, w_009_1361, w_009_1362, w_009_1363, w_009_1364, w_009_1365, w_009_1366, w_009_1367, w_009_1368, w_009_1370, w_009_1373, w_009_1374, w_009_1375, w_009_1376, w_009_1377, w_009_1378, w_009_1379, w_009_1380, w_009_1381, w_009_1382, w_009_1383, w_009_1384, w_009_1385, w_009_1386, w_009_1387, w_009_1388, w_009_1389, w_009_1390, w_009_1391, w_009_1392, w_009_1393, w_009_1395, w_009_1396, w_009_1397, w_009_1398, w_009_1400, w_009_1401, w_009_1402, w_009_1403, w_009_1404, w_009_1405, w_009_1406, w_009_1407, w_009_1408, w_009_1409, w_009_1410, w_009_1411, w_009_1412, w_009_1413, w_009_1414, w_009_1415, w_009_1416, w_009_1417, w_009_1418, w_009_1419, w_009_1420, w_009_1421, w_009_1422, w_009_1423, w_009_1424, w_009_1425, w_009_1426, w_009_1427, w_009_1428, w_009_1429, w_009_1430, w_009_1431, w_009_1432, w_009_1433, w_009_1435, w_009_1436, w_009_1437, w_009_1438, w_009_1439, w_009_1440, w_009_1441, w_009_1442, w_009_1443, w_009_1444, w_009_1445, w_009_1446, w_009_1447, w_009_1448, w_009_1449, w_009_1450, w_009_1451, w_009_1452, w_009_1453, w_009_1454, w_009_1455, w_009_1456, w_009_1457, w_009_1458, w_009_1459, w_009_1460, w_009_1461, w_009_1462, w_009_1463, w_009_1464, w_009_1465, w_009_1466, w_009_1467, w_009_1468, w_009_1469, w_009_1470, w_009_1471, w_009_1472, w_009_1473, w_009_1474, w_009_1475, w_009_1476, w_009_1477, w_009_1478, w_009_1479, w_009_1481, w_009_1482, w_009_1483, w_009_1484, w_009_1485, w_009_1486, w_009_1488, w_009_1489, w_009_1490, w_009_1491, w_009_1492, w_009_1493, w_009_1494, w_009_1495, w_009_1496, w_009_1497, w_009_1498, w_009_1499, w_009_1500, w_009_1501, w_009_1502, w_009_1503, w_009_1504, w_009_1505, w_009_1506, w_009_1507, w_009_1508, w_009_1509, w_009_1510, w_009_1511, w_009_1512, w_009_1513, w_009_1514, w_009_1515, w_009_1516, w_009_1517, w_009_1518, w_009_1520, w_009_1521, w_009_1522, w_009_1523, w_009_1524, w_009_1525, w_009_1526, w_009_1527, w_009_1528, w_009_1529, w_009_1530, w_009_1531, w_009_1532, w_009_1533, w_009_1534, w_009_1535, w_009_1536, w_009_1537, w_009_1538, w_009_1539, w_009_1540, w_009_1542, w_009_1543, w_009_1544, w_009_1545, w_009_1546, w_009_1547, w_009_1548, w_009_1549, w_009_1550, w_009_1551, w_009_1552, w_009_1553, w_009_1555, w_009_1556, w_009_1557, w_009_1558, w_009_1559, w_009_1560, w_009_1561, w_009_1562, w_009_1563, w_009_1564, w_009_1565, w_009_1566, w_009_1567, w_009_1568, w_009_1569, w_009_1570, w_009_1572, w_009_1573, w_009_1574, w_009_1575, w_009_1576, w_009_1577, w_009_1578, w_009_1579, w_009_1580, w_009_1581, w_009_1583, w_009_1584, w_009_1585, w_009_1586, w_009_1587, w_009_1588, w_009_1589, w_009_1590, w_009_1591, w_009_1592, w_009_1593, w_009_1594, w_009_1595, w_009_1596, w_009_1598, w_009_1599, w_009_1600, w_009_1601, w_009_1602, w_009_1603, w_009_1604, w_009_1605, w_009_1606, w_009_1607, w_009_1608, w_009_1609, w_009_1610, w_009_1611, w_009_1612, w_009_1613, w_009_1614, w_009_1615, w_009_1617, w_009_1618, w_009_1619, w_009_1620, w_009_1621, w_009_1622, w_009_1623, w_009_1624, w_009_1625, w_009_1626, w_009_1627, w_009_1628, w_009_1629, w_009_1630, w_009_1631, w_009_1632, w_009_1634, w_009_1635, w_009_1636, w_009_1637, w_009_1638, w_009_1639, w_009_1640, w_009_1641, w_009_1642, w_009_1643, w_009_1644, w_009_1645, w_009_1646, w_009_1647, w_009_1648, w_009_1649, w_009_1650, w_009_1651, w_009_1652, w_009_1653, w_009_1654, w_009_1655, w_009_1656, w_009_1657, w_009_1658, w_009_1659, w_009_1660, w_009_1661, w_009_1662, w_009_1663, w_009_1664, w_009_1665, w_009_1666, w_009_1667, w_009_1669, w_009_1670, w_009_1671, w_009_1672, w_009_1673, w_009_1674, w_009_1675, w_009_1676, w_009_1677, w_009_1678, w_009_1679, w_009_1680, w_009_1681, w_009_1682, w_009_1683, w_009_1684, w_009_1685, w_009_1686, w_009_1687, w_009_1688, w_009_1689, w_009_1690, w_009_1691, w_009_1692, w_009_1693, w_009_1694, w_009_1695, w_009_1696, w_009_1697, w_009_1698, w_009_1699, w_009_1700, w_009_1701, w_009_1702, w_009_1703, w_009_1704, w_009_1705, w_009_1706, w_009_1708, w_009_1709, w_009_1710, w_009_1711, w_009_1712, w_009_1713, w_009_1714, w_009_1715, w_009_1716, w_009_1717, w_009_1718, w_009_1719, w_009_1720, w_009_1721, w_009_1722, w_009_1723, w_009_1724, w_009_1725, w_009_1726, w_009_1727, w_009_1728, w_009_1729, w_009_1730, w_009_1731, w_009_1732, w_009_1733, w_009_1734, w_009_1735, w_009_1736, w_009_1737, w_009_1738, w_009_1739, w_009_1740, w_009_1741, w_009_1742, w_009_1743, w_009_1744, w_009_1745, w_009_1747, w_009_1749, w_009_1750, w_009_1751, w_009_1752, w_009_1753, w_009_1754, w_009_1755, w_009_1756, w_009_1757, w_009_1758, w_009_1759, w_009_1760, w_009_1761, w_009_1762, w_009_1763, w_009_1764, w_009_1765, w_009_1766, w_009_1767, w_009_1768, w_009_1769, w_009_1770, w_009_1771, w_009_1772, w_009_1773, w_009_1774, w_009_1775, w_009_1776, w_009_1777, w_009_1779, w_009_1780, w_009_1781, w_009_1782, w_009_1783, w_009_1784, w_009_1785, w_009_1786, w_009_1787, w_009_1788, w_009_1789, w_009_1790, w_009_1791, w_009_1792, w_009_1793, w_009_1794, w_009_1795, w_009_1796, w_009_1797, w_009_1800, w_009_1801, w_009_1803, w_009_1804, w_009_1805, w_009_1806, w_009_1808, w_009_1809, w_009_1810, w_009_1811, w_009_1812, w_009_1813, w_009_1814, w_009_1815, w_009_1816, w_009_1817, w_009_1818, w_009_1820, w_009_1821, w_009_1822, w_009_1823, w_009_1824, w_009_1825, w_009_1826, w_009_1827, w_009_1828, w_009_1830, w_009_1831, w_009_1832, w_009_1833, w_009_1834, w_009_1835, w_009_1836, w_009_1837, w_009_1838, w_009_1839, w_009_1840, w_009_1841, w_009_1842, w_009_1843, w_009_1844, w_009_1845, w_009_1846, w_009_1847, w_009_1848, w_009_1849, w_009_1850, w_009_1851, w_009_1852, w_009_1853, w_009_1854, w_009_1855, w_009_1856, w_009_1857, w_009_1858, w_009_1859, w_009_1860, w_009_1861, w_009_1862, w_009_1864, w_009_1865, w_009_1866, w_009_1867, w_009_1869, w_009_1870, w_009_1871, w_009_1872, w_009_1873, w_009_1875, w_009_1876, w_009_1877, w_009_1878, w_009_1879, w_009_1880, w_009_1881, w_009_1882, w_009_1883, w_009_1885, w_009_1886, w_009_1887, w_009_1888, w_009_1889, w_009_1890, w_009_1891, w_009_1892, w_009_1893, w_009_1894, w_009_1895, w_009_1896, w_009_1897, w_009_1898, w_009_1899, w_009_1900, w_009_1901, w_009_1902, w_009_1903, w_009_1904, w_009_1905, w_009_1906, w_009_1907, w_009_1908, w_009_1909, w_009_1910, w_009_1911, w_009_1912, w_009_1913, w_009_1914, w_009_1915, w_009_1916, w_009_1917, w_009_1918, w_009_1919, w_009_1920, w_009_1921, w_009_1922, w_009_1923, w_009_1924, w_009_1925, w_009_1926, w_009_1927, w_009_1928, w_009_1929, w_009_1930, w_009_1931, w_009_1932, w_009_1933, w_009_1935, w_009_1936, w_009_1937, w_009_1938, w_009_1939, w_009_1940, w_009_1941, w_009_1942, w_009_1943, w_009_1944, w_009_1945, w_009_1946, w_009_1947, w_009_1948, w_009_1950, w_009_1951, w_009_1952, w_009_1953, w_009_1954, w_009_1955, w_009_1956, w_009_1957, w_009_1958, w_009_1959, w_009_1960, w_009_1961, w_009_1962, w_009_1963, w_009_1965, w_009_1966, w_009_1967, w_009_1969, w_009_1970, w_009_1971, w_009_1972, w_009_1973, w_009_1974, w_009_1975, w_009_1976, w_009_1977, w_009_1978, w_009_1979, w_009_1980, w_009_1981, w_009_1982, w_009_1983, w_009_1984, w_009_1985, w_009_1986, w_009_1987, w_009_1988, w_009_1989, w_009_1990, w_009_1991, w_009_1992, w_009_1993, w_009_1994, w_009_1996, w_009_1997, w_009_1998, w_009_1999, w_009_2000, w_009_2001, w_009_2002, w_009_2003, w_009_2004, w_009_2005, w_009_2006, w_009_2007, w_009_2008, w_009_2010, w_009_2011, w_009_2012, w_009_2013, w_009_2014, w_009_2015, w_009_2016, w_009_2017, w_009_2018, w_009_2019, w_009_2020, w_009_2021, w_009_2022, w_009_2023, w_009_2024, w_009_2025, w_009_2026, w_009_2027, w_009_2028, w_009_2030, w_009_2031, w_009_2032, w_009_2033, w_009_2034, w_009_2035, w_009_2036, w_009_2037, w_009_2038, w_009_2039, w_009_2040, w_009_2041, w_009_2042, w_009_2043, w_009_2044, w_009_2045, w_009_2046, w_009_2047, w_009_2048, w_009_2049, w_009_2050, w_009_2051, w_009_2052, w_009_2053, w_009_2054, w_009_2055, w_009_2056, w_009_2057, w_009_2058, w_009_2059, w_009_2060, w_009_2063, w_009_2064, w_009_2065, w_009_2066, w_009_2067, w_009_2068, w_009_2069, w_009_2070, w_009_2071, w_009_2072, w_009_2073, w_009_2074, w_009_2075, w_009_2077, w_009_2078, w_009_2079, w_009_2080, w_009_2081, w_009_2082, w_009_2083, w_009_2084, w_009_2085, w_009_2086, w_009_2087, w_009_2088, w_009_2089, w_009_2090, w_009_2091, w_009_2092, w_009_2093, w_009_2095, w_009_2096, w_009_2097, w_009_2098, w_009_2099, w_009_2100, w_009_2101, w_009_2102, w_009_2103, w_009_2105, w_009_2106, w_009_2107, w_009_2108, w_009_2110, w_009_2111, w_009_2112, w_009_2113, w_009_2114, w_009_2115, w_009_2116, w_009_2117, w_009_2118, w_009_2119, w_009_2120, w_009_2121, w_009_2122, w_009_2123, w_009_2124, w_009_2125, w_009_2126, w_009_2127, w_009_2128, w_009_2129, w_009_2130, w_009_2131, w_009_2132, w_009_2133, w_009_2134, w_009_2135, w_009_2136, w_009_2137, w_009_2138, w_009_2139, w_009_2141, w_009_2142, w_009_2143, w_009_2144, w_009_2145, w_009_2146, w_009_2147, w_009_2148, w_009_2149, w_009_2150, w_009_2151, w_009_2152, w_009_2153, w_009_2154, w_009_2155, w_009_2156, w_009_2157, w_009_2158, w_009_2160, w_009_2161, w_009_2162, w_009_2163, w_009_2164, w_009_2165, w_009_2166, w_009_2167, w_009_2168, w_009_2169, w_009_2170, w_009_2171, w_009_2172, w_009_2173, w_009_2174, w_009_2175, w_009_2176, w_009_2177, w_009_2178, w_009_2179, w_009_2180, w_009_2181, w_009_2182, w_009_2183, w_009_2184, w_009_2185, w_009_2186, w_009_2187, w_009_2188, w_009_2189, w_009_2190, w_009_2191, w_009_2192, w_009_2193, w_009_2194, w_009_2195, w_009_2196, w_009_2197, w_009_2199, w_009_2200, w_009_2201, w_009_2202, w_009_2203, w_009_2204, w_009_2205, w_009_2206, w_009_2208, w_009_2209, w_009_2210, w_009_2211, w_009_2212, w_009_2213, w_009_2214, w_009_2215, w_009_2216, w_009_2217, w_009_2218, w_009_2219, w_009_2220, w_009_2221, w_009_2222, w_009_2223, w_009_2224, w_009_2225, w_009_2226, w_009_2227, w_009_2228, w_009_2229, w_009_2230, w_009_2231, w_009_2232, w_009_2233, w_009_2235, w_009_2236, w_009_2237, w_009_2238, w_009_2239, w_009_2240, w_009_2241, w_009_2242, w_009_2243, w_009_2244, w_009_2245, w_009_2246, w_009_2247, w_009_2248, w_009_2249, w_009_2250, w_009_2251, w_009_2252, w_009_2253, w_009_2254, w_009_2255, w_009_2256, w_009_2257, w_009_2258, w_009_2259, w_009_2260, w_009_2261, w_009_2262, w_009_2263, w_009_2264, w_009_2265, w_009_2266, w_009_2267, w_009_2268, w_009_2269, w_009_2270, w_009_2271, w_009_2272, w_009_2273, w_009_2274, w_009_2275, w_009_2276, w_009_2277, w_009_2278, w_009_2279, w_009_2280, w_009_2281, w_009_2282, w_009_2283, w_009_2284, w_009_2285, w_009_2286, w_009_2287, w_009_2288, w_009_2289, w_009_2290, w_009_2292, w_009_2294, w_009_2295, w_009_2296, w_009_2297, w_009_2298, w_009_2299, w_009_2300, w_009_2301, w_009_2302, w_009_2303, w_009_2304, w_009_2305, w_009_2306, w_009_2307, w_009_2308, w_009_2309, w_009_2310, w_009_2311, w_009_2312, w_009_2313, w_009_2314, w_009_2315, w_009_2316, w_009_2317, w_009_2318, w_009_2319, w_009_2321, w_009_2323, w_009_2324, w_009_2325, w_009_2326, w_009_2327, w_009_2328, w_009_2329, w_009_2330, w_009_2331, w_009_2332, w_009_2333, w_009_2334, w_009_2335, w_009_2336, w_009_2337, w_009_2338, w_009_2339, w_009_2340, w_009_2341, w_009_2342, w_009_2343, w_009_2344, w_009_2345, w_009_2346, w_009_2347, w_009_2348, w_009_2349, w_009_2350, w_009_2351, w_009_2352, w_009_2353, w_009_2354, w_009_2355, w_009_2356, w_009_2357, w_009_2358, w_009_2359, w_009_2360, w_009_2361, w_009_2362, w_009_2363, w_009_2364, w_009_2365, w_009_2366, w_009_2367, w_009_2368, w_009_2369, w_009_2370, w_009_2371, w_009_2372, w_009_2373, w_009_2374, w_009_2375, w_009_2376, w_009_2377, w_009_2378, w_009_2379, w_009_2380, w_009_2381, w_009_2382, w_009_2383, w_009_2385, w_009_2386, w_009_2387, w_009_2389, w_009_2390, w_009_2391, w_009_2392, w_009_2393, w_009_2394, w_009_2395, w_009_2396, w_009_2397, w_009_2398, w_009_2399, w_009_2400, w_009_2401, w_009_2402, w_009_2403, w_009_2404, w_009_2405, w_009_2406, w_009_2407, w_009_2408, w_009_2409, w_009_2410, w_009_2411, w_009_2412, w_009_2413, w_009_2414, w_009_2415, w_009_2416, w_009_2417, w_009_2418, w_009_2419, w_009_2420, w_009_2421, w_009_2422, w_009_2423, w_009_2424, w_009_2425, w_009_2426, w_009_2427, w_009_2429, w_009_2430, w_009_2431, w_009_2432, w_009_2433, w_009_2434, w_009_2435, w_009_2436, w_009_2437, w_009_2438, w_009_2439, w_009_2440, w_009_2441, w_009_2442, w_009_2443, w_009_2444, w_009_2445, w_009_2446, w_009_2447, w_009_2448, w_009_2449, w_009_2450, w_009_2451, w_009_2452, w_009_2453, w_009_2454, w_009_2455, w_009_2456, w_009_2457, w_009_2458, w_009_2459, w_009_2460, w_009_2462, w_009_2463, w_009_2464, w_009_2465, w_009_2466, w_009_2467, w_009_2468, w_009_2469, w_009_2471, w_009_2472, w_009_2473, w_009_2474, w_009_2475, w_009_2476, w_009_2477, w_009_2478, w_009_2479, w_009_2480, w_009_2481, w_009_2482, w_009_2483, w_009_2484, w_009_2485, w_009_2486, w_009_2487, w_009_2489, w_009_2490, w_009_2491, w_009_2492, w_009_2493, w_009_2494, w_009_2495, w_009_2496, w_009_2497, w_009_2498, w_009_2499, w_009_2500, w_009_2501, w_009_2502, w_009_2503, w_009_2504, w_009_2505, w_009_2506, w_009_2507, w_009_2508, w_009_2509, w_009_2510, w_009_2511, w_009_2512, w_009_2513, w_009_2514, w_009_2515, w_009_2516, w_009_2517, w_009_2518, w_009_2519, w_009_2520, w_009_2521, w_009_2522, w_009_2523, w_009_2524, w_009_2525, w_009_2526, w_009_2527, w_009_2528, w_009_2529, w_009_2530, w_009_2531, w_009_2532, w_009_2533, w_009_2534, w_009_2535, w_009_2536, w_009_2537, w_009_2538, w_009_2539, w_009_2541, w_009_2542, w_009_2543, w_009_2544, w_009_2545, w_009_2546, w_009_2547, w_009_2548, w_009_2549, w_009_2550, w_009_2551, w_009_2552, w_009_2553, w_009_2554, w_009_2555, w_009_2556, w_009_2557, w_009_2558, w_009_2559, w_009_2560, w_009_2561, w_009_2562, w_009_2563, w_009_2564, w_009_2565, w_009_2567, w_009_2568, w_009_2569, w_009_2570, w_009_2571, w_009_2572, w_009_2573, w_009_2574, w_009_2575, w_009_2576, w_009_2577, w_009_2578, w_009_2579, w_009_2580, w_009_2581, w_009_2582, w_009_2583, w_009_2585, w_009_2586, w_009_2587, w_009_2588, w_009_2589, w_009_2590, w_009_2591, w_009_2593, w_009_2594, w_009_2595, w_009_2596, w_009_2597, w_009_2598, w_009_2599, w_009_2600, w_009_2601, w_009_2602, w_009_2603, w_009_2604, w_009_2605, w_009_2606, w_009_2607, w_009_2608, w_009_2609, w_009_2610, w_009_2611, w_009_2612, w_009_2613, w_009_2614, w_009_2615, w_009_2616, w_009_2617, w_009_2618, w_009_2619, w_009_2620, w_009_2621, w_009_2622, w_009_2623, w_009_2624, w_009_2625, w_009_2626, w_009_2627, w_009_2628, w_009_2629, w_009_2630, w_009_2631, w_009_2632, w_009_2633, w_009_2634, w_009_2635, w_009_2636, w_009_2637, w_009_2638, w_009_2639, w_009_2640, w_009_2641, w_009_2642, w_009_2643, w_009_2644, w_009_2646, w_009_2647, w_009_2648, w_009_2649, w_009_2650, w_009_2651, w_009_2652, w_009_2653, w_009_2654, w_009_2655, w_009_2656, w_009_2657, w_009_2658, w_009_2659, w_009_2660, w_009_2661, w_009_2662, w_009_2663, w_009_2664, w_009_2665, w_009_2666, w_009_2667, w_009_2668, w_009_2669, w_009_2670, w_009_2671, w_009_2672, w_009_2673, w_009_2674, w_009_2675, w_009_2676, w_009_2677, w_009_2678, w_009_2679, w_009_2680, w_009_2681, w_009_2682, w_009_2683, w_009_2684, w_009_2686, w_009_2687, w_009_2688, w_009_2689, w_009_2690, w_009_2691, w_009_2692, w_009_2693, w_009_2694, w_009_2696, w_009_2697, w_009_2698, w_009_2699, w_009_2700, w_009_2701, w_009_2703, w_009_2704, w_009_2705, w_009_2708, w_009_2709, w_009_2710, w_009_2711, w_009_2712, w_009_2713, w_009_2714, w_009_2715, w_009_2716, w_009_2717, w_009_2718, w_009_2719, w_009_2720, w_009_2721, w_009_2722, w_009_2723, w_009_2724, w_009_2725, w_009_2726, w_009_2727, w_009_2728, w_009_2729, w_009_2730, w_009_2731, w_009_2732, w_009_2733, w_009_2734, w_009_2735, w_009_2736, w_009_2737, w_009_2738, w_009_2739, w_009_2740, w_009_2741, w_009_2742, w_009_2743, w_009_2744, w_009_2745, w_009_2746, w_009_2747, w_009_2748, w_009_2749, w_009_2750, w_009_2751, w_009_2752, w_009_2753, w_009_2754, w_009_2755, w_009_2756, w_009_2758, w_009_2759, w_009_2760, w_009_2761, w_009_2762, w_009_2763, w_009_2764, w_009_2765, w_009_2766, w_009_2767, w_009_2768, w_009_2769, w_009_2770, w_009_2771, w_009_2772, w_009_2773, w_009_2774, w_009_2776, w_009_2777, w_009_2778, w_009_2779, w_009_2781, w_009_2782, w_009_2783, w_009_2784, w_009_2785, w_009_2786, w_009_2787, w_009_2788, w_009_2789, w_009_2790, w_009_2791, w_009_2792, w_009_2793, w_009_2795, w_009_2796, w_009_2797, w_009_2798, w_009_2799, w_009_2800, w_009_2801, w_009_2802, w_009_2803, w_009_2804, w_009_2805, w_009_2806, w_009_2807, w_009_2808, w_009_2809, w_009_2810, w_009_2811, w_009_2812, w_009_2813, w_009_2814, w_009_2815, w_009_2816, w_009_2817, w_009_2818, w_009_2819, w_009_2820, w_009_2821, w_009_2822, w_009_2823, w_009_2824, w_009_2825, w_009_2826, w_009_2827, w_009_2828, w_009_2829, w_009_2830, w_009_2831, w_009_2832, w_009_2833, w_009_2834, w_009_2835, w_009_2836, w_009_2837, w_009_2838, w_009_2840, w_009_2841, w_009_2842, w_009_2843, w_009_2844, w_009_2845, w_009_2846, w_009_2847, w_009_2848, w_009_2849, w_009_2850, w_009_2851, w_009_2852, w_009_2853, w_009_2854, w_009_2855, w_009_2856, w_009_2857, w_009_2858, w_009_2859, w_009_2860, w_009_2861, w_009_2862, w_009_2863, w_009_2864, w_009_2865, w_009_2866, w_009_2867, w_009_2868, w_009_2869, w_009_2870, w_009_2871, w_009_2872, w_009_2873, w_009_2874, w_009_2875, w_009_2876, w_009_2877, w_009_2878, w_009_2879, w_009_2880, w_009_2881, w_009_2883, w_009_2884, w_009_2885, w_009_2886, w_009_2887, w_009_2888, w_009_2889, w_009_2890, w_009_2891, w_009_2892, w_009_2893, w_009_2894, w_009_2896, w_009_2897, w_009_2900, w_009_2901, w_009_2902, w_009_2903, w_009_2904, w_009_2905, w_009_2906, w_009_2907, w_009_2908, w_009_2909, w_009_2910, w_009_2911, w_009_2912, w_009_2913, w_009_2914, w_009_2915, w_009_2916, w_009_2917, w_009_2918, w_009_2919, w_009_2920, w_009_2921, w_009_2922, w_009_2923, w_009_2924, w_009_2925, w_009_2926, w_009_2927, w_009_2928, w_009_2929, w_009_2930, w_009_2931, w_009_2932, w_009_2933, w_009_2934, w_009_2935, w_009_2936, w_009_2937, w_009_2938, w_009_2939, w_009_2940, w_009_2941, w_009_2942, w_009_2943, w_009_2944, w_009_2945, w_009_2946, w_009_2947, w_009_2948, w_009_2949, w_009_2950, w_009_2951, w_009_2953, w_009_2954, w_009_2955, w_009_2956, w_009_2957, w_009_2958, w_009_2959, w_009_2960, w_009_2961, w_009_2962, w_009_2963, w_009_2964, w_009_2965, w_009_2966, w_009_2967, w_009_2968, w_009_2969, w_009_2971, w_009_2972, w_009_2973, w_009_2974, w_009_2975, w_009_2976, w_009_2977, w_009_2978, w_009_2979, w_009_2980, w_009_2981, w_009_2982, w_009_2983, w_009_2984, w_009_2985, w_009_2986, w_009_2987, w_009_2988, w_009_2990, w_009_2991, w_009_2992, w_009_2993, w_009_2994, w_009_2995, w_009_2996, w_009_2997, w_009_2998, w_009_2999, w_009_3000, w_009_3001, w_009_3002, w_009_3003, w_009_3004, w_009_3005, w_009_3006, w_009_3007, w_009_3008, w_009_3009, w_009_3010, w_009_3011, w_009_3012, w_009_3013, w_009_3014, w_009_3015, w_009_3016, w_009_3017, w_009_3019, w_009_3020, w_009_3021, w_009_3022, w_009_3023, w_009_3024, w_009_3026, w_009_3027, w_009_3028, w_009_3029, w_009_3030, w_009_3031, w_009_3032, w_009_3033, w_009_3034, w_009_3035, w_009_3036, w_009_3037, w_009_3038, w_009_3039, w_009_3040, w_009_3041, w_009_3042, w_009_3043, w_009_3044, w_009_3045, w_009_3046, w_009_3047, w_009_3049, w_009_3050, w_009_3052, w_009_3053, w_009_3054, w_009_3055, w_009_3056, w_009_3057, w_009_3058, w_009_3059, w_009_3060, w_009_3061, w_009_3062, w_009_3063, w_009_3064, w_009_3065, w_009_3066, w_009_3067, w_009_3069, w_009_3070, w_009_3071, w_009_3073, w_009_3074, w_009_3075, w_009_3076, w_009_3077, w_009_3078, w_009_3079, w_009_3080, w_009_3081, w_009_3082, w_009_3083, w_009_3084, w_009_3085, w_009_3086, w_009_3087, w_009_3088, w_009_3089, w_009_3090, w_009_3091, w_009_3092, w_009_3093, w_009_3094, w_009_3095, w_009_3096, w_009_3097, w_009_3098, w_009_3099, w_009_3100, w_009_3102, w_009_3103, w_009_3104, w_009_3105, w_009_3107, w_009_3109, w_009_3110, w_009_3111, w_009_3112, w_009_3113, w_009_3115, w_009_3116, w_009_3117, w_009_3118, w_009_3119, w_009_3120, w_009_3121, w_009_3122, w_009_3123, w_009_3124, w_009_3125, w_009_3126, w_009_3127, w_009_3128, w_009_3129, w_009_3130, w_009_3131, w_009_3132, w_009_3133, w_009_3134, w_009_3136, w_009_3137, w_009_3138, w_009_3139, w_009_3140, w_009_3141, w_009_3142, w_009_3143, w_009_3144, w_009_3145, w_009_3146, w_009_3147, w_009_3148, w_009_3149, w_009_3150, w_009_3151, w_009_3152, w_009_3153, w_009_3154, w_009_3155, w_009_3156, w_009_3157, w_009_3158, w_009_3159, w_009_3160, w_009_3161, w_009_3162, w_009_3163, w_009_3164, w_009_3165, w_009_3166, w_009_3167, w_009_3168, w_009_3169, w_009_3170, w_009_3171, w_009_3172, w_009_3173, w_009_3174, w_009_3175, w_009_3176, w_009_3177, w_009_3178, w_009_3179, w_009_3180, w_009_3181, w_009_3182, w_009_3183, w_009_3184, w_009_3185, w_009_3186, w_009_3187, w_009_3188, w_009_3189, w_009_3190, w_009_3191, w_009_3192, w_009_3193, w_009_3194, w_009_3195, w_009_3196, w_009_3197, w_009_3198, w_009_3199, w_009_3200, w_009_3201, w_009_3202, w_009_3203, w_009_3204, w_009_3205, w_009_3206, w_009_3207, w_009_3208, w_009_3209, w_009_3210, w_009_3211, w_009_3212, w_009_3213, w_009_3214, w_009_3215, w_009_3216, w_009_3217, w_009_3218, w_009_3219, w_009_3220, w_009_3221, w_009_3222, w_009_3223, w_009_3224, w_009_3225, w_009_3226, w_009_3227, w_009_3228, w_009_3230, w_009_3232, w_009_3233, w_009_3234, w_009_3235, w_009_3236, w_009_3237, w_009_3238, w_009_3239, w_009_3240, w_009_3241, w_009_3242, w_009_3243, w_009_3244, w_009_3245, w_009_3247, w_009_3248, w_009_3249, w_009_3250, w_009_3251, w_009_3252, w_009_3253, w_009_3254, w_009_3255, w_009_3256, w_009_3257, w_009_3258, w_009_3259, w_009_3260, w_009_3261, w_009_3262, w_009_3263, w_009_3264, w_009_3265, w_009_3266, w_009_3267, w_009_3268, w_009_3269, w_009_3270, w_009_3271, w_009_3273, w_009_3274, w_009_3275, w_009_3276, w_009_3277, w_009_3278, w_009_3279, w_009_3280, w_009_3281, w_009_3282, w_009_3283, w_009_3284, w_009_3285, w_009_3287, w_009_3288, w_009_3289, w_009_3290, w_009_3291, w_009_3292, w_009_3293, w_009_3294, w_009_3295, w_009_3296, w_009_3297, w_009_3299, w_009_3300, w_009_3301, w_009_3302, w_009_3303, w_009_3304, w_009_3305, w_009_3306, w_009_3307, w_009_3308, w_009_3309, w_009_3311, w_009_3312, w_009_3313, w_009_3314, w_009_3315, w_009_3316, w_009_3317, w_009_3318, w_009_3319, w_009_3320, w_009_3321, w_009_3322, w_009_3323, w_009_3324, w_009_3325, w_009_3326, w_009_3327, w_009_3328, w_009_3329, w_009_3330, w_009_3331, w_009_3333, w_009_3335, w_009_3336, w_009_3337, w_009_3338, w_009_3339, w_009_3340, w_009_3342, w_009_3343, w_009_3344, w_009_3345, w_009_3346, w_009_3347, w_009_3348, w_009_3350, w_009_3351, w_009_3352, w_009_3353, w_009_3354, w_009_3355, w_009_3356, w_009_3357, w_009_3358, w_009_3359, w_009_3360, w_009_3361, w_009_3362, w_009_3363, w_009_3364, w_009_3365, w_009_3367, w_009_3368, w_009_3369, w_009_3370, w_009_3371, w_009_3372, w_009_3373, w_009_3374, w_009_3375, w_009_3376, w_009_3377, w_009_3378, w_009_3379, w_009_3380, w_009_3381, w_009_3382, w_009_3383, w_009_3385, w_009_3386, w_009_3387, w_009_3388, w_009_3389, w_009_3390, w_009_3391, w_009_3392, w_009_3393, w_009_3394, w_009_3395, w_009_3396, w_009_3397, w_009_3398, w_009_3399, w_009_3400, w_009_3401, w_009_3402, w_009_3403, w_009_3404, w_009_3405, w_009_3406, w_009_3407, w_009_3408, w_009_3409, w_009_3410, w_009_3411, w_009_3412, w_009_3413, w_009_3414, w_009_3415, w_009_3416, w_009_3417, w_009_3418, w_009_3419, w_009_3420, w_009_3421, w_009_3422, w_009_3423, w_009_3424, w_009_3425, w_009_3426, w_009_3427, w_009_3428, w_009_3429, w_009_3430, w_009_3431, w_009_3432, w_009_3433, w_009_3434, w_009_3436, w_009_3437, w_009_3438, w_009_3439, w_009_3440, w_009_3442, w_009_3444, w_009_3445, w_009_3446, w_009_3447, w_009_3448, w_009_3449, w_009_3450, w_009_3451, w_009_3452, w_009_3453, w_009_3454, w_009_3455, w_009_3456, w_009_3457, w_009_3458, w_009_3459, w_009_3460, w_009_3461, w_009_3462, w_009_3463, w_009_3464, w_009_3465, w_009_3466, w_009_3467, w_009_3468, w_009_3469, w_009_3470, w_009_3471, w_009_3472, w_009_3473, w_009_3474, w_009_3476, w_009_3477, w_009_3478, w_009_3479, w_009_3480, w_009_3481, w_009_3482, w_009_3483, w_009_3484, w_009_3485, w_009_3486, w_009_3488, w_009_3489, w_009_3490, w_009_3491, w_009_3492, w_009_3493, w_009_3494, w_009_3495, w_009_3496, w_009_3497, w_009_3498, w_009_3500, w_009_3501, w_009_3502, w_009_3503, w_009_3504, w_009_3505, w_009_3506, w_009_3507, w_009_3508, w_009_3509, w_009_3510, w_009_3511, w_009_3512, w_009_3513, w_009_3514, w_009_3515, w_009_3516, w_009_3517, w_009_3518, w_009_3519, w_009_3520, w_009_3521, w_009_3522, w_009_3523, w_009_3524, w_009_3525, w_009_3526, w_009_3527, w_009_3528, w_009_3529, w_009_3530, w_009_3531, w_009_3532, w_009_3533, w_009_3534, w_009_3536, w_009_3537, w_009_3538, w_009_3539, w_009_3540, w_009_3542, w_009_3543, w_009_3544, w_009_3546, w_009_3547, w_009_3548, w_009_3549, w_009_3550, w_009_3551, w_009_3553, w_009_3554, w_009_3555, w_009_3556, w_009_3557, w_009_3558, w_009_3559, w_009_3561, w_009_3562, w_009_3563, w_009_3564, w_009_3565, w_009_3566, w_009_3567, w_009_3568, w_009_3569, w_009_3570, w_009_3571, w_009_3572, w_009_3573, w_009_3574, w_009_3575, w_009_3576, w_009_3577, w_009_3578, w_009_3581, w_009_3582, w_009_3583, w_009_3584, w_009_3585, w_009_3586, w_009_3587, w_009_3588, w_009_3589, w_009_3590, w_009_3591, w_009_3592, w_009_3593, w_009_3594, w_009_3595, w_009_3596, w_009_3597, w_009_3598, w_009_3599, w_009_3600, w_009_3601, w_009_3602, w_009_3603, w_009_3604, w_009_3605, w_009_3606, w_009_3607, w_009_3608, w_009_3609, w_009_3610, w_009_3611, w_009_3612, w_009_3613, w_009_3614, w_009_3615, w_009_3617, w_009_3618, w_009_3619, w_009_3620, w_009_3621, w_009_3622, w_009_3623, w_009_3625, w_009_3626, w_009_3627, w_009_3628, w_009_3629, w_009_3630, w_009_3631, w_009_3632, w_009_3633, w_009_3634, w_009_3635, w_009_3636, w_009_3637, w_009_3638, w_009_3639, w_009_3640, w_009_3641, w_009_3642, w_009_3643, w_009_3645, w_009_3646, w_009_3648, w_009_3649, w_009_3650, w_009_3651, w_009_3652, w_009_3654, w_009_3655, w_009_3656, w_009_3657, w_009_3658, w_009_3659, w_009_3660, w_009_3661, w_009_3662, w_009_3663, w_009_3664, w_009_3665, w_009_3667, w_009_3668, w_009_3669, w_009_3670, w_009_3671, w_009_3672, w_009_3673, w_009_3674, w_009_3675, w_009_3676, w_009_3677, w_009_3679, w_009_3680, w_009_3681, w_009_3683, w_009_3684, w_009_3685, w_009_3686, w_009_3687, w_009_3688, w_009_3689, w_009_3690, w_009_3691, w_009_3692, w_009_3694, w_009_3695, w_009_3696, w_009_3697, w_009_3698, w_009_3699, w_009_3700, w_009_3701, w_009_3702, w_009_3703, w_009_3704, w_009_3705, w_009_3706, w_009_3707, w_009_3708, w_009_3709, w_009_3710, w_009_3711, w_009_3712, w_009_3713, w_009_3714, w_009_3715, w_009_3716, w_009_3717, w_009_3718, w_009_3719, w_009_3720, w_009_3721, w_009_3722, w_009_3723, w_009_3724, w_009_3725, w_009_3726, w_009_3727, w_009_3728, w_009_3729, w_009_3730, w_009_3731, w_009_3732, w_009_3733, w_009_3734, w_009_3735, w_009_3736, w_009_3737, w_009_3738, w_009_3739, w_009_3740, w_009_3741, w_009_3742, w_009_3743, w_009_3744, w_009_3745, w_009_3746, w_009_3747, w_009_3749, w_009_3750, w_009_3751, w_009_3752, w_009_3754, w_009_3755, w_009_3756, w_009_3757, w_009_3758, w_009_3759, w_009_3760, w_009_3761, w_009_3763, w_009_3764, w_009_3765, w_009_3766, w_009_3767, w_009_3768, w_009_3769, w_009_3770, w_009_3771, w_009_3772, w_009_3773, w_009_3774, w_009_3775, w_009_3776, w_009_3777, w_009_3778, w_009_3779, w_009_3780, w_009_3781, w_009_3782, w_009_3783, w_009_3784, w_009_3785, w_009_3786, w_009_3787, w_009_3788, w_009_3789, w_009_3791, w_009_3792, w_009_3793, w_009_3794, w_009_3795, w_009_3796, w_009_3797, w_009_3798, w_009_3799, w_009_3800, w_009_3801, w_009_3802, w_009_3803, w_009_3804, w_009_3805, w_009_3806, w_009_3807, w_009_3809, w_009_3810, w_009_3811, w_009_3812, w_009_3813, w_009_3814, w_009_3815, w_009_3816, w_009_3817, w_009_3818, w_009_3819, w_009_3820, w_009_3821, w_009_3822, w_009_3823, w_009_3824, w_009_3825, w_009_3826, w_009_3827, w_009_3828, w_009_3829, w_009_3830, w_009_3832, w_009_3833, w_009_3834, w_009_3835, w_009_3836, w_009_3837, w_009_3838, w_009_3839, w_009_3840, w_009_3841, w_009_3842, w_009_3843, w_009_3844, w_009_3845, w_009_3846, w_009_3847, w_009_3848, w_009_3849, w_009_3850, w_009_3851, w_009_3852, w_009_3853, w_009_3854, w_009_3855, w_009_3856, w_009_3857, w_009_3858, w_009_3859, w_009_3860, w_009_3861, w_009_3862, w_009_3863, w_009_3864, w_009_3865, w_009_3866, w_009_3867, w_009_3868, w_009_3869, w_009_3870, w_009_3871, w_009_3872, w_009_3873, w_009_3874, w_009_3875, w_009_3876, w_009_3877, w_009_3878, w_009_3879, w_009_3880, w_009_3882, w_009_3883, w_009_3884, w_009_3885, w_009_3886, w_009_3887, w_009_3888, w_009_3889, w_009_3890, w_009_3891, w_009_3892, w_009_3894, w_009_3895, w_009_3896, w_009_3897, w_009_3898, w_009_3899, w_009_3900, w_009_3901, w_009_3902, w_009_3903, w_009_3904, w_009_3905, w_009_3906, w_009_3907, w_009_3908, w_009_3909, w_009_3910, w_009_3911, w_009_3912, w_009_3913, w_009_3914, w_009_3915, w_009_3916, w_009_3917, w_009_3918, w_009_3919, w_009_3920, w_009_3921, w_009_3922, w_009_3923, w_009_3924, w_009_3925, w_009_3926, w_009_3927, w_009_3928, w_009_3929, w_009_3930, w_009_3931, w_009_3932, w_009_3933, w_009_3934, w_009_3935, w_009_3936, w_009_3937, w_009_3938, w_009_3939, w_009_3940, w_009_3942, w_009_3943, w_009_3944, w_009_3945, w_009_3946, w_009_3947, w_009_3948, w_009_3949, w_009_3950, w_009_3951, w_009_3952, w_009_3953, w_009_3954, w_009_3955, w_009_3956, w_009_3957, w_009_3959, w_009_3960, w_009_3961, w_009_3962, w_009_3963, w_009_3964, w_009_3965, w_009_3967, w_009_3968, w_009_3969, w_009_3970, w_009_3971, w_009_3972, w_009_3973, w_009_3974, w_009_3975, w_009_3976, w_009_3977, w_009_3978, w_009_3979, w_009_3980, w_009_3981, w_009_3982, w_009_3983, w_009_3984, w_009_3985, w_009_3986, w_009_3987, w_009_3988, w_009_3989, w_009_3990, w_009_3991, w_009_3992, w_009_3993, w_009_3994, w_009_3995, w_009_3996, w_009_3997, w_009_3998, w_009_3999, w_009_4000, w_009_4001, w_009_4002, w_009_4003, w_009_4004, w_009_4005, w_009_4006, w_009_4007, w_009_4008, w_009_4009, w_009_4010, w_009_4011, w_009_4012, w_009_4013, w_009_4014, w_009_4015, w_009_4016, w_009_4017, w_009_4018, w_009_4019, w_009_4021, w_009_4022, w_009_4023, w_009_4024, w_009_4025, w_009_4026, w_009_4027, w_009_4028, w_009_4029, w_009_4030, w_009_4031, w_009_4032, w_009_4033, w_009_4034, w_009_4035, w_009_4036, w_009_4037, w_009_4038, w_009_4039, w_009_4040, w_009_4041, w_009_4042, w_009_4043, w_009_4045, w_009_4046, w_009_4048, w_009_4049, w_009_4050, w_009_4051, w_009_4052, w_009_4053, w_009_4054, w_009_4055, w_009_4056, w_009_4057, w_009_4058, w_009_4059, w_009_4060, w_009_4061, w_009_4062, w_009_4063, w_009_4064, w_009_4065, w_009_4066, w_009_4067, w_009_4068, w_009_4069, w_009_4070, w_009_4071, w_009_4072, w_009_4073, w_009_4074, w_009_4075, w_009_4076, w_009_4077, w_009_4078, w_009_4079, w_009_4080, w_009_4081, w_009_4082, w_009_4083, w_009_4084, w_009_4085, w_009_4086, w_009_4087, w_009_4088, w_009_4089, w_009_4090, w_009_4091, w_009_4092, w_009_4093, w_009_4095, w_009_4096, w_009_4097, w_009_4098, w_009_4099, w_009_4100, w_009_4101, w_009_4102, w_009_4103, w_009_4104, w_009_4105, w_009_4106, w_009_4107, w_009_4108, w_009_4109, w_009_4110, w_009_4111, w_009_4112, w_009_4113, w_009_4114, w_009_4115, w_009_4116, w_009_4118, w_009_4119, w_009_4120, w_009_4122, w_009_4123, w_009_4124, w_009_4125, w_009_4126, w_009_4127, w_009_4128, w_009_4129, w_009_4130, w_009_4131, w_009_4132, w_009_4133, w_009_4134, w_009_4135, w_009_4136, w_009_4137, w_009_4138, w_009_4139, w_009_4140, w_009_4141, w_009_4142, w_009_4143, w_009_4144, w_009_4145, w_009_4146, w_009_4147, w_009_4148, w_009_4149, w_009_4150, w_009_4151, w_009_4152, w_009_4153, w_009_4154, w_009_4155, w_009_4156, w_009_4157, w_009_4158, w_009_4159, w_009_4160, w_009_4161, w_009_4162, w_009_4163, w_009_4164, w_009_4165, w_009_4166, w_009_4167, w_009_4168, w_009_4169, w_009_4170, w_009_4171, w_009_4172, w_009_4173, w_009_4174, w_009_4176, w_009_4177, w_009_4179, w_009_4180, w_009_4181, w_009_4182, w_009_4183, w_009_4184, w_009_4185, w_009_4186, w_009_4187, w_009_4188, w_009_4189, w_009_4190, w_009_4191, w_009_4192, w_009_4193, w_009_4194, w_009_4195, w_009_4196, w_009_4197, w_009_4198, w_009_4199, w_009_4200, w_009_4201, w_009_4202, w_009_4203, w_009_4204, w_009_4205, w_009_4206, w_009_4207, w_009_4208, w_009_4209, w_009_4210, w_009_4211, w_009_4213, w_009_4214, w_009_4215, w_009_4216, w_009_4217, w_009_4218, w_009_4219, w_009_4220, w_009_4221, w_009_4222, w_009_4223, w_009_4224, w_009_4225, w_009_4226, w_009_4227, w_009_4228, w_009_4229, w_009_4230, w_009_4231, w_009_4232, w_009_4233, w_009_4234, w_009_4235, w_009_4236, w_009_4237, w_009_4238, w_009_4239, w_009_4240, w_009_4241, w_009_4242, w_009_4243, w_009_4244, w_009_4245, w_009_4246, w_009_4247, w_009_4248, w_009_4249, w_009_4250, w_009_4251, w_009_4252, w_009_4253, w_009_4254, w_009_4255, w_009_4256, w_009_4257, w_009_4258, w_009_4259, w_009_4260, w_009_4261, w_009_4262, w_009_4263, w_009_4264, w_009_4265, w_009_4266, w_009_4267, w_009_4268, w_009_4269, w_009_4270, w_009_4271, w_009_4272, w_009_4273, w_009_4274, w_009_4275, w_009_4276, w_009_4277, w_009_4278, w_009_4279, w_009_4280, w_009_4281, w_009_4282, w_009_4283, w_009_4284, w_009_4285, w_009_4286, w_009_4287, w_009_4288, w_009_4289, w_009_4290, w_009_4291, w_009_4293, w_009_4294, w_009_4295, w_009_4296, w_009_4297, w_009_4298, w_009_4299, w_009_4300, w_009_4301, w_009_4302, w_009_4303, w_009_4304, w_009_4305, w_009_4306, w_009_4307, w_009_4308, w_009_4309, w_009_4310, w_009_4311, w_009_4313, w_009_4314, w_009_4315, w_009_4316, w_009_4317, w_009_4318, w_009_4319, w_009_4320, w_009_4321, w_009_4322, w_009_4323, w_009_4324, w_009_4325, w_009_4326, w_009_4327, w_009_4328, w_009_4329, w_009_4330, w_009_4331, w_009_4332, w_009_4333, w_009_4334, w_009_4335, w_009_4336, w_009_4337, w_009_4338, w_009_4339, w_009_4340, w_009_4342, w_009_4343, w_009_4344, w_009_4345, w_009_4346, w_009_4347, w_009_4348, w_009_4349, w_009_4351, w_009_4352, w_009_4353, w_009_4354, w_009_4355, w_009_4356, w_009_4357, w_009_4358, w_009_4359, w_009_4360, w_009_4361, w_009_4362, w_009_4363, w_009_4364, w_009_4365, w_009_4366, w_009_4367, w_009_4368, w_009_4369, w_009_4370, w_009_4371, w_009_4372, w_009_4373, w_009_4374, w_009_4375, w_009_4376, w_009_4377, w_009_4378, w_009_4379, w_009_4380, w_009_4381, w_009_4382, w_009_4383, w_009_4384, w_009_4385, w_009_4387, w_009_4388, w_009_4389, w_009_4390, w_009_4391, w_009_4392, w_009_4393, w_009_4394, w_009_4395, w_009_4396, w_009_4397, w_009_4398, w_009_4399, w_009_4400, w_009_4401, w_009_4402, w_009_4403, w_009_4404, w_009_4405, w_009_4406, w_009_4407, w_009_4408, w_009_4409, w_009_4410, w_009_4411, w_009_4412, w_009_4413, w_009_4414, w_009_4416, w_009_4417, w_009_4418, w_009_4419, w_009_4420, w_009_4421, w_009_4422, w_009_4423, w_009_4424, w_009_4425, w_009_4426, w_009_4427, w_009_4428, w_009_4429, w_009_4430, w_009_4431, w_009_4432, w_009_4433, w_009_4434, w_009_4435, w_009_4436, w_009_4437, w_009_4438, w_009_4439, w_009_4440, w_009_4441, w_009_4442, w_009_4443, w_009_4444, w_009_4445, w_009_4446, w_009_4447, w_009_4448, w_009_4450, w_009_4451, w_009_4452, w_009_4453, w_009_4454, w_009_4455, w_009_4456, w_009_4457, w_009_4458, w_009_4459, w_009_4460, w_009_4461, w_009_4462, w_009_4463, w_009_4464, w_009_4465, w_009_4466, w_009_4467, w_009_4468, w_009_4469, w_009_4470, w_009_4472, w_009_4473, w_009_4474, w_009_4475, w_009_4476, w_009_4477, w_009_4478, w_009_4479, w_009_4480, w_009_4481, w_009_4482, w_009_4483, w_009_4484, w_009_4485, w_009_4487, w_009_4489, w_009_4490, w_009_4491, w_009_4492, w_009_4493, w_009_4494, w_009_4495, w_009_4496, w_009_4497, w_009_4498, w_009_4499, w_009_4500, w_009_4501, w_009_4502, w_009_4503, w_009_4504, w_009_4505, w_009_4506, w_009_4507, w_009_4508, w_009_4510, w_009_4511, w_009_4512, w_009_4513, w_009_4514, w_009_4515, w_009_4516, w_009_4517, w_009_4518, w_009_4520, w_009_4521, w_009_4522, w_009_4523, w_009_4524, w_009_4526, w_009_4527, w_009_4528, w_009_4529, w_009_4530, w_009_4531, w_009_4532, w_009_4533, w_009_4534, w_009_4535, w_009_4536, w_009_4537, w_009_4538, w_009_4539, w_009_4540, w_009_4541, w_009_4542, w_009_4543, w_009_4544;
  wire w_010_000, w_010_001, w_010_002, w_010_003, w_010_004, w_010_005, w_010_006, w_010_007, w_010_009, w_010_010, w_010_011, w_010_012, w_010_013, w_010_014, w_010_015, w_010_016, w_010_017, w_010_018, w_010_019, w_010_020, w_010_021, w_010_022, w_010_023, w_010_024, w_010_025, w_010_026, w_010_027, w_010_028, w_010_029, w_010_030, w_010_031, w_010_032, w_010_033, w_010_034, w_010_035, w_010_036, w_010_037, w_010_039, w_010_040, w_010_041, w_010_042, w_010_043, w_010_044, w_010_045, w_010_046, w_010_047, w_010_048, w_010_049, w_010_050, w_010_051, w_010_052, w_010_053, w_010_054, w_010_055, w_010_056, w_010_057, w_010_058, w_010_059, w_010_060, w_010_061, w_010_062, w_010_063, w_010_064, w_010_065, w_010_066, w_010_067, w_010_068, w_010_069, w_010_070, w_010_071, w_010_072, w_010_073, w_010_074, w_010_076, w_010_077, w_010_078, w_010_080, w_010_081, w_010_082, w_010_083, w_010_084, w_010_085, w_010_086, w_010_087, w_010_088, w_010_089, w_010_091, w_010_092, w_010_094, w_010_095, w_010_096, w_010_097, w_010_098, w_010_099, w_010_100, w_010_101, w_010_102, w_010_103, w_010_104, w_010_105, w_010_106, w_010_107, w_010_108, w_010_109, w_010_110, w_010_111, w_010_112, w_010_113, w_010_114, w_010_115, w_010_116, w_010_117, w_010_118, w_010_119, w_010_120, w_010_121, w_010_122, w_010_123, w_010_124, w_010_125, w_010_126, w_010_127, w_010_128, w_010_129, w_010_130, w_010_131, w_010_132, w_010_133, w_010_134, w_010_135, w_010_136, w_010_137, w_010_138, w_010_139, w_010_140, w_010_141, w_010_142, w_010_143, w_010_144, w_010_145, w_010_146, w_010_147, w_010_148, w_010_149, w_010_150, w_010_151, w_010_152, w_010_153, w_010_154, w_010_155, w_010_156, w_010_157, w_010_158, w_010_159, w_010_160, w_010_161, w_010_162, w_010_163, w_010_166, w_010_167, w_010_168, w_010_169, w_010_170, w_010_171, w_010_172, w_010_173, w_010_174, w_010_175, w_010_176, w_010_178, w_010_179, w_010_180, w_010_181, w_010_183, w_010_184, w_010_185, w_010_187, w_010_188, w_010_189, w_010_190, w_010_191, w_010_192, w_010_193, w_010_194, w_010_195, w_010_196, w_010_197, w_010_198, w_010_199, w_010_200, w_010_201, w_010_202, w_010_203, w_010_204, w_010_205, w_010_206, w_010_207, w_010_208, w_010_209, w_010_211, w_010_212, w_010_213, w_010_214, w_010_215, w_010_216, w_010_217, w_010_218, w_010_219, w_010_220, w_010_221, w_010_222, w_010_223, w_010_224, w_010_225, w_010_226, w_010_227, w_010_228, w_010_229, w_010_230, w_010_231, w_010_232, w_010_233, w_010_234, w_010_235, w_010_236, w_010_238, w_010_239, w_010_240, w_010_242, w_010_243, w_010_244, w_010_245, w_010_246, w_010_247, w_010_248, w_010_250, w_010_251, w_010_252, w_010_253, w_010_254, w_010_255, w_010_256, w_010_257, w_010_258, w_010_259, w_010_260, w_010_262, w_010_263, w_010_264, w_010_265, w_010_266, w_010_267, w_010_268, w_010_269, w_010_271, w_010_272, w_010_273, w_010_274, w_010_275, w_010_276, w_010_277, w_010_278, w_010_279, w_010_280, w_010_281, w_010_282, w_010_283, w_010_284, w_010_285, w_010_286, w_010_287, w_010_288, w_010_289, w_010_290, w_010_291, w_010_292, w_010_293, w_010_294, w_010_295, w_010_296, w_010_297, w_010_298, w_010_299, w_010_300, w_010_302, w_010_303, w_010_304, w_010_305, w_010_308, w_010_309, w_010_310, w_010_311, w_010_312, w_010_313, w_010_314, w_010_315, w_010_316, w_010_317, w_010_318, w_010_319, w_010_320, w_010_321, w_010_322, w_010_323, w_010_324, w_010_326, w_010_327, w_010_328, w_010_329, w_010_330, w_010_331, w_010_332, w_010_333, w_010_334, w_010_335, w_010_336, w_010_339, w_010_340, w_010_341, w_010_342, w_010_343, w_010_344, w_010_345, w_010_346, w_010_347, w_010_349, w_010_350, w_010_351, w_010_352, w_010_353, w_010_354, w_010_355, w_010_356, w_010_357, w_010_358, w_010_359, w_010_360, w_010_362, w_010_363, w_010_364, w_010_365, w_010_366, w_010_367, w_010_368, w_010_369, w_010_371, w_010_372, w_010_373, w_010_374, w_010_375, w_010_376, w_010_377, w_010_378, w_010_380, w_010_381, w_010_382, w_010_384, w_010_385, w_010_387, w_010_388, w_010_389, w_010_390, w_010_391, w_010_392, w_010_393, w_010_394, w_010_395, w_010_396, w_010_397, w_010_398, w_010_399, w_010_400, w_010_401, w_010_402, w_010_403, w_010_404, w_010_406, w_010_407, w_010_408, w_010_409, w_010_410, w_010_411, w_010_413, w_010_414, w_010_415, w_010_416, w_010_417, w_010_419, w_010_420, w_010_421, w_010_422, w_010_423, w_010_424, w_010_425, w_010_426, w_010_427, w_010_428, w_010_429, w_010_430, w_010_431, w_010_432, w_010_433, w_010_435, w_010_436, w_010_437, w_010_438, w_010_439, w_010_440, w_010_441, w_010_442, w_010_443, w_010_444, w_010_445, w_010_446, w_010_447, w_010_448, w_010_449, w_010_450, w_010_451, w_010_452, w_010_453, w_010_454, w_010_455, w_010_456, w_010_457, w_010_458, w_010_459, w_010_460, w_010_461, w_010_462, w_010_463, w_010_464, w_010_465, w_010_466, w_010_467, w_010_468, w_010_469, w_010_470, w_010_471, w_010_472, w_010_473, w_010_474, w_010_476, w_010_477, w_010_478, w_010_479, w_010_480, w_010_481, w_010_482, w_010_483, w_010_484, w_010_485, w_010_487, w_010_488, w_010_489, w_010_490, w_010_491, w_010_492, w_010_493, w_010_494, w_010_495, w_010_496, w_010_497, w_010_498, w_010_500, w_010_502, w_010_503, w_010_504, w_010_505, w_010_506, w_010_507, w_010_508, w_010_509, w_010_510, w_010_511, w_010_512, w_010_513, w_010_514, w_010_515, w_010_516, w_010_517, w_010_518, w_010_519, w_010_521, w_010_522, w_010_523, w_010_524, w_010_525, w_010_526, w_010_528, w_010_529, w_010_530, w_010_531, w_010_532, w_010_533, w_010_534, w_010_535, w_010_536, w_010_537, w_010_538, w_010_539, w_010_540, w_010_541, w_010_542, w_010_543, w_010_544, w_010_545, w_010_547, w_010_548, w_010_549, w_010_550, w_010_551, w_010_552, w_010_553, w_010_554, w_010_555, w_010_556, w_010_557, w_010_558, w_010_559, w_010_560, w_010_561, w_010_563, w_010_564, w_010_565, w_010_566, w_010_567, w_010_568, w_010_569, w_010_571, w_010_572, w_010_573, w_010_574, w_010_575, w_010_576, w_010_577, w_010_578, w_010_579, w_010_580, w_010_581, w_010_582, w_010_583, w_010_584, w_010_586, w_010_587, w_010_588, w_010_589, w_010_590, w_010_591, w_010_592, w_010_593, w_010_594, w_010_595, w_010_596, w_010_597, w_010_598, w_010_599, w_010_600, w_010_601, w_010_602, w_010_603, w_010_604, w_010_605, w_010_606, w_010_607, w_010_608, w_010_609, w_010_610, w_010_611, w_010_612, w_010_613, w_010_615, w_010_616, w_010_617, w_010_618, w_010_619, w_010_620, w_010_621, w_010_622, w_010_623, w_010_624, w_010_625, w_010_626, w_010_628, w_010_629, w_010_630, w_010_631, w_010_632, w_010_633, w_010_635, w_010_636, w_010_637, w_010_638, w_010_639, w_010_640, w_010_641, w_010_642, w_010_643, w_010_644, w_010_645, w_010_646, w_010_647, w_010_648, w_010_649, w_010_650, w_010_651, w_010_652, w_010_653, w_010_654, w_010_655, w_010_656, w_010_657, w_010_658, w_010_659, w_010_660, w_010_661, w_010_662, w_010_663, w_010_664, w_010_665, w_010_666, w_010_667, w_010_668, w_010_669, w_010_670, w_010_671, w_010_672, w_010_673, w_010_674, w_010_675, w_010_676, w_010_677, w_010_678, w_010_679, w_010_680, w_010_682, w_010_683, w_010_684, w_010_685, w_010_686, w_010_687, w_010_688, w_010_689, w_010_690, w_010_691, w_010_693, w_010_694, w_010_695, w_010_696, w_010_697, w_010_698, w_010_699, w_010_700, w_010_701, w_010_702, w_010_703, w_010_704, w_010_705, w_010_706, w_010_707, w_010_708, w_010_709, w_010_710, w_010_711, w_010_712, w_010_713, w_010_714, w_010_715, w_010_716, w_010_718, w_010_719, w_010_721, w_010_722, w_010_723, w_010_724, w_010_726, w_010_727, w_010_728, w_010_729, w_010_730, w_010_731, w_010_732, w_010_733, w_010_734, w_010_735, w_010_736, w_010_737, w_010_738, w_010_739, w_010_741, w_010_742, w_010_743, w_010_744, w_010_745, w_010_747, w_010_749, w_010_751, w_010_752, w_010_753, w_010_754, w_010_755, w_010_756, w_010_757, w_010_758, w_010_759, w_010_760, w_010_761, w_010_762, w_010_763, w_010_764, w_010_765, w_010_766, w_010_767, w_010_768, w_010_769, w_010_770, w_010_771, w_010_772, w_010_773, w_010_774, w_010_775, w_010_776, w_010_777, w_010_778, w_010_779, w_010_780, w_010_781, w_010_782, w_010_783, w_010_784, w_010_785, w_010_786, w_010_787, w_010_788, w_010_789, w_010_790, w_010_791, w_010_792, w_010_793, w_010_794, w_010_795, w_010_796, w_010_797, w_010_798, w_010_799, w_010_800, w_010_801, w_010_802, w_010_803, w_010_804, w_010_805, w_010_806, w_010_807, w_010_808, w_010_809, w_010_810, w_010_811, w_010_812, w_010_813, w_010_814, w_010_815, w_010_816, w_010_817, w_010_818, w_010_819, w_010_820, w_010_821, w_010_822, w_010_823, w_010_824, w_010_825, w_010_826, w_010_827, w_010_828, w_010_829, w_010_830, w_010_831, w_010_832, w_010_833, w_010_834, w_010_835, w_010_836, w_010_838, w_010_840, w_010_841, w_010_842, w_010_844, w_010_845, w_010_846, w_010_847, w_010_848, w_010_849, w_010_850, w_010_851, w_010_853, w_010_854, w_010_855, w_010_856, w_010_857, w_010_858, w_010_859, w_010_860, w_010_861, w_010_862, w_010_863, w_010_864, w_010_865, w_010_866, w_010_867, w_010_868, w_010_869, w_010_870, w_010_871, w_010_872, w_010_873, w_010_874, w_010_875, w_010_876, w_010_877, w_010_878, w_010_879, w_010_880, w_010_881, w_010_882, w_010_883, w_010_884, w_010_885, w_010_886, w_010_887, w_010_888, w_010_889, w_010_890, w_010_891, w_010_892, w_010_894, w_010_895, w_010_896, w_010_897, w_010_898, w_010_899, w_010_900, w_010_902, w_010_903, w_010_904, w_010_905, w_010_906, w_010_907, w_010_908, w_010_909, w_010_910, w_010_911, w_010_912, w_010_913, w_010_915, w_010_916, w_010_917, w_010_918, w_010_920, w_010_921, w_010_922, w_010_923, w_010_924, w_010_925, w_010_926, w_010_927, w_010_928, w_010_929, w_010_930, w_010_932, w_010_933, w_010_934, w_010_935, w_010_936, w_010_937, w_010_938, w_010_939, w_010_940, w_010_941, w_010_942, w_010_943, w_010_944, w_010_945, w_010_947, w_010_948, w_010_949, w_010_950, w_010_951, w_010_952, w_010_953, w_010_954, w_010_955, w_010_956, w_010_957, w_010_958, w_010_959, w_010_960, w_010_961, w_010_962, w_010_963, w_010_964, w_010_965, w_010_966, w_010_967, w_010_968, w_010_969, w_010_970, w_010_971, w_010_972, w_010_973, w_010_974, w_010_975, w_010_976, w_010_977, w_010_978, w_010_979, w_010_980, w_010_981, w_010_982, w_010_983, w_010_984, w_010_985, w_010_986, w_010_987, w_010_988, w_010_989, w_010_990, w_010_991, w_010_992, w_010_993, w_010_994, w_010_995, w_010_996, w_010_997, w_010_998, w_010_999, w_010_1000, w_010_1001, w_010_1002, w_010_1003, w_010_1004, w_010_1005, w_010_1006, w_010_1007, w_010_1008, w_010_1009, w_010_1010, w_010_1011, w_010_1012, w_010_1013, w_010_1014, w_010_1015, w_010_1016, w_010_1017, w_010_1018, w_010_1019, w_010_1022, w_010_1023, w_010_1024, w_010_1025, w_010_1026, w_010_1027, w_010_1028, w_010_1029, w_010_1030, w_010_1032, w_010_1034, w_010_1035, w_010_1036, w_010_1037, w_010_1038, w_010_1039, w_010_1040, w_010_1041, w_010_1042, w_010_1043, w_010_1044, w_010_1045, w_010_1046, w_010_1047, w_010_1048, w_010_1049, w_010_1050, w_010_1051, w_010_1052, w_010_1053, w_010_1054, w_010_1055, w_010_1056, w_010_1057, w_010_1058, w_010_1059, w_010_1060, w_010_1061, w_010_1062, w_010_1063, w_010_1064, w_010_1065, w_010_1067, w_010_1068, w_010_1069, w_010_1071, w_010_1072, w_010_1073, w_010_1074, w_010_1075, w_010_1076, w_010_1077, w_010_1078, w_010_1079, w_010_1080, w_010_1081, w_010_1082, w_010_1083, w_010_1084, w_010_1085, w_010_1086, w_010_1088, w_010_1089, w_010_1090, w_010_1091, w_010_1092, w_010_1093, w_010_1094, w_010_1095, w_010_1096, w_010_1097, w_010_1098, w_010_1099, w_010_1100, w_010_1101, w_010_1102, w_010_1103, w_010_1104, w_010_1105, w_010_1106, w_010_1107, w_010_1108, w_010_1109, w_010_1110, w_010_1111, w_010_1112, w_010_1113, w_010_1114, w_010_1115, w_010_1117, w_010_1118, w_010_1120, w_010_1121, w_010_1122, w_010_1123, w_010_1124, w_010_1125, w_010_1126, w_010_1127, w_010_1128, w_010_1129, w_010_1130, w_010_1131, w_010_1132, w_010_1133, w_010_1134, w_010_1135, w_010_1136, w_010_1137, w_010_1138, w_010_1139, w_010_1140, w_010_1141, w_010_1142, w_010_1143, w_010_1144, w_010_1145, w_010_1146, w_010_1147, w_010_1148, w_010_1149, w_010_1150, w_010_1151, w_010_1152, w_010_1153, w_010_1154, w_010_1156, w_010_1157, w_010_1158, w_010_1159, w_010_1160, w_010_1162, w_010_1163, w_010_1164, w_010_1165, w_010_1166, w_010_1167, w_010_1168, w_010_1169, w_010_1170, w_010_1171, w_010_1172, w_010_1173, w_010_1175, w_010_1176, w_010_1177, w_010_1178, w_010_1179, w_010_1180, w_010_1181, w_010_1182, w_010_1183, w_010_1184, w_010_1185, w_010_1186, w_010_1187, w_010_1188, w_010_1189, w_010_1190, w_010_1191, w_010_1192, w_010_1193, w_010_1194, w_010_1195, w_010_1196, w_010_1197, w_010_1198, w_010_1199, w_010_1200, w_010_1201, w_010_1202, w_010_1203, w_010_1204, w_010_1205, w_010_1206, w_010_1207, w_010_1208, w_010_1209, w_010_1210, w_010_1211, w_010_1212, w_010_1213, w_010_1214, w_010_1215, w_010_1216, w_010_1217, w_010_1218, w_010_1219, w_010_1220, w_010_1221, w_010_1222, w_010_1223, w_010_1224, w_010_1225, w_010_1226, w_010_1227, w_010_1228, w_010_1229, w_010_1230, w_010_1231, w_010_1232, w_010_1234, w_010_1236, w_010_1238, w_010_1239, w_010_1240, w_010_1241, w_010_1242, w_010_1243, w_010_1244, w_010_1245, w_010_1246, w_010_1247, w_010_1248, w_010_1249, w_010_1250, w_010_1251, w_010_1252, w_010_1253, w_010_1254, w_010_1255, w_010_1256, w_010_1257, w_010_1258, w_010_1259, w_010_1260, w_010_1261, w_010_1263, w_010_1264, w_010_1265, w_010_1266, w_010_1267, w_010_1268, w_010_1269, w_010_1270, w_010_1271, w_010_1272, w_010_1273, w_010_1274, w_010_1275, w_010_1276, w_010_1277, w_010_1278, w_010_1279, w_010_1280, w_010_1281, w_010_1282, w_010_1283, w_010_1284, w_010_1285, w_010_1286, w_010_1287, w_010_1288, w_010_1289, w_010_1290, w_010_1291, w_010_1292, w_010_1293, w_010_1294, w_010_1296, w_010_1297, w_010_1298, w_010_1299, w_010_1300, w_010_1301, w_010_1302, w_010_1303, w_010_1304, w_010_1305, w_010_1306, w_010_1307, w_010_1308, w_010_1309, w_010_1310, w_010_1311, w_010_1312, w_010_1313, w_010_1314, w_010_1315, w_010_1316, w_010_1317, w_010_1318, w_010_1319, w_010_1320, w_010_1321, w_010_1322, w_010_1323, w_010_1324, w_010_1325, w_010_1326, w_010_1327, w_010_1328, w_010_1329, w_010_1330, w_010_1331, w_010_1332, w_010_1333, w_010_1335, w_010_1336, w_010_1338, w_010_1339, w_010_1340, w_010_1341, w_010_1342, w_010_1343, w_010_1344, w_010_1345, w_010_1346, w_010_1347, w_010_1348, w_010_1349, w_010_1350, w_010_1351, w_010_1352, w_010_1353, w_010_1354, w_010_1355, w_010_1356, w_010_1358, w_010_1359, w_010_1360, w_010_1361, w_010_1362, w_010_1363, w_010_1364, w_010_1365, w_010_1366, w_010_1367, w_010_1369, w_010_1371, w_010_1372, w_010_1373, w_010_1374, w_010_1375, w_010_1376, w_010_1377, w_010_1378, w_010_1379, w_010_1380, w_010_1381, w_010_1382, w_010_1383, w_010_1384, w_010_1385, w_010_1386, w_010_1387, w_010_1388, w_010_1389, w_010_1390, w_010_1391, w_010_1392, w_010_1393, w_010_1394, w_010_1395, w_010_1396, w_010_1397, w_010_1398, w_010_1399, w_010_1400, w_010_1401, w_010_1402, w_010_1403, w_010_1404, w_010_1405, w_010_1406, w_010_1407, w_010_1408, w_010_1409, w_010_1410, w_010_1411, w_010_1412, w_010_1413, w_010_1415, w_010_1416, w_010_1417, w_010_1418, w_010_1419, w_010_1421, w_010_1422, w_010_1423, w_010_1424, w_010_1425, w_010_1426, w_010_1427, w_010_1428, w_010_1429, w_010_1430, w_010_1431, w_010_1432, w_010_1433, w_010_1434, w_010_1435, w_010_1436, w_010_1437, w_010_1438, w_010_1439, w_010_1440, w_010_1441, w_010_1442, w_010_1443, w_010_1444, w_010_1445, w_010_1446, w_010_1447, w_010_1448, w_010_1449, w_010_1450, w_010_1451, w_010_1452, w_010_1454, w_010_1455, w_010_1456, w_010_1457, w_010_1458, w_010_1459, w_010_1460, w_010_1461, w_010_1462, w_010_1463, w_010_1464, w_010_1465, w_010_1466, w_010_1468, w_010_1469, w_010_1470, w_010_1471, w_010_1472, w_010_1473, w_010_1474, w_010_1475, w_010_1476, w_010_1477, w_010_1478, w_010_1479, w_010_1480, w_010_1481, w_010_1483, w_010_1484, w_010_1485, w_010_1487, w_010_1488, w_010_1489, w_010_1490, w_010_1491, w_010_1493, w_010_1494, w_010_1495, w_010_1496, w_010_1497, w_010_1498, w_010_1500, w_010_1501, w_010_1502, w_010_1503, w_010_1504, w_010_1505, w_010_1507, w_010_1508, w_010_1509, w_010_1510, w_010_1511, w_010_1512, w_010_1513, w_010_1514, w_010_1516, w_010_1517, w_010_1518, w_010_1519, w_010_1520, w_010_1522, w_010_1523, w_010_1524, w_010_1525, w_010_1526, w_010_1527, w_010_1528, w_010_1529, w_010_1530, w_010_1531, w_010_1532, w_010_1533, w_010_1534, w_010_1535, w_010_1536, w_010_1537, w_010_1538, w_010_1539, w_010_1540, w_010_1541, w_010_1542, w_010_1543, w_010_1545, w_010_1546, w_010_1548, w_010_1549, w_010_1550, w_010_1551, w_010_1552, w_010_1553, w_010_1554, w_010_1555, w_010_1556, w_010_1557, w_010_1559, w_010_1560, w_010_1561, w_010_1562, w_010_1563, w_010_1564, w_010_1565, w_010_1566, w_010_1567, w_010_1568, w_010_1569, w_010_1570, w_010_1571, w_010_1572, w_010_1573, w_010_1575, w_010_1576, w_010_1577, w_010_1578, w_010_1579, w_010_1580, w_010_1581, w_010_1582, w_010_1583, w_010_1584, w_010_1585, w_010_1586, w_010_1587, w_010_1588, w_010_1589, w_010_1590, w_010_1591, w_010_1592, w_010_1593, w_010_1594, w_010_1595, w_010_1596, w_010_1597, w_010_1598, w_010_1599, w_010_1600, w_010_1601, w_010_1602, w_010_1603, w_010_1604, w_010_1605, w_010_1606, w_010_1607, w_010_1608, w_010_1609, w_010_1610, w_010_1611, w_010_1612, w_010_1613, w_010_1614, w_010_1615, w_010_1616, w_010_1617, w_010_1618, w_010_1619, w_010_1620, w_010_1621, w_010_1623, w_010_1624, w_010_1625, w_010_1626, w_010_1627, w_010_1628, w_010_1629, w_010_1630, w_010_1631, w_010_1632, w_010_1633, w_010_1634, w_010_1635, w_010_1636, w_010_1637, w_010_1638, w_010_1639, w_010_1640, w_010_1641, w_010_1642, w_010_1643, w_010_1644, w_010_1645, w_010_1646, w_010_1647, w_010_1648, w_010_1649, w_010_1650, w_010_1651, w_010_1652, w_010_1653, w_010_1654, w_010_1656, w_010_1657, w_010_1658, w_010_1659, w_010_1660, w_010_1661, w_010_1662, w_010_1663, w_010_1664, w_010_1665, w_010_1666, w_010_1668, w_010_1669, w_010_1671, w_010_1672, w_010_1673, w_010_1675, w_010_1676, w_010_1677, w_010_1678, w_010_1680, w_010_1681, w_010_1682, w_010_1683, w_010_1684, w_010_1685, w_010_1686, w_010_1687, w_010_1688, w_010_1690, w_010_1691, w_010_1692, w_010_1693, w_010_1694, w_010_1695, w_010_1696, w_010_1697, w_010_1698, w_010_1700, w_010_1701, w_010_1702, w_010_1703, w_010_1704, w_010_1705, w_010_1706, w_010_1707, w_010_1708, w_010_1709, w_010_1710, w_010_1712, w_010_1713, w_010_1714, w_010_1715, w_010_1716, w_010_1717, w_010_1718, w_010_1719, w_010_1720, w_010_1721, w_010_1722, w_010_1723, w_010_1724, w_010_1725, w_010_1726, w_010_1727, w_010_1728, w_010_1729, w_010_1730, w_010_1731, w_010_1732, w_010_1733, w_010_1734, w_010_1735, w_010_1736, w_010_1737, w_010_1738, w_010_1739, w_010_1740, w_010_1741, w_010_1742, w_010_1743, w_010_1744, w_010_1745, w_010_1746, w_010_1747, w_010_1748, w_010_1749, w_010_1750, w_010_1751, w_010_1752, w_010_1753, w_010_1754, w_010_1755, w_010_1756, w_010_1757, w_010_1758, w_010_1760, w_010_1761, w_010_1762, w_010_1763, w_010_1764, w_010_1765, w_010_1766, w_010_1767, w_010_1769, w_010_1770, w_010_1771, w_010_1772, w_010_1773, w_010_1774, w_010_1775, w_010_1776, w_010_1778, w_010_1779, w_010_1780, w_010_1782, w_010_1783, w_010_1784, w_010_1785, w_010_1786, w_010_1787, w_010_1788, w_010_1789, w_010_1790, w_010_1791, w_010_1792, w_010_1793, w_010_1794, w_010_1795, w_010_1796, w_010_1797, w_010_1798, w_010_1799, w_010_1801, w_010_1802, w_010_1803, w_010_1804, w_010_1805, w_010_1806, w_010_1807, w_010_1808, w_010_1809, w_010_1810, w_010_1811, w_010_1812, w_010_1813, w_010_1814, w_010_1815, w_010_1817, w_010_1818, w_010_1819, w_010_1820, w_010_1821, w_010_1822, w_010_1823, w_010_1824, w_010_1825, w_010_1826, w_010_1827, w_010_1828, w_010_1829, w_010_1830, w_010_1831, w_010_1832, w_010_1833, w_010_1834, w_010_1835, w_010_1837, w_010_1838, w_010_1839, w_010_1840, w_010_1841, w_010_1842, w_010_1843, w_010_1844, w_010_1845, w_010_1846, w_010_1848, w_010_1849, w_010_1850, w_010_1851, w_010_1852, w_010_1853, w_010_1854, w_010_1855, w_010_1856, w_010_1857, w_010_1858, w_010_1859, w_010_1860, w_010_1861, w_010_1862, w_010_1863, w_010_1864, w_010_1865, w_010_1866, w_010_1867, w_010_1871, w_010_1872, w_010_1873, w_010_1874, w_010_1875, w_010_1876, w_010_1877, w_010_1878, w_010_1879, w_010_1880, w_010_1881, w_010_1882, w_010_1883, w_010_1884, w_010_1885, w_010_1886, w_010_1887, w_010_1888, w_010_1889, w_010_1890, w_010_1891, w_010_1892, w_010_1893, w_010_1894, w_010_1895, w_010_1896, w_010_1897, w_010_1898, w_010_1899, w_010_1900, w_010_1902, w_010_1903, w_010_1905, w_010_1906, w_010_1907, w_010_1908, w_010_1909, w_010_1910, w_010_1911, w_010_1912, w_010_1913, w_010_1914, w_010_1915, w_010_1916, w_010_1917, w_010_1918, w_010_1919, w_010_1920, w_010_1921, w_010_1922, w_010_1923, w_010_1924, w_010_1925, w_010_1926, w_010_1927, w_010_1928, w_010_1929, w_010_1930, w_010_1931, w_010_1932, w_010_1933, w_010_1934, w_010_1935, w_010_1936, w_010_1937, w_010_1938, w_010_1939, w_010_1940, w_010_1941, w_010_1942, w_010_1943, w_010_1944, w_010_1945, w_010_1946, w_010_1947, w_010_1948, w_010_1949, w_010_1951, w_010_1952, w_010_1953, w_010_1955, w_010_1956, w_010_1957, w_010_1958, w_010_1959, w_010_1960, w_010_1961, w_010_1962, w_010_1963, w_010_1966, w_010_1967, w_010_1968, w_010_1969, w_010_1970, w_010_1971, w_010_1972, w_010_1973, w_010_1974, w_010_1975, w_010_1976, w_010_1977, w_010_1978, w_010_1979, w_010_1980, w_010_1981, w_010_1982, w_010_1983, w_010_1984, w_010_1985, w_010_1986, w_010_1987, w_010_1988, w_010_1989, w_010_1990, w_010_1991, w_010_1992, w_010_1993, w_010_1994, w_010_1995, w_010_1996, w_010_1997, w_010_1998, w_010_1999, w_010_2000, w_010_2001, w_010_2002, w_010_2003, w_010_2004, w_010_2005, w_010_2006, w_010_2007, w_010_2008, w_010_2009, w_010_2010, w_010_2011, w_010_2012, w_010_2013, w_010_2014, w_010_2015, w_010_2016, w_010_2017, w_010_2018, w_010_2019, w_010_2020, w_010_2021, w_010_2022, w_010_2023, w_010_2024, w_010_2025, w_010_2026, w_010_2027, w_010_2028, w_010_2029, w_010_2030, w_010_2031, w_010_2032, w_010_2033, w_010_2034, w_010_2035, w_010_2036, w_010_2037, w_010_2038, w_010_2039, w_010_2040, w_010_2041, w_010_2042, w_010_2043, w_010_2044, w_010_2045, w_010_2046, w_010_2047, w_010_2048, w_010_2050, w_010_2051, w_010_2052, w_010_2053, w_010_2054, w_010_2055, w_010_2056, w_010_2057, w_010_2058, w_010_2059, w_010_2060, w_010_2061, w_010_2062, w_010_2063, w_010_2065, w_010_2066, w_010_2067, w_010_2068, w_010_2069, w_010_2070, w_010_2071, w_010_2072, w_010_2073, w_010_2074, w_010_2075, w_010_2076, w_010_2077, w_010_2078, w_010_2079, w_010_2080, w_010_2081, w_010_2082, w_010_2083, w_010_2084, w_010_2085, w_010_2086, w_010_2087, w_010_2089, w_010_2090, w_010_2091, w_010_2093, w_010_2094, w_010_2095, w_010_2096, w_010_2097, w_010_2098, w_010_2099, w_010_2100, w_010_2101, w_010_2102, w_010_2103, w_010_2104, w_010_2105, w_010_2106, w_010_2107, w_010_2108, w_010_2109, w_010_2110, w_010_2111, w_010_2112, w_010_2113, w_010_2114, w_010_2115, w_010_2116, w_010_2117, w_010_2118, w_010_2119, w_010_2120, w_010_2121, w_010_2122, w_010_2123, w_010_2124, w_010_2125, w_010_2126, w_010_2127, w_010_2128, w_010_2129, w_010_2130, w_010_2131, w_010_2132, w_010_2133, w_010_2134, w_010_2135, w_010_2136, w_010_2137, w_010_2138, w_010_2139, w_010_2140, w_010_2141, w_010_2142, w_010_2143, w_010_2144, w_010_2145, w_010_2146, w_010_2147, w_010_2148, w_010_2149, w_010_2150, w_010_2151, w_010_2152, w_010_2153, w_010_2154, w_010_2155, w_010_2156, w_010_2159, w_010_2160, w_010_2161, w_010_2162, w_010_2163, w_010_2164, w_010_2165, w_010_2166, w_010_2167, w_010_2168, w_010_2169, w_010_2171, w_010_2173, w_010_2174, w_010_2175, w_010_2176, w_010_2177, w_010_2178, w_010_2180, w_010_2181, w_010_2182, w_010_2183, w_010_2184, w_010_2185, w_010_2186, w_010_2187, w_010_2188, w_010_2189, w_010_2190, w_010_2191, w_010_2192, w_010_2193, w_010_2195, w_010_2196, w_010_2197, w_010_2198, w_010_2199, w_010_2200, w_010_2201, w_010_2202, w_010_2203, w_010_2204, w_010_2205, w_010_2206, w_010_2207, w_010_2208, w_010_2209, w_010_2210, w_010_2211, w_010_2212, w_010_2213, w_010_2216, w_010_2217, w_010_2218, w_010_2219, w_010_2220, w_010_2221, w_010_2222, w_010_2223, w_010_2224, w_010_2225, w_010_2227, w_010_2228, w_010_2229, w_010_2230, w_010_2231, w_010_2232, w_010_2233, w_010_2234, w_010_2235, w_010_2236, w_010_2237, w_010_2238, w_010_2239, w_010_2240, w_010_2241, w_010_2242, w_010_2243, w_010_2244, w_010_2245, w_010_2246, w_010_2247, w_010_2248, w_010_2249, w_010_2250, w_010_2251, w_010_2252, w_010_2253, w_010_2255, w_010_2256, w_010_2257, w_010_2258, w_010_2259, w_010_2260, w_010_2261, w_010_2262, w_010_2263, w_010_2264, w_010_2265, w_010_2266, w_010_2267, w_010_2268, w_010_2269, w_010_2270, w_010_2271, w_010_2272, w_010_2273, w_010_2274, w_010_2275, w_010_2276, w_010_2278, w_010_2279, w_010_2280, w_010_2281, w_010_2282, w_010_2284, w_010_2285, w_010_2286, w_010_2287, w_010_2288, w_010_2289, w_010_2290, w_010_2291, w_010_2292, w_010_2293, w_010_2294, w_010_2295, w_010_2296, w_010_2297, w_010_2298, w_010_2299, w_010_2300, w_010_2301, w_010_2302, w_010_2303, w_010_2304, w_010_2305, w_010_2306, w_010_2307, w_010_2309, w_010_2310, w_010_2311, w_010_2312, w_010_2313, w_010_2314, w_010_2315, w_010_2316, w_010_2317, w_010_2318, w_010_2319, w_010_2320, w_010_2321, w_010_2322, w_010_2323, w_010_2324, w_010_2325, w_010_2327, w_010_2328, w_010_2329, w_010_2330, w_010_2331, w_010_2332, w_010_2333, w_010_2334, w_010_2335, w_010_2336, w_010_2337, w_010_2338, w_010_2340, w_010_2341, w_010_2342, w_010_2343, w_010_2344, w_010_2345, w_010_2346, w_010_2347, w_010_2348, w_010_2349, w_010_2350, w_010_2351, w_010_2352, w_010_2353, w_010_2354, w_010_2356, w_010_2357, w_010_2358, w_010_2359, w_010_2360, w_010_2361, w_010_2363, w_010_2364, w_010_2365, w_010_2366, w_010_2367, w_010_2370, w_010_2371, w_010_2372, w_010_2373, w_010_2374, w_010_2375, w_010_2376, w_010_2377, w_010_2378, w_010_2379, w_010_2380, w_010_2381, w_010_2382, w_010_2383, w_010_2384, w_010_2385, w_010_2386, w_010_2387, w_010_2388, w_010_2389, w_010_2390, w_010_2391, w_010_2392, w_010_2393, w_010_2394, w_010_2395, w_010_2396, w_010_2397, w_010_2398, w_010_2399, w_010_2400, w_010_2401, w_010_2402, w_010_2403, w_010_2404, w_010_2405, w_010_2406, w_010_2407, w_010_2408, w_010_2409, w_010_2410, w_010_2411, w_010_2412, w_010_2413, w_010_2414, w_010_2415, w_010_2416, w_010_2417, w_010_2418, w_010_2419, w_010_2420, w_010_2421, w_010_2422, w_010_2423, w_010_2424, w_010_2425, w_010_2426, w_010_2428, w_010_2429, w_010_2430, w_010_2431, w_010_2432, w_010_2433, w_010_2434, w_010_2435, w_010_2436, w_010_2437, w_010_2438, w_010_2439, w_010_2440, w_010_2441, w_010_2442, w_010_2443, w_010_2444, w_010_2445, w_010_2446, w_010_2447, w_010_2448, w_010_2449, w_010_2450, w_010_2451, w_010_2452, w_010_2453, w_010_2454, w_010_2455, w_010_2456, w_010_2457, w_010_2458, w_010_2459, w_010_2460, w_010_2461, w_010_2462, w_010_2463, w_010_2464, w_010_2465, w_010_2466, w_010_2467, w_010_2469, w_010_2470, w_010_2471, w_010_2472, w_010_2473, w_010_2474, w_010_2475, w_010_2476, w_010_2477, w_010_2478, w_010_2479, w_010_2480, w_010_2481, w_010_2482, w_010_2483, w_010_2484, w_010_2485, w_010_2486, w_010_2487, w_010_2488, w_010_2489, w_010_2490, w_010_2491, w_010_2492, w_010_2493, w_010_2494, w_010_2495, w_010_2496, w_010_2497, w_010_2498, w_010_2499, w_010_2500, w_010_2501, w_010_2502, w_010_2503, w_010_2504, w_010_2505, w_010_2506, w_010_2507, w_010_2508, w_010_2509, w_010_2510, w_010_2511, w_010_2512, w_010_2513, w_010_2514, w_010_2516, w_010_2517, w_010_2518, w_010_2519, w_010_2520, w_010_2521, w_010_2522, w_010_2523, w_010_2524, w_010_2525, w_010_2526, w_010_2527, w_010_2528, w_010_2529, w_010_2530, w_010_2531, w_010_2532, w_010_2533, w_010_2534, w_010_2535, w_010_2536, w_010_2537, w_010_2538, w_010_2539, w_010_2540, w_010_2541, w_010_2542, w_010_2543, w_010_2544, w_010_2545, w_010_2546, w_010_2547, w_010_2548, w_010_2549, w_010_2550, w_010_2551, w_010_2552, w_010_2553, w_010_2554, w_010_2555, w_010_2556, w_010_2557, w_010_2558, w_010_2559, w_010_2560, w_010_2561, w_010_2562, w_010_2563, w_010_2564, w_010_2565, w_010_2566, w_010_2567, w_010_2568, w_010_2569, w_010_2570, w_010_2571, w_010_2572, w_010_2573, w_010_2574, w_010_2575, w_010_2576, w_010_2577, w_010_2578, w_010_2579, w_010_2580, w_010_2581, w_010_2582, w_010_2583, w_010_2584, w_010_2585, w_010_2586, w_010_2587, w_010_2588, w_010_2590, w_010_2591, w_010_2592, w_010_2593, w_010_2594, w_010_2595, w_010_2596, w_010_2597, w_010_2598, w_010_2599, w_010_2601, w_010_2602, w_010_2603, w_010_2604, w_010_2605, w_010_2606, w_010_2607, w_010_2608, w_010_2609, w_010_2610, w_010_2611, w_010_2612, w_010_2613, w_010_2616, w_010_2617, w_010_2618, w_010_2619, w_010_2620, w_010_2621, w_010_2623, w_010_2624, w_010_2625, w_010_2626, w_010_2627, w_010_2628, w_010_2629, w_010_2630, w_010_2631, w_010_2632, w_010_2633, w_010_2634, w_010_2635, w_010_2636, w_010_2637, w_010_2638, w_010_2639, w_010_2640, w_010_2642, w_010_2643, w_010_2645, w_010_2646, w_010_2647, w_010_2648, w_010_2649, w_010_2650, w_010_2651, w_010_2652, w_010_2653, w_010_2654, w_010_2655, w_010_2657, w_010_2658, w_010_2659, w_010_2660, w_010_2661, w_010_2662, w_010_2663, w_010_2664, w_010_2665, w_010_2666, w_010_2667, w_010_2668, w_010_2669, w_010_2671, w_010_2672, w_010_2674, w_010_2675, w_010_2676, w_010_2677, w_010_2678, w_010_2680, w_010_2681, w_010_2682, w_010_2683, w_010_2684, w_010_2685, w_010_2686, w_010_2688, w_010_2689, w_010_2690, w_010_2692, w_010_2693, w_010_2694, w_010_2696, w_010_2697, w_010_2698, w_010_2699, w_010_2700, w_010_2701, w_010_2702, w_010_2703, w_010_2704, w_010_2705, w_010_2706, w_010_2707, w_010_2708, w_010_2709, w_010_2710, w_010_2711, w_010_2712, w_010_2713, w_010_2714, w_010_2715, w_010_2717, w_010_2718, w_010_2719, w_010_2720, w_010_2721, w_010_2722, w_010_2723, w_010_2724, w_010_2725, w_010_2726, w_010_2727, w_010_2728, w_010_2729, w_010_2730, w_010_2731, w_010_2732, w_010_2734, w_010_2735, w_010_2736, w_010_2737, w_010_2738, w_010_2739, w_010_2740, w_010_2741, w_010_2742, w_010_2743, w_010_2744, w_010_2745, w_010_2746, w_010_2747, w_010_2748, w_010_2749, w_010_2750, w_010_2751, w_010_2752, w_010_2753, w_010_2754, w_010_2755, w_010_2756, w_010_2757, w_010_2758, w_010_2759, w_010_2761, w_010_2762, w_010_2763, w_010_2764, w_010_2765, w_010_2766, w_010_2767, w_010_2768, w_010_2769, w_010_2770, w_010_2771, w_010_2772, w_010_2773, w_010_2774, w_010_2776, w_010_2777, w_010_2779, w_010_2780, w_010_2781, w_010_2782, w_010_2783, w_010_2784, w_010_2785, w_010_2786, w_010_2787, w_010_2788, w_010_2789, w_010_2790, w_010_2791, w_010_2792, w_010_2793, w_010_2794, w_010_2795, w_010_2796, w_010_2797, w_010_2798, w_010_2799, w_010_2800, w_010_2801, w_010_2802, w_010_2803, w_010_2804, w_010_2805, w_010_2806, w_010_2807, w_010_2808, w_010_2809, w_010_2810, w_010_2811, w_010_2812, w_010_2813, w_010_2815, w_010_2816, w_010_2817, w_010_2818, w_010_2819, w_010_2820, w_010_2821, w_010_2822, w_010_2823, w_010_2824, w_010_2825, w_010_2826, w_010_2827, w_010_2828, w_010_2829, w_010_2830, w_010_2831, w_010_2832, w_010_2833, w_010_2834, w_010_2835, w_010_2836, w_010_2837, w_010_2838, w_010_2839, w_010_2840, w_010_2841, w_010_2842, w_010_2843, w_010_2844, w_010_2845, w_010_2846, w_010_2847, w_010_2848, w_010_2849, w_010_2850, w_010_2851, w_010_2852, w_010_2854, w_010_2855, w_010_2856, w_010_2857, w_010_2858, w_010_2859, w_010_2860, w_010_2861, w_010_2862, w_010_2863, w_010_2864, w_010_2865, w_010_2866, w_010_2867, w_010_2868, w_010_2869, w_010_2870, w_010_2871, w_010_2872, w_010_2873, w_010_2874, w_010_2875, w_010_2876, w_010_2877, w_010_2878, w_010_2879, w_010_2880, w_010_2881, w_010_2882, w_010_2883, w_010_2884, w_010_2885, w_010_2886, w_010_2888, w_010_2889, w_010_2890, w_010_2891, w_010_2892, w_010_2893, w_010_2894, w_010_2895, w_010_2896, w_010_2897, w_010_2898, w_010_2899, w_010_2901, w_010_2902, w_010_2904, w_010_2905, w_010_2906, w_010_2907, w_010_2908, w_010_2909, w_010_2910, w_010_2911, w_010_2912, w_010_2913, w_010_2916, w_010_2917, w_010_2918, w_010_2919, w_010_2920, w_010_2921, w_010_2922, w_010_2923, w_010_2924, w_010_2925, w_010_2926, w_010_2928, w_010_2929, w_010_2930, w_010_2932, w_010_2933, w_010_2934, w_010_2937, w_010_2938, w_010_2939, w_010_2940, w_010_2941, w_010_2942, w_010_2943, w_010_2944, w_010_2945, w_010_2946, w_010_2947, w_010_2948, w_010_2949, w_010_2950, w_010_2951, w_010_2952, w_010_2953, w_010_2954, w_010_2955, w_010_2956, w_010_2958, w_010_2959, w_010_2960, w_010_2961, w_010_2962, w_010_2963, w_010_2964, w_010_2965, w_010_2966, w_010_2968, w_010_2969, w_010_2971, w_010_2972, w_010_2973, w_010_2974, w_010_2975, w_010_2976, w_010_2977, w_010_2978, w_010_2980, w_010_2981, w_010_2982, w_010_2983, w_010_2984, w_010_2985, w_010_2986, w_010_2987, w_010_2988, w_010_2989, w_010_2990, w_010_2991, w_010_2992, w_010_2993, w_010_2994, w_010_2995, w_010_2996, w_010_2997, w_010_2998, w_010_2999, w_010_3000, w_010_3001, w_010_3002, w_010_3003, w_010_3004, w_010_3005, w_010_3006, w_010_3007, w_010_3008, w_010_3009, w_010_3010, w_010_3011, w_010_3013, w_010_3014, w_010_3015, w_010_3016, w_010_3017, w_010_3018, w_010_3019, w_010_3020, w_010_3021, w_010_3022, w_010_3023, w_010_3024, w_010_3025, w_010_3026, w_010_3027, w_010_3029, w_010_3030, w_010_3031, w_010_3032, w_010_3033, w_010_3034, w_010_3035, w_010_3036, w_010_3037, w_010_3038, w_010_3039, w_010_3040, w_010_3041, w_010_3043, w_010_3044, w_010_3045, w_010_3046, w_010_3047, w_010_3048, w_010_3049, w_010_3050, w_010_3051, w_010_3052, w_010_3053, w_010_3054, w_010_3055, w_010_3056, w_010_3057, w_010_3058, w_010_3059, w_010_3060, w_010_3061, w_010_3062, w_010_3063, w_010_3064, w_010_3065, w_010_3066, w_010_3067, w_010_3068, w_010_3069, w_010_3070, w_010_3071, w_010_3072, w_010_3073, w_010_3074, w_010_3075, w_010_3076, w_010_3077, w_010_3078, w_010_3079, w_010_3080, w_010_3081, w_010_3082, w_010_3083, w_010_3084, w_010_3085, w_010_3086, w_010_3087, w_010_3088, w_010_3090, w_010_3091, w_010_3092, w_010_3093, w_010_3094, w_010_3095, w_010_3096, w_010_3097, w_010_3098, w_010_3099, w_010_3100, w_010_3101, w_010_3102, w_010_3103, w_010_3104, w_010_3105, w_010_3106, w_010_3107, w_010_3108, w_010_3109, w_010_3110, w_010_3111, w_010_3112, w_010_3113, w_010_3114, w_010_3115, w_010_3116, w_010_3117, w_010_3118, w_010_3119, w_010_3120, w_010_3121, w_010_3122, w_010_3123, w_010_3124, w_010_3125, w_010_3126, w_010_3127, w_010_3128, w_010_3129, w_010_3130, w_010_3131, w_010_3132, w_010_3133, w_010_3134, w_010_3135, w_010_3136, w_010_3137, w_010_3139, w_010_3140, w_010_3141, w_010_3142, w_010_3143, w_010_3144, w_010_3145, w_010_3146, w_010_3147, w_010_3148, w_010_3150, w_010_3151, w_010_3152, w_010_3153, w_010_3154, w_010_3155, w_010_3156, w_010_3157, w_010_3158, w_010_3159, w_010_3160, w_010_3161, w_010_3162, w_010_3163, w_010_3164, w_010_3165, w_010_3166, w_010_3167, w_010_3168, w_010_3169, w_010_3170, w_010_3171, w_010_3172, w_010_3173, w_010_3174, w_010_3175, w_010_3177, w_010_3179, w_010_3180, w_010_3181, w_010_3182, w_010_3183, w_010_3184, w_010_3185, w_010_3186, w_010_3187, w_010_3188, w_010_3189, w_010_3190, w_010_3191, w_010_3192, w_010_3193, w_010_3194, w_010_3195, w_010_3196, w_010_3197, w_010_3198, w_010_3200, w_010_3201, w_010_3202, w_010_3203, w_010_3205, w_010_3206, w_010_3207, w_010_3208, w_010_3209, w_010_3210, w_010_3211, w_010_3212, w_010_3214, w_010_3215, w_010_3216, w_010_3217, w_010_3218, w_010_3219, w_010_3220, w_010_3221, w_010_3222, w_010_3224, w_010_3225, w_010_3226, w_010_3227, w_010_3228, w_010_3229, w_010_3232, w_010_3233, w_010_3234, w_010_3235, w_010_3236, w_010_3238, w_010_3239, w_010_3240, w_010_3241, w_010_3242, w_010_3243, w_010_3244, w_010_3245, w_010_3246, w_010_3247, w_010_3248, w_010_3249, w_010_3250, w_010_3251, w_010_3252, w_010_3253, w_010_3254, w_010_3255, w_010_3256, w_010_3257, w_010_3258, w_010_3259, w_010_3260, w_010_3261, w_010_3262, w_010_3264, w_010_3265, w_010_3266, w_010_3267, w_010_3269, w_010_3271, w_010_3272, w_010_3273, w_010_3274, w_010_3275, w_010_3276, w_010_3277, w_010_3278, w_010_3279, w_010_3280, w_010_3281, w_010_3282, w_010_3284, w_010_3285, w_010_3286, w_010_3287, w_010_3288, w_010_3289, w_010_3290, w_010_3291, w_010_3292, w_010_3293, w_010_3294, w_010_3295, w_010_3296, w_010_3297, w_010_3298, w_010_3299, w_010_3300, w_010_3301, w_010_3302, w_010_3303, w_010_3304, w_010_3305, w_010_3306, w_010_3307, w_010_3308, w_010_3309, w_010_3310, w_010_3312, w_010_3313, w_010_3314, w_010_3315, w_010_3316, w_010_3317, w_010_3318, w_010_3319, w_010_3320, w_010_3321, w_010_3322, w_010_3323, w_010_3324, w_010_3325, w_010_3326, w_010_3327, w_010_3328, w_010_3329, w_010_3330, w_010_3331, w_010_3332, w_010_3333, w_010_3334, w_010_3335, w_010_3336, w_010_3337, w_010_3338, w_010_3339, w_010_3341, w_010_3342, w_010_3343, w_010_3344, w_010_3345, w_010_3346, w_010_3347, w_010_3348, w_010_3349, w_010_3350, w_010_3351, w_010_3352, w_010_3353, w_010_3354, w_010_3355, w_010_3356, w_010_3357, w_010_3358, w_010_3359, w_010_3360, w_010_3361, w_010_3362, w_010_3363, w_010_3364, w_010_3365, w_010_3366, w_010_3367, w_010_3368, w_010_3369, w_010_3370, w_010_3371, w_010_3372, w_010_3373, w_010_3374, w_010_3375, w_010_3377, w_010_3378, w_010_3379, w_010_3380, w_010_3382, w_010_3383, w_010_3384, w_010_3385, w_010_3386, w_010_3387, w_010_3388, w_010_3389, w_010_3390, w_010_3391, w_010_3395, w_010_3396, w_010_3397, w_010_3399, w_010_3400, w_010_3401, w_010_3402, w_010_3403, w_010_3405, w_010_3406, w_010_3407, w_010_3408, w_010_3409, w_010_3410, w_010_3411, w_010_3412, w_010_3413, w_010_3414, w_010_3415, w_010_3416, w_010_3417, w_010_3418, w_010_3419, w_010_3420, w_010_3421, w_010_3422, w_010_3423, w_010_3424, w_010_3425, w_010_3426, w_010_3428, w_010_3429, w_010_3430, w_010_3431, w_010_3432, w_010_3433, w_010_3434, w_010_3435, w_010_3436, w_010_3437, w_010_3438, w_010_3439, w_010_3440, w_010_3441, w_010_3442, w_010_3443, w_010_3444, w_010_3445, w_010_3446, w_010_3447, w_010_3448, w_010_3449, w_010_3450, w_010_3451, w_010_3452, w_010_3453, w_010_3454, w_010_3455, w_010_3456, w_010_3457, w_010_3458, w_010_3459, w_010_3460, w_010_3461, w_010_3462, w_010_3463, w_010_3464, w_010_3465, w_010_3467, w_010_3468, w_010_3469, w_010_3470, w_010_3471, w_010_3472, w_010_3473, w_010_3474, w_010_3475, w_010_3476, w_010_3477, w_010_3478, w_010_3479, w_010_3480, w_010_3482, w_010_3484, w_010_3485, w_010_3486, w_010_3487, w_010_3488, w_010_3489, w_010_3490, w_010_3491, w_010_3492, w_010_3493, w_010_3495, w_010_3496, w_010_3497, w_010_3498, w_010_3499, w_010_3500, w_010_3501, w_010_3502, w_010_3503, w_010_3504, w_010_3505, w_010_3506, w_010_3507, w_010_3508, w_010_3509, w_010_3510, w_010_3511, w_010_3512, w_010_3513, w_010_3514, w_010_3515, w_010_3516, w_010_3517, w_010_3518, w_010_3519, w_010_3520, w_010_3521, w_010_3522, w_010_3523, w_010_3524, w_010_3526, w_010_3527, w_010_3528, w_010_3529, w_010_3530, w_010_3531, w_010_3532, w_010_3533, w_010_3534, w_010_3535, w_010_3536, w_010_3537, w_010_3538, w_010_3539, w_010_3540, w_010_3541, w_010_3542, w_010_3543, w_010_3544, w_010_3545, w_010_3546, w_010_3547, w_010_3548, w_010_3549, w_010_3550, w_010_3551, w_010_3552, w_010_3553, w_010_3554, w_010_3555, w_010_3556, w_010_3557, w_010_3558, w_010_3559, w_010_3560, w_010_3561, w_010_3562, w_010_3563, w_010_3564, w_010_3565, w_010_3566, w_010_3567, w_010_3568, w_010_3569, w_010_3570, w_010_3571, w_010_3572, w_010_3573, w_010_3574, w_010_3575, w_010_3576, w_010_3577, w_010_3578, w_010_3579, w_010_3580, w_010_3581, w_010_3582, w_010_3584, w_010_3585, w_010_3586, w_010_3587, w_010_3588, w_010_3589, w_010_3590, w_010_3591, w_010_3592, w_010_3593, w_010_3595, w_010_3597, w_010_3598, w_010_3599, w_010_3600, w_010_3601, w_010_3602, w_010_3603, w_010_3604, w_010_3606, w_010_3607, w_010_3608, w_010_3609, w_010_3610, w_010_3611, w_010_3612, w_010_3613, w_010_3614, w_010_3615, w_010_3616, w_010_3618, w_010_3619, w_010_3620, w_010_3621, w_010_3622, w_010_3623, w_010_3624, w_010_3625, w_010_3626, w_010_3627, w_010_3628, w_010_3629, w_010_3630, w_010_3631, w_010_3632, w_010_3633, w_010_3634, w_010_3635, w_010_3636, w_010_3637, w_010_3638, w_010_3639, w_010_3641, w_010_3642, w_010_3643, w_010_3644, w_010_3645, w_010_3646, w_010_3647, w_010_3648, w_010_3649, w_010_3651, w_010_3652, w_010_3653, w_010_3655, w_010_3656, w_010_3657, w_010_3658, w_010_3659, w_010_3660, w_010_3662, w_010_3663, w_010_3664, w_010_3665, w_010_3666, w_010_3667, w_010_3668, w_010_3669, w_010_3670, w_010_3671, w_010_3672, w_010_3673, w_010_3674, w_010_3675, w_010_3676, w_010_3677, w_010_3678, w_010_3679, w_010_3680, w_010_3681, w_010_3682, w_010_3683, w_010_3684, w_010_3685, w_010_3686, w_010_3687, w_010_3688, w_010_3689, w_010_3690, w_010_3691, w_010_3693, w_010_3694, w_010_3695, w_010_3696, w_010_3697, w_010_3698, w_010_3699, w_010_3700, w_010_3701, w_010_3702, w_010_3703, w_010_3704, w_010_3705, w_010_3706, w_010_3708, w_010_3709, w_010_3710, w_010_3711, w_010_3712, w_010_3713, w_010_3714, w_010_3715, w_010_3716, w_010_3717, w_010_3718, w_010_3719, w_010_3720, w_010_3721, w_010_3722, w_010_3723, w_010_3724, w_010_3725, w_010_3726, w_010_3727, w_010_3728, w_010_3729, w_010_3730, w_010_3731, w_010_3732, w_010_3733, w_010_3734, w_010_3735, w_010_3736, w_010_3737, w_010_3738, w_010_3739, w_010_3740, w_010_3741, w_010_3742, w_010_3743, w_010_3744, w_010_3745, w_010_3746, w_010_3747, w_010_3748, w_010_3749, w_010_3750, w_010_3751, w_010_3752, w_010_3753, w_010_3754, w_010_3755, w_010_3756, w_010_3757, w_010_3758, w_010_3759, w_010_3760, w_010_3761, w_010_3762, w_010_3763, w_010_3764, w_010_3765, w_010_3766, w_010_3767, w_010_3768, w_010_3769, w_010_3770, w_010_3771, w_010_3772, w_010_3773, w_010_3774, w_010_3775, w_010_3776, w_010_3777, w_010_3778, w_010_3779, w_010_3781, w_010_3782, w_010_3783, w_010_3784, w_010_3785, w_010_3786, w_010_3787, w_010_3788, w_010_3789, w_010_3790, w_010_3791, w_010_3792, w_010_3793, w_010_3794, w_010_3795, w_010_3796, w_010_3797, w_010_3798, w_010_3799, w_010_3800, w_010_3801, w_010_3802, w_010_3803, w_010_3804, w_010_3805, w_010_3806, w_010_3807, w_010_3808, w_010_3809, w_010_3810, w_010_3811, w_010_3812, w_010_3813, w_010_3814, w_010_3815, w_010_3816, w_010_3818, w_010_3819, w_010_3820, w_010_3821, w_010_3822, w_010_3823, w_010_3824, w_010_3825, w_010_3826, w_010_3827, w_010_3831, w_010_3832, w_010_3833, w_010_3834, w_010_3835, w_010_3836, w_010_3837, w_010_3838, w_010_3839, w_010_3840, w_010_3841, w_010_3842, w_010_3844, w_010_3845, w_010_3846, w_010_3848, w_010_3849, w_010_3850, w_010_3851, w_010_3852, w_010_3853, w_010_3854, w_010_3855, w_010_3856, w_010_3857, w_010_3858, w_010_3859, w_010_3860, w_010_3861, w_010_3862, w_010_3863, w_010_3864, w_010_3865, w_010_3866, w_010_3867, w_010_3868, w_010_3869, w_010_3870, w_010_3871, w_010_3872, w_010_3873, w_010_3875, w_010_3876, w_010_3877, w_010_3878, w_010_3879, w_010_3880, w_010_3881, w_010_3882, w_010_3883, w_010_3884, w_010_3885, w_010_3886, w_010_3887, w_010_3888, w_010_3889, w_010_3890, w_010_3891, w_010_3892, w_010_3893, w_010_3894, w_010_3895, w_010_3896, w_010_3897, w_010_3898, w_010_3900, w_010_3901, w_010_3902, w_010_3903, w_010_3904, w_010_3905, w_010_3906, w_010_3907, w_010_3908, w_010_3909, w_010_3910, w_010_3911, w_010_3912, w_010_3913, w_010_3915, w_010_3916, w_010_3917, w_010_3918, w_010_3919, w_010_3920, w_010_3921, w_010_3922, w_010_3923, w_010_3924, w_010_3925, w_010_3926, w_010_3927, w_010_3928, w_010_3929, w_010_3930, w_010_3931, w_010_3932, w_010_3933, w_010_3934, w_010_3935, w_010_3936, w_010_3937, w_010_3938, w_010_3940, w_010_3941, w_010_3942, w_010_3943, w_010_3944, w_010_3945, w_010_3946, w_010_3949, w_010_3950, w_010_3952, w_010_3953, w_010_3954, w_010_3955, w_010_3956, w_010_3958, w_010_3959, w_010_3960, w_010_3961, w_010_3962, w_010_3963, w_010_3964, w_010_3965, w_010_3966, w_010_3967, w_010_3968, w_010_3969, w_010_3970, w_010_3971, w_010_3972, w_010_3973, w_010_3974, w_010_3975, w_010_3976, w_010_3977, w_010_3978, w_010_3979, w_010_3980, w_010_3981, w_010_3982, w_010_3983, w_010_3984, w_010_3985, w_010_3986, w_010_3987, w_010_3988, w_010_3989, w_010_3990, w_010_3991, w_010_3992, w_010_3993, w_010_3994, w_010_3995, w_010_3996, w_010_3997, w_010_3998, w_010_3999, w_010_4000, w_010_4001, w_010_4002, w_010_4003, w_010_4004, w_010_4005, w_010_4006, w_010_4007, w_010_4008, w_010_4009, w_010_4010, w_010_4011, w_010_4012, w_010_4013, w_010_4014, w_010_4015, w_010_4016, w_010_4017, w_010_4018, w_010_4019, w_010_4020, w_010_4021, w_010_4022, w_010_4023, w_010_4024, w_010_4025, w_010_4026, w_010_4027, w_010_4028, w_010_4030, w_010_4031, w_010_4032, w_010_4033, w_010_4034, w_010_4035, w_010_4036, w_010_4037, w_010_4038, w_010_4039, w_010_4040, w_010_4041, w_010_4042, w_010_4044, w_010_4045, w_010_4046, w_010_4047, w_010_4048, w_010_4050, w_010_4051, w_010_4052, w_010_4054, w_010_4056, w_010_4057, w_010_4058, w_010_4059, w_010_4060, w_010_4061, w_010_4062, w_010_4063, w_010_4064, w_010_4065, w_010_4066, w_010_4067, w_010_4068, w_010_4069, w_010_4070, w_010_4071, w_010_4072, w_010_4073, w_010_4074, w_010_4075, w_010_4076, w_010_4077, w_010_4078, w_010_4079, w_010_4080, w_010_4081, w_010_4082, w_010_4083, w_010_4084, w_010_4085, w_010_4086, w_010_4087, w_010_4089, w_010_4090, w_010_4091, w_010_4092, w_010_4093, w_010_4094, w_010_4095, w_010_4096, w_010_4097, w_010_4098, w_010_4099, w_010_4100, w_010_4101, w_010_4102, w_010_4103, w_010_4104, w_010_4105, w_010_4106, w_010_4107, w_010_4108, w_010_4109, w_010_4110, w_010_4112, w_010_4113, w_010_4114, w_010_4115, w_010_4116, w_010_4117, w_010_4118, w_010_4119, w_010_4120, w_010_4121, w_010_4122, w_010_4123, w_010_4124, w_010_4125, w_010_4126, w_010_4127, w_010_4128, w_010_4129, w_010_4131, w_010_4132, w_010_4133, w_010_4134, w_010_4135, w_010_4136, w_010_4137, w_010_4138, w_010_4139, w_010_4140, w_010_4141, w_010_4142, w_010_4143, w_010_4144, w_010_4145, w_010_4146, w_010_4147, w_010_4148, w_010_4149, w_010_4150, w_010_4151, w_010_4152, w_010_4153, w_010_4154, w_010_4155, w_010_4156, w_010_4157, w_010_4158, w_010_4159, w_010_4160, w_010_4161, w_010_4163, w_010_4164, w_010_4165, w_010_4166, w_010_4167, w_010_4168, w_010_4169, w_010_4170, w_010_4171, w_010_4172, w_010_4173, w_010_4174, w_010_4175, w_010_4176, w_010_4177, w_010_4178, w_010_4179, w_010_4181, w_010_4182, w_010_4183, w_010_4186, w_010_4187, w_010_4188, w_010_4189, w_010_4190, w_010_4191, w_010_4192, w_010_4193, w_010_4194, w_010_4195, w_010_4196, w_010_4197, w_010_4198, w_010_4199, w_010_4200, w_010_4201, w_010_4202, w_010_4203, w_010_4204, w_010_4205, w_010_4206, w_010_4207, w_010_4208, w_010_4209, w_010_4210, w_010_4211, w_010_4212, w_010_4213, w_010_4214, w_010_4215, w_010_4216, w_010_4217, w_010_4218, w_010_4219, w_010_4220, w_010_4221, w_010_4222, w_010_4223, w_010_4224, w_010_4225, w_010_4226, w_010_4227, w_010_4228, w_010_4229, w_010_4230, w_010_4231, w_010_4232, w_010_4233, w_010_4236, w_010_4237, w_010_4238, w_010_4239, w_010_4240, w_010_4242, w_010_4243, w_010_4244, w_010_4245, w_010_4246, w_010_4247, w_010_4248, w_010_4249, w_010_4250, w_010_4251, w_010_4252, w_010_4253, w_010_4254, w_010_4255, w_010_4256, w_010_4257, w_010_4258, w_010_4259, w_010_4260, w_010_4261, w_010_4262, w_010_4263, w_010_4264, w_010_4265, w_010_4266, w_010_4267, w_010_4268, w_010_4269, w_010_4271, w_010_4272, w_010_4273, w_010_4274, w_010_4276, w_010_4277, w_010_4278, w_010_4279, w_010_4280, w_010_4281, w_010_4282, w_010_4283, w_010_4284, w_010_4285, w_010_4286, w_010_4287, w_010_4288, w_010_4289, w_010_4290, w_010_4291, w_010_4292, w_010_4293, w_010_4294, w_010_4296, w_010_4297, w_010_4298, w_010_4300, w_010_4301, w_010_4302, w_010_4303, w_010_4304, w_010_4305, w_010_4307, w_010_4308, w_010_4309, w_010_4311, w_010_4312, w_010_4313, w_010_4314, w_010_4315, w_010_4316, w_010_4317, w_010_4318, w_010_4319, w_010_4320, w_010_4321, w_010_4322, w_010_4323, w_010_4324, w_010_4325, w_010_4326, w_010_4328, w_010_4329, w_010_4330, w_010_4331, w_010_4332, w_010_4333, w_010_4334, w_010_4335, w_010_4336, w_010_4337, w_010_4338, w_010_4339, w_010_4340, w_010_4342, w_010_4343, w_010_4344, w_010_4345, w_010_4346, w_010_4347, w_010_4349, w_010_4350, w_010_4351, w_010_4352, w_010_4353, w_010_4354, w_010_4355, w_010_4356, w_010_4357, w_010_4358, w_010_4359, w_010_4360, w_010_4361, w_010_4362, w_010_4363, w_010_4364, w_010_4365, w_010_4367, w_010_4368, w_010_4369, w_010_4370, w_010_4371, w_010_4372, w_010_4373, w_010_4374, w_010_4375, w_010_4376, w_010_4377, w_010_4378, w_010_4379, w_010_4380, w_010_4381, w_010_4382, w_010_4383, w_010_4384, w_010_4385, w_010_4386, w_010_4387, w_010_4388, w_010_4389, w_010_4390, w_010_4391, w_010_4392, w_010_4393, w_010_4394, w_010_4395, w_010_4397, w_010_4398, w_010_4399, w_010_4400, w_010_4401, w_010_4402, w_010_4403, w_010_4404, w_010_4405, w_010_4406, w_010_4407, w_010_4408, w_010_4409, w_010_4410, w_010_4411, w_010_4412, w_010_4413, w_010_4414, w_010_4415, w_010_4416, w_010_4417, w_010_4419, w_010_4420, w_010_4421, w_010_4422, w_010_4423, w_010_4424, w_010_4425, w_010_4426, w_010_4427, w_010_4428, w_010_4429, w_010_4430, w_010_4431, w_010_4432, w_010_4433, w_010_4434, w_010_4435, w_010_4436, w_010_4437, w_010_4438, w_010_4439, w_010_4440, w_010_4441, w_010_4442, w_010_4443, w_010_4445, w_010_4446, w_010_4447, w_010_4448, w_010_4449, w_010_4450, w_010_4451, w_010_4452, w_010_4453, w_010_4454, w_010_4456, w_010_4457, w_010_4458, w_010_4460, w_010_4461, w_010_4462, w_010_4463, w_010_4464, w_010_4465, w_010_4466, w_010_4467, w_010_4468, w_010_4469, w_010_4470, w_010_4471, w_010_4472, w_010_4473, w_010_4474, w_010_4476, w_010_4477, w_010_4478, w_010_4479, w_010_4480, w_010_4481, w_010_4482, w_010_4483, w_010_4485, w_010_4486, w_010_4487, w_010_4488, w_010_4489, w_010_4490, w_010_4492, w_010_4493, w_010_4494, w_010_4495, w_010_4496, w_010_4497, w_010_4499, w_010_4500, w_010_4501, w_010_4502, w_010_4503, w_010_4504, w_010_4505, w_010_4506, w_010_4507, w_010_4508, w_010_4509, w_010_4510, w_010_4511, w_010_4512, w_010_4514, w_010_4515, w_010_4516, w_010_4517, w_010_4518, w_010_4519, w_010_4520, w_010_4521, w_010_4522, w_010_4523, w_010_4524, w_010_4525, w_010_4526, w_010_4527, w_010_4528, w_010_4529, w_010_4530, w_010_4531, w_010_4532, w_010_4533, w_010_4534, w_010_4535, w_010_4536, w_010_4537, w_010_4538, w_010_4539, w_010_4540, w_010_4541, w_010_4542, w_010_4543, w_010_4544, w_010_4546, w_010_4547, w_010_4548, w_010_4549, w_010_4550, w_010_4551, w_010_4552, w_010_4553, w_010_4554, w_010_4555, w_010_4556, w_010_4557, w_010_4558, w_010_4559, w_010_4560, w_010_4561, w_010_4562, w_010_4563, w_010_4564, w_010_4565, w_010_4566, w_010_4567, w_010_4568, w_010_4569, w_010_4570, w_010_4571, w_010_4573, w_010_4574, w_010_4575, w_010_4576, w_010_4577, w_010_4578, w_010_4579, w_010_4580, w_010_4581, w_010_4582, w_010_4583, w_010_4584, w_010_4585, w_010_4586, w_010_4587, w_010_4588, w_010_4589, w_010_4590, w_010_4592, w_010_4593, w_010_4595, w_010_4596, w_010_4597, w_010_4600, w_010_4601, w_010_4602, w_010_4603, w_010_4604, w_010_4605, w_010_4606, w_010_4607, w_010_4608, w_010_4609, w_010_4610, w_010_4611, w_010_4612, w_010_4613, w_010_4614, w_010_4615, w_010_4616, w_010_4617, w_010_4619, w_010_4620, w_010_4621, w_010_4622, w_010_4623, w_010_4625, w_010_4627, w_010_4628, w_010_4629, w_010_4630, w_010_4631, w_010_4632, w_010_4633, w_010_4635, w_010_4636, w_010_4637, w_010_4638, w_010_4639, w_010_4641, w_010_4642, w_010_4643, w_010_4644, w_010_4645, w_010_4646, w_010_4647, w_010_4648, w_010_4649, w_010_4650, w_010_4651, w_010_4652, w_010_4653, w_010_4654, w_010_4655, w_010_4656, w_010_4657, w_010_4658, w_010_4659, w_010_4660, w_010_4661, w_010_4662, w_010_4663, w_010_4664, w_010_4665, w_010_4666, w_010_4668, w_010_4669, w_010_4670, w_010_4671, w_010_4672, w_010_4673, w_010_4674, w_010_4675, w_010_4677, w_010_4678, w_010_4679, w_010_4680, w_010_4681, w_010_4682, w_010_4683, w_010_4684, w_010_4685, w_010_4686, w_010_4688, w_010_4689, w_010_4690, w_010_4691, w_010_4692, w_010_4693, w_010_4695, w_010_4696, w_010_4697, w_010_4698, w_010_4699, w_010_4700, w_010_4701, w_010_4702, w_010_4703, w_010_4704, w_010_4705, w_010_4708, w_010_4709, w_010_4711, w_010_4712, w_010_4713, w_010_4714, w_010_4717, w_010_4718, w_010_4719, w_010_4721, w_010_4722, w_010_4724, w_010_4725, w_010_4726, w_010_4727, w_010_4728, w_010_4729, w_010_4731, w_010_4734, w_010_4737, w_010_4738, w_010_4740, w_010_4741, w_010_4742, w_010_4744, w_010_4746, w_010_4747, w_010_4748, w_010_4749, w_010_4750, w_010_4752, w_010_4753, w_010_4754, w_010_4756, w_010_4757, w_010_4758, w_010_4759, w_010_4761, w_010_4762, w_010_4763, w_010_4764, w_010_4765, w_010_4767, w_010_4768, w_010_4770, w_010_4771, w_010_4772, w_010_4773, w_010_4774, w_010_4775, w_010_4776, w_010_4780, w_010_4781, w_010_4783, w_010_4784, w_010_4785, w_010_4786, w_010_4787, w_010_4788, w_010_4790, w_010_4794, w_010_4795, w_010_4796, w_010_4797, w_010_4798, w_010_4799, w_010_4800, w_010_4801, w_010_4802, w_010_4803, w_010_4804, w_010_4805, w_010_4806, w_010_4807, w_010_4808, w_010_4809, w_010_4810, w_010_4812, w_010_4813, w_010_4816, w_010_4820, w_010_4821, w_010_4822, w_010_4824, w_010_4826, w_010_4827, w_010_4828, w_010_4829, w_010_4830, w_010_4831, w_010_4832, w_010_4833, w_010_4834, w_010_4835, w_010_4836, w_010_4837, w_010_4839, w_010_4840, w_010_4841, w_010_4843, w_010_4845, w_010_4846, w_010_4847, w_010_4848, w_010_4849, w_010_4851, w_010_4853, w_010_4854, w_010_4856, w_010_4857, w_010_4859, w_010_4861, w_010_4862, w_010_4863, w_010_4865, w_010_4866, w_010_4867, w_010_4868, w_010_4870, w_010_4871, w_010_4872, w_010_4873, w_010_4875, w_010_4877, w_010_4878, w_010_4879, w_010_4882, w_010_4885, w_010_4887, w_010_4888, w_010_4889, w_010_4890, w_010_4891, w_010_4894, w_010_4895, w_010_4896, w_010_4900, w_010_4901, w_010_4902, w_010_4904, w_010_4905, w_010_4906, w_010_4907, w_010_4910, w_010_4911, w_010_4912, w_010_4913, w_010_4914, w_010_4915, w_010_4917, w_010_4918, w_010_4919, w_010_4920, w_010_4921, w_010_4922, w_010_4923, w_010_4924, w_010_4926, w_010_4927, w_010_4928, w_010_4930, w_010_4931, w_010_4932, w_010_4933, w_010_4934, w_010_4936, w_010_4937, w_010_4941, w_010_4942, w_010_4946, w_010_4948, w_010_4949, w_010_4950, w_010_4951, w_010_4952, w_010_4953, w_010_4954, w_010_4955, w_010_4956, w_010_4957, w_010_4958, w_010_4959, w_010_4960, w_010_4961, w_010_4962, w_010_4963, w_010_4964, w_010_4965, w_010_4966, w_010_4967, w_010_4968, w_010_4969, w_010_4970, w_010_4971, w_010_4972, w_010_4973, w_010_4974, w_010_4975, w_010_4977, w_010_4979, w_010_4980, w_010_4981, w_010_4983, w_010_4984, w_010_4985, w_010_4987, w_010_4988, w_010_4989, w_010_4993, w_010_4994, w_010_4996, w_010_4997, w_010_4999, w_010_5000, w_010_5001, w_010_5002, w_010_5003, w_010_5004, w_010_5006, w_010_5007, w_010_5008, w_010_5009, w_010_5010, w_010_5011, w_010_5012, w_010_5014, w_010_5016, w_010_5017, w_010_5018, w_010_5019, w_010_5020, w_010_5022, w_010_5025, w_010_5026, w_010_5027, w_010_5028, w_010_5029, w_010_5030, w_010_5031, w_010_5032, w_010_5034, w_010_5035, w_010_5036, w_010_5037, w_010_5039, w_010_5040, w_010_5041, w_010_5042, w_010_5043, w_010_5044, w_010_5045, w_010_5047, w_010_5048, w_010_5049, w_010_5050, w_010_5051, w_010_5052, w_010_5053, w_010_5054, w_010_5055, w_010_5056, w_010_5057, w_010_5058, w_010_5059, w_010_5060, w_010_5061, w_010_5063, w_010_5064, w_010_5065, w_010_5066, w_010_5068, w_010_5069, w_010_5071, w_010_5072, w_010_5073, w_010_5074, w_010_5075, w_010_5076, w_010_5077, w_010_5080, w_010_5081, w_010_5082, w_010_5083, w_010_5084, w_010_5085, w_010_5088, w_010_5089, w_010_5090, w_010_5091, w_010_5094, w_010_5095, w_010_5096, w_010_5097, w_010_5098, w_010_5100, w_010_5101, w_010_5103, w_010_5104, w_010_5105, w_010_5109, w_010_5110, w_010_5113, w_010_5115, w_010_5116, w_010_5118, w_010_5119, w_010_5120, w_010_5121, w_010_5122, w_010_5124, w_010_5125, w_010_5126, w_010_5127, w_010_5128, w_010_5129, w_010_5131, w_010_5132, w_010_5133, w_010_5138, w_010_5139, w_010_5140, w_010_5141, w_010_5142, w_010_5143, w_010_5144, w_010_5145, w_010_5147, w_010_5148, w_010_5149, w_010_5150, w_010_5151, w_010_5152, w_010_5153, w_010_5154, w_010_5155, w_010_5156, w_010_5158, w_010_5160, w_010_5161, w_010_5162, w_010_5164, w_010_5166, w_010_5167, w_010_5168, w_010_5169, w_010_5170, w_010_5173, w_010_5174, w_010_5175, w_010_5177, w_010_5178, w_010_5179, w_010_5180, w_010_5182, w_010_5183, w_010_5184, w_010_5185, w_010_5186, w_010_5189, w_010_5190, w_010_5191, w_010_5192, w_010_5193, w_010_5194, w_010_5195, w_010_5196, w_010_5198, w_010_5199, w_010_5200, w_010_5201, w_010_5202, w_010_5203, w_010_5204, w_010_5205, w_010_5206, w_010_5207, w_010_5208, w_010_5210, w_010_5211, w_010_5212, w_010_5213, w_010_5214, w_010_5215, w_010_5216, w_010_5217, w_010_5218, w_010_5219, w_010_5220, w_010_5222, w_010_5223, w_010_5224, w_010_5225, w_010_5226, w_010_5228, w_010_5229, w_010_5231, w_010_5232, w_010_5233, w_010_5234, w_010_5235, w_010_5236, w_010_5237, w_010_5238, w_010_5239, w_010_5240, w_010_5241, w_010_5242, w_010_5243, w_010_5244, w_010_5245, w_010_5246, w_010_5247, w_010_5249, w_010_5250, w_010_5252, w_010_5255, w_010_5256, w_010_5257, w_010_5258, w_010_5260, w_010_5261, w_010_5264, w_010_5265, w_010_5266, w_010_5267, w_010_5268, w_010_5269, w_010_5270, w_010_5271, w_010_5273, w_010_5274, w_010_5275, w_010_5276, w_010_5277, w_010_5280, w_010_5282, w_010_5283, w_010_5285, w_010_5286, w_010_5287, w_010_5288, w_010_5289, w_010_5290, w_010_5291, w_010_5292, w_010_5294, w_010_5295, w_010_5296, w_010_5297, w_010_5300, w_010_5301, w_010_5302, w_010_5303, w_010_5304, w_010_5305, w_010_5307, w_010_5308, w_010_5309, w_010_5311, w_010_5312, w_010_5314, w_010_5315, w_010_5316, w_010_5317, w_010_5318, w_010_5319, w_010_5320, w_010_5321, w_010_5322, w_010_5323;
  wire w_011_000, w_011_001, w_011_002, w_011_003, w_011_004, w_011_005, w_011_006, w_011_007, w_011_008, w_011_009, w_011_010, w_011_011, w_011_012, w_011_014, w_011_015, w_011_016, w_011_017, w_011_018, w_011_019, w_011_020, w_011_021, w_011_022, w_011_023, w_011_024, w_011_025, w_011_027, w_011_028, w_011_029, w_011_030, w_011_031, w_011_032, w_011_033, w_011_034, w_011_035, w_011_036, w_011_037, w_011_039, w_011_041, w_011_042, w_011_043, w_011_044, w_011_046, w_011_047, w_011_048, w_011_049, w_011_050, w_011_052, w_011_054, w_011_055, w_011_056, w_011_057, w_011_058, w_011_059, w_011_061, w_011_062, w_011_063, w_011_064, w_011_065, w_011_066, w_011_067, w_011_068, w_011_070, w_011_071, w_011_072, w_011_073, w_011_074, w_011_075, w_011_076, w_011_077, w_011_078, w_011_079, w_011_080, w_011_081, w_011_082, w_011_083, w_011_084, w_011_085, w_011_086, w_011_087, w_011_088, w_011_089, w_011_090, w_011_091, w_011_092, w_011_093, w_011_094, w_011_095, w_011_096, w_011_097, w_011_098, w_011_099, w_011_100, w_011_101, w_011_102, w_011_103, w_011_104, w_011_106, w_011_107, w_011_108, w_011_109, w_011_110, w_011_111, w_011_112, w_011_113, w_011_114, w_011_115, w_011_116, w_011_117, w_011_119, w_011_120, w_011_122, w_011_123, w_011_124, w_011_126, w_011_127, w_011_128, w_011_129, w_011_130, w_011_131, w_011_132, w_011_133, w_011_134, w_011_135, w_011_136, w_011_137, w_011_138, w_011_140, w_011_141, w_011_142, w_011_143, w_011_144, w_011_145, w_011_146, w_011_147, w_011_148, w_011_149, w_011_150, w_011_151, w_011_152, w_011_153, w_011_154, w_011_155, w_011_157, w_011_158, w_011_159, w_011_160, w_011_161, w_011_163, w_011_164, w_011_165, w_011_166, w_011_167, w_011_171, w_011_173, w_011_174, w_011_175, w_011_176, w_011_177, w_011_178, w_011_179, w_011_180, w_011_181, w_011_182, w_011_183, w_011_184, w_011_185, w_011_186, w_011_187, w_011_188, w_011_189, w_011_190, w_011_191, w_011_192, w_011_193, w_011_194, w_011_195, w_011_196, w_011_198, w_011_199, w_011_200, w_011_202, w_011_203, w_011_204, w_011_205, w_011_206, w_011_207, w_011_208, w_011_209, w_011_210, w_011_211, w_011_212, w_011_213, w_011_214, w_011_215, w_011_216, w_011_217, w_011_218, w_011_219, w_011_220, w_011_221, w_011_222, w_011_224, w_011_225, w_011_226, w_011_227, w_011_228, w_011_229, w_011_230, w_011_231, w_011_232, w_011_233, w_011_234, w_011_235, w_011_236, w_011_238, w_011_239, w_011_240, w_011_241, w_011_242, w_011_243, w_011_244, w_011_245, w_011_246, w_011_248, w_011_249, w_011_250, w_011_251, w_011_252, w_011_253, w_011_254, w_011_255, w_011_256, w_011_257, w_011_258, w_011_259, w_011_260, w_011_261, w_011_262, w_011_263, w_011_264, w_011_265, w_011_266, w_011_267, w_011_268, w_011_270, w_011_271, w_011_272, w_011_273, w_011_274, w_011_275, w_011_276, w_011_277, w_011_279, w_011_280, w_011_281, w_011_282, w_011_283, w_011_284, w_011_285, w_011_286, w_011_287, w_011_288, w_011_289, w_011_290, w_011_291, w_011_292, w_011_293, w_011_294, w_011_295, w_011_296, w_011_297, w_011_298, w_011_299, w_011_301, w_011_302, w_011_303, w_011_304, w_011_305, w_011_306, w_011_308, w_011_309, w_011_310, w_011_311, w_011_313, w_011_314, w_011_315, w_011_316, w_011_318, w_011_319, w_011_320, w_011_321, w_011_322, w_011_323, w_011_324, w_011_325, w_011_326, w_011_327, w_011_328, w_011_329, w_011_330, w_011_331, w_011_332, w_011_333, w_011_334, w_011_335, w_011_336, w_011_338, w_011_339, w_011_340, w_011_341, w_011_342, w_011_343, w_011_344, w_011_345, w_011_346, w_011_347, w_011_348, w_011_349, w_011_350, w_011_351, w_011_352, w_011_353, w_011_354, w_011_355, w_011_356, w_011_357, w_011_358, w_011_359, w_011_360, w_011_361, w_011_362, w_011_363, w_011_364, w_011_366, w_011_367, w_011_369, w_011_370, w_011_371, w_011_372, w_011_373, w_011_374, w_011_375, w_011_376, w_011_377, w_011_378, w_011_379, w_011_380, w_011_381, w_011_382, w_011_383, w_011_384, w_011_385, w_011_386, w_011_387, w_011_388, w_011_389, w_011_390, w_011_391, w_011_393, w_011_394, w_011_395, w_011_396, w_011_397, w_011_398, w_011_399, w_011_400, w_011_401, w_011_402, w_011_403, w_011_404, w_011_406, w_011_407, w_011_408, w_011_409, w_011_410, w_011_411, w_011_412, w_011_413, w_011_414, w_011_415, w_011_416, w_011_417, w_011_418, w_011_419, w_011_420, w_011_421, w_011_422, w_011_423, w_011_424, w_011_425, w_011_426, w_011_427, w_011_428, w_011_429, w_011_430, w_011_431, w_011_432, w_011_434, w_011_435, w_011_436, w_011_437, w_011_438, w_011_439, w_011_441, w_011_442, w_011_443, w_011_444, w_011_445, w_011_446, w_011_447, w_011_448, w_011_449, w_011_450, w_011_451, w_011_452, w_011_453, w_011_454, w_011_455, w_011_457, w_011_458, w_011_459, w_011_460, w_011_461, w_011_462, w_011_463, w_011_464, w_011_465, w_011_466, w_011_467, w_011_468, w_011_469, w_011_470, w_011_471, w_011_472, w_011_473, w_011_474, w_011_475, w_011_476, w_011_477, w_011_479, w_011_480, w_011_482, w_011_483, w_011_484, w_011_485, w_011_486, w_011_487, w_011_488, w_011_489, w_011_491, w_011_492, w_011_493, w_011_494, w_011_495, w_011_496, w_011_497, w_011_498, w_011_499, w_011_500, w_011_502, w_011_503, w_011_504, w_011_505, w_011_506, w_011_507, w_011_508, w_011_509, w_011_510, w_011_511, w_011_512, w_011_513, w_011_514, w_011_515, w_011_516, w_011_517, w_011_518, w_011_519, w_011_520, w_011_521, w_011_522, w_011_523, w_011_524, w_011_525, w_011_526, w_011_528, w_011_530, w_011_531, w_011_532, w_011_533, w_011_534, w_011_535, w_011_536, w_011_537, w_011_539, w_011_540, w_011_541, w_011_542, w_011_543, w_011_544, w_011_545, w_011_546, w_011_547, w_011_548, w_011_549, w_011_550, w_011_551, w_011_552, w_011_553, w_011_554, w_011_555, w_011_556, w_011_557, w_011_558, w_011_559, w_011_560, w_011_561, w_011_562, w_011_563, w_011_564, w_011_565, w_011_566, w_011_567, w_011_568, w_011_569, w_011_571, w_011_572, w_011_573, w_011_574, w_011_575, w_011_576, w_011_577, w_011_578, w_011_579, w_011_580, w_011_581, w_011_582, w_011_583, w_011_584, w_011_585, w_011_586, w_011_587, w_011_589, w_011_590, w_011_591, w_011_592, w_011_596, w_011_597, w_011_598, w_011_599, w_011_600, w_011_601, w_011_602, w_011_603, w_011_604, w_011_605, w_011_606, w_011_607, w_011_608, w_011_609, w_011_610, w_011_611, w_011_612, w_011_613, w_011_614, w_011_615, w_011_616, w_011_617, w_011_618, w_011_619, w_011_620, w_011_622, w_011_623, w_011_624, w_011_625, w_011_626, w_011_627, w_011_628, w_011_629, w_011_630, w_011_631, w_011_632, w_011_633, w_011_634, w_011_635, w_011_636, w_011_637, w_011_638, w_011_639, w_011_640, w_011_641, w_011_642, w_011_643, w_011_644, w_011_645, w_011_646, w_011_648, w_011_649, w_011_652, w_011_653, w_011_654, w_011_655, w_011_656, w_011_657, w_011_658, w_011_659, w_011_660, w_011_661, w_011_662, w_011_663, w_011_664, w_011_665, w_011_666, w_011_667, w_011_670, w_011_671, w_011_672, w_011_673, w_011_674, w_011_675, w_011_676, w_011_677, w_011_678, w_011_679, w_011_680, w_011_681, w_011_682, w_011_684, w_011_685, w_011_687, w_011_688, w_011_689, w_011_690, w_011_691, w_011_692, w_011_693, w_011_696, w_011_697, w_011_698, w_011_699, w_011_700, w_011_701, w_011_702, w_011_703, w_011_704, w_011_705, w_011_706, w_011_707, w_011_708, w_011_709, w_011_710, w_011_712, w_011_713, w_011_715, w_011_716, w_011_718, w_011_719, w_011_720, w_011_721, w_011_722, w_011_723, w_011_726, w_011_727, w_011_728, w_011_729, w_011_730, w_011_731, w_011_732, w_011_733, w_011_735, w_011_736, w_011_737, w_011_738, w_011_739, w_011_740, w_011_741, w_011_742, w_011_743, w_011_744, w_011_745, w_011_746, w_011_747, w_011_748, w_011_749, w_011_750, w_011_751, w_011_752, w_011_753, w_011_754, w_011_755, w_011_756, w_011_757, w_011_758, w_011_759, w_011_760, w_011_761, w_011_763, w_011_764, w_011_765, w_011_767, w_011_768, w_011_769, w_011_770, w_011_771, w_011_772, w_011_773, w_011_774, w_011_775, w_011_776, w_011_777, w_011_778, w_011_779, w_011_780, w_011_781, w_011_782, w_011_783, w_011_784, w_011_786, w_011_787, w_011_788, w_011_789, w_011_790, w_011_791, w_011_792, w_011_793, w_011_794, w_011_795, w_011_796, w_011_797, w_011_798, w_011_799, w_011_800, w_011_802, w_011_803, w_011_804, w_011_805, w_011_806, w_011_807, w_011_809, w_011_811, w_011_812, w_011_813, w_011_814, w_011_815, w_011_816, w_011_817, w_011_818, w_011_819, w_011_820, w_011_821, w_011_822, w_011_823, w_011_824, w_011_825, w_011_826, w_011_827, w_011_828, w_011_829, w_011_830, w_011_831, w_011_832, w_011_833, w_011_834, w_011_835, w_011_836, w_011_837, w_011_838, w_011_839, w_011_840, w_011_841, w_011_843, w_011_844, w_011_845, w_011_846, w_011_847, w_011_848, w_011_851, w_011_852, w_011_854, w_011_855, w_011_856, w_011_860, w_011_861, w_011_862, w_011_863, w_011_866, w_011_867, w_011_868, w_011_869, w_011_870, w_011_871, w_011_872, w_011_873, w_011_874, w_011_875, w_011_877, w_011_878, w_011_879, w_011_880, w_011_881, w_011_882, w_011_884, w_011_885, w_011_886, w_011_889, w_011_890, w_011_892, w_011_894, w_011_897, w_011_898, w_011_899, w_011_900, w_011_901, w_011_903, w_011_904, w_011_905, w_011_908, w_011_910, w_011_911, w_011_913, w_011_914, w_011_915, w_011_916, w_011_918, w_011_921, w_011_922, w_011_923, w_011_924, w_011_925, w_011_926, w_011_927, w_011_928, w_011_929, w_011_930, w_011_931, w_011_933, w_011_935, w_011_936, w_011_937, w_011_938, w_011_939, w_011_940, w_011_941, w_011_943, w_011_944, w_011_945, w_011_946, w_011_947, w_011_948, w_011_949, w_011_951, w_011_952, w_011_953, w_011_954, w_011_955, w_011_956, w_011_957, w_011_958, w_011_959, w_011_961, w_011_962, w_011_963, w_011_964, w_011_965, w_011_967, w_011_968, w_011_969, w_011_970, w_011_972, w_011_973, w_011_974, w_011_975, w_011_976, w_011_980, w_011_981, w_011_982, w_011_983, w_011_985, w_011_986, w_011_987, w_011_988, w_011_989, w_011_990, w_011_991, w_011_993, w_011_994, w_011_995, w_011_996, w_011_997, w_011_998, w_011_999, w_011_1001, w_011_1002, w_011_1005, w_011_1006, w_011_1007, w_011_1009, w_011_1011, w_011_1013, w_011_1014, w_011_1015, w_011_1017, w_011_1019, w_011_1021, w_011_1023, w_011_1024, w_011_1026, w_011_1027, w_011_1028, w_011_1030, w_011_1032, w_011_1033, w_011_1036, w_011_1037, w_011_1038, w_011_1039, w_011_1042, w_011_1043, w_011_1045, w_011_1046, w_011_1048, w_011_1049, w_011_1050, w_011_1051, w_011_1052, w_011_1054, w_011_1055, w_011_1056, w_011_1057, w_011_1058, w_011_1059, w_011_1060, w_011_1062, w_011_1063, w_011_1064, w_011_1065, w_011_1066, w_011_1067, w_011_1068, w_011_1069, w_011_1070, w_011_1072, w_011_1073, w_011_1074, w_011_1076, w_011_1077, w_011_1079, w_011_1080, w_011_1081, w_011_1082, w_011_1083, w_011_1084, w_011_1085, w_011_1086, w_011_1087, w_011_1088, w_011_1090, w_011_1091, w_011_1092, w_011_1093, w_011_1095, w_011_1097, w_011_1098, w_011_1099, w_011_1100, w_011_1101, w_011_1102, w_011_1103, w_011_1104, w_011_1105, w_011_1106, w_011_1108, w_011_1109, w_011_1110, w_011_1112, w_011_1113, w_011_1114, w_011_1115, w_011_1116, w_011_1117, w_011_1119, w_011_1120, w_011_1121, w_011_1123, w_011_1124, w_011_1125, w_011_1126, w_011_1127, w_011_1128, w_011_1129, w_011_1130, w_011_1131, w_011_1132, w_011_1133, w_011_1134, w_011_1135, w_011_1137, w_011_1138, w_011_1139, w_011_1140, w_011_1141, w_011_1142, w_011_1143, w_011_1144, w_011_1145, w_011_1146, w_011_1147, w_011_1149, w_011_1152, w_011_1154, w_011_1155, w_011_1156, w_011_1157, w_011_1158, w_011_1161, w_011_1164, w_011_1165, w_011_1169, w_011_1171, w_011_1172, w_011_1173, w_011_1174, w_011_1178, w_011_1180, w_011_1185, w_011_1186, w_011_1187, w_011_1188, w_011_1189, w_011_1191, w_011_1192, w_011_1193, w_011_1194, w_011_1196, w_011_1197, w_011_1199, w_011_1202, w_011_1203, w_011_1204, w_011_1209, w_011_1210, w_011_1212, w_011_1214, w_011_1216, w_011_1217, w_011_1219, w_011_1220, w_011_1223, w_011_1226, w_011_1227, w_011_1228, w_011_1229, w_011_1230, w_011_1231, w_011_1232, w_011_1234, w_011_1235, w_011_1236, w_011_1237, w_011_1238, w_011_1239, w_011_1240, w_011_1242, w_011_1243, w_011_1247, w_011_1250, w_011_1251, w_011_1252, w_011_1253, w_011_1255, w_011_1256, w_011_1258, w_011_1260, w_011_1262, w_011_1263, w_011_1264, w_011_1265, w_011_1266, w_011_1267, w_011_1268, w_011_1271, w_011_1274, w_011_1275, w_011_1276, w_011_1277, w_011_1278, w_011_1279, w_011_1281, w_011_1282, w_011_1283, w_011_1284, w_011_1286, w_011_1288, w_011_1289, w_011_1291, w_011_1293, w_011_1294, w_011_1296, w_011_1298, w_011_1299, w_011_1300, w_011_1301, w_011_1302, w_011_1304, w_011_1306, w_011_1308, w_011_1309, w_011_1310, w_011_1311, w_011_1312, w_011_1313, w_011_1314, w_011_1316, w_011_1317, w_011_1318, w_011_1319, w_011_1320, w_011_1321, w_011_1322, w_011_1323, w_011_1324, w_011_1327, w_011_1329, w_011_1331, w_011_1332, w_011_1333, w_011_1334, w_011_1335, w_011_1337, w_011_1338, w_011_1339, w_011_1340, w_011_1341, w_011_1343, w_011_1344, w_011_1345, w_011_1346, w_011_1347, w_011_1348, w_011_1350, w_011_1352, w_011_1353, w_011_1354, w_011_1356, w_011_1357, w_011_1358, w_011_1359, w_011_1361, w_011_1364, w_011_1365, w_011_1366, w_011_1367, w_011_1368, w_011_1369, w_011_1372, w_011_1373, w_011_1374, w_011_1375, w_011_1376, w_011_1377, w_011_1378, w_011_1379, w_011_1380, w_011_1381, w_011_1385, w_011_1386, w_011_1388, w_011_1389, w_011_1391, w_011_1392, w_011_1394, w_011_1395, w_011_1397, w_011_1398, w_011_1399, w_011_1400, w_011_1402, w_011_1403, w_011_1405, w_011_1406, w_011_1408, w_011_1410, w_011_1411, w_011_1414, w_011_1416, w_011_1417, w_011_1418, w_011_1420, w_011_1421, w_011_1422, w_011_1423, w_011_1424, w_011_1425, w_011_1426, w_011_1427, w_011_1429, w_011_1430, w_011_1431, w_011_1432, w_011_1434, w_011_1435, w_011_1437, w_011_1439, w_011_1440, w_011_1441, w_011_1442, w_011_1444, w_011_1445, w_011_1446, w_011_1447, w_011_1448, w_011_1449, w_011_1453, w_011_1454, w_011_1455, w_011_1456, w_011_1457, w_011_1458, w_011_1459, w_011_1460, w_011_1461, w_011_1462, w_011_1463, w_011_1464, w_011_1465, w_011_1466, w_011_1468, w_011_1471, w_011_1473, w_011_1474, w_011_1475, w_011_1476, w_011_1477, w_011_1478, w_011_1479, w_011_1480, w_011_1481, w_011_1482, w_011_1483, w_011_1484, w_011_1485, w_011_1486, w_011_1487, w_011_1488, w_011_1489, w_011_1490, w_011_1491, w_011_1492, w_011_1493, w_011_1496, w_011_1497, w_011_1498, w_011_1499, w_011_1500, w_011_1501, w_011_1502, w_011_1504, w_011_1508, w_011_1509, w_011_1512, w_011_1513, w_011_1514, w_011_1516, w_011_1517, w_011_1518, w_011_1519, w_011_1520, w_011_1521, w_011_1522, w_011_1523, w_011_1524, w_011_1525, w_011_1526, w_011_1527, w_011_1528, w_011_1529, w_011_1530, w_011_1531, w_011_1533, w_011_1534, w_011_1535, w_011_1538, w_011_1539, w_011_1540, w_011_1541, w_011_1542, w_011_1543, w_011_1545, w_011_1546, w_011_1550, w_011_1551, w_011_1552, w_011_1554, w_011_1555, w_011_1556, w_011_1558, w_011_1559, w_011_1561, w_011_1562, w_011_1564, w_011_1565, w_011_1566, w_011_1567, w_011_1569, w_011_1571, w_011_1572, w_011_1573, w_011_1574, w_011_1575, w_011_1576, w_011_1577, w_011_1580, w_011_1582, w_011_1583, w_011_1584, w_011_1587, w_011_1588, w_011_1589, w_011_1591, w_011_1593, w_011_1594, w_011_1596, w_011_1597, w_011_1598, w_011_1600, w_011_1601, w_011_1602, w_011_1603, w_011_1604, w_011_1605, w_011_1606, w_011_1607, w_011_1609, w_011_1611, w_011_1612, w_011_1613, w_011_1615, w_011_1617, w_011_1619, w_011_1621, w_011_1622, w_011_1623, w_011_1626, w_011_1627, w_011_1629, w_011_1633, w_011_1634, w_011_1635, w_011_1636, w_011_1637, w_011_1638, w_011_1640, w_011_1641, w_011_1642, w_011_1644, w_011_1646, w_011_1649, w_011_1650, w_011_1651, w_011_1652, w_011_1654, w_011_1657, w_011_1658, w_011_1659, w_011_1660, w_011_1661, w_011_1664, w_011_1666, w_011_1667, w_011_1668, w_011_1672, w_011_1673, w_011_1674, w_011_1675, w_011_1676, w_011_1677, w_011_1678, w_011_1679, w_011_1681, w_011_1682, w_011_1683, w_011_1684, w_011_1685, w_011_1686, w_011_1687, w_011_1689, w_011_1690, w_011_1692, w_011_1695, w_011_1696, w_011_1698, w_011_1699, w_011_1700, w_011_1701, w_011_1704, w_011_1705, w_011_1706, w_011_1708, w_011_1711, w_011_1713, w_011_1714, w_011_1715, w_011_1716, w_011_1717, w_011_1718, w_011_1719, w_011_1722, w_011_1723, w_011_1724, w_011_1725, w_011_1726, w_011_1730, w_011_1732, w_011_1733, w_011_1735, w_011_1736, w_011_1737, w_011_1739, w_011_1740, w_011_1742, w_011_1745, w_011_1747, w_011_1748, w_011_1749, w_011_1750, w_011_1751, w_011_1754, w_011_1755, w_011_1756, w_011_1757, w_011_1758, w_011_1759, w_011_1760, w_011_1763, w_011_1764, w_011_1765, w_011_1767, w_011_1768, w_011_1770, w_011_1771, w_011_1773, w_011_1774, w_011_1776, w_011_1777, w_011_1778, w_011_1780, w_011_1781, w_011_1783, w_011_1784, w_011_1785, w_011_1786, w_011_1787, w_011_1788, w_011_1789, w_011_1791, w_011_1792, w_011_1793, w_011_1794, w_011_1795, w_011_1796, w_011_1798, w_011_1799, w_011_1802, w_011_1805, w_011_1807, w_011_1808, w_011_1809, w_011_1810, w_011_1811, w_011_1812, w_011_1813, w_011_1814, w_011_1815, w_011_1816, w_011_1818, w_011_1819, w_011_1821, w_011_1823, w_011_1824, w_011_1826, w_011_1827, w_011_1830, w_011_1831, w_011_1832, w_011_1833, w_011_1834, w_011_1836, w_011_1837, w_011_1838, w_011_1839, w_011_1840, w_011_1841, w_011_1842, w_011_1844, w_011_1845, w_011_1847, w_011_1848, w_011_1851, w_011_1852, w_011_1855, w_011_1856, w_011_1858, w_011_1859, w_011_1860, w_011_1861, w_011_1862, w_011_1863, w_011_1864, w_011_1865, w_011_1867, w_011_1868, w_011_1870, w_011_1872, w_011_1873, w_011_1874, w_011_1876, w_011_1877, w_011_1878, w_011_1879, w_011_1882, w_011_1883, w_011_1884, w_011_1885, w_011_1886, w_011_1889, w_011_1891, w_011_1892, w_011_1893, w_011_1894, w_011_1895, w_011_1896, w_011_1897, w_011_1898, w_011_1899, w_011_1900, w_011_1903, w_011_1904, w_011_1905, w_011_1906, w_011_1907, w_011_1908, w_011_1909, w_011_1910, w_011_1911, w_011_1912, w_011_1913, w_011_1915, w_011_1917, w_011_1918, w_011_1919, w_011_1920, w_011_1921, w_011_1922, w_011_1923, w_011_1924, w_011_1925, w_011_1927, w_011_1928, w_011_1933, w_011_1934, w_011_1935, w_011_1936, w_011_1937, w_011_1940, w_011_1942, w_011_1943, w_011_1945, w_011_1946, w_011_1947, w_011_1949, w_011_1950, w_011_1953, w_011_1954, w_011_1955, w_011_1956, w_011_1957, w_011_1958, w_011_1959, w_011_1960, w_011_1961, w_011_1962, w_011_1963, w_011_1964, w_011_1965, w_011_1966, w_011_1967, w_011_1968, w_011_1969, w_011_1970, w_011_1971, w_011_1972, w_011_1973, w_011_1975, w_011_1976, w_011_1977, w_011_1978, w_011_1979, w_011_1981, w_011_1982, w_011_1983, w_011_1984, w_011_1985, w_011_1986, w_011_1987, w_011_1988, w_011_1990, w_011_1991, w_011_1993, w_011_1995, w_011_2000, w_011_2001, w_011_2002, w_011_2003, w_011_2004, w_011_2005, w_011_2006, w_011_2007, w_011_2010, w_011_2013, w_011_2014, w_011_2015, w_011_2017, w_011_2019, w_011_2020, w_011_2021, w_011_2022, w_011_2023, w_011_2024, w_011_2027, w_011_2028, w_011_2029, w_011_2031, w_011_2035, w_011_2037, w_011_2040, w_011_2042, w_011_2043, w_011_2045, w_011_2047, w_011_2048, w_011_2049, w_011_2050, w_011_2051, w_011_2053, w_011_2054, w_011_2056, w_011_2061, w_011_2062, w_011_2063, w_011_2066, w_011_2067, w_011_2068, w_011_2071, w_011_2073, w_011_2075, w_011_2079, w_011_2080, w_011_2081, w_011_2082, w_011_2083, w_011_2084, w_011_2085, w_011_2086, w_011_2088, w_011_2089, w_011_2090, w_011_2092, w_011_2093, w_011_2094, w_011_2095, w_011_2097, w_011_2099, w_011_2100, w_011_2102, w_011_2103, w_011_2105, w_011_2107, w_011_2108, w_011_2110, w_011_2112, w_011_2114, w_011_2115, w_011_2116, w_011_2117, w_011_2120, w_011_2121, w_011_2123, w_011_2124, w_011_2125, w_011_2127, w_011_2128, w_011_2129, w_011_2130, w_011_2131, w_011_2132, w_011_2133, w_011_2134, w_011_2135, w_011_2136, w_011_2137, w_011_2139, w_011_2142, w_011_2144, w_011_2146, w_011_2147, w_011_2150, w_011_2151, w_011_2155, w_011_2157, w_011_2158, w_011_2159, w_011_2160, w_011_2161, w_011_2162, w_011_2163, w_011_2166, w_011_2167, w_011_2169, w_011_2170, w_011_2171, w_011_2172, w_011_2173, w_011_2175, w_011_2178, w_011_2181, w_011_2183, w_011_2185, w_011_2186, w_011_2187, w_011_2188, w_011_2189, w_011_2190, w_011_2191, w_011_2192, w_011_2193, w_011_2194, w_011_2195, w_011_2196, w_011_2197, w_011_2198, w_011_2199, w_011_2200, w_011_2201, w_011_2203, w_011_2204, w_011_2205, w_011_2206, w_011_2207, w_011_2208, w_011_2209, w_011_2210, w_011_2211, w_011_2213, w_011_2215, w_011_2216, w_011_2217, w_011_2218, w_011_2219, w_011_2220, w_011_2221, w_011_2222, w_011_2223, w_011_2224, w_011_2227, w_011_2228, w_011_2229, w_011_2230, w_011_2233, w_011_2234, w_011_2235, w_011_2237, w_011_2238, w_011_2239, w_011_2240, w_011_2241, w_011_2242, w_011_2243, w_011_2244, w_011_2245, w_011_2246, w_011_2247, w_011_2248, w_011_2249, w_011_2250, w_011_2251, w_011_2252, w_011_2253, w_011_2254, w_011_2256, w_011_2258, w_011_2259, w_011_2261, w_011_2262, w_011_2263, w_011_2264, w_011_2267, w_011_2269, w_011_2270, w_011_2272, w_011_2273, w_011_2274, w_011_2276, w_011_2277, w_011_2278, w_011_2281, w_011_2282, w_011_2284, w_011_2287, w_011_2289, w_011_2291, w_011_2292, w_011_2293, w_011_2294, w_011_2297, w_011_2298, w_011_2299, w_011_2300, w_011_2301, w_011_2303, w_011_2304, w_011_2305, w_011_2307, w_011_2308, w_011_2309, w_011_2310, w_011_2311, w_011_2314, w_011_2315, w_011_2316, w_011_2317, w_011_2318, w_011_2319, w_011_2320, w_011_2323, w_011_2324, w_011_2325, w_011_2326, w_011_2327, w_011_2330, w_011_2331, w_011_2332, w_011_2333, w_011_2334, w_011_2335, w_011_2336, w_011_2337, w_011_2339, w_011_2340, w_011_2341, w_011_2342, w_011_2344, w_011_2345, w_011_2348, w_011_2350, w_011_2351, w_011_2352, w_011_2353, w_011_2355, w_011_2356, w_011_2357, w_011_2359, w_011_2362, w_011_2363, w_011_2365, w_011_2366, w_011_2367, w_011_2368, w_011_2369, w_011_2372, w_011_2374, w_011_2376, w_011_2377, w_011_2378, w_011_2379, w_011_2382, w_011_2384, w_011_2385, w_011_2386, w_011_2387, w_011_2388, w_011_2390, w_011_2391, w_011_2392, w_011_2393, w_011_2394, w_011_2395, w_011_2398, w_011_2399, w_011_2400, w_011_2401, w_011_2402, w_011_2403, w_011_2404, w_011_2408, w_011_2410, w_011_2411, w_011_2413, w_011_2414, w_011_2415, w_011_2417, w_011_2420, w_011_2421, w_011_2422, w_011_2423, w_011_2424, w_011_2425, w_011_2426, w_011_2428, w_011_2429, w_011_2430, w_011_2431, w_011_2432, w_011_2433, w_011_2435, w_011_2438, w_011_2439, w_011_2440, w_011_2441, w_011_2443, w_011_2444, w_011_2446, w_011_2447, w_011_2448, w_011_2449, w_011_2451, w_011_2452, w_011_2453, w_011_2454, w_011_2455, w_011_2456, w_011_2457, w_011_2458, w_011_2459, w_011_2460, w_011_2462, w_011_2463, w_011_2464, w_011_2465, w_011_2466, w_011_2467, w_011_2469, w_011_2470, w_011_2471, w_011_2472, w_011_2474, w_011_2475, w_011_2476, w_011_2479, w_011_2481, w_011_2482, w_011_2484, w_011_2485, w_011_2486, w_011_2487, w_011_2488, w_011_2490, w_011_2493, w_011_2496, w_011_2497, w_011_2498, w_011_2499, w_011_2500, w_011_2501, w_011_2502, w_011_2503, w_011_2504, w_011_2505, w_011_2506, w_011_2509, w_011_2510, w_011_2511, w_011_2512, w_011_2513, w_011_2514, w_011_2515, w_011_2516, w_011_2517, w_011_2518, w_011_2519, w_011_2520, w_011_2521, w_011_2522, w_011_2523, w_011_2524, w_011_2525, w_011_2526, w_011_2527, w_011_2528, w_011_2530, w_011_2531, w_011_2532, w_011_2533, w_011_2535, w_011_2536, w_011_2537, w_011_2538, w_011_2540, w_011_2541, w_011_2542, w_011_2543, w_011_2544, w_011_2545, w_011_2546, w_011_2547, w_011_2548, w_011_2549, w_011_2550, w_011_2551, w_011_2552, w_011_2553, w_011_2554, w_011_2555, w_011_2556, w_011_2558, w_011_2559, w_011_2560, w_011_2561, w_011_2563, w_011_2565, w_011_2566, w_011_2567, w_011_2568, w_011_2569, w_011_2571, w_011_2573, w_011_2574, w_011_2575, w_011_2576, w_011_2577, w_011_2578, w_011_2579, w_011_2580, w_011_2581, w_011_2582, w_011_2583, w_011_2584, w_011_2586, w_011_2587, w_011_2588, w_011_2589, w_011_2590, w_011_2592, w_011_2593, w_011_2597, w_011_2599, w_011_2600, w_011_2601, w_011_2602, w_011_2603, w_011_2604, w_011_2605, w_011_2607, w_011_2608, w_011_2610, w_011_2613, w_011_2615, w_011_2617, w_011_2619, w_011_2621, w_011_2622, w_011_2624, w_011_2625, w_011_2626, w_011_2627, w_011_2628, w_011_2629, w_011_2630, w_011_2632, w_011_2634, w_011_2635, w_011_2638, w_011_2639, w_011_2642, w_011_2643, w_011_2644, w_011_2645, w_011_2646, w_011_2647, w_011_2649, w_011_2650, w_011_2651, w_011_2652, w_011_2655, w_011_2660, w_011_2661, w_011_2662, w_011_2663, w_011_2665, w_011_2666, w_011_2667, w_011_2668, w_011_2672, w_011_2674, w_011_2675, w_011_2676, w_011_2679, w_011_2680, w_011_2681, w_011_2682, w_011_2683, w_011_2687, w_011_2689, w_011_2690, w_011_2691, w_011_2692, w_011_2693, w_011_2695, w_011_2696, w_011_2697, w_011_2699, w_011_2701, w_011_2702, w_011_2703, w_011_2705, w_011_2706, w_011_2711, w_011_2712, w_011_2713, w_011_2714, w_011_2715, w_011_2716, w_011_2717, w_011_2718, w_011_2719, w_011_2722, w_011_2723, w_011_2724, w_011_2725, w_011_2726, w_011_2727, w_011_2730, w_011_2731, w_011_2733, w_011_2734, w_011_2735, w_011_2738, w_011_2740, w_011_2741, w_011_2742, w_011_2743, w_011_2744, w_011_2748, w_011_2749, w_011_2750, w_011_2752, w_011_2753, w_011_2754, w_011_2755, w_011_2756, w_011_2757, w_011_2758, w_011_2759, w_011_2760, w_011_2764, w_011_2766, w_011_2767, w_011_2769, w_011_2770, w_011_2771, w_011_2772, w_011_2773, w_011_2774, w_011_2775, w_011_2776, w_011_2777, w_011_2779, w_011_2780, w_011_2781, w_011_2783, w_011_2784, w_011_2785, w_011_2787, w_011_2788, w_011_2789, w_011_2790, w_011_2791, w_011_2792, w_011_2793, w_011_2795, w_011_2796, w_011_2797, w_011_2798, w_011_2799, w_011_2800, w_011_2802, w_011_2803, w_011_2804, w_011_2805, w_011_2807, w_011_2808, w_011_2810, w_011_2811, w_011_2812, w_011_2813, w_011_2814, w_011_2815, w_011_2816, w_011_2817, w_011_2818, w_011_2819, w_011_2820, w_011_2823, w_011_2824, w_011_2825, w_011_2828, w_011_2829, w_011_2830, w_011_2831, w_011_2833, w_011_2834, w_011_2835, w_011_2836, w_011_2838, w_011_2839, w_011_2840, w_011_2841, w_011_2844, w_011_2845, w_011_2846, w_011_2849, w_011_2850, w_011_2851, w_011_2852, w_011_2853, w_011_2854, w_011_2855, w_011_2857, w_011_2860, w_011_2863, w_011_2864, w_011_2865, w_011_2868, w_011_2869, w_011_2870, w_011_2871, w_011_2874, w_011_2875, w_011_2876, w_011_2877, w_011_2879, w_011_2881, w_011_2882, w_011_2883, w_011_2884, w_011_2885, w_011_2887, w_011_2888, w_011_2890, w_011_2893, w_011_2894, w_011_2895, w_011_2896, w_011_2898, w_011_2899, w_011_2900, w_011_2901, w_011_2902, w_011_2903, w_011_2904, w_011_2905, w_011_2907, w_011_2909, w_011_2911, w_011_2912, w_011_2913, w_011_2914, w_011_2915, w_011_2916, w_011_2917, w_011_2918, w_011_2919, w_011_2920, w_011_2921, w_011_2922, w_011_2923, w_011_2924, w_011_2928, w_011_2930, w_011_2933, w_011_2934, w_011_2935, w_011_2936, w_011_2937, w_011_2938, w_011_2941, w_011_2942, w_011_2943, w_011_2944, w_011_2945, w_011_2949, w_011_2950, w_011_2951, w_011_2952, w_011_2955, w_011_2956, w_011_2960, w_011_2961, w_011_2963, w_011_2964, w_011_2965, w_011_2968, w_011_2969, w_011_2970, w_011_2972, w_011_2973, w_011_2974, w_011_2976, w_011_2977, w_011_2980, w_011_2981, w_011_2983, w_011_2984, w_011_2987, w_011_2989, w_011_2990, w_011_2991, w_011_2992, w_011_2993, w_011_2994, w_011_2995, w_011_2996, w_011_2998, w_011_2999, w_011_3001, w_011_3003, w_011_3005, w_011_3006, w_011_3007, w_011_3009, w_011_3010, w_011_3013, w_011_3015, w_011_3016, w_011_3017, w_011_3018, w_011_3019, w_011_3020, w_011_3021, w_011_3022, w_011_3023, w_011_3024, w_011_3025, w_011_3026, w_011_3027, w_011_3032, w_011_3033, w_011_3034, w_011_3035, w_011_3037, w_011_3039, w_011_3040, w_011_3041, w_011_3044, w_011_3045, w_011_3048, w_011_3049, w_011_3051, w_011_3052, w_011_3053, w_011_3055, w_011_3059, w_011_3060, w_011_3062, w_011_3063, w_011_3064, w_011_3065, w_011_3067, w_011_3068, w_011_3070, w_011_3072, w_011_3073, w_011_3075, w_011_3076, w_011_3077, w_011_3078, w_011_3080, w_011_3081, w_011_3082, w_011_3084, w_011_3086, w_011_3087, w_011_3090, w_011_3091, w_011_3092, w_011_3093, w_011_3095, w_011_3097, w_011_3098, w_011_3099, w_011_3101, w_011_3102, w_011_3105, w_011_3106, w_011_3107, w_011_3108, w_011_3109, w_011_3110, w_011_3111, w_011_3113, w_011_3115, w_011_3116, w_011_3118, w_011_3119, w_011_3120, w_011_3121, w_011_3122, w_011_3124, w_011_3126, w_011_3127, w_011_3128, w_011_3129, w_011_3130, w_011_3131, w_011_3132, w_011_3135, w_011_3136, w_011_3137, w_011_3138, w_011_3139, w_011_3140, w_011_3141, w_011_3142, w_011_3143, w_011_3144, w_011_3145, w_011_3146, w_011_3147, w_011_3148, w_011_3149, w_011_3151, w_011_3152, w_011_3154, w_011_3156, w_011_3158, w_011_3159, w_011_3160, w_011_3161, w_011_3164, w_011_3168, w_011_3169, w_011_3171, w_011_3172, w_011_3173, w_011_3174, w_011_3178, w_011_3179, w_011_3180, w_011_3181, w_011_3183, w_011_3184, w_011_3185, w_011_3186, w_011_3188, w_011_3189, w_011_3190, w_011_3191, w_011_3194, w_011_3195, w_011_3196, w_011_3197, w_011_3198, w_011_3199, w_011_3200, w_011_3206, w_011_3207, w_011_3208, w_011_3209, w_011_3210, w_011_3211, w_011_3212, w_011_3213, w_011_3214, w_011_3216, w_011_3217, w_011_3218, w_011_3219, w_011_3220, w_011_3221, w_011_3223, w_011_3225, w_011_3226, w_011_3227, w_011_3228, w_011_3230, w_011_3231, w_011_3232, w_011_3234, w_011_3235, w_011_3238, w_011_3239, w_011_3240, w_011_3241, w_011_3246, w_011_3247, w_011_3248, w_011_3250, w_011_3251, w_011_3253, w_011_3254, w_011_3255, w_011_3257, w_011_3258, w_011_3261, w_011_3264, w_011_3267, w_011_3269, w_011_3271, w_011_3272, w_011_3273, w_011_3274, w_011_3275, w_011_3276, w_011_3277, w_011_3279, w_011_3280, w_011_3281, w_011_3282, w_011_3284, w_011_3286, w_011_3287, w_011_3289, w_011_3290, w_011_3291, w_011_3292, w_011_3293, w_011_3294, w_011_3295, w_011_3296, w_011_3297, w_011_3298, w_011_3299, w_011_3301, w_011_3302, w_011_3303, w_011_3307, w_011_3309, w_011_3311, w_011_3312, w_011_3313, w_011_3317, w_011_3321, w_011_3322, w_011_3323, w_011_3324, w_011_3325, w_011_3328, w_011_3329, w_011_3332, w_011_3334, w_011_3335, w_011_3336, w_011_3337, w_011_3338, w_011_3340, w_011_3341, w_011_3343, w_011_3344, w_011_3345, w_011_3348, w_011_3350, w_011_3352, w_011_3353, w_011_3354, w_011_3355, w_011_3357, w_011_3358, w_011_3360, w_011_3362, w_011_3363, w_011_3364, w_011_3365, w_011_3366, w_011_3367, w_011_3369, w_011_3370, w_011_3371, w_011_3372, w_011_3373, w_011_3375, w_011_3377, w_011_3379, w_011_3380, w_011_3381, w_011_3382, w_011_3384, w_011_3385, w_011_3387, w_011_3388, w_011_3390, w_011_3391, w_011_3392, w_011_3395, w_011_3396, w_011_3397, w_011_3402, w_011_3403, w_011_3404, w_011_3405, w_011_3406, w_011_3407, w_011_3410, w_011_3411, w_011_3412, w_011_3413, w_011_3414, w_011_3415, w_011_3416, w_011_3417, w_011_3418, w_011_3419, w_011_3420, w_011_3422, w_011_3423, w_011_3424, w_011_3426, w_011_3429, w_011_3430, w_011_3431, w_011_3433, w_011_3434, w_011_3435, w_011_3438, w_011_3439, w_011_3440, w_011_3441, w_011_3443, w_011_3444, w_011_3445, w_011_3446, w_011_3447, w_011_3448, w_011_3449, w_011_3450, w_011_3451, w_011_3452, w_011_3453, w_011_3454, w_011_3455, w_011_3456, w_011_3457, w_011_3459, w_011_3460, w_011_3461, w_011_3463, w_011_3465, w_011_3466, w_011_3467, w_011_3468, w_011_3470, w_011_3471, w_011_3473, w_011_3475, w_011_3476, w_011_3477, w_011_3478, w_011_3480, w_011_3481, w_011_3482, w_011_3483, w_011_3485, w_011_3486, w_011_3487, w_011_3488, w_011_3489, w_011_3490, w_011_3492, w_011_3493, w_011_3497, w_011_3498, w_011_3499, w_011_3500, w_011_3501, w_011_3503, w_011_3504, w_011_3505, w_011_3506, w_011_3507, w_011_3509, w_011_3510, w_011_3511, w_011_3513, w_011_3514, w_011_3515, w_011_3516, w_011_3517, w_011_3519, w_011_3520, w_011_3522, w_011_3523, w_011_3524, w_011_3526, w_011_3527, w_011_3529, w_011_3530, w_011_3531, w_011_3532, w_011_3533, w_011_3534, w_011_3535, w_011_3537, w_011_3538, w_011_3540, w_011_3541, w_011_3542, w_011_3543, w_011_3544, w_011_3545, w_011_3546, w_011_3547, w_011_3549, w_011_3550, w_011_3551, w_011_3552, w_011_3553, w_011_3554, w_011_3555, w_011_3556, w_011_3558, w_011_3559, w_011_3561, w_011_3562, w_011_3563, w_011_3564, w_011_3565, w_011_3567, w_011_3569, w_011_3571, w_011_3574, w_011_3577, w_011_3578, w_011_3580, w_011_3581, w_011_3582, w_011_3584, w_011_3585, w_011_3586, w_011_3587, w_011_3588, w_011_3589, w_011_3590, w_011_3591, w_011_3593, w_011_3594, w_011_3595, w_011_3596, w_011_3598, w_011_3599, w_011_3600, w_011_3601, w_011_3604, w_011_3605, w_011_3607, w_011_3609, w_011_3610, w_011_3611, w_011_3612, w_011_3613, w_011_3614, w_011_3615, w_011_3616, w_011_3617, w_011_3618, w_011_3619, w_011_3620, w_011_3622, w_011_3623, w_011_3624, w_011_3625, w_011_3626, w_011_3628, w_011_3629, w_011_3630, w_011_3632, w_011_3636, w_011_3638, w_011_3639, w_011_3641, w_011_3642, w_011_3644, w_011_3645, w_011_3646, w_011_3651, w_011_3652, w_011_3654, w_011_3655, w_011_3656, w_011_3657, w_011_3658, w_011_3660, w_011_3661, w_011_3663, w_011_3665, w_011_3666, w_011_3668, w_011_3670, w_011_3671, w_011_3672, w_011_3673, w_011_3674, w_011_3676, w_011_3677, w_011_3680, w_011_3682, w_011_3683, w_011_3684, w_011_3685, w_011_3686, w_011_3687, w_011_3688, w_011_3690, w_011_3691, w_011_3693, w_011_3695, w_011_3697, w_011_3698, w_011_3699, w_011_3700, w_011_3701, w_011_3702, w_011_3703, w_011_3704, w_011_3705, w_011_3706, w_011_3707, w_011_3709, w_011_3711, w_011_3712, w_011_3714, w_011_3715, w_011_3718, w_011_3719, w_011_3721, w_011_3722, w_011_3723, w_011_3725, w_011_3726, w_011_3727, w_011_3728, w_011_3729, w_011_3730, w_011_3731, w_011_3732, w_011_3733, w_011_3734, w_011_3735, w_011_3736, w_011_3737, w_011_3738, w_011_3739, w_011_3741, w_011_3742, w_011_3743, w_011_3744, w_011_3745, w_011_3746, w_011_3747, w_011_3748, w_011_3749, w_011_3750, w_011_3755, w_011_3756, w_011_3758, w_011_3759, w_011_3760, w_011_3761, w_011_3762, w_011_3763, w_011_3765, w_011_3767, w_011_3768, w_011_3769, w_011_3770, w_011_3771, w_011_3772, w_011_3774, w_011_3775, w_011_3776, w_011_3777, w_011_3779, w_011_3780, w_011_3781, w_011_3783, w_011_3784, w_011_3786, w_011_3787, w_011_3788, w_011_3789, w_011_3791, w_011_3792, w_011_3793, w_011_3794, w_011_3797, w_011_3798, w_011_3799, w_011_3801, w_011_3803, w_011_3804, w_011_3805, w_011_3806, w_011_3807, w_011_3808, w_011_3809, w_011_3810, w_011_3813, w_011_3814, w_011_3815, w_011_3816, w_011_3817, w_011_3818, w_011_3819, w_011_3820, w_011_3821, w_011_3823, w_011_3824, w_011_3825, w_011_3826, w_011_3829, w_011_3830, w_011_3832, w_011_3833, w_011_3834, w_011_3835, w_011_3836, w_011_3838, w_011_3839, w_011_3840, w_011_3842, w_011_3843, w_011_3844, w_011_3845, w_011_3846, w_011_3848, w_011_3849, w_011_3850, w_011_3851, w_011_3852, w_011_3853, w_011_3855, w_011_3857, w_011_3859, w_011_3860, w_011_3861, w_011_3863, w_011_3865, w_011_3867, w_011_3868, w_011_3869, w_011_3870, w_011_3873, w_011_3874, w_011_3875, w_011_3876, w_011_3877, w_011_3879, w_011_3880, w_011_3881, w_011_3882, w_011_3883, w_011_3884, w_011_3886, w_011_3888, w_011_3892, w_011_3894, w_011_3895, w_011_3897, w_011_3899, w_011_3900, w_011_3901, w_011_3902, w_011_3904, w_011_3905, w_011_3906, w_011_3907, w_011_3908, w_011_3909, w_011_3910, w_011_3911, w_011_3914, w_011_3915, w_011_3916, w_011_3917, w_011_3918, w_011_3919, w_011_3920, w_011_3921, w_011_3922, w_011_3923, w_011_3924, w_011_3925, w_011_3926, w_011_3927, w_011_3928, w_011_3929, w_011_3930, w_011_3931, w_011_3933, w_011_3934, w_011_3935, w_011_3936, w_011_3937, w_011_3938, w_011_3940, w_011_3942, w_011_3944, w_011_3945, w_011_3946, w_011_3947, w_011_3950, w_011_3951, w_011_3952, w_011_3953, w_011_3954, w_011_3955, w_011_3956, w_011_3957, w_011_3958, w_011_3959, w_011_3961, w_011_3962, w_011_3965, w_011_3966, w_011_3967, w_011_3968, w_011_3969, w_011_3970, w_011_3971, w_011_3972, w_011_3973, w_011_3977, w_011_3978, w_011_3979, w_011_3981, w_011_3982, w_011_3983, w_011_3984, w_011_3986, w_011_3987, w_011_3988, w_011_3989, w_011_3991, w_011_3992, w_011_3995, w_011_3997, w_011_3999, w_011_4001, w_011_4004, w_011_4008, w_011_4009, w_011_4010, w_011_4011, w_011_4012, w_011_4013, w_011_4014, w_011_4015, w_011_4016, w_011_4018, w_011_4020, w_011_4021, w_011_4022, w_011_4023, w_011_4024, w_011_4025, w_011_4026, w_011_4028, w_011_4031, w_011_4032, w_011_4033, w_011_4034, w_011_4035, w_011_4036, w_011_4037, w_011_4038, w_011_4039, w_011_4040, w_011_4044, w_011_4046, w_011_4047, w_011_4049, w_011_4050, w_011_4052, w_011_4053, w_011_4054, w_011_4056, w_011_4057, w_011_4058, w_011_4060, w_011_4061, w_011_4062, w_011_4063, w_011_4064, w_011_4067, w_011_4068, w_011_4070, w_011_4071, w_011_4074, w_011_4075, w_011_4078, w_011_4081, w_011_4082, w_011_4083, w_011_4084, w_011_4085, w_011_4086, w_011_4087, w_011_4088, w_011_4089, w_011_4091, w_011_4094, w_011_4096, w_011_4097, w_011_4098, w_011_4099, w_011_4100, w_011_4102, w_011_4104, w_011_4105, w_011_4107, w_011_4109, w_011_4111, w_011_4112, w_011_4114, w_011_4117, w_011_4118, w_011_4119, w_011_4120, w_011_4121, w_011_4122, w_011_4123, w_011_4124, w_011_4125, w_011_4126, w_011_4128, w_011_4129, w_011_4130, w_011_4131, w_011_4132, w_011_4133, w_011_4134, w_011_4135, w_011_4141, w_011_4142, w_011_4143, w_011_4145, w_011_4146, w_011_4147, w_011_4148, w_011_4149, w_011_4150, w_011_4151, w_011_4152, w_011_4154, w_011_4155, w_011_4156, w_011_4157, w_011_4159, w_011_4160, w_011_4161, w_011_4162, w_011_4169, w_011_4171, w_011_4173, w_011_4175, w_011_4176, w_011_4177, w_011_4180, w_011_4181, w_011_4182, w_011_4183, w_011_4186, w_011_4187, w_011_4188, w_011_4189, w_011_4191, w_011_4193, w_011_4194, w_011_4195, w_011_4196, w_011_4197, w_011_4198, w_011_4199, w_011_4200, w_011_4201, w_011_4202, w_011_4203, w_011_4206, w_011_4209, w_011_4210, w_011_4211, w_011_4212, w_011_4213, w_011_4215, w_011_4217, w_011_4218, w_011_4219, w_011_4220, w_011_4221, w_011_4222, w_011_4223, w_011_4230, w_011_4231, w_011_4232, w_011_4234, w_011_4237, w_011_4238, w_011_4239, w_011_4240, w_011_4242, w_011_4243, w_011_4245, w_011_4247, w_011_4248, w_011_4249, w_011_4254, w_011_4255, w_011_4257, w_011_4258, w_011_4259, w_011_4261, w_011_4264, w_011_4265, w_011_4266, w_011_4269, w_011_4271, w_011_4274, w_011_4275, w_011_4276, w_011_4278, w_011_4279, w_011_4281, w_011_4282, w_011_4284, w_011_4285, w_011_4289, w_011_4290, w_011_4291, w_011_4292, w_011_4294, w_011_4295, w_011_4296, w_011_4297, w_011_4298, w_011_4299, w_011_4300, w_011_4301, w_011_4302, w_011_4303, w_011_4304, w_011_4306, w_011_4308, w_011_4309, w_011_4310, w_011_4311, w_011_4314, w_011_4315, w_011_4317, w_011_4318, w_011_4319, w_011_4320, w_011_4322, w_011_4323, w_011_4324, w_011_4326, w_011_4327, w_011_4328, w_011_4329, w_011_4331, w_011_4334, w_011_4335, w_011_4336, w_011_4338, w_011_4339, w_011_4340, w_011_4342, w_011_4343, w_011_4344, w_011_4345, w_011_4346, w_011_4348, w_011_4350, w_011_4353, w_011_4354, w_011_4356, w_011_4357, w_011_4358, w_011_4359, w_011_4361, w_011_4362, w_011_4363, w_011_4364, w_011_4365, w_011_4366, w_011_4368, w_011_4369, w_011_4370, w_011_4372, w_011_4374, w_011_4375, w_011_4377, w_011_4379, w_011_4381, w_011_4382, w_011_4383, w_011_4384, w_011_4385, w_011_4386, w_011_4387, w_011_4391, w_011_4392, w_011_4394, w_011_4396, w_011_4397, w_011_4398, w_011_4400, w_011_4402, w_011_4403, w_011_4404, w_011_4405, w_011_4406, w_011_4407, w_011_4408, w_011_4412, w_011_4413, w_011_4414, w_011_4415, w_011_4416, w_011_4417, w_011_4418, w_011_4420, w_011_4421, w_011_4422, w_011_4423, w_011_4424, w_011_4425, w_011_4426, w_011_4427, w_011_4428, w_011_4429, w_011_4430, w_011_4431, w_011_4432, w_011_4433, w_011_4434, w_011_4435, w_011_4437, w_011_4438, w_011_4440, w_011_4441, w_011_4442, w_011_4443, w_011_4444, w_011_4445, w_011_4449, w_011_4452, w_011_4453, w_011_4454, w_011_4455, w_011_4456, w_011_4457, w_011_4458, w_011_4459, w_011_4460, w_011_4461, w_011_4462, w_011_4463, w_011_4464, w_011_4465, w_011_4467, w_011_4469, w_011_4470, w_011_4472, w_011_4473, w_011_4474, w_011_4475, w_011_4476, w_011_4477, w_011_4478, w_011_4479, w_011_4481, w_011_4482, w_011_4483, w_011_4484, w_011_4487, w_011_4489, w_011_4490, w_011_4491, w_011_4492, w_011_4493, w_011_4495, w_011_4496, w_011_4497, w_011_4498, w_011_4499, w_011_4502, w_011_4503, w_011_4505, w_011_4506, w_011_4507, w_011_4508, w_011_4509, w_011_4511, w_011_4512, w_011_4514, w_011_4515, w_011_4517, w_011_4518, w_011_4519, w_011_4520, w_011_4521, w_011_4523, w_011_4524, w_011_4525, w_011_4526, w_011_4527, w_011_4530, w_011_4531, w_011_4532, w_011_4534, w_011_4537, w_011_4538, w_011_4539, w_011_4540, w_011_4542, w_011_4543, w_011_4544, w_011_4545, w_011_4546, w_011_4547, w_011_4548, w_011_4549, w_011_4552, w_011_4554, w_011_4556, w_011_4558, w_011_4560, w_011_4563, w_011_4564, w_011_4565, w_011_4566, w_011_4567, w_011_4570, w_011_4571, w_011_4572, w_011_4573, w_011_4574, w_011_4575, w_011_4577, w_011_4580, w_011_4581, w_011_4582, w_011_4588, w_011_4589, w_011_4590, w_011_4591, w_011_4593, w_011_4594, w_011_4595, w_011_4596, w_011_4597, w_011_4598, w_011_4599, w_011_4603, w_011_4604, w_011_4605, w_011_4606, w_011_4608, w_011_4610, w_011_4611, w_011_4613, w_011_4615, w_011_4616, w_011_4618, w_011_4621, w_011_4622, w_011_4624, w_011_4626, w_011_4627, w_011_4628, w_011_4629, w_011_4631, w_011_4632, w_011_4634, w_011_4636, w_011_4637, w_011_4638, w_011_4639, w_011_4641, w_011_4642, w_011_4643, w_011_4644, w_011_4645, w_011_4646, w_011_4647, w_011_4648, w_011_4649, w_011_4650, w_011_4651, w_011_4653, w_011_4654, w_011_4655, w_011_4657, w_011_4658, w_011_4659, w_011_4660, w_011_4661, w_011_4663, w_011_4664, w_011_4665, w_011_4666, w_011_4668, w_011_4669, w_011_4670, w_011_4671, w_011_4673, w_011_4675, w_011_4676, w_011_4677, w_011_4678, w_011_4679, w_011_4680, w_011_4681, w_011_4682, w_011_4683, w_011_4684, w_011_4685, w_011_4687, w_011_4688, w_011_4689, w_011_4691, w_011_4692, w_011_4694, w_011_4695, w_011_4697, w_011_4698, w_011_4699, w_011_4700, w_011_4701, w_011_4703, w_011_4705, w_011_4710, w_011_4711, w_011_4712, w_011_4713, w_011_4714, w_011_4715, w_011_4716, w_011_4717, w_011_4718, w_011_4719, w_011_4720, w_011_4722, w_011_4723, w_011_4724, w_011_4725, w_011_4726, w_011_4727, w_011_4728, w_011_4729, w_011_4733, w_011_4735, w_011_4736, w_011_4737, w_011_4739, w_011_4740, w_011_4742, w_011_4743, w_011_4744, w_011_4747, w_011_4748, w_011_4749, w_011_4750, w_011_4751, w_011_4752, w_011_4753, w_011_4754, w_011_4755, w_011_4757, w_011_4758, w_011_4759, w_011_4760, w_011_4761, w_011_4763, w_011_4764, w_011_4765, w_011_4766, w_011_4767, w_011_4768, w_011_4772, w_011_4773, w_011_4774, w_011_4775, w_011_4776, w_011_4778, w_011_4779, w_011_4780, w_011_4781, w_011_4784, w_011_4785, w_011_4786, w_011_4787, w_011_4788, w_011_4789, w_011_4790, w_011_4791, w_011_4793, w_011_4794, w_011_4795, w_011_4796, w_011_4797, w_011_4798, w_011_4799, w_011_4801, w_011_4803, w_011_4804, w_011_4805, w_011_4806, w_011_4807, w_011_4810, w_011_4812, w_011_4813, w_011_4814, w_011_4815, w_011_4816, w_011_4817, w_011_4818, w_011_4819, w_011_4820, w_011_4821, w_011_4823, w_011_4824, w_011_4825, w_011_4826, w_011_4827, w_011_4828, w_011_4829, w_011_4832, w_011_4833, w_011_4834, w_011_4837, w_011_4838, w_011_4839, w_011_4840, w_011_4841, w_011_4844, w_011_4845, w_011_4846, w_011_4847, w_011_4848, w_011_4849, w_011_4850, w_011_4851, w_011_4852, w_011_4853, w_011_4854, w_011_4855, w_011_4856, w_011_4859, w_011_4861, w_011_4862, w_011_4864, w_011_4865, w_011_4866, w_011_4867, w_011_4868, w_011_4869, w_011_4870, w_011_4871, w_011_4873, w_011_4874, w_011_4876, w_011_4877, w_011_4878, w_011_4879, w_011_4880, w_011_4881, w_011_4882, w_011_4883, w_011_4884, w_011_4886, w_011_4889, w_011_4890, w_011_4891, w_011_4892, w_011_4893, w_011_4894, w_011_4896, w_011_4897, w_011_4898, w_011_4899, w_011_4900, w_011_4901, w_011_4902, w_011_4904, w_011_4906, w_011_4907, w_011_4908, w_011_4911, w_011_4912, w_011_4915, w_011_4916, w_011_4917, w_011_4918, w_011_4919, w_011_4920, w_011_4921, w_011_4922, w_011_4923, w_011_4924, w_011_4925, w_011_4927, w_011_4928, w_011_4929, w_011_4930, w_011_4931, w_011_4932, w_011_4933, w_011_4935, w_011_4936, w_011_4938, w_011_4939, w_011_4940, w_011_4941, w_011_4944, w_011_4945, w_011_4947, w_011_4949, w_011_4951, w_011_4952, w_011_4954, w_011_4955, w_011_4959, w_011_4960, w_011_4963, w_011_4965, w_011_4966, w_011_4967, w_011_4968, w_011_4969, w_011_4970, w_011_4971, w_011_4974, w_011_4975, w_011_4976, w_011_4977, w_011_4978, w_011_4979, w_011_4980, w_011_4981, w_011_4983, w_011_4984, w_011_4985, w_011_4987, w_011_4989, w_011_4990, w_011_4991, w_011_4993, w_011_4994, w_011_4995, w_011_4996, w_011_4998, w_011_4999, w_011_5001, w_011_5002, w_011_5003, w_011_5004, w_011_5005, w_011_5007, w_011_5008, w_011_5009, w_011_5010, w_011_5012, w_011_5013, w_011_5014, w_011_5015, w_011_5016, w_011_5017, w_011_5019, w_011_5020, w_011_5021, w_011_5022, w_011_5023, w_011_5024, w_011_5025, w_011_5029, w_011_5031, w_011_5032, w_011_5034, w_011_5035, w_011_5036, w_011_5037, w_011_5038, w_011_5039, w_011_5040, w_011_5041, w_011_5042, w_011_5043, w_011_5044, w_011_5046, w_011_5047, w_011_5049, w_011_5050, w_011_5051, w_011_5053, w_011_5054, w_011_5055, w_011_5056, w_011_5057, w_011_5058, w_011_5059, w_011_5060, w_011_5061, w_011_5062, w_011_5063, w_011_5064, w_011_5065, w_011_5066, w_011_5070, w_011_5073, w_011_5074, w_011_5077, w_011_5078, w_011_5080, w_011_5081, w_011_5082, w_011_5083, w_011_5085, w_011_5086, w_011_5087, w_011_5089, w_011_5090, w_011_5091, w_011_5092, w_011_5093, w_011_5094, w_011_5095, w_011_5097, w_011_5100, w_011_5101, w_011_5102, w_011_5103, w_011_5104, w_011_5105, w_011_5106, w_011_5107, w_011_5108, w_011_5109, w_011_5110, w_011_5111, w_011_5112, w_011_5113, w_011_5116, w_011_5117, w_011_5118, w_011_5119, w_011_5121, w_011_5123, w_011_5124, w_011_5127, w_011_5128, w_011_5130, w_011_5131, w_011_5132, w_011_5136, w_011_5138, w_011_5141, w_011_5142, w_011_5143, w_011_5144, w_011_5145, w_011_5146, w_011_5147, w_011_5148, w_011_5150, w_011_5153, w_011_5155, w_011_5156, w_011_5159, w_011_5161, w_011_5162, w_011_5165, w_011_5166, w_011_5168, w_011_5169, w_011_5170, w_011_5172, w_011_5173, w_011_5174, w_011_5176, w_011_5177, w_011_5178, w_011_5179, w_011_5182, w_011_5183, w_011_5184, w_011_5185, w_011_5186, w_011_5187, w_011_5189, w_011_5190, w_011_5191, w_011_5192, w_011_5193, w_011_5194, w_011_5196, w_011_5197, w_011_5198, w_011_5200, w_011_5201, w_011_5202, w_011_5204, w_011_5207, w_011_5208, w_011_5210, w_011_5212, w_011_5213, w_011_5214, w_011_5215, w_011_5216, w_011_5217, w_011_5218, w_011_5219, w_011_5220, w_011_5221, w_011_5223, w_011_5224, w_011_5225, w_011_5226, w_011_5227, w_011_5231, w_011_5232, w_011_5233, w_011_5235, w_011_5236, w_011_5237, w_011_5238, w_011_5239, w_011_5240, w_011_5242, w_011_5243, w_011_5246, w_011_5247, w_011_5248, w_011_5249, w_011_5251, w_011_5252, w_011_5253, w_011_5254, w_011_5255, w_011_5256, w_011_5257, w_011_5259, w_011_5263, w_011_5264, w_011_5265, w_011_5266, w_011_5269, w_011_5271, w_011_5272, w_011_5274, w_011_5276, w_011_5278, w_011_5281, w_011_5282, w_011_5283, w_011_5284, w_011_5285, w_011_5286, w_011_5287, w_011_5288, w_011_5290, w_011_5291, w_011_5292, w_011_5293, w_011_5294, w_011_5295, w_011_5296, w_011_5297, w_011_5298, w_011_5299, w_011_5301, w_011_5302, w_011_5303, w_011_5304, w_011_5305, w_011_5307, w_011_5309, w_011_5310, w_011_5313, w_011_5314, w_011_5315, w_011_5317, w_011_5318, w_011_5322, w_011_5323, w_011_5324, w_011_5326, w_011_5328, w_011_5330, w_011_5331, w_011_5332, w_011_5334, w_011_5335, w_011_5336, w_011_5337, w_011_5338, w_011_5339, w_011_5340, w_011_5342, w_011_5343, w_011_5344, w_011_5345, w_011_5347, w_011_5349, w_011_5351, w_011_5352, w_011_5353, w_011_5354, w_011_5355, w_011_5356, w_011_5357, w_011_5358, w_011_5359, w_011_5360, w_011_5361, w_011_5363, w_011_5365, w_011_5366, w_011_5367, w_011_5368, w_011_5369, w_011_5370, w_011_5374, w_011_5375, w_011_5376, w_011_5379, w_011_5380, w_011_5381, w_011_5382, w_011_5383, w_011_5385, w_011_5386, w_011_5387, w_011_5389, w_011_5391, w_011_5393, w_011_5394, w_011_5396, w_011_5397, w_011_5399, w_011_5400, w_011_5401, w_011_5402, w_011_5404, w_011_5409, w_011_5410, w_011_5411, w_011_5413, w_011_5414, w_011_5416, w_011_5417, w_011_5419, w_011_5420, w_011_5421, w_011_5422, w_011_5423, w_011_5424, w_011_5429, w_011_5430, w_011_5431, w_011_5433, w_011_5434, w_011_5435, w_011_5436, w_011_5437, w_011_5438, w_011_5439, w_011_5440, w_011_5441, w_011_5442, w_011_5443, w_011_5445, w_011_5446, w_011_5447, w_011_5448, w_011_5449, w_011_5451, w_011_5452, w_011_5453, w_011_5454, w_011_5455, w_011_5456, w_011_5457, w_011_5458, w_011_5459, w_011_5460, w_011_5462, w_011_5464, w_011_5465, w_011_5467, w_011_5468, w_011_5469, w_011_5470, w_011_5471, w_011_5472, w_011_5473, w_011_5475, w_011_5476, w_011_5477, w_011_5479, w_011_5480, w_011_5481, w_011_5482, w_011_5484, w_011_5487, w_011_5488, w_011_5489, w_011_5490, w_011_5491, w_011_5494, w_011_5495, w_011_5500, w_011_5502, w_011_5503, w_011_5504, w_011_5506, w_011_5507, w_011_5508, w_011_5509, w_011_5510, w_011_5512, w_011_5513, w_011_5514, w_011_5515, w_011_5516, w_011_5517, w_011_5520, w_011_5522, w_011_5524, w_011_5525, w_011_5526, w_011_5528, w_011_5529, w_011_5530, w_011_5531, w_011_5532, w_011_5533, w_011_5534, w_011_5535, w_011_5537, w_011_5538, w_011_5539, w_011_5540, w_011_5541, w_011_5542, w_011_5544, w_011_5546, w_011_5547, w_011_5550, w_011_5551, w_011_5552, w_011_5553, w_011_5554, w_011_5555, w_011_5558, w_011_5560, w_011_5561, w_011_5563, w_011_5564, w_011_5565, w_011_5566, w_011_5567, w_011_5568, w_011_5569, w_011_5570, w_011_5575, w_011_5576, w_011_5580, w_011_5581, w_011_5584, w_011_5585, w_011_5587, w_011_5589, w_011_5591, w_011_5592, w_011_5593, w_011_5594, w_011_5596, w_011_5599, w_011_5600, w_011_5601, w_011_5602, w_011_5603, w_011_5604, w_011_5605, w_011_5606, w_011_5608, w_011_5609, w_011_5611, w_011_5612, w_011_5616, w_011_5617, w_011_5618, w_011_5619, w_011_5620, w_011_5622, w_011_5623, w_011_5624, w_011_5625, w_011_5626, w_011_5627, w_011_5628, w_011_5630, w_011_5632, w_011_5633, w_011_5634, w_011_5635, w_011_5637, w_011_5638, w_011_5639, w_011_5640, w_011_5642, w_011_5644, w_011_5645, w_011_5646, w_011_5647, w_011_5649, w_011_5650, w_011_5651, w_011_5652, w_011_5655, w_011_5658, w_011_5659, w_011_5660, w_011_5661, w_011_5662, w_011_5663, w_011_5665, w_011_5667, w_011_5668, w_011_5669, w_011_5670, w_011_5671, w_011_5672, w_011_5673, w_011_5674, w_011_5675, w_011_5677, w_011_5679, w_011_5680, w_011_5681, w_011_5682, w_011_5683, w_011_5684, w_011_5685, w_011_5686, w_011_5687, w_011_5688, w_011_5690, w_011_5691, w_011_5692, w_011_5693, w_011_5694, w_011_5695, w_011_5697, w_011_5698, w_011_5699, w_011_5700, w_011_5701, w_011_5702, w_011_5704, w_011_5706, w_011_5707, w_011_5708, w_011_5709, w_011_5710, w_011_5711, w_011_5712, w_011_5713, w_011_5714, w_011_5715, w_011_5716, w_011_5717, w_011_5718, w_011_5719, w_011_5720, w_011_5722, w_011_5724, w_011_5727, w_011_5728, w_011_5730, w_011_5732, w_011_5733, w_011_5737, w_011_5741, w_011_5742, w_011_5743, w_011_5744, w_011_5745, w_011_5747, w_011_5748, w_011_5749, w_011_5750, w_011_5751, w_011_5752, w_011_5753, w_011_5755, w_011_5757, w_011_5758, w_011_5759, w_011_5760, w_011_5761, w_011_5764, w_011_5765, w_011_5767, w_011_5768, w_011_5769, w_011_5771, w_011_5772, w_011_5773, w_011_5774, w_011_5775, w_011_5776, w_011_5777, w_011_5778, w_011_5779, w_011_5780, w_011_5782, w_011_5783, w_011_5784, w_011_5787, w_011_5788, w_011_5789, w_011_5790, w_011_5793, w_011_5794, w_011_5795, w_011_5796, w_011_5797, w_011_5798, w_011_5799, w_011_5800, w_011_5802, w_011_5804, w_011_5805, w_011_5806, w_011_5809, w_011_5810, w_011_5811, w_011_5812, w_011_5813, w_011_5814, w_011_5815, w_011_5816, w_011_5817, w_011_5818, w_011_5819, w_011_5820, w_011_5821, w_011_5822, w_011_5823, w_011_5825, w_011_5826, w_011_5828, w_011_5829, w_011_5830, w_011_5831, w_011_5832, w_011_5833, w_011_5835, w_011_5836, w_011_5837, w_011_5840, w_011_5845, w_011_5846, w_011_5847, w_011_5848, w_011_5849, w_011_5850, w_011_5851, w_011_5852, w_011_5853, w_011_5854, w_011_5855, w_011_5857, w_011_5858, w_011_5859, w_011_5860, w_011_5861, w_011_5862, w_011_5864, w_011_5865, w_011_5866, w_011_5867, w_011_5868, w_011_5870, w_011_5871, w_011_5873, w_011_5875, w_011_5876, w_011_5877, w_011_5878, w_011_5879, w_011_5881, w_011_5882, w_011_5883, w_011_5884, w_011_5885, w_011_5888, w_011_5890, w_011_5891, w_011_5893, w_011_5894, w_011_5896, w_011_5900, w_011_5901, w_011_5902, w_011_5903, w_011_5904, w_011_5906, w_011_5907, w_011_5908, w_011_5909, w_011_5911, w_011_5912, w_011_5913, w_011_5915, w_011_5916, w_011_5919, w_011_5921, w_011_5924, w_011_5925, w_011_5926, w_011_5927, w_011_5929, w_011_5930, w_011_5933, w_011_5934, w_011_5935, w_011_5936, w_011_5937, w_011_5938, w_011_5941, w_011_5942, w_011_5943, w_011_5944, w_011_5945, w_011_5946, w_011_5947, w_011_5948, w_011_5949, w_011_5950, w_011_5952, w_011_5955, w_011_5956, w_011_5957, w_011_5958, w_011_5959, w_011_5960, w_011_5961, w_011_5962, w_011_5963, w_011_5964, w_011_5965, w_011_5967, w_011_5969, w_011_5970, w_011_5972, w_011_5973, w_011_5974, w_011_5975, w_011_5976, w_011_5980, w_011_5981, w_011_5983, w_011_5985, w_011_5986, w_011_5987, w_011_5988, w_011_5990, w_011_5991, w_011_5992, w_011_5993, w_011_5994, w_011_5995, w_011_5996, w_011_5997, w_011_5998, w_011_5999, w_011_6000, w_011_6001, w_011_6002, w_011_6005, w_011_6007, w_011_6008, w_011_6011, w_011_6012, w_011_6013, w_011_6014, w_011_6016, w_011_6017, w_011_6019, w_011_6021, w_011_6022, w_011_6023, w_011_6024, w_011_6025, w_011_6029, w_011_6030, w_011_6032, w_011_6033, w_011_6034, w_011_6035, w_011_6036, w_011_6038, w_011_6039, w_011_6040, w_011_6041, w_011_6042, w_011_6044, w_011_6045, w_011_6046, w_011_6047, w_011_6048, w_011_6050, w_011_6051, w_011_6053, w_011_6054, w_011_6055, w_011_6056, w_011_6057, w_011_6060, w_011_6061, w_011_6062, w_011_6067, w_011_6069, w_011_6070, w_011_6071, w_011_6072, w_011_6073, w_011_6074, w_011_6075, w_011_6076, w_011_6077, w_011_6078, w_011_6079, w_011_6080, w_011_6081, w_011_6082, w_011_6083, w_011_6084, w_011_6085, w_011_6086, w_011_6087, w_011_6089, w_011_6090, w_011_6092, w_011_6095, w_011_6097, w_011_6098, w_011_6100, w_011_6101, w_011_6103, w_011_6104, w_011_6105, w_011_6106, w_011_6108, w_011_6110, w_011_6111, w_011_6112, w_011_6116, w_011_6117, w_011_6118, w_011_6120, w_011_6122, w_011_6123, w_011_6124, w_011_6125, w_011_6126, w_011_6132, w_011_6133, w_011_6134, w_011_6135, w_011_6136, w_011_6137, w_011_6138, w_011_6139, w_011_6140, w_011_6141, w_011_6142, w_011_6143, w_011_6145, w_011_6146, w_011_6147, w_011_6148, w_011_6149, w_011_6151, w_011_6153, w_011_6157, w_011_6159, w_011_6161, w_011_6162, w_011_6163, w_011_6164, w_011_6165, w_011_6166, w_011_6167, w_011_6168, w_011_6169, w_011_6170, w_011_6171, w_011_6172, w_011_6173, w_011_6174, w_011_6175, w_011_6176, w_011_6178, w_011_6179, w_011_6181, w_011_6182, w_011_6183, w_011_6185, w_011_6187, w_011_6189, w_011_6190, w_011_6191, w_011_6192, w_011_6194, w_011_6197, w_011_6198, w_011_6199, w_011_6200, w_011_6201, w_011_6203, w_011_6205, w_011_6206, w_011_6208, w_011_6210, w_011_6211, w_011_6212, w_011_6214, w_011_6215, w_011_6216, w_011_6217, w_011_6218, w_011_6219, w_011_6220, w_011_6221, w_011_6223, w_011_6224, w_011_6225, w_011_6227, w_011_6228, w_011_6229, w_011_6230, w_011_6231, w_011_6232, w_011_6233, w_011_6234, w_011_6235, w_011_6238, w_011_6239, w_011_6240, w_011_6241, w_011_6243, w_011_6244, w_011_6245, w_011_6246, w_011_6247, w_011_6249, w_011_6250, w_011_6252, w_011_6253, w_011_6254, w_011_6255, w_011_6256, w_011_6257, w_011_6258, w_011_6260, w_011_6261, w_011_6262, w_011_6263, w_011_6264, w_011_6265, w_011_6266, w_011_6268, w_011_6270, w_011_6272, w_011_6273, w_011_6274, w_011_6275, w_011_6276, w_011_6278, w_011_6279, w_011_6280, w_011_6282, w_011_6283, w_011_6285, w_011_6288, w_011_6289, w_011_6290, w_011_6291, w_011_6294, w_011_6296, w_011_6297, w_011_6298, w_011_6299, w_011_6300, w_011_6302, w_011_6303, w_011_6304, w_011_6305, w_011_6308, w_011_6309, w_011_6310, w_011_6311, w_011_6312, w_011_6313, w_011_6317, w_011_6318, w_011_6320, w_011_6321, w_011_6322, w_011_6323, w_011_6324, w_011_6325, w_011_6326, w_011_6327, w_011_6328, w_011_6329, w_011_6330, w_011_6331, w_011_6332, w_011_6334, w_011_6336, w_011_6337, w_011_6338, w_011_6340, w_011_6341, w_011_6342, w_011_6343, w_011_6344, w_011_6346, w_011_6348, w_011_6349, w_011_6350, w_011_6351, w_011_6352, w_011_6353, w_011_6354, w_011_6355, w_011_6356, w_011_6357, w_011_6358, w_011_6361, w_011_6363, w_011_6365, w_011_6366, w_011_6373, w_011_6375, w_011_6376, w_011_6377, w_011_6380, w_011_6381, w_011_6382, w_011_6383, w_011_6384, w_011_6385, w_011_6386, w_011_6387, w_011_6389, w_011_6390, w_011_6392, w_011_6394, w_011_6395, w_011_6397, w_011_6398, w_011_6401, w_011_6403, w_011_6404, w_011_6405, w_011_6406, w_011_6407, w_011_6408, w_011_6409, w_011_6410, w_011_6414, w_011_6415, w_011_6416, w_011_6417, w_011_6418, w_011_6419, w_011_6422, w_011_6423, w_011_6424, w_011_6425, w_011_6427, w_011_6428, w_011_6431, w_011_6432, w_011_6434, w_011_6438, w_011_6439, w_011_6440, w_011_6441, w_011_6444, w_011_6445, w_011_6446, w_011_6447, w_011_6448, w_011_6449, w_011_6451, w_011_6453, w_011_6454, w_011_6455, w_011_6456, w_011_6458, w_011_6459, w_011_6460, w_011_6461, w_011_6462, w_011_6463, w_011_6464, w_011_6465, w_011_6466, w_011_6467, w_011_6468, w_011_6469, w_011_6470, w_011_6471, w_011_6472, w_011_6474, w_011_6475, w_011_6476, w_011_6478, w_011_6479, w_011_6481, w_011_6482, w_011_6483, w_011_6484, w_011_6486, w_011_6487, w_011_6488, w_011_6489, w_011_6491, w_011_6492, w_011_6493, w_011_6494, w_011_6495, w_011_6496, w_011_6497, w_011_6499, w_011_6501, w_011_6502, w_011_6504, w_011_6505, w_011_6506, w_011_6507, w_011_6508, w_011_6509, w_011_6510, w_011_6511, w_011_6512, w_011_6513, w_011_6514, w_011_6515, w_011_6519, w_011_6522, w_011_6523, w_011_6524, w_011_6525, w_011_6526, w_011_6527, w_011_6528, w_011_6529, w_011_6531, w_011_6532, w_011_6533, w_011_6539, w_011_6540, w_011_6541, w_011_6542, w_011_6543, w_011_6544, w_011_6545, w_011_6546, w_011_6547, w_011_6548, w_011_6550, w_011_6552, w_011_6554, w_011_6555, w_011_6556, w_011_6557, w_011_6558, w_011_6561, w_011_6562, w_011_6563, w_011_6564, w_011_6565, w_011_6567, w_011_6568, w_011_6569, w_011_6570, w_011_6571, w_011_6573, w_011_6576, w_011_6577, w_011_6578, w_011_6579, w_011_6582, w_011_6583, w_011_6584, w_011_6585, w_011_6586, w_011_6587, w_011_6588, w_011_6590, w_011_6591, w_011_6592, w_011_6593, w_011_6594, w_011_6595, w_011_6598, w_011_6599, w_011_6600, w_011_6604, w_011_6605, w_011_6606, w_011_6607, w_011_6609, w_011_6610, w_011_6611, w_011_6612, w_011_6613, w_011_6616, w_011_6617, w_011_6618, w_011_6619, w_011_6620, w_011_6622, w_011_6623, w_011_6625, w_011_6626, w_011_6627, w_011_6628, w_011_6629, w_011_6630, w_011_6631, w_011_6632, w_011_6633, w_011_6635, w_011_6636, w_011_6637, w_011_6638, w_011_6639, w_011_6640, w_011_6641, w_011_6644, w_011_6645, w_011_6647, w_011_6648, w_011_6649, w_011_6650, w_011_6651, w_011_6652, w_011_6656, w_011_6657, w_011_6658, w_011_6661, w_011_6664, w_011_6665, w_011_6666, w_011_6667, w_011_6669, w_011_6670, w_011_6671, w_011_6673, w_011_6674, w_011_6675, w_011_6676, w_011_6677, w_011_6678, w_011_6679, w_011_6680, w_011_6682, w_011_6683, w_011_6684, w_011_6685, w_011_6687, w_011_6690, w_011_6692, w_011_6693, w_011_6694, w_011_6695, w_011_6697, w_011_6698, w_011_6699, w_011_6701, w_011_6702, w_011_6703, w_011_6704, w_011_6705, w_011_6707, w_011_6708, w_011_6709, w_011_6710, w_011_6712, w_011_6714, w_011_6715, w_011_6716, w_011_6718, w_011_6719, w_011_6720, w_011_6721, w_011_6722, w_011_6723, w_011_6724, w_011_6725, w_011_6726, w_011_6727, w_011_6728, w_011_6730, w_011_6731, w_011_6735, w_011_6736, w_011_6737, w_011_6738, w_011_6739, w_011_6740, w_011_6741, w_011_6742, w_011_6743, w_011_6744, w_011_6745, w_011_6747, w_011_6748, w_011_6749, w_011_6750, w_011_6751, w_011_6752, w_011_6753, w_011_6754, w_011_6755, w_011_6756, w_011_6758, w_011_6759, w_011_6760, w_011_6762, w_011_6764, w_011_6765, w_011_6767, w_011_6768, w_011_6769, w_011_6771, w_011_6772, w_011_6773, w_011_6774, w_011_6775, w_011_6776, w_011_6777, w_011_6779, w_011_6780, w_011_6782, w_011_6784, w_011_6789, w_011_6790, w_011_6792, w_011_6793, w_011_6795, w_011_6796, w_011_6797, w_011_6798, w_011_6799, w_011_6800, w_011_6801, w_011_6805, w_011_6807, w_011_6808, w_011_6809, w_011_6810, w_011_6811, w_011_6814, w_011_6815, w_011_6816, w_011_6817, w_011_6818, w_011_6819, w_011_6820, w_011_6821, w_011_6822, w_011_6823, w_011_6824, w_011_6825, w_011_6826, w_011_6827, w_011_6828, w_011_6830, w_011_6831, w_011_6832, w_011_6833, w_011_6834, w_011_6838, w_011_6839, w_011_6840, w_011_6843, w_011_6844, w_011_6846, w_011_6847, w_011_6848, w_011_6851, w_011_6853, w_011_6854, w_011_6855, w_011_6857, w_011_6858, w_011_6859, w_011_6862, w_011_6863, w_011_6864, w_011_6865, w_011_6866, w_011_6867, w_011_6868, w_011_6869, w_011_6870, w_011_6872, w_011_6875, w_011_6876, w_011_6877, w_011_6878, w_011_6879, w_011_6880, w_011_6881, w_011_6882, w_011_6884, w_011_6885, w_011_6886, w_011_6887, w_011_6888, w_011_6890, w_011_6891, w_011_6893, w_011_6894, w_011_6895, w_011_6898, w_011_6899, w_011_6901, w_011_6902, w_011_6903, w_011_6904, w_011_6906, w_011_6908, w_011_6911, w_011_6912, w_011_6914, w_011_6915, w_011_6916, w_011_6917, w_011_6918, w_011_6920, w_011_6921, w_011_6922, w_011_6923, w_011_6924, w_011_6925, w_011_6927, w_011_6929, w_011_6930, w_011_6931, w_011_6932, w_011_6933, w_011_6934, w_011_6935, w_011_6936, w_011_6937, w_011_6938, w_011_6939, w_011_6941, w_011_6943, w_011_6944, w_011_6945, w_011_6946, w_011_6947, w_011_6948, w_011_6949, w_011_6950, w_011_6952, w_011_6953, w_011_6954, w_011_6955, w_011_6956, w_011_6957, w_011_6958, w_011_6959, w_011_6960, w_011_6961, w_011_6962, w_011_6963, w_011_6964, w_011_6965, w_011_6966, w_011_6967, w_011_6969, w_011_6971, w_011_6972, w_011_6973, w_011_6974, w_011_6975, w_011_6977, w_011_6979, w_011_6980, w_011_6982, w_011_6983, w_011_6984, w_011_6986, w_011_6987, w_011_6988, w_011_6990, w_011_6991, w_011_6992, w_011_6994, w_011_6995, w_011_6996, w_011_6998, w_011_6999, w_011_7000, w_011_7001, w_011_7002, w_011_7003, w_011_7004, w_011_7006, w_011_7007, w_011_7009, w_011_7011, w_011_7013, w_011_7015, w_011_7017, w_011_7018, w_011_7019, w_011_7020, w_011_7021, w_011_7022, w_011_7023, w_011_7024, w_011_7025, w_011_7026, w_011_7027, w_011_7028, w_011_7029, w_011_7030, w_011_7031, w_011_7032, w_011_7033, w_011_7035, w_011_7037, w_011_7038, w_011_7039, w_011_7040, w_011_7041, w_011_7042, w_011_7043, w_011_7044, w_011_7046, w_011_7047, w_011_7048, w_011_7049, w_011_7050, w_011_7051, w_011_7052, w_011_7053, w_011_7054, w_011_7055, w_011_7058, w_011_7059, w_011_7060, w_011_7061, w_011_7062, w_011_7063, w_011_7064, w_011_7066, w_011_7069, w_011_7070, w_011_7072, w_011_7074, w_011_7075, w_011_7080, w_011_7081, w_011_7082, w_011_7083, w_011_7084, w_011_7085, w_011_7086, w_011_7087, w_011_7088, w_011_7089, w_011_7090, w_011_7091, w_011_7092, w_011_7093, w_011_7094, w_011_7095, w_011_7098, w_011_7101, w_011_7103, w_011_7104, w_011_7106, w_011_7107, w_011_7108, w_011_7109, w_011_7110, w_011_7111, w_011_7112, w_011_7113, w_011_7114, w_011_7115, w_011_7116, w_011_7117, w_011_7118, w_011_7119, w_011_7121, w_011_7122, w_011_7123, w_011_7124, w_011_7125, w_011_7126, w_011_7127, w_011_7129, w_011_7131, w_011_7132, w_011_7133, w_011_7134, w_011_7137, w_011_7138, w_011_7139, w_011_7142, w_011_7143, w_011_7144, w_011_7146, w_011_7148, w_011_7149, w_011_7150, w_011_7151, w_011_7152, w_011_7153, w_011_7154, w_011_7155, w_011_7156, w_011_7157, w_011_7159, w_011_7160, w_011_7162, w_011_7164, w_011_7165, w_011_7166, w_011_7172, w_011_7173, w_011_7174, w_011_7175, w_011_7176, w_011_7179, w_011_7180, w_011_7181, w_011_7182, w_011_7183, w_011_7184, w_011_7186, w_011_7187, w_011_7188, w_011_7191, w_011_7194, w_011_7196, w_011_7198, w_011_7199, w_011_7201, w_011_7202, w_011_7203, w_011_7206, w_011_7208, w_011_7209, w_011_7211, w_011_7213, w_011_7216, w_011_7217, w_011_7218, w_011_7219, w_011_7220, w_011_7221, w_011_7222, w_011_7223, w_011_7224, w_011_7225, w_011_7226, w_011_7228, w_011_7229, w_011_7230, w_011_7231, w_011_7232, w_011_7234, w_011_7235, w_011_7236, w_011_7238, w_011_7242, w_011_7243, w_011_7244, w_011_7245, w_011_7246, w_011_7247, w_011_7249, w_011_7250, w_011_7251, w_011_7252, w_011_7253, w_011_7254, w_011_7255, w_011_7256, w_011_7257, w_011_7258, w_011_7259, w_011_7261, w_011_7262, w_011_7263, w_011_7264, w_011_7265, w_011_7266, w_011_7268, w_011_7270, w_011_7271, w_011_7272, w_011_7274, w_011_7275, w_011_7277, w_011_7278, w_011_7279, w_011_7280, w_011_7281, w_011_7284, w_011_7286, w_011_7288, w_011_7289, w_011_7290, w_011_7291, w_011_7292, w_011_7293, w_011_7294, w_011_7295, w_011_7297, w_011_7298, w_011_7299, w_011_7300, w_011_7301, w_011_7305, w_011_7306, w_011_7307, w_011_7308, w_011_7309, w_011_7311, w_011_7312, w_011_7313, w_011_7314, w_011_7315, w_011_7316, w_011_7318, w_011_7319, w_011_7321, w_011_7322, w_011_7323, w_011_7324, w_011_7329, w_011_7330, w_011_7331, w_011_7332, w_011_7333, w_011_7334, w_011_7335, w_011_7336, w_011_7337, w_011_7338, w_011_7339, w_011_7342, w_011_7344, w_011_7345, w_011_7346, w_011_7347, w_011_7348, w_011_7349, w_011_7350, w_011_7351, w_011_7352, w_011_7354, w_011_7355, w_011_7357, w_011_7358, w_011_7360, w_011_7361, w_011_7362, w_011_7363, w_011_7366, w_011_7367, w_011_7368, w_011_7369, w_011_7373, w_011_7374, w_011_7376, w_011_7378, w_011_7379, w_011_7380, w_011_7383, w_011_7384, w_011_7385, w_011_7389, w_011_7390, w_011_7391, w_011_7392, w_011_7393, w_011_7395, w_011_7397, w_011_7398, w_011_7401, w_011_7406, w_011_7407, w_011_7411, w_011_7412, w_011_7416, w_011_7417, w_011_7418, w_011_7420, w_011_7421, w_011_7423, w_011_7424, w_011_7425, w_011_7426, w_011_7427, w_011_7428, w_011_7429, w_011_7431, w_011_7432, w_011_7433, w_011_7435, w_011_7436, w_011_7437, w_011_7438, w_011_7440, w_011_7441, w_011_7443, w_011_7444, w_011_7447, w_011_7454, w_011_7456, w_011_7457, w_011_7459, w_011_7461, w_011_7462, w_011_7470, w_011_7471, w_011_7472, w_011_7473, w_011_7475, w_011_7477, w_011_7478, w_011_7479, w_011_7480, w_011_7481, w_011_7482, w_011_7483, w_011_7485, w_011_7486, w_011_7487, w_011_7488, w_011_7489, w_011_7490, w_011_7495, w_011_7496, w_011_7497, w_011_7498, w_011_7499, w_011_7500, w_011_7501, w_011_7503, w_011_7504, w_011_7506, w_011_7507, w_011_7509, w_011_7510, w_011_7511, w_011_7512, w_011_7513, w_011_7515, w_011_7517, w_011_7519, w_011_7520, w_011_7521, w_011_7522, w_011_7523, w_011_7524, w_011_7525, w_011_7526, w_011_7527, w_011_7528, w_011_7529, w_011_7530, w_011_7531, w_011_7532, w_011_7533, w_011_7534, w_011_7536, w_011_7537, w_011_7539, w_011_7541, w_011_7542, w_011_7543, w_011_7544, w_011_7545, w_011_7548, w_011_7549, w_011_7551, w_011_7552, w_011_7553, w_011_7554, w_011_7556, w_011_7557, w_011_7558, w_011_7559, w_011_7560, w_011_7563, w_011_7565, w_011_7566, w_011_7567, w_011_7568, w_011_7571, w_011_7573, w_011_7574, w_011_7576, w_011_7578, w_011_7580, w_011_7583, w_011_7584, w_011_7585, w_011_7588, w_011_7589, w_011_7590, w_011_7594, w_011_7595, w_011_7596, w_011_7597, w_011_7598, w_011_7599, w_011_7601, w_011_7602, w_011_7603, w_011_7604, w_011_7605, w_011_7606, w_011_7608, w_011_7609, w_011_7610, w_011_7611, w_011_7612, w_011_7614, w_011_7615, w_011_7616, w_011_7617, w_011_7619, w_011_7620, w_011_7621, w_011_7623, w_011_7624, w_011_7626, w_011_7629, w_011_7630, w_011_7632, w_011_7633, w_011_7635, w_011_7636, w_011_7638, w_011_7639, w_011_7641, w_011_7642, w_011_7646, w_011_7647, w_011_7652, w_011_7653, w_011_7654, w_011_7655, w_011_7656, w_011_7657, w_011_7659, w_011_7660, w_011_7661, w_011_7663, w_011_7664, w_011_7665, w_011_7666, w_011_7667, w_011_7668, w_011_7669, w_011_7671, w_011_7672, w_011_7674, w_011_7675, w_011_7676, w_011_7677, w_011_7678, w_011_7679, w_011_7680, w_011_7681, w_011_7682, w_011_7683, w_011_7684, w_011_7685, w_011_7688, w_011_7689, w_011_7692, w_011_7693, w_011_7694, w_011_7695, w_011_7696, w_011_7698, w_011_7699, w_011_7700, w_011_7702, w_011_7703, w_011_7704, w_011_7705, w_011_7706, w_011_7707, w_011_7708, w_011_7709, w_011_7711, w_011_7714, w_011_7715, w_011_7716, w_011_7717, w_011_7718, w_011_7720, w_011_7721, w_011_7722, w_011_7723, w_011_7724, w_011_7725, w_011_7726, w_011_7727, w_011_7729, w_011_7730, w_011_7731, w_011_7732, w_011_7733, w_011_7736, w_011_7737, w_011_7738, w_011_7739, w_011_7741, w_011_7743, w_011_7744, w_011_7746, w_011_7747, w_011_7748, w_011_7749, w_011_7750, w_011_7751, w_011_7752, w_011_7753, w_011_7755, w_011_7756, w_011_7758, w_011_7759, w_011_7762, w_011_7766, w_011_7767, w_011_7768, w_011_7770, w_011_7771, w_011_7773, w_011_7774, w_011_7775, w_011_7777, w_011_7778, w_011_7779, w_011_7780, w_011_7781, w_011_7782, w_011_7783, w_011_7784, w_011_7786, w_011_7787, w_011_7788, w_011_7789, w_011_7790, w_011_7792, w_011_7793, w_011_7794, w_011_7796, w_011_7799, w_011_7800, w_011_7802, w_011_7805, w_011_7806, w_011_7807, w_011_7809, w_011_7813, w_011_7815, w_011_7816, w_011_7817, w_011_7819, w_011_7821, w_011_7823, w_011_7824, w_011_7825, w_011_7826, w_011_7827, w_011_7831, w_011_7833, w_011_7834, w_011_7835, w_011_7837, w_011_7838, w_011_7839, w_011_7840, w_011_7841, w_011_7842, w_011_7843, w_011_7845, w_011_7847, w_011_7848, w_011_7849, w_011_7850, w_011_7851, w_011_7852, w_011_7853, w_011_7854, w_011_7855, w_011_7857, w_011_7858, w_011_7859, w_011_7860, w_011_7861, w_011_7862, w_011_7863, w_011_7865, w_011_7867, w_011_7868, w_011_7869, w_011_7870, w_011_7871, w_011_7872, w_011_7873, w_011_7874, w_011_7875, w_011_7876, w_011_7877, w_011_7882, w_011_7883, w_011_7885, w_011_7886, w_011_7887, w_011_7888, w_011_7889, w_011_7890, w_011_7892, w_011_7893, w_011_7894, w_011_7895, w_011_7896, w_011_7898, w_011_7899, w_011_7900, w_011_7901, w_011_7903, w_011_7904, w_011_7908, w_011_7909, w_011_7910, w_011_7912, w_011_7913, w_011_7914, w_011_7915, w_011_7917, w_011_7918, w_011_7919, w_011_7920, w_011_7921, w_011_7922, w_011_7923, w_011_7924, w_011_7925, w_011_7926, w_011_7927, w_011_7928, w_011_7929, w_011_7930, w_011_7933, w_011_7934, w_011_7935, w_011_7939, w_011_7940, w_011_7941, w_011_7942, w_011_7943, w_011_7944, w_011_7945, w_011_7947, w_011_7948, w_011_7949, w_011_7950, w_011_7951, w_011_7952, w_011_7955, w_011_7956, w_011_7957, w_011_7958, w_011_7959, w_011_7961, w_011_7962, w_011_7963, w_011_7964, w_011_7967, w_011_7968, w_011_7969, w_011_7970, w_011_7972, w_011_7973, w_011_7974, w_011_7975, w_011_7976, w_011_7978, w_011_7979, w_011_7980, w_011_7984, w_011_7985, w_011_7986, w_011_7987, w_011_7988, w_011_7989, w_011_7991, w_011_7992, w_011_7993, w_011_7994, w_011_7995, w_011_7996, w_011_7998, w_011_7999, w_011_8000, w_011_8002, w_011_8003, w_011_8004, w_011_8005, w_011_8007, w_011_8009, w_011_8010, w_011_8011, w_011_8012, w_011_8013, w_011_8015, w_011_8016, w_011_8017, w_011_8018, w_011_8019, w_011_8020, w_011_8021, w_011_8022, w_011_8023, w_011_8024, w_011_8025, w_011_8027, w_011_8029, w_011_8032, w_011_8035, w_011_8036, w_011_8038, w_011_8039, w_011_8040, w_011_8041, w_011_8043, w_011_8044, w_011_8045, w_011_8046, w_011_8047, w_011_8048, w_011_8049, w_011_8050, w_011_8052, w_011_8053, w_011_8054, w_011_8055, w_011_8058, w_011_8061, w_011_8062, w_011_8063, w_011_8065, w_011_8067, w_011_8068, w_011_8069, w_011_8071, w_011_8072, w_011_8073, w_011_8074, w_011_8075, w_011_8080, w_011_8081, w_011_8082, w_011_8083, w_011_8085, w_011_8087, w_011_8089, w_011_8091, w_011_8092, w_011_8093, w_011_8094, w_011_8095, w_011_8098, w_011_8100, w_011_8101, w_011_8103, w_011_8104, w_011_8105, w_011_8106, w_011_8107, w_011_8109, w_011_8110, w_011_8111, w_011_8112, w_011_8115, w_011_8117, w_011_8118, w_011_8120, w_011_8122, w_011_8123, w_011_8124, w_011_8125, w_011_8126, w_011_8127, w_011_8128, w_011_8129, w_011_8130, w_011_8131, w_011_8134, w_011_8135, w_011_8136, w_011_8137, w_011_8138, w_011_8141, w_011_8144, w_011_8145, w_011_8146, w_011_8147, w_011_8148, w_011_8149, w_011_8150, w_011_8151, w_011_8152, w_011_8154, w_011_8155, w_011_8156, w_011_8157, w_011_8158, w_011_8159, w_011_8160, w_011_8161, w_011_8162, w_011_8163, w_011_8164, w_011_8165, w_011_8166, w_011_8167, w_011_8168, w_011_8169, w_011_8170, w_011_8173, w_011_8174, w_011_8176, w_011_8177, w_011_8178, w_011_8179, w_011_8180, w_011_8181, w_011_8182, w_011_8183, w_011_8185, w_011_8186, w_011_8187, w_011_8189, w_011_8190, w_011_8192, w_011_8193, w_011_8194, w_011_8195, w_011_8198, w_011_8202, w_011_8203, w_011_8204, w_011_8205, w_011_8206, w_011_8208, w_011_8210, w_011_8211, w_011_8212, w_011_8213, w_011_8214, w_011_8215, w_011_8216, w_011_8217, w_011_8220, w_011_8221, w_011_8222, w_011_8225, w_011_8226, w_011_8230, w_011_8232, w_011_8233, w_011_8234, w_011_8236, w_011_8237, w_011_8238, w_011_8239, w_011_8240, w_011_8241, w_011_8243, w_011_8245, w_011_8246, w_011_8247, w_011_8248, w_011_8249, w_011_8251, w_011_8252, w_011_8253, w_011_8254, w_011_8255, w_011_8256, w_011_8257, w_011_8259, w_011_8260, w_011_8261, w_011_8262, w_011_8263, w_011_8264, w_011_8265, w_011_8266, w_011_8268, w_011_8269, w_011_8270, w_011_8271, w_011_8272, w_011_8274, w_011_8275, w_011_8277, w_011_8278, w_011_8279, w_011_8280, w_011_8282, w_011_8284, w_011_8285, w_011_8286, w_011_8288, w_011_8289, w_011_8290, w_011_8292, w_011_8293, w_011_8294, w_011_8295, w_011_8296, w_011_8297, w_011_8300, w_011_8301, w_011_8302, w_011_8303, w_011_8306, w_011_8307, w_011_8308, w_011_8309, w_011_8310, w_011_8311, w_011_8312, w_011_8316, w_011_8317, w_011_8318, w_011_8319, w_011_8322, w_011_8324, w_011_8325, w_011_8328, w_011_8329, w_011_8330, w_011_8331, w_011_8332, w_011_8333, w_011_8337, w_011_8338, w_011_8339, w_011_8340, w_011_8341, w_011_8342, w_011_8343, w_011_8344, w_011_8345, w_011_8346, w_011_8348, w_011_8350, w_011_8352, w_011_8353, w_011_8354, w_011_8356, w_011_8358, w_011_8359, w_011_8362, w_011_8363, w_011_8364, w_011_8366, w_011_8367, w_011_8368, w_011_8370, w_011_8371, w_011_8374, w_011_8376, w_011_8377, w_011_8378, w_011_8381, w_011_8382, w_011_8383, w_011_8384, w_011_8385, w_011_8386, w_011_8387, w_011_8388, w_011_8389, w_011_8390, w_011_8391, w_011_8392, w_011_8393, w_011_8394, w_011_8395, w_011_8396, w_011_8397, w_011_8398, w_011_8399, w_011_8400, w_011_8402, w_011_8403, w_011_8404, w_011_8405, w_011_8406, w_011_8407, w_011_8409, w_011_8414, w_011_8415, w_011_8417, w_011_8418, w_011_8419, w_011_8420, w_011_8421, w_011_8422, w_011_8425, w_011_8426, w_011_8427, w_011_8428, w_011_8429, w_011_8430, w_011_8431, w_011_8433, w_011_8434, w_011_8436, w_011_8437, w_011_8439, w_011_8440, w_011_8441, w_011_8444, w_011_8446, w_011_8447, w_011_8448, w_011_8449, w_011_8450, w_011_8452, w_011_8453, w_011_8456, w_011_8457, w_011_8458, w_011_8459, w_011_8460, w_011_8461, w_011_8462, w_011_8463, w_011_8466, w_011_8469, w_011_8470, w_011_8471, w_011_8472, w_011_8473, w_011_8474, w_011_8476, w_011_8477, w_011_8478, w_011_8481, w_011_8483, w_011_8484, w_011_8485, w_011_8487, w_011_8488, w_011_8490, w_011_8491, w_011_8492, w_011_8493, w_011_8494, w_011_8495, w_011_8496, w_011_8497, w_011_8498, w_011_8499, w_011_8501, w_011_8502, w_011_8503, w_011_8504, w_011_8505, w_011_8508, w_011_8509, w_011_8510, w_011_8511, w_011_8512, w_011_8513, w_011_8514, w_011_8515, w_011_8517, w_011_8522, w_011_8523, w_011_8524, w_011_8525, w_011_8526, w_011_8527, w_011_8528, w_011_8529, w_011_8531, w_011_8534, w_011_8535, w_011_8536, w_011_8537, w_011_8538, w_011_8539, w_011_8540, w_011_8541, w_011_8542, w_011_8544, w_011_8545, w_011_8546, w_011_8547, w_011_8548, w_011_8549, w_011_8550, w_011_8551, w_011_8552, w_011_8554, w_011_8555, w_011_8556, w_011_8557, w_011_8558, w_011_8559, w_011_8561, w_011_8566, w_011_8567, w_011_8568, w_011_8569, w_011_8570, w_011_8571, w_011_8572, w_011_8573, w_011_8574, w_011_8575, w_011_8576, w_011_8577, w_011_8578, w_011_8581, w_011_8583, w_011_8584, w_011_8586, w_011_8587, w_011_8588, w_011_8589, w_011_8590, w_011_8592, w_011_8594, w_011_8598, w_011_8600, w_011_8601, w_011_8604, w_011_8606, w_011_8609, w_011_8610, w_011_8611, w_011_8612, w_011_8613, w_011_8614, w_011_8616, w_011_8617, w_011_8618, w_011_8619, w_011_8620, w_011_8622, w_011_8623, w_011_8624, w_011_8625, w_011_8626, w_011_8628, w_011_8629, w_011_8633, w_011_8634, w_011_8635, w_011_8637, w_011_8638, w_011_8639, w_011_8640, w_011_8641, w_011_8643, w_011_8644, w_011_8645, w_011_8646, w_011_8647, w_011_8649, w_011_8651, w_011_8652, w_011_8654, w_011_8655, w_011_8656, w_011_8657, w_011_8658, w_011_8659, w_011_8660, w_011_8661, w_011_8662, w_011_8663, w_011_8665, w_011_8667, w_011_8668, w_011_8669, w_011_8670, w_011_8672, w_011_8674, w_011_8675, w_011_8676, w_011_8677, w_011_8678, w_011_8679, w_011_8680, w_011_8682, w_011_8683, w_011_8684, w_011_8685, w_011_8688, w_011_8689, w_011_8690, w_011_8691, w_011_8692, w_011_8693, w_011_8694, w_011_8695, w_011_8696, w_011_8698, w_011_8699, w_011_8700, w_011_8701, w_011_8704, w_011_8705, w_011_8706, w_011_8708, w_011_8709, w_011_8710, w_011_8711, w_011_8712, w_011_8713, w_011_8715, w_011_8716, w_011_8717, w_011_8718, w_011_8719, w_011_8722, w_011_8723, w_011_8724, w_011_8726, w_011_8727, w_011_8728, w_011_8732, w_011_8733, w_011_8736, w_011_8737, w_011_8740, w_011_8742, w_011_8743, w_011_8744, w_011_8745, w_011_8747, w_011_8748, w_011_8750, w_011_8751, w_011_8753, w_011_8755, w_011_8756, w_011_8757, w_011_8758, w_011_8759, w_011_8760, w_011_8761, w_011_8765, w_011_8766, w_011_8767, w_011_8768, w_011_8771, w_011_8772, w_011_8773, w_011_8774, w_011_8775, w_011_8776, w_011_8777, w_011_8778, w_011_8779, w_011_8780, w_011_8781, w_011_8782, w_011_8783, w_011_8786, w_011_8787, w_011_8788, w_011_8789, w_011_8790, w_011_8793, w_011_8794, w_011_8795, w_011_8796, w_011_8797, w_011_8799, w_011_8800, w_011_8801, w_011_8802, w_011_8803, w_011_8805, w_011_8806, w_011_8807, w_011_8808, w_011_8809, w_011_8810, w_011_8811, w_011_8813, w_011_8814, w_011_8815, w_011_8817, w_011_8818, w_011_8819, w_011_8820, w_011_8821, w_011_8824, w_011_8825, w_011_8826, w_011_8827, w_011_8828, w_011_8830, w_011_8831, w_011_8832, w_011_8833, w_011_8835, w_011_8836, w_011_8837, w_011_8838, w_011_8839, w_011_8840, w_011_8841, w_011_8842, w_011_8845, w_011_8847, w_011_8848, w_011_8849, w_011_8851, w_011_8852, w_011_8856, w_011_8858, w_011_8859, w_011_8860, w_011_8861, w_011_8862, w_011_8865, w_011_8866, w_011_8867, w_011_8868, w_011_8869, w_011_8870, w_011_8871, w_011_8872, w_011_8874, w_011_8875, w_011_8876, w_011_8877, w_011_8878, w_011_8879, w_011_8880, w_011_8881, w_011_8884, w_011_8885, w_011_8887, w_011_8888, w_011_8890, w_011_8891, w_011_8892, w_011_8893, w_011_8896, w_011_8897, w_011_8898, w_011_8901, w_011_8902, w_011_8903, w_011_8905, w_011_8906, w_011_8910, w_011_8912, w_011_8913, w_011_8914, w_011_8915, w_011_8917, w_011_8918, w_011_8919, w_011_8921, w_011_8922, w_011_8923, w_011_8924, w_011_8925, w_011_8926, w_011_8927, w_011_8928, w_011_8929, w_011_8930, w_011_8931, w_011_8932, w_011_8933, w_011_8934, w_011_8935, w_011_8936, w_011_8937, w_011_8942, w_011_8947, w_011_8949, w_011_8950, w_011_8951, w_011_8952, w_011_8953, w_011_8954, w_011_8955, w_011_8956, w_011_8957, w_011_8958, w_011_8960, w_011_8962, w_011_8963, w_011_8964, w_011_8965, w_011_8966, w_011_8967, w_011_8971, w_011_8972, w_011_8973, w_011_8974, w_011_8976, w_011_8979, w_011_8981, w_011_8982, w_011_8983, w_011_8984, w_011_8985, w_011_8986, w_011_8987, w_011_8988, w_011_8991, w_011_8992, w_011_8993, w_011_8994, w_011_8995, w_011_8996, w_011_8998, w_011_8999, w_011_9000, w_011_9001, w_011_9003, w_011_9004, w_011_9007, w_011_9008, w_011_9009, w_011_9010, w_011_9011, w_011_9012, w_011_9013, w_011_9014, w_011_9015, w_011_9016, w_011_9017, w_011_9018, w_011_9019, w_011_9021, w_011_9022, w_011_9023, w_011_9025, w_011_9026, w_011_9028, w_011_9029, w_011_9030, w_011_9031, w_011_9032, w_011_9033, w_011_9034, w_011_9035, w_011_9036, w_011_9037, w_011_9038, w_011_9039, w_011_9040, w_011_9041, w_011_9042, w_011_9044, w_011_9045, w_011_9046, w_011_9047, w_011_9048, w_011_9049, w_011_9050, w_011_9051, w_011_9054, w_011_9055, w_011_9056, w_011_9057, w_011_9058, w_011_9059, w_011_9060, w_011_9061, w_011_9063, w_011_9065, w_011_9066, w_011_9067, w_011_9069, w_011_9070, w_011_9074, w_011_9076, w_011_9077, w_011_9078, w_011_9079, w_011_9080, w_011_9081, w_011_9082, w_011_9083, w_011_9084, w_011_9085, w_011_9086, w_011_9087, w_011_9088, w_011_9089, w_011_9090, w_011_9091, w_011_9093, w_011_9094, w_011_9095, w_011_9096, w_011_9098, w_011_9099, w_011_9100, w_011_9101, w_011_9102, w_011_9103, w_011_9105, w_011_9106, w_011_9107, w_011_9108, w_011_9109, w_011_9110, w_011_9111, w_011_9113, w_011_9114, w_011_9115, w_011_9117, w_011_9118, w_011_9119, w_011_9120, w_011_9121, w_011_9124, w_011_9125, w_011_9127, w_011_9129, w_011_9130, w_011_9131, w_011_9132, w_011_9134, w_011_9135, w_011_9136, w_011_9137, w_011_9138, w_011_9139, w_011_9142, w_011_9143, w_011_9144, w_011_9146, w_011_9148, w_011_9149, w_011_9150, w_011_9151, w_011_9152, w_011_9153, w_011_9154, w_011_9155, w_011_9156, w_011_9157;
  wire w_012_000, w_012_001, w_012_002, w_012_003, w_012_004, w_012_005, w_012_006, w_012_007, w_012_008, w_012_009, w_012_010, w_012_011, w_012_012, w_012_013, w_012_014, w_012_015, w_012_016, w_012_017, w_012_018, w_012_019, w_012_020, w_012_021, w_012_022, w_012_023, w_012_024, w_012_025, w_012_026, w_012_027, w_012_028, w_012_029, w_012_030, w_012_031, w_012_032, w_012_033, w_012_034, w_012_035, w_012_036, w_012_037, w_012_038, w_012_039, w_012_040, w_012_041, w_012_042, w_012_043, w_012_044, w_012_045, w_012_046, w_012_047, w_012_048, w_012_049, w_012_050, w_012_051, w_012_052, w_012_053, w_012_054, w_012_055, w_012_056, w_012_057, w_012_058, w_012_059, w_012_060, w_012_061, w_012_062, w_012_063, w_012_064, w_012_065, w_012_066, w_012_067, w_012_068, w_012_069, w_012_070, w_012_071, w_012_072, w_012_073, w_012_074, w_012_075, w_012_076, w_012_077, w_012_078, w_012_079, w_012_080, w_012_081, w_012_082, w_012_083, w_012_084, w_012_085, w_012_086, w_012_087, w_012_088, w_012_089, w_012_091, w_012_092, w_012_093, w_012_094, w_012_095, w_012_096, w_012_097, w_012_098, w_012_099, w_012_100, w_012_101, w_012_102, w_012_103, w_012_104, w_012_105, w_012_106, w_012_107, w_012_108, w_012_109, w_012_110, w_012_111, w_012_112, w_012_113, w_012_114, w_012_115, w_012_116, w_012_117, w_012_118, w_012_119, w_012_120, w_012_121, w_012_122, w_012_123, w_012_124, w_012_125, w_012_126, w_012_127, w_012_128, w_012_129, w_012_130, w_012_131, w_012_132, w_012_133, w_012_134, w_012_135, w_012_136, w_012_137, w_012_138, w_012_139, w_012_140, w_012_141, w_012_142, w_012_143, w_012_144, w_012_145, w_012_146, w_012_147, w_012_148, w_012_149, w_012_150, w_012_151, w_012_152, w_012_153, w_012_154, w_012_155, w_012_156, w_012_157, w_012_158, w_012_159, w_012_160, w_012_161, w_012_162, w_012_163, w_012_164, w_012_165, w_012_166, w_012_167, w_012_168, w_012_169, w_012_170, w_012_171, w_012_172, w_012_173, w_012_174, w_012_175, w_012_176, w_012_177, w_012_178, w_012_179, w_012_180, w_012_181, w_012_182, w_012_183, w_012_184, w_012_185, w_012_186, w_012_187, w_012_188, w_012_189, w_012_190, w_012_191, w_012_192, w_012_193, w_012_194, w_012_195, w_012_196, w_012_197, w_012_198, w_012_199, w_012_200, w_012_201, w_012_202, w_012_203, w_012_204, w_012_206, w_012_207, w_012_208, w_012_209, w_012_210, w_012_211, w_012_212, w_012_213, w_012_214, w_012_215, w_012_216, w_012_217, w_012_218, w_012_219, w_012_220, w_012_221, w_012_222, w_012_223, w_012_224, w_012_225, w_012_226, w_012_227, w_012_228, w_012_229, w_012_230, w_012_231, w_012_232, w_012_233, w_012_234, w_012_235, w_012_236, w_012_237, w_012_238, w_012_239, w_012_240, w_012_241, w_012_242, w_012_243, w_012_244, w_012_245, w_012_246, w_012_247, w_012_248, w_012_249, w_012_250, w_012_251, w_012_252, w_012_253, w_012_254, w_012_255, w_012_256, w_012_257, w_012_258, w_012_259, w_012_260, w_012_261, w_012_262, w_012_263, w_012_264, w_012_265, w_012_266, w_012_267, w_012_268, w_012_269, w_012_270, w_012_271, w_012_272, w_012_273, w_012_274, w_012_275, w_012_276, w_012_277, w_012_278, w_012_279, w_012_280, w_012_281, w_012_282, w_012_283, w_012_284, w_012_285, w_012_286, w_012_287, w_012_288, w_012_289, w_012_290, w_012_291, w_012_292, w_012_293, w_012_294, w_012_295, w_012_296, w_012_297, w_012_298, w_012_299, w_012_300, w_012_301, w_012_302, w_012_303, w_012_304, w_012_305, w_012_306, w_012_307, w_012_308, w_012_309, w_012_310, w_012_311, w_012_312, w_012_313, w_012_314, w_012_315, w_012_316, w_012_317, w_012_318, w_012_319, w_012_320, w_012_321, w_012_322, w_012_323, w_012_324, w_012_325, w_012_326, w_012_327, w_012_328, w_012_329, w_012_330, w_012_331, w_012_332, w_012_333, w_012_334, w_012_335, w_012_336, w_012_337, w_012_338, w_012_339, w_012_340, w_012_341, w_012_342, w_012_343, w_012_344, w_012_345, w_012_346, w_012_347, w_012_348, w_012_349, w_012_350, w_012_351, w_012_352, w_012_353, w_012_354, w_012_355, w_012_356, w_012_357, w_012_358, w_012_359, w_012_360, w_012_361, w_012_362, w_012_363, w_012_364, w_012_365, w_012_366, w_012_367, w_012_368, w_012_369, w_012_370, w_012_371, w_012_372, w_012_373, w_012_374, w_012_375, w_012_376, w_012_377, w_012_378, w_012_379, w_012_380, w_012_381, w_012_382, w_012_383, w_012_384, w_012_385, w_012_386, w_012_387, w_012_388, w_012_389, w_012_390, w_012_391, w_012_392, w_012_393, w_012_394, w_012_395, w_012_396, w_012_397, w_012_398, w_012_399, w_012_400, w_012_401, w_012_402, w_012_403, w_012_404, w_012_405, w_012_406, w_012_407, w_012_408, w_012_409, w_012_410, w_012_411, w_012_412, w_012_413, w_012_414, w_012_415, w_012_416, w_012_417, w_012_418, w_012_419, w_012_420, w_012_421, w_012_422, w_012_423, w_012_424, w_012_425, w_012_426, w_012_427, w_012_428, w_012_429, w_012_430, w_012_431, w_012_432, w_012_433, w_012_434, w_012_435, w_012_436, w_012_437, w_012_438, w_012_439, w_012_440, w_012_441, w_012_442, w_012_443, w_012_444, w_012_445, w_012_446, w_012_447, w_012_448, w_012_449, w_012_450, w_012_451, w_012_452, w_012_453, w_012_454, w_012_455, w_012_456, w_012_457, w_012_458, w_012_459, w_012_460, w_012_461, w_012_462, w_012_463, w_012_464, w_012_465, w_012_466, w_012_467, w_012_468, w_012_469, w_012_470, w_012_471, w_012_472, w_012_473, w_012_474, w_012_475, w_012_476, w_012_477, w_012_478, w_012_479, w_012_480, w_012_481, w_012_482, w_012_483, w_012_484, w_012_485, w_012_486, w_012_487, w_012_488, w_012_489, w_012_490, w_012_491, w_012_492, w_012_493, w_012_494, w_012_495, w_012_496, w_012_497, w_012_498, w_012_499, w_012_500, w_012_501, w_012_502, w_012_503, w_012_504, w_012_505, w_012_506, w_012_507, w_012_508, w_012_509, w_012_510, w_012_511, w_012_512, w_012_513, w_012_514, w_012_515, w_012_516, w_012_517, w_012_518, w_012_519, w_012_520, w_012_521, w_012_522, w_012_523, w_012_524, w_012_525, w_012_526, w_012_527, w_012_528, w_012_529, w_012_530, w_012_531, w_012_532, w_012_533, w_012_534, w_012_535, w_012_536, w_012_537, w_012_538, w_012_539, w_012_540, w_012_541, w_012_542, w_012_543, w_012_544, w_012_545, w_012_546, w_012_547, w_012_548, w_012_549, w_012_550, w_012_551, w_012_552, w_012_553, w_012_554, w_012_555, w_012_556, w_012_557, w_012_558, w_012_559, w_012_560, w_012_561, w_012_562, w_012_563, w_012_564, w_012_565, w_012_566, w_012_567, w_012_568, w_012_569, w_012_570, w_012_571, w_012_572, w_012_573, w_012_574, w_012_575, w_012_576, w_012_577, w_012_578, w_012_579, w_012_580, w_012_581, w_012_582, w_012_583, w_012_584, w_012_585, w_012_586, w_012_587, w_012_588, w_012_589, w_012_590, w_012_591, w_012_592, w_012_593, w_012_594, w_012_595, w_012_596, w_012_597, w_012_598, w_012_599, w_012_600, w_012_601, w_012_602, w_012_603, w_012_604, w_012_605, w_012_606, w_012_607, w_012_608, w_012_609, w_012_610, w_012_611, w_012_612, w_012_613, w_012_614, w_012_615, w_012_616, w_012_617, w_012_618, w_012_619, w_012_620, w_012_621, w_012_622, w_012_623, w_012_624, w_012_625, w_012_626, w_012_627, w_012_628, w_012_629, w_012_630, w_012_631, w_012_632, w_012_633, w_012_634, w_012_635, w_012_636, w_012_637, w_012_638, w_012_639, w_012_640, w_012_641, w_012_642, w_012_644, w_012_645, w_012_646, w_012_647, w_012_648, w_012_649, w_012_650, w_012_651, w_012_652, w_012_653, w_012_654, w_012_655, w_012_656, w_012_657, w_012_658, w_012_659, w_012_660, w_012_661, w_012_662, w_012_663, w_012_664, w_012_665, w_012_666, w_012_667, w_012_668, w_012_669, w_012_670, w_012_671, w_012_672, w_012_673, w_012_674, w_012_675, w_012_676, w_012_677, w_012_678, w_012_679, w_012_680, w_012_681, w_012_682, w_012_683, w_012_684, w_012_685, w_012_686, w_012_687, w_012_688, w_012_689, w_012_690, w_012_691, w_012_692, w_012_693, w_012_694, w_012_695, w_012_696, w_012_697, w_012_698, w_012_699, w_012_700, w_012_701, w_012_702, w_012_703, w_012_704, w_012_705, w_012_706, w_012_707, w_012_708, w_012_709, w_012_710, w_012_711, w_012_712, w_012_713, w_012_714, w_012_715, w_012_717, w_012_718, w_012_719, w_012_720, w_012_721, w_012_722, w_012_723, w_012_724, w_012_725, w_012_726, w_012_727, w_012_728, w_012_729, w_012_730, w_012_731, w_012_732, w_012_733, w_012_734, w_012_735, w_012_736, w_012_737, w_012_738, w_012_739, w_012_740, w_012_741, w_012_742, w_012_743, w_012_744, w_012_745, w_012_746, w_012_747, w_012_748, w_012_749, w_012_750, w_012_751, w_012_752, w_012_753, w_012_754, w_012_755, w_012_756, w_012_757, w_012_758, w_012_759, w_012_760, w_012_761, w_012_762, w_012_763, w_012_764, w_012_766, w_012_767, w_012_768, w_012_770, w_012_771, w_012_772, w_012_773, w_012_774, w_012_776, w_012_777, w_012_778, w_012_779, w_012_780, w_012_781, w_012_782, w_012_783, w_012_784, w_012_785, w_012_786, w_012_787, w_012_788, w_012_789, w_012_790, w_012_792, w_012_793, w_012_795, w_012_796, w_012_797, w_012_798, w_012_799, w_012_800, w_012_801, w_012_802, w_012_803, w_012_804, w_012_805, w_012_806, w_012_807, w_012_808, w_012_809, w_012_810, w_012_811, w_012_812, w_012_813, w_012_814, w_012_815, w_012_816, w_012_817, w_012_818, w_012_819, w_012_820, w_012_821, w_012_822, w_012_823, w_012_824, w_012_825, w_012_826, w_012_827, w_012_828, w_012_829, w_012_830, w_012_831, w_012_832, w_012_833, w_012_834, w_012_835, w_012_836, w_012_837, w_012_838, w_012_839, w_012_840, w_012_841, w_012_842, w_012_843, w_012_844, w_012_845, w_012_846, w_012_847, w_012_848, w_012_849, w_012_850, w_012_851, w_012_852, w_012_853, w_012_854, w_012_855, w_012_856, w_012_857, w_012_858, w_012_859, w_012_860, w_012_861, w_012_862, w_012_863, w_012_864, w_012_865, w_012_866, w_012_867, w_012_868, w_012_869, w_012_870, w_012_871, w_012_872, w_012_873, w_012_874, w_012_875, w_012_876, w_012_877, w_012_878, w_012_879, w_012_880, w_012_881, w_012_882, w_012_883, w_012_884, w_012_885, w_012_886, w_012_887, w_012_888, w_012_889, w_012_890, w_012_891, w_012_892, w_012_893, w_012_894, w_012_895, w_012_896, w_012_897, w_012_898, w_012_899, w_012_900, w_012_901, w_012_902, w_012_903, w_012_904, w_012_905, w_012_906, w_012_907, w_012_908, w_012_909, w_012_910, w_012_911, w_012_912, w_012_913, w_012_914, w_012_915, w_012_916, w_012_917, w_012_918, w_012_919, w_012_920, w_012_921, w_012_922, w_012_923, w_012_924, w_012_925, w_012_926, w_012_927, w_012_928, w_012_929, w_012_930, w_012_931, w_012_932, w_012_933, w_012_934, w_012_935, w_012_936, w_012_937, w_012_938, w_012_939, w_012_940, w_012_941, w_012_942, w_012_943, w_012_944, w_012_945, w_012_946, w_012_947, w_012_948, w_012_949, w_012_950, w_012_951, w_012_952, w_012_953, w_012_954, w_012_955, w_012_956, w_012_957, w_012_958, w_012_959, w_012_960, w_012_961, w_012_962, w_012_963, w_012_964, w_012_965, w_012_966, w_012_967, w_012_968, w_012_969, w_012_970, w_012_971, w_012_972, w_012_974, w_012_975, w_012_976, w_012_977, w_012_978, w_012_979, w_012_980, w_012_981, w_012_982, w_012_983, w_012_984, w_012_985, w_012_986, w_012_987, w_012_988, w_012_989, w_012_990, w_012_991, w_012_992, w_012_993, w_012_994, w_012_995, w_012_996, w_012_997, w_012_998, w_012_999, w_012_1000, w_012_1001, w_012_1002, w_012_1003, w_012_1004, w_012_1005, w_012_1006, w_012_1007, w_012_1008, w_012_1009, w_012_1010, w_012_1011, w_012_1012, w_012_1013, w_012_1014, w_012_1015, w_012_1016, w_012_1017, w_012_1018, w_012_1019, w_012_1020, w_012_1021, w_012_1022, w_012_1023, w_012_1024, w_012_1025, w_012_1026, w_012_1028, w_012_1029, w_012_1030, w_012_1031, w_012_1032, w_012_1033, w_012_1034, w_012_1035, w_012_1036, w_012_1037, w_012_1038, w_012_1039, w_012_1040, w_012_1041, w_012_1042, w_012_1043, w_012_1044, w_012_1045, w_012_1046, w_012_1047, w_012_1048, w_012_1049, w_012_1050, w_012_1051, w_012_1052, w_012_1053, w_012_1054, w_012_1055, w_012_1056, w_012_1057, w_012_1058, w_012_1059, w_012_1060, w_012_1061, w_012_1062, w_012_1063, w_012_1064, w_012_1065, w_012_1066, w_012_1067, w_012_1068, w_012_1069, w_012_1070, w_012_1071, w_012_1072, w_012_1073, w_012_1074, w_012_1075, w_012_1076, w_012_1077, w_012_1078, w_012_1079, w_012_1080, w_012_1081, w_012_1082, w_012_1083, w_012_1084, w_012_1085, w_012_1086, w_012_1087, w_012_1088, w_012_1089, w_012_1090, w_012_1091, w_012_1092, w_012_1093, w_012_1094, w_012_1095, w_012_1096, w_012_1097, w_012_1098, w_012_1099, w_012_1100, w_012_1101, w_012_1102, w_012_1103, w_012_1104, w_012_1105, w_012_1106, w_012_1107, w_012_1108, w_012_1109, w_012_1110, w_012_1111, w_012_1112, w_012_1113, w_012_1114, w_012_1115, w_012_1116, w_012_1117, w_012_1118, w_012_1119, w_012_1120, w_012_1121, w_012_1122, w_012_1123, w_012_1124, w_012_1125, w_012_1126, w_012_1127, w_012_1128, w_012_1129, w_012_1130, w_012_1131, w_012_1132, w_012_1133, w_012_1134, w_012_1135, w_012_1136, w_012_1137, w_012_1138, w_012_1139, w_012_1140, w_012_1141, w_012_1142, w_012_1143, w_012_1144, w_012_1145, w_012_1147, w_012_1148, w_012_1149, w_012_1150, w_012_1151, w_012_1152, w_012_1153, w_012_1154, w_012_1155, w_012_1156, w_012_1157, w_012_1158, w_012_1160, w_012_1161, w_012_1162, w_012_1163, w_012_1164, w_012_1165, w_012_1166, w_012_1167, w_012_1168, w_012_1169, w_012_1170, w_012_1171, w_012_1172, w_012_1173, w_012_1174, w_012_1175, w_012_1176, w_012_1177, w_012_1178, w_012_1179, w_012_1180, w_012_1181, w_012_1182, w_012_1183, w_012_1184, w_012_1185, w_012_1187, w_012_1188, w_012_1189, w_012_1190, w_012_1191, w_012_1192, w_012_1193, w_012_1194, w_012_1195, w_012_1196, w_012_1197, w_012_1198, w_012_1199, w_012_1200, w_012_1201, w_012_1202, w_012_1203, w_012_1204, w_012_1205, w_012_1206, w_012_1207, w_012_1208, w_012_1209, w_012_1210, w_012_1211, w_012_1212, w_012_1213, w_012_1214, w_012_1215, w_012_1216, w_012_1217, w_012_1218, w_012_1219, w_012_1220, w_012_1221, w_012_1222, w_012_1223, w_012_1224, w_012_1225, w_012_1226, w_012_1227, w_012_1228, w_012_1229, w_012_1230, w_012_1231, w_012_1232, w_012_1233, w_012_1234, w_012_1235, w_012_1236, w_012_1237, w_012_1238, w_012_1239, w_012_1240, w_012_1241, w_012_1242, w_012_1243, w_012_1244, w_012_1245, w_012_1246, w_012_1247, w_012_1248, w_012_1249, w_012_1250, w_012_1251, w_012_1252, w_012_1253, w_012_1254, w_012_1255, w_012_1256, w_012_1257, w_012_1258, w_012_1259, w_012_1260, w_012_1261, w_012_1262, w_012_1263, w_012_1264, w_012_1265, w_012_1266, w_012_1267, w_012_1268, w_012_1269, w_012_1270, w_012_1271, w_012_1272, w_012_1274, w_012_1275, w_012_1276, w_012_1277, w_012_1278, w_012_1279, w_012_1280, w_012_1281, w_012_1282, w_012_1283, w_012_1284, w_012_1285, w_012_1286, w_012_1287, w_012_1288, w_012_1289, w_012_1290, w_012_1291, w_012_1292, w_012_1293, w_012_1294, w_012_1295, w_012_1296, w_012_1297, w_012_1298, w_012_1299, w_012_1300, w_012_1301, w_012_1302, w_012_1303, w_012_1304, w_012_1305, w_012_1306, w_012_1307, w_012_1308, w_012_1309, w_012_1310, w_012_1311, w_012_1312, w_012_1313, w_012_1314, w_012_1315, w_012_1316, w_012_1317, w_012_1318, w_012_1319, w_012_1320, w_012_1322, w_012_1323, w_012_1324, w_012_1325, w_012_1326, w_012_1327, w_012_1328, w_012_1329, w_012_1330, w_012_1331, w_012_1332, w_012_1334, w_012_1335, w_012_1336, w_012_1337, w_012_1338, w_012_1339, w_012_1340, w_012_1341, w_012_1342, w_012_1343, w_012_1344, w_012_1345, w_012_1346, w_012_1347, w_012_1348, w_012_1349, w_012_1350, w_012_1351, w_012_1352, w_012_1353, w_012_1354, w_012_1355, w_012_1356, w_012_1357, w_012_1358, w_012_1359, w_012_1360, w_012_1361, w_012_1362, w_012_1363, w_012_1364, w_012_1365, w_012_1366, w_012_1367, w_012_1368, w_012_1369, w_012_1370, w_012_1371, w_012_1372, w_012_1373, w_012_1374, w_012_1375, w_012_1376, w_012_1377, w_012_1378, w_012_1379, w_012_1380, w_012_1381, w_012_1382, w_012_1383, w_012_1384, w_012_1385, w_012_1386, w_012_1387, w_012_1388, w_012_1389, w_012_1390, w_012_1391, w_012_1392, w_012_1393, w_012_1394, w_012_1395, w_012_1396, w_012_1397, w_012_1398, w_012_1399, w_012_1400, w_012_1401, w_012_1402, w_012_1403, w_012_1404, w_012_1405, w_012_1406, w_012_1407, w_012_1408, w_012_1409, w_012_1410, w_012_1411, w_012_1412, w_012_1413, w_012_1414, w_012_1415, w_012_1416, w_012_1417, w_012_1418, w_012_1419, w_012_1420, w_012_1421, w_012_1422, w_012_1423, w_012_1424, w_012_1425, w_012_1426, w_012_1427, w_012_1428, w_012_1429, w_012_1430, w_012_1431, w_012_1432, w_012_1433, w_012_1435, w_012_1436, w_012_1437, w_012_1438, w_012_1439, w_012_1440, w_012_1441, w_012_1442, w_012_1443, w_012_1444, w_012_1445, w_012_1446, w_012_1447, w_012_1448, w_012_1449, w_012_1450, w_012_1451, w_012_1452, w_012_1453, w_012_1454, w_012_1455, w_012_1456, w_012_1457, w_012_1458, w_012_1459, w_012_1460, w_012_1461, w_012_1462, w_012_1463, w_012_1464, w_012_1465, w_012_1466, w_012_1467, w_012_1468, w_012_1469, w_012_1471, w_012_1472, w_012_1473, w_012_1474, w_012_1475, w_012_1476, w_012_1477, w_012_1479, w_012_1480, w_012_1481, w_012_1482, w_012_1483, w_012_1484, w_012_1485, w_012_1486, w_012_1487, w_012_1488, w_012_1489, w_012_1490, w_012_1491, w_012_1492, w_012_1494, w_012_1495, w_012_1496, w_012_1497, w_012_1498, w_012_1499, w_012_1500, w_012_1501, w_012_1502, w_012_1503, w_012_1504, w_012_1505, w_012_1506, w_012_1507, w_012_1508, w_012_1509, w_012_1510, w_012_1511, w_012_1512, w_012_1513, w_012_1514, w_012_1515, w_012_1516, w_012_1517, w_012_1519, w_012_1520, w_012_1521, w_012_1522, w_012_1523, w_012_1524, w_012_1525, w_012_1526, w_012_1527, w_012_1528, w_012_1529, w_012_1530, w_012_1531, w_012_1532, w_012_1533, w_012_1534, w_012_1535, w_012_1536, w_012_1537, w_012_1538, w_012_1539, w_012_1540, w_012_1541, w_012_1542, w_012_1543, w_012_1544, w_012_1545, w_012_1546, w_012_1547, w_012_1548, w_012_1549, w_012_1550, w_012_1551, w_012_1552, w_012_1553, w_012_1554, w_012_1555, w_012_1556, w_012_1557, w_012_1558, w_012_1559, w_012_1561, w_012_1562, w_012_1563, w_012_1565, w_012_1566, w_012_1567, w_012_1568, w_012_1569, w_012_1570, w_012_1571, w_012_1572, w_012_1574, w_012_1575, w_012_1576, w_012_1577, w_012_1578, w_012_1579, w_012_1580, w_012_1581, w_012_1582, w_012_1583, w_012_1584, w_012_1585, w_012_1586, w_012_1588, w_012_1589, w_012_1590, w_012_1591, w_012_1592, w_012_1593, w_012_1594, w_012_1595, w_012_1596, w_012_1597, w_012_1598, w_012_1599, w_012_1600, w_012_1601, w_012_1602, w_012_1603, w_012_1604, w_012_1605, w_012_1606, w_012_1607, w_012_1608, w_012_1609, w_012_1610, w_012_1611, w_012_1612, w_012_1613, w_012_1614, w_012_1615, w_012_1616, w_012_1617, w_012_1618, w_012_1619, w_012_1620, w_012_1621, w_012_1622, w_012_1623, w_012_1624, w_012_1625, w_012_1626, w_012_1627, w_012_1628, w_012_1630, w_012_1631, w_012_1633, w_012_1634, w_012_1635, w_012_1636, w_012_1637, w_012_1638, w_012_1639, w_012_1640, w_012_1641, w_012_1642, w_012_1643, w_012_1644, w_012_1645, w_012_1646, w_012_1647, w_012_1648, w_012_1649, w_012_1650, w_012_1651, w_012_1652, w_012_1653, w_012_1654, w_012_1655, w_012_1656, w_012_1657, w_012_1658, w_012_1659, w_012_1660, w_012_1661, w_012_1662, w_012_1663, w_012_1664, w_012_1665, w_012_1666, w_012_1667, w_012_1668, w_012_1669, w_012_1670, w_012_1671, w_012_1672, w_012_1673, w_012_1674, w_012_1675, w_012_1676, w_012_1677, w_012_1678, w_012_1679, w_012_1680, w_012_1681, w_012_1682, w_012_1683, w_012_1684, w_012_1685, w_012_1686, w_012_1687, w_012_1688, w_012_1689, w_012_1690, w_012_1691, w_012_1692, w_012_1693, w_012_1694, w_012_1695, w_012_1696, w_012_1697, w_012_1698, w_012_1699, w_012_1700, w_012_1701, w_012_1702, w_012_1703, w_012_1704, w_012_1705, w_012_1706, w_012_1707, w_012_1708, w_012_1709, w_012_1710, w_012_1711, w_012_1712, w_012_1713, w_012_1714, w_012_1715, w_012_1716, w_012_1717, w_012_1718, w_012_1719, w_012_1720, w_012_1721, w_012_1722, w_012_1723, w_012_1724, w_012_1725, w_012_1726, w_012_1727, w_012_1728, w_012_1729, w_012_1730, w_012_1731, w_012_1732, w_012_1733, w_012_1734, w_012_1735, w_012_1736, w_012_1737, w_012_1738, w_012_1740, w_012_1741, w_012_1742, w_012_1743, w_012_1744, w_012_1745, w_012_1746, w_012_1747, w_012_1748, w_012_1749, w_012_1750, w_012_1751, w_012_1752, w_012_1753, w_012_1754, w_012_1755, w_012_1756, w_012_1757, w_012_1758, w_012_1759, w_012_1760, w_012_1761, w_012_1762, w_012_1763, w_012_1764, w_012_1765, w_012_1766, w_012_1767, w_012_1768, w_012_1769, w_012_1770, w_012_1771, w_012_1772, w_012_1773, w_012_1774, w_012_1775, w_012_1776, w_012_1777, w_012_1778, w_012_1779, w_012_1780, w_012_1781, w_012_1782, w_012_1783, w_012_1784, w_012_1785, w_012_1786, w_012_1787, w_012_1788, w_012_1789, w_012_1790, w_012_1791, w_012_1792, w_012_1793, w_012_1794, w_012_1795, w_012_1796, w_012_1797, w_012_1798, w_012_1799, w_012_1800, w_012_1801, w_012_1802, w_012_1803, w_012_1804, w_012_1805, w_012_1806, w_012_1807, w_012_1808, w_012_1809, w_012_1810, w_012_1811, w_012_1812, w_012_1813, w_012_1814, w_012_1815, w_012_1816, w_012_1817, w_012_1818, w_012_1819, w_012_1820, w_012_1821, w_012_1822, w_012_1823, w_012_1824, w_012_1825, w_012_1826, w_012_1827, w_012_1828, w_012_1829, w_012_1831, w_012_1832, w_012_1833, w_012_1834, w_012_1835, w_012_1836, w_012_1837, w_012_1838, w_012_1839, w_012_1840, w_012_1841, w_012_1842, w_012_1843, w_012_1844, w_012_1845, w_012_1846, w_012_1847, w_012_1848, w_012_1849, w_012_1850, w_012_1851, w_012_1852, w_012_1853, w_012_1854, w_012_1855, w_012_1857, w_012_1858, w_012_1859, w_012_1860, w_012_1861, w_012_1862, w_012_1863, w_012_1864, w_012_1865, w_012_1866, w_012_1867, w_012_1868, w_012_1869, w_012_1870, w_012_1871, w_012_1873, w_012_1874, w_012_1875, w_012_1876, w_012_1877, w_012_1878, w_012_1879, w_012_1880, w_012_1881, w_012_1882, w_012_1883, w_012_1884, w_012_1885, w_012_1886, w_012_1887, w_012_1888, w_012_1889, w_012_1890, w_012_1891, w_012_1892, w_012_1893, w_012_1894, w_012_1895, w_012_1896, w_012_1897, w_012_1898, w_012_1899, w_012_1900, w_012_1901, w_012_1902, w_012_1903, w_012_1905, w_012_1906, w_012_1907, w_012_1908, w_012_1909, w_012_1910, w_012_1911, w_012_1912, w_012_1913, w_012_1914, w_012_1915, w_012_1916, w_012_1917, w_012_1918, w_012_1919, w_012_1920, w_012_1921, w_012_1922, w_012_1923, w_012_1924, w_012_1925, w_012_1926, w_012_1927, w_012_1928, w_012_1929, w_012_1930, w_012_1931, w_012_1932, w_012_1933, w_012_1934, w_012_1936, w_012_1937, w_012_1938, w_012_1939, w_012_1940, w_012_1941, w_012_1943, w_012_1944, w_012_1945, w_012_1946, w_012_1947, w_012_1948, w_012_1949, w_012_1950, w_012_1951, w_012_1952, w_012_1953, w_012_1954, w_012_1955, w_012_1956, w_012_1957, w_012_1958, w_012_1959, w_012_1960, w_012_1961, w_012_1962, w_012_1963, w_012_1964, w_012_1965, w_012_1966, w_012_1967, w_012_1968, w_012_1969, w_012_1970, w_012_1971, w_012_1972, w_012_1973, w_012_1974, w_012_1975, w_012_1976, w_012_1977, w_012_1978, w_012_1979, w_012_1980, w_012_1981, w_012_1982, w_012_1983, w_012_1984, w_012_1985, w_012_1986, w_012_1987, w_012_1988, w_012_1989, w_012_1990, w_012_1991, w_012_1992, w_012_1993, w_012_1994, w_012_1995, w_012_1996, w_012_1997, w_012_1999, w_012_2000, w_012_2001, w_012_2002, w_012_2003, w_012_2004, w_012_2005, w_012_2006, w_012_2007, w_012_2008, w_012_2009, w_012_2010, w_012_2011, w_012_2012, w_012_2013, w_012_2014, w_012_2015, w_012_2016, w_012_2017, w_012_2018, w_012_2019, w_012_2020, w_012_2021, w_012_2022, w_012_2023, w_012_2024, w_012_2025, w_012_2026, w_012_2027, w_012_2028, w_012_2029, w_012_2030, w_012_2031, w_012_2032, w_012_2033, w_012_2034, w_012_2035, w_012_2036, w_012_2037, w_012_2038, w_012_2039, w_012_2040, w_012_2041, w_012_2042, w_012_2043, w_012_2044, w_012_2045, w_012_2046, w_012_2047, w_012_2048, w_012_2049, w_012_2050, w_012_2051, w_012_2052, w_012_2053, w_012_2054, w_012_2055, w_012_2056, w_012_2057, w_012_2058, w_012_2059, w_012_2060, w_012_2061, w_012_2062, w_012_2063, w_012_2064, w_012_2065, w_012_2066, w_012_2067, w_012_2068, w_012_2069, w_012_2070, w_012_2071, w_012_2072, w_012_2073, w_012_2074, w_012_2075, w_012_2076, w_012_2077, w_012_2078, w_012_2080, w_012_2081, w_012_2082, w_012_2084, w_012_2085, w_012_2086, w_012_2087, w_012_2088, w_012_2089, w_012_2090, w_012_2091, w_012_2092, w_012_2093, w_012_2094, w_012_2095, w_012_2096, w_012_2097, w_012_2098, w_012_2099, w_012_2100, w_012_2101, w_012_2102, w_012_2103, w_012_2104, w_012_2105, w_012_2106, w_012_2107, w_012_2108, w_012_2109, w_012_2110, w_012_2111, w_012_2112, w_012_2113, w_012_2114, w_012_2115, w_012_2116, w_012_2117, w_012_2118, w_012_2119, w_012_2120, w_012_2121, w_012_2122, w_012_2123, w_012_2124, w_012_2125, w_012_2126, w_012_2127, w_012_2128, w_012_2129, w_012_2130, w_012_2131, w_012_2132, w_012_2133, w_012_2134, w_012_2135, w_012_2136, w_012_2137, w_012_2138, w_012_2139, w_012_2140, w_012_2141, w_012_2142, w_012_2143, w_012_2144, w_012_2145, w_012_2146, w_012_2147, w_012_2148, w_012_2149, w_012_2150, w_012_2151, w_012_2152, w_012_2153, w_012_2154, w_012_2155, w_012_2156, w_012_2157, w_012_2158, w_012_2159, w_012_2160, w_012_2161, w_012_2162, w_012_2163, w_012_2164, w_012_2165, w_012_2166, w_012_2167, w_012_2168, w_012_2169, w_012_2170, w_012_2171, w_012_2172, w_012_2173, w_012_2174, w_012_2175, w_012_2176, w_012_2177, w_012_2178, w_012_2179, w_012_2181, w_012_2182, w_012_2183, w_012_2184, w_012_2185, w_012_2186, w_012_2187, w_012_2188, w_012_2189, w_012_2190, w_012_2191, w_012_2192, w_012_2193, w_012_2194, w_012_2195, w_012_2196, w_012_2197, w_012_2198, w_012_2199, w_012_2200, w_012_2201, w_012_2202, w_012_2203, w_012_2204, w_012_2205, w_012_2206, w_012_2207, w_012_2208, w_012_2209, w_012_2210, w_012_2211, w_012_2212, w_012_2213, w_012_2214, w_012_2215, w_012_2216, w_012_2217, w_012_2218, w_012_2219, w_012_2220, w_012_2221, w_012_2222, w_012_2223, w_012_2224, w_012_2225, w_012_2226, w_012_2227, w_012_2228, w_012_2229, w_012_2230, w_012_2231, w_012_2232, w_012_2233, w_012_2234, w_012_2235, w_012_2236, w_012_2237, w_012_2238, w_012_2239, w_012_2240, w_012_2241, w_012_2242, w_012_2243, w_012_2244, w_012_2246, w_012_2247, w_012_2248, w_012_2249, w_012_2250, w_012_2252, w_012_2253, w_012_2254, w_012_2255, w_012_2256, w_012_2257, w_012_2258, w_012_2259, w_012_2260, w_012_2261, w_012_2262, w_012_2263, w_012_2264, w_012_2265, w_012_2266, w_012_2267, w_012_2268, w_012_2269, w_012_2270, w_012_2271, w_012_2272, w_012_2273, w_012_2274, w_012_2275, w_012_2276, w_012_2277, w_012_2278, w_012_2279, w_012_2280, w_012_2281, w_012_2282, w_012_2283, w_012_2284, w_012_2285, w_012_2286, w_012_2287, w_012_2288, w_012_2289, w_012_2290, w_012_2292, w_012_2293, w_012_2294, w_012_2295, w_012_2296, w_012_2297, w_012_2298, w_012_2299, w_012_2300, w_012_2301, w_012_2302, w_012_2303, w_012_2304, w_012_2305, w_012_2306, w_012_2307, w_012_2308, w_012_2309, w_012_2310, w_012_2311, w_012_2312, w_012_2313, w_012_2314, w_012_2315, w_012_2316, w_012_2317, w_012_2318, w_012_2319, w_012_2320, w_012_2321, w_012_2322, w_012_2323, w_012_2324, w_012_2325, w_012_2326, w_012_2327, w_012_2328, w_012_2329, w_012_2330, w_012_2331, w_012_2332, w_012_2333, w_012_2334, w_012_2335, w_012_2336, w_012_2337, w_012_2338, w_012_2339, w_012_2340, w_012_2341, w_012_2342, w_012_2343, w_012_2344, w_012_2345, w_012_2346, w_012_2347, w_012_2348, w_012_2349, w_012_2350, w_012_2351, w_012_2352, w_012_2353, w_012_2354, w_012_2355, w_012_2356, w_012_2358, w_012_2359, w_012_2360, w_012_2361, w_012_2362, w_012_2363, w_012_2364, w_012_2365, w_012_2366, w_012_2367, w_012_2368, w_012_2369, w_012_2370, w_012_2371, w_012_2372, w_012_2373, w_012_2374, w_012_2375, w_012_2376, w_012_2377, w_012_2378, w_012_2379, w_012_2380, w_012_2381, w_012_2382, w_012_2383, w_012_2384, w_012_2385, w_012_2386, w_012_2387, w_012_2388, w_012_2389, w_012_2390, w_012_2392, w_012_2393, w_012_2394, w_012_2395, w_012_2396, w_012_2397, w_012_2398, w_012_2399, w_012_2400, w_012_2401, w_012_2402, w_012_2403, w_012_2404, w_012_2405, w_012_2406, w_012_2407, w_012_2408, w_012_2409, w_012_2410, w_012_2411, w_012_2412, w_012_2413, w_012_2414, w_012_2415, w_012_2416, w_012_2417, w_012_2418, w_012_2419, w_012_2420, w_012_2421, w_012_2422, w_012_2423, w_012_2424, w_012_2425, w_012_2426, w_012_2427, w_012_2428, w_012_2429, w_012_2430, w_012_2431, w_012_2432, w_012_2433, w_012_2434, w_012_2435, w_012_2436, w_012_2438, w_012_2439, w_012_2440, w_012_2441, w_012_2442, w_012_2443, w_012_2444, w_012_2445, w_012_2446, w_012_2447, w_012_2448, w_012_2449, w_012_2450, w_012_2451, w_012_2452, w_012_2454, w_012_2455, w_012_2456, w_012_2457, w_012_2458, w_012_2459, w_012_2460, w_012_2461, w_012_2462, w_012_2463, w_012_2464, w_012_2465, w_012_2466, w_012_2467, w_012_2468, w_012_2469, w_012_2470, w_012_2471, w_012_2472, w_012_2473, w_012_2474, w_012_2475, w_012_2476, w_012_2477, w_012_2478, w_012_2479, w_012_2480, w_012_2481, w_012_2483, w_012_2484, w_012_2485, w_012_2486, w_012_2487, w_012_2488, w_012_2489, w_012_2490, w_012_2491, w_012_2492, w_012_2493, w_012_2494, w_012_2495, w_012_2496, w_012_2497, w_012_2498, w_012_2499, w_012_2500, w_012_2501, w_012_2502, w_012_2504, w_012_2505, w_012_2506, w_012_2507, w_012_2508, w_012_2509, w_012_2510, w_012_2511, w_012_2512, w_012_2513, w_012_2514, w_012_2515, w_012_2516, w_012_2517, w_012_2518, w_012_2519, w_012_2520, w_012_2521, w_012_2522, w_012_2523, w_012_2524, w_012_2525, w_012_2526, w_012_2527, w_012_2528, w_012_2529, w_012_2530, w_012_2531, w_012_2532, w_012_2533, w_012_2535, w_012_2536, w_012_2537, w_012_2538, w_012_2539, w_012_2540, w_012_2541, w_012_2542, w_012_2543, w_012_2545, w_012_2546, w_012_2547, w_012_2549, w_012_2550, w_012_2551, w_012_2552, w_012_2553, w_012_2554, w_012_2555, w_012_2556, w_012_2557, w_012_2558, w_012_2559, w_012_2560, w_012_2561, w_012_2562, w_012_2563, w_012_2564, w_012_2565, w_012_2566, w_012_2567, w_012_2568, w_012_2569, w_012_2570, w_012_2571, w_012_2572, w_012_2573, w_012_2574, w_012_2575, w_012_2576, w_012_2577, w_012_2578, w_012_2579, w_012_2580, w_012_2581, w_012_2582, w_012_2583, w_012_2584, w_012_2585, w_012_2586, w_012_2587, w_012_2588, w_012_2589, w_012_2590, w_012_2591, w_012_2592, w_012_2593, w_012_2594, w_012_2595, w_012_2596, w_012_2597, w_012_2598, w_012_2599, w_012_2600, w_012_2601, w_012_2602, w_012_2603, w_012_2604, w_012_2605, w_012_2606, w_012_2607, w_012_2608, w_012_2609, w_012_2610, w_012_2611, w_012_2612, w_012_2613, w_012_2614, w_012_2615, w_012_2616, w_012_2617, w_012_2618, w_012_2619, w_012_2620, w_012_2621, w_012_2622, w_012_2623, w_012_2624, w_012_2625, w_012_2626, w_012_2627, w_012_2628, w_012_2629, w_012_2630, w_012_2631, w_012_2632, w_012_2633, w_012_2634, w_012_2635, w_012_2636, w_012_2637, w_012_2638, w_012_2639, w_012_2640, w_012_2641, w_012_2642, w_012_2643, w_012_2644, w_012_2645, w_012_2646, w_012_2647, w_012_2648, w_012_2649, w_012_2650, w_012_2651, w_012_2652, w_012_2653, w_012_2654, w_012_2655, w_012_2656, w_012_2657, w_012_2658, w_012_2659, w_012_2660, w_012_2661, w_012_2662, w_012_2663, w_012_2664, w_012_2665, w_012_2666, w_012_2668, w_012_2669, w_012_2670, w_012_2671, w_012_2672, w_012_2673, w_012_2674, w_012_2675, w_012_2676, w_012_2677, w_012_2678, w_012_2679, w_012_2680, w_012_2681, w_012_2682, w_012_2683, w_012_2684, w_012_2685, w_012_2686, w_012_2687, w_012_2688, w_012_2689, w_012_2690, w_012_2691, w_012_2692, w_012_2693, w_012_2694, w_012_2695, w_012_2696, w_012_2697, w_012_2698, w_012_2699, w_012_2700, w_012_2701, w_012_2702, w_012_2703, w_012_2704, w_012_2705, w_012_2706, w_012_2707, w_012_2708, w_012_2709, w_012_2710, w_012_2711, w_012_2712, w_012_2713, w_012_2714, w_012_2715, w_012_2716, w_012_2717, w_012_2718, w_012_2719, w_012_2720, w_012_2721, w_012_2722, w_012_2723, w_012_2724, w_012_2725, w_012_2726, w_012_2727, w_012_2728, w_012_2729, w_012_2730, w_012_2731, w_012_2732, w_012_2733, w_012_2734, w_012_2735, w_012_2736, w_012_2737, w_012_2738, w_012_2739, w_012_2740, w_012_2741, w_012_2742, w_012_2743, w_012_2744, w_012_2745, w_012_2746, w_012_2747, w_012_2749, w_012_2750, w_012_2751, w_012_2752, w_012_2753, w_012_2754, w_012_2755, w_012_2756, w_012_2757, w_012_2758, w_012_2759, w_012_2760, w_012_2761, w_012_2762, w_012_2763, w_012_2764, w_012_2765, w_012_2766, w_012_2767, w_012_2768, w_012_2769, w_012_2770, w_012_2771, w_012_2772, w_012_2773, w_012_2774, w_012_2775, w_012_2776, w_012_2777, w_012_2778, w_012_2779, w_012_2780, w_012_2781, w_012_2782, w_012_2783, w_012_2784, w_012_2785, w_012_2786, w_012_2787, w_012_2788, w_012_2789, w_012_2790, w_012_2791, w_012_2792, w_012_2793, w_012_2794, w_012_2795, w_012_2796, w_012_2797, w_012_2798, w_012_2799, w_012_2800, w_012_2801, w_012_2802, w_012_2803, w_012_2804, w_012_2805, w_012_2806, w_012_2807, w_012_2808, w_012_2809, w_012_2810, w_012_2811, w_012_2812, w_012_2813, w_012_2814, w_012_2815, w_012_2816, w_012_2817, w_012_2818, w_012_2819, w_012_2820, w_012_2821, w_012_2822, w_012_2823, w_012_2824, w_012_2825, w_012_2826, w_012_2827, w_012_2828, w_012_2829, w_012_2830, w_012_2831, w_012_2832, w_012_2833, w_012_2834, w_012_2835, w_012_2836, w_012_2837, w_012_2838, w_012_2839, w_012_2840, w_012_2843, w_012_2844, w_012_2845, w_012_2846, w_012_2847, w_012_2848, w_012_2849, w_012_2850, w_012_2851, w_012_2852, w_012_2853, w_012_2854, w_012_2855, w_012_2856, w_012_2857, w_012_2858, w_012_2859, w_012_2860, w_012_2861, w_012_2862, w_012_2863, w_012_2864, w_012_2865, w_012_2866, w_012_2867, w_012_2868, w_012_2869, w_012_2870, w_012_2872, w_012_2873, w_012_2874, w_012_2875, w_012_2876, w_012_2877, w_012_2878, w_012_2879, w_012_2880, w_012_2881, w_012_2882, w_012_2883, w_012_2884, w_012_2885, w_012_2886, w_012_2887, w_012_2888, w_012_2889, w_012_2890, w_012_2891, w_012_2892, w_012_2893, w_012_2894, w_012_2895, w_012_2896, w_012_2897, w_012_2898, w_012_2899, w_012_2900, w_012_2901, w_012_2902, w_012_2903, w_012_2904, w_012_2905, w_012_2906, w_012_2907, w_012_2908, w_012_2909, w_012_2910, w_012_2911, w_012_2912, w_012_2913, w_012_2914, w_012_2915, w_012_2916, w_012_2917, w_012_2918, w_012_2919, w_012_2920, w_012_2921, w_012_2922, w_012_2923, w_012_2924, w_012_2925, w_012_2926, w_012_2927, w_012_2928, w_012_2929, w_012_2930, w_012_2931, w_012_2932, w_012_2933, w_012_2934, w_012_2935, w_012_2936, w_012_2937, w_012_2938, w_012_2939, w_012_2940, w_012_2941, w_012_2942, w_012_2943, w_012_2944, w_012_2945, w_012_2946, w_012_2947, w_012_2948, w_012_2950, w_012_2951, w_012_2952, w_012_2953, w_012_2954, w_012_2955, w_012_2956, w_012_2957, w_012_2958, w_012_2959, w_012_2960, w_012_2961, w_012_2962, w_012_2963, w_012_2964, w_012_2965, w_012_2966, w_012_2967, w_012_2968, w_012_2969, w_012_2970, w_012_2971, w_012_2972, w_012_2973, w_012_2974, w_012_2975, w_012_2976, w_012_2977, w_012_2978, w_012_2979, w_012_2980, w_012_2981, w_012_2982, w_012_2983, w_012_2984, w_012_2985, w_012_2986, w_012_2987, w_012_2988, w_012_2989, w_012_2990, w_012_2991, w_012_2992, w_012_2993, w_012_2994, w_012_2995, w_012_2996, w_012_2997, w_012_2998, w_012_2999, w_012_3000, w_012_3001, w_012_3002, w_012_3003, w_012_3004, w_012_3005, w_012_3006, w_012_3007, w_012_3008, w_012_3009, w_012_3010, w_012_3011, w_012_3012, w_012_3013, w_012_3014, w_012_3015, w_012_3016, w_012_3017, w_012_3018, w_012_3019, w_012_3020, w_012_3021, w_012_3022, w_012_3023, w_012_3024, w_012_3025, w_012_3026, w_012_3027, w_012_3028, w_012_3029, w_012_3030, w_012_3031, w_012_3032, w_012_3033, w_012_3034, w_012_3035, w_012_3036, w_012_3037, w_012_3038, w_012_3039, w_012_3040, w_012_3041, w_012_3042, w_012_3043, w_012_3044, w_012_3045, w_012_3046, w_012_3047, w_012_3048, w_012_3049, w_012_3050, w_012_3051, w_012_3052, w_012_3053, w_012_3054, w_012_3055, w_012_3056, w_012_3057, w_012_3058, w_012_3059, w_012_3060, w_012_3061, w_012_3062, w_012_3063, w_012_3064, w_012_3065, w_012_3066, w_012_3067, w_012_3068, w_012_3069, w_012_3070, w_012_3071, w_012_3072, w_012_3073, w_012_3074, w_012_3075, w_012_3076, w_012_3077, w_012_3078, w_012_3079, w_012_3081, w_012_3082, w_012_3083, w_012_3084, w_012_3085, w_012_3086, w_012_3087, w_012_3088, w_012_3089, w_012_3090, w_012_3091, w_012_3092, w_012_3093, w_012_3094, w_012_3095, w_012_3096, w_012_3097, w_012_3098, w_012_3099, w_012_3100, w_012_3101, w_012_3102, w_012_3103, w_012_3104, w_012_3105, w_012_3106, w_012_3107, w_012_3108, w_012_3109, w_012_3110, w_012_3111, w_012_3112, w_012_3113, w_012_3114, w_012_3115, w_012_3116, w_012_3117, w_012_3118, w_012_3119, w_012_3120, w_012_3121, w_012_3122, w_012_3123, w_012_3124, w_012_3125, w_012_3126, w_012_3127, w_012_3128, w_012_3129, w_012_3130, w_012_3131, w_012_3132, w_012_3133, w_012_3134, w_012_3135, w_012_3136, w_012_3137, w_012_3138, w_012_3139, w_012_3140, w_012_3141, w_012_3142, w_012_3143, w_012_3144, w_012_3145, w_012_3146;
  wire w_013_002, w_013_003, w_013_004, w_013_005, w_013_007, w_013_008, w_013_009, w_013_010, w_013_011, w_013_012, w_013_013, w_013_014, w_013_015, w_013_016, w_013_017, w_013_018, w_013_019, w_013_020, w_013_021, w_013_022, w_013_023, w_013_024, w_013_025, w_013_026, w_013_027, w_013_028, w_013_029, w_013_030, w_013_031, w_013_033, w_013_034, w_013_035, w_013_036, w_013_037, w_013_038, w_013_039, w_013_041, w_013_042, w_013_043, w_013_044, w_013_045, w_013_046, w_013_047, w_013_048, w_013_049, w_013_050, w_013_051, w_013_052, w_013_053, w_013_054, w_013_056, w_013_058, w_013_059, w_013_060, w_013_062, w_013_063, w_013_064, w_013_065, w_013_066, w_013_067, w_013_068, w_013_069, w_013_070, w_013_072, w_013_073, w_013_075, w_013_076, w_013_077, w_013_078, w_013_079, w_013_080, w_013_081, w_013_082, w_013_083, w_013_084, w_013_085, w_013_086, w_013_087, w_013_088, w_013_089, w_013_090, w_013_091, w_013_092, w_013_093, w_013_094, w_013_095, w_013_096, w_013_097, w_013_098, w_013_099, w_013_100, w_013_101, w_013_103, w_013_104, w_013_106, w_013_108, w_013_109, w_013_110, w_013_111, w_013_112, w_013_113, w_013_114, w_013_115, w_013_117, w_013_118, w_013_119, w_013_120, w_013_121, w_013_122, w_013_123, w_013_124, w_013_125, w_013_126, w_013_127, w_013_129, w_013_130, w_013_132, w_013_133, w_013_134, w_013_135, w_013_136, w_013_137, w_013_138, w_013_139, w_013_140, w_013_141, w_013_142, w_013_143, w_013_144, w_013_146, w_013_147, w_013_148, w_013_149, w_013_150, w_013_152, w_013_153, w_013_154, w_013_155, w_013_156, w_013_157, w_013_158, w_013_159, w_013_160, w_013_161, w_013_162, w_013_163, w_013_164, w_013_165, w_013_166, w_013_167, w_013_168, w_013_169, w_013_171, w_013_173, w_013_174, w_013_176, w_013_177, w_013_178, w_013_179, w_013_180, w_013_181, w_013_182, w_013_183, w_013_184, w_013_185, w_013_186, w_013_187, w_013_188, w_013_189, w_013_190, w_013_191, w_013_192, w_013_193, w_013_194, w_013_196, w_013_197, w_013_198, w_013_199, w_013_200, w_013_201, w_013_203, w_013_204, w_013_205, w_013_206, w_013_207, w_013_208, w_013_209, w_013_210, w_013_211, w_013_212, w_013_213, w_013_214, w_013_215, w_013_216, w_013_217, w_013_219, w_013_220, w_013_221, w_013_222, w_013_223, w_013_225, w_013_226, w_013_227, w_013_228, w_013_229, w_013_231, w_013_232, w_013_233, w_013_234, w_013_235, w_013_236, w_013_237, w_013_238, w_013_239, w_013_240, w_013_241, w_013_242, w_013_243, w_013_244, w_013_245, w_013_246, w_013_247, w_013_248, w_013_249, w_013_251, w_013_252, w_013_253, w_013_254, w_013_255, w_013_256, w_013_257, w_013_258, w_013_259, w_013_260, w_013_261, w_013_262, w_013_263, w_013_264, w_013_265, w_013_266, w_013_267, w_013_268, w_013_269, w_013_270, w_013_271, w_013_273, w_013_274, w_013_276, w_013_277, w_013_278, w_013_280, w_013_281, w_013_282, w_013_283, w_013_284, w_013_286, w_013_287, w_013_288, w_013_289, w_013_290, w_013_291, w_013_292, w_013_293, w_013_294, w_013_295, w_013_296, w_013_297, w_013_298, w_013_299, w_013_300, w_013_301, w_013_302, w_013_303, w_013_304, w_013_305, w_013_306, w_013_308, w_013_309, w_013_310, w_013_311, w_013_312, w_013_313, w_013_314, w_013_315, w_013_316, w_013_317, w_013_318, w_013_319, w_013_320, w_013_321, w_013_322, w_013_323, w_013_324, w_013_325, w_013_326, w_013_327, w_013_328, w_013_329, w_013_330, w_013_331, w_013_332, w_013_333, w_013_334, w_013_335, w_013_336, w_013_337, w_013_338, w_013_339, w_013_340, w_013_341, w_013_342, w_013_343, w_013_345, w_013_347, w_013_349, w_013_353, w_013_354, w_013_355, w_013_356, w_013_357, w_013_358, w_013_359, w_013_360, w_013_361, w_013_362, w_013_363, w_013_364, w_013_365, w_013_366, w_013_367, w_013_368, w_013_370, w_013_371, w_013_372, w_013_374, w_013_375, w_013_376, w_013_377, w_013_378, w_013_379, w_013_380, w_013_381, w_013_383, w_013_384, w_013_385, w_013_386, w_013_387, w_013_388, w_013_389, w_013_390, w_013_391, w_013_392, w_013_393, w_013_394, w_013_395, w_013_396, w_013_397, w_013_398, w_013_399, w_013_400, w_013_401, w_013_402, w_013_403, w_013_404, w_013_405, w_013_406, w_013_407, w_013_408, w_013_409, w_013_410, w_013_411, w_013_412, w_013_413, w_013_414, w_013_415, w_013_416, w_013_417, w_013_418, w_013_419, w_013_420, w_013_421, w_013_422, w_013_423, w_013_426, w_013_428, w_013_429, w_013_430, w_013_431, w_013_432, w_013_433, w_013_434, w_013_435, w_013_436, w_013_437, w_013_439, w_013_440, w_013_441, w_013_442, w_013_443, w_013_444, w_013_445, w_013_446, w_013_447, w_013_448, w_013_449, w_013_451, w_013_452, w_013_453, w_013_454, w_013_455, w_013_456, w_013_457, w_013_458, w_013_459, w_013_460, w_013_461, w_013_462, w_013_463, w_013_464, w_013_465, w_013_466, w_013_467, w_013_468, w_013_469, w_013_470, w_013_471, w_013_472, w_013_473, w_013_474, w_013_476, w_013_477, w_013_478, w_013_479, w_013_480, w_013_481, w_013_482, w_013_483, w_013_484, w_013_485, w_013_486, w_013_487, w_013_488, w_013_489, w_013_490, w_013_491, w_013_492, w_013_493, w_013_494, w_013_495, w_013_496, w_013_497, w_013_498, w_013_500, w_013_501, w_013_502, w_013_503, w_013_504, w_013_505, w_013_506, w_013_507, w_013_508, w_013_509, w_013_510, w_013_512, w_013_513, w_013_514, w_013_515, w_013_516, w_013_517, w_013_518, w_013_519, w_013_522, w_013_523, w_013_524, w_013_525, w_013_526, w_013_527, w_013_528, w_013_529, w_013_530, w_013_531, w_013_533, w_013_534, w_013_535, w_013_537, w_013_538, w_013_540, w_013_541, w_013_542, w_013_543, w_013_544, w_013_545, w_013_546, w_013_547, w_013_548, w_013_549, w_013_551, w_013_552, w_013_553, w_013_554, w_013_555, w_013_557, w_013_558, w_013_559, w_013_560, w_013_561, w_013_563, w_013_564, w_013_565, w_013_566, w_013_567, w_013_568, w_013_569, w_013_570, w_013_571, w_013_572, w_013_573, w_013_574, w_013_575, w_013_576, w_013_577, w_013_579, w_013_580, w_013_581, w_013_582, w_013_585, w_013_586, w_013_587, w_013_588, w_013_589, w_013_591, w_013_592, w_013_593, w_013_594, w_013_595, w_013_597, w_013_598, w_013_599, w_013_600, w_013_601, w_013_602, w_013_603, w_013_604, w_013_605, w_013_606, w_013_607, w_013_608, w_013_609, w_013_610, w_013_611, w_013_612, w_013_613, w_013_614, w_013_615, w_013_619, w_013_620, w_013_621, w_013_622, w_013_623, w_013_624, w_013_625, w_013_626, w_013_628, w_013_629, w_013_630, w_013_631, w_013_632, w_013_633, w_013_634, w_013_635, w_013_636, w_013_637, w_013_638, w_013_639, w_013_640, w_013_641, w_013_642, w_013_644, w_013_645, w_013_646, w_013_647, w_013_648, w_013_649, w_013_650, w_013_651, w_013_652, w_013_653, w_013_654, w_013_655, w_013_656, w_013_657, w_013_658, w_013_659, w_013_661, w_013_662, w_013_664, w_013_665, w_013_666, w_013_667, w_013_668, w_013_669, w_013_670, w_013_671, w_013_672, w_013_673, w_013_674, w_013_675, w_013_676, w_013_677, w_013_678, w_013_679, w_013_680, w_013_681, w_013_682, w_013_683, w_013_684, w_013_685, w_013_686, w_013_687, w_013_688, w_013_689, w_013_690, w_013_691, w_013_692, w_013_693, w_013_694, w_013_695, w_013_696, w_013_697, w_013_698, w_013_699, w_013_700, w_013_701, w_013_702, w_013_703, w_013_704, w_013_705, w_013_706, w_013_707, w_013_708, w_013_709, w_013_710, w_013_711, w_013_712, w_013_713, w_013_714, w_013_715, w_013_716, w_013_717, w_013_718, w_013_719, w_013_720, w_013_721, w_013_722, w_013_723, w_013_724, w_013_725, w_013_726, w_013_727, w_013_728, w_013_729, w_013_730, w_013_731, w_013_732, w_013_733, w_013_734, w_013_735, w_013_736, w_013_737, w_013_738, w_013_739, w_013_740, w_013_741, w_013_742, w_013_743, w_013_744, w_013_746, w_013_748, w_013_750, w_013_752, w_013_753, w_013_754, w_013_755, w_013_757, w_013_758, w_013_760, w_013_761, w_013_762, w_013_763, w_013_764, w_013_765, w_013_766, w_013_767, w_013_768, w_013_769, w_013_770, w_013_771, w_013_772, w_013_773, w_013_774, w_013_775, w_013_776, w_013_777, w_013_778, w_013_779, w_013_780, w_013_781, w_013_782, w_013_783, w_013_785, w_013_786, w_013_787, w_013_788, w_013_789, w_013_790, w_013_791, w_013_792, w_013_793, w_013_794, w_013_795, w_013_796, w_013_797, w_013_799, w_013_800, w_013_801, w_013_802, w_013_803, w_013_804, w_013_805, w_013_806, w_013_807, w_013_808, w_013_809, w_013_810, w_013_811, w_013_812, w_013_813, w_013_814, w_013_818, w_013_819, w_013_820, w_013_821, w_013_822, w_013_823, w_013_825, w_013_826, w_013_827, w_013_828, w_013_829, w_013_830, w_013_831, w_013_832, w_013_833, w_013_834, w_013_835, w_013_836, w_013_837, w_013_839, w_013_840, w_013_841, w_013_842, w_013_843, w_013_844, w_013_845, w_013_846, w_013_847, w_013_848, w_013_850, w_013_851, w_013_852, w_013_853, w_013_854, w_013_855, w_013_856, w_013_857, w_013_858, w_013_859, w_013_860, w_013_861, w_013_862, w_013_863, w_013_864, w_013_866, w_013_867, w_013_868, w_013_869, w_013_870, w_013_872, w_013_873, w_013_874, w_013_875, w_013_876, w_013_877, w_013_878, w_013_879, w_013_881, w_013_882, w_013_883, w_013_884, w_013_885, w_013_886, w_013_887, w_013_888, w_013_889, w_013_890, w_013_891, w_013_892, w_013_893, w_013_894, w_013_895, w_013_896, w_013_897, w_013_898, w_013_899, w_013_900, w_013_901, w_013_902, w_013_904, w_013_905, w_013_906, w_013_907, w_013_908, w_013_909, w_013_910, w_013_911, w_013_912, w_013_913, w_013_914, w_013_915, w_013_916, w_013_917, w_013_918, w_013_919, w_013_920, w_013_921, w_013_922, w_013_924, w_013_925, w_013_926, w_013_927, w_013_928, w_013_930, w_013_931, w_013_932, w_013_933, w_013_934, w_013_935, w_013_936, w_013_937, w_013_938, w_013_939, w_013_940, w_013_941, w_013_943, w_013_944, w_013_945, w_013_946, w_013_947, w_013_948, w_013_949, w_013_950, w_013_951, w_013_952, w_013_953, w_013_954, w_013_955, w_013_956, w_013_957, w_013_958, w_013_959, w_013_961, w_013_962, w_013_963, w_013_964, w_013_965, w_013_966, w_013_967, w_013_968, w_013_969, w_013_970, w_013_971, w_013_972, w_013_973, w_013_974, w_013_975, w_013_976, w_013_977, w_013_978, w_013_979, w_013_980, w_013_981, w_013_983, w_013_984, w_013_985, w_013_986, w_013_987, w_013_988, w_013_989, w_013_990, w_013_991, w_013_992, w_013_993, w_013_994, w_013_995, w_013_997, w_013_999, w_013_1000, w_013_1001, w_013_1002, w_013_1003, w_013_1004, w_013_1006, w_013_1007, w_013_1008, w_013_1009, w_013_1010, w_013_1011, w_013_1013, w_013_1014, w_013_1015, w_013_1017, w_013_1018, w_013_1019, w_013_1020, w_013_1022, w_013_1024, w_013_1025, w_013_1027, w_013_1028, w_013_1029, w_013_1030, w_013_1031, w_013_1032, w_013_1033, w_013_1034, w_013_1035, w_013_1036, w_013_1037, w_013_1038, w_013_1039, w_013_1040, w_013_1041, w_013_1042, w_013_1043, w_013_1044, w_013_1045, w_013_1046, w_013_1047, w_013_1048, w_013_1049, w_013_1050, w_013_1051, w_013_1052, w_013_1054, w_013_1057, w_013_1059, w_013_1060, w_013_1061, w_013_1062, w_013_1063, w_013_1064, w_013_1065, w_013_1066, w_013_1067, w_013_1068, w_013_1069, w_013_1071, w_013_1072, w_013_1073, w_013_1075, w_013_1076, w_013_1077, w_013_1078, w_013_1079, w_013_1081, w_013_1082, w_013_1083, w_013_1084, w_013_1085, w_013_1086, w_013_1087, w_013_1088, w_013_1089, w_013_1090, w_013_1092, w_013_1095, w_013_1096, w_013_1097, w_013_1098, w_013_1099, w_013_1100, w_013_1101, w_013_1102, w_013_1103, w_013_1104, w_013_1105, w_013_1106, w_013_1107, w_013_1108, w_013_1109, w_013_1110, w_013_1111, w_013_1112, w_013_1113, w_013_1114, w_013_1115, w_013_1116, w_013_1117, w_013_1118, w_013_1119, w_013_1120, w_013_1121, w_013_1122, w_013_1123, w_013_1124, w_013_1125, w_013_1126, w_013_1127, w_013_1128, w_013_1129, w_013_1130, w_013_1131, w_013_1132, w_013_1134, w_013_1135, w_013_1136, w_013_1137, w_013_1139, w_013_1140, w_013_1141, w_013_1142, w_013_1143, w_013_1144, w_013_1146, w_013_1147, w_013_1148, w_013_1149, w_013_1150, w_013_1151, w_013_1152, w_013_1153, w_013_1154, w_013_1155, w_013_1156, w_013_1157, w_013_1158, w_013_1159, w_013_1160, w_013_1161, w_013_1162, w_013_1163, w_013_1164, w_013_1165, w_013_1166, w_013_1167, w_013_1168, w_013_1169, w_013_1170, w_013_1171, w_013_1172, w_013_1173, w_013_1175, w_013_1176, w_013_1177, w_013_1178, w_013_1179, w_013_1180, w_013_1181, w_013_1182, w_013_1183, w_013_1185, w_013_1186, w_013_1187, w_013_1188, w_013_1189, w_013_1190, w_013_1192, w_013_1193, w_013_1194, w_013_1195, w_013_1197, w_013_1198, w_013_1199, w_013_1200, w_013_1201, w_013_1202, w_013_1203, w_013_1204, w_013_1205, w_013_1206, w_013_1208, w_013_1209, w_013_1210, w_013_1211, w_013_1212, w_013_1213, w_013_1214, w_013_1215, w_013_1216, w_013_1217, w_013_1218, w_013_1219, w_013_1220, w_013_1221, w_013_1222, w_013_1223, w_013_1224, w_013_1225, w_013_1226, w_013_1228, w_013_1229, w_013_1230, w_013_1231, w_013_1232, w_013_1233, w_013_1235, w_013_1236, w_013_1237, w_013_1238, w_013_1239, w_013_1240, w_013_1241, w_013_1242, w_013_1243, w_013_1244, w_013_1245, w_013_1246, w_013_1247, w_013_1248, w_013_1249, w_013_1250, w_013_1251, w_013_1252, w_013_1253, w_013_1254, w_013_1255, w_013_1256, w_013_1257, w_013_1259, w_013_1260, w_013_1261, w_013_1262, w_013_1263, w_013_1265, w_013_1267, w_013_1268, w_013_1269, w_013_1270, w_013_1272, w_013_1273, w_013_1274, w_013_1275, w_013_1276, w_013_1277, w_013_1279, w_013_1280, w_013_1281, w_013_1282, w_013_1283, w_013_1284, w_013_1285, w_013_1286, w_013_1287, w_013_1288, w_013_1289, w_013_1290, w_013_1291, w_013_1292, w_013_1293, w_013_1294, w_013_1295, w_013_1296, w_013_1297, w_013_1298, w_013_1299, w_013_1300, w_013_1301, w_013_1302, w_013_1303, w_013_1304, w_013_1305, w_013_1306, w_013_1307, w_013_1308, w_013_1309, w_013_1310, w_013_1311, w_013_1312, w_013_1313, w_013_1314, w_013_1316, w_013_1317, w_013_1318, w_013_1319, w_013_1321, w_013_1322, w_013_1323, w_013_1324, w_013_1325, w_013_1326, w_013_1328, w_013_1330, w_013_1331, w_013_1332, w_013_1333, w_013_1334, w_013_1335, w_013_1336, w_013_1337, w_013_1338, w_013_1339, w_013_1341, w_013_1342, w_013_1343, w_013_1344, w_013_1345, w_013_1347, w_013_1348, w_013_1349, w_013_1351, w_013_1352, w_013_1353, w_013_1354, w_013_1356, w_013_1357, w_013_1358, w_013_1359, w_013_1361, w_013_1363, w_013_1364, w_013_1365, w_013_1366, w_013_1367, w_013_1368, w_013_1369, w_013_1370, w_013_1371, w_013_1372, w_013_1373, w_013_1374, w_013_1375, w_013_1376, w_013_1377, w_013_1378, w_013_1379, w_013_1380, w_013_1381, w_013_1382, w_013_1383, w_013_1384, w_013_1385, w_013_1386, w_013_1387, w_013_1388, w_013_1389, w_013_1390, w_013_1391, w_013_1392, w_013_1393, w_013_1394, w_013_1395, w_013_1396, w_013_1397, w_013_1399, w_013_1400, w_013_1401, w_013_1402, w_013_1403, w_013_1404, w_013_1405, w_013_1407, w_013_1408, w_013_1409, w_013_1412, w_013_1413, w_013_1414, w_013_1415, w_013_1416, w_013_1417, w_013_1418, w_013_1419, w_013_1420, w_013_1421, w_013_1422, w_013_1423, w_013_1424, w_013_1425, w_013_1426, w_013_1427, w_013_1428, w_013_1429, w_013_1430, w_013_1431, w_013_1432, w_013_1434, w_013_1435, w_013_1436, w_013_1437, w_013_1439, w_013_1441, w_013_1442, w_013_1443, w_013_1444, w_013_1445, w_013_1446, w_013_1447, w_013_1448, w_013_1449, w_013_1450, w_013_1451, w_013_1452, w_013_1453, w_013_1455, w_013_1456, w_013_1457, w_013_1458, w_013_1459, w_013_1460, w_013_1461, w_013_1462, w_013_1463, w_013_1464, w_013_1465, w_013_1466, w_013_1467, w_013_1468, w_013_1469, w_013_1470, w_013_1471, w_013_1472, w_013_1473, w_013_1474, w_013_1476, w_013_1477, w_013_1479, w_013_1480, w_013_1481, w_013_1482, w_013_1483, w_013_1484, w_013_1485, w_013_1486, w_013_1487, w_013_1488, w_013_1489, w_013_1490, w_013_1491, w_013_1492, w_013_1493, w_013_1494, w_013_1495, w_013_1496, w_013_1497, w_013_1498, w_013_1499, w_013_1502, w_013_1503, w_013_1504, w_013_1505, w_013_1508, w_013_1509, w_013_1510, w_013_1511, w_013_1512, w_013_1513, w_013_1514, w_013_1515, w_013_1516, w_013_1518, w_013_1519, w_013_1520, w_013_1521, w_013_1522, w_013_1523, w_013_1524, w_013_1525, w_013_1527, w_013_1528, w_013_1529, w_013_1530, w_013_1531, w_013_1532, w_013_1534, w_013_1535, w_013_1536, w_013_1537, w_013_1538, w_013_1540, w_013_1541, w_013_1542, w_013_1543, w_013_1544, w_013_1545, w_013_1547, w_013_1548, w_013_1549, w_013_1550, w_013_1551, w_013_1552, w_013_1553, w_013_1554, w_013_1555, w_013_1556, w_013_1557, w_013_1558, w_013_1559, w_013_1560, w_013_1561, w_013_1562, w_013_1563, w_013_1564, w_013_1565, w_013_1566, w_013_1567, w_013_1568, w_013_1570, w_013_1571, w_013_1572, w_013_1573, w_013_1574, w_013_1575, w_013_1576, w_013_1577, w_013_1578, w_013_1579, w_013_1580, w_013_1581, w_013_1582, w_013_1583, w_013_1584, w_013_1585, w_013_1586, w_013_1588, w_013_1589, w_013_1590, w_013_1591, w_013_1592, w_013_1593, w_013_1594, w_013_1597, w_013_1598, w_013_1599, w_013_1600, w_013_1601, w_013_1602, w_013_1603, w_013_1604, w_013_1605, w_013_1606, w_013_1607, w_013_1609, w_013_1610, w_013_1611, w_013_1612, w_013_1613, w_013_1614, w_013_1615, w_013_1616, w_013_1617, w_013_1618, w_013_1619, w_013_1620, w_013_1621, w_013_1622, w_013_1623, w_013_1626, w_013_1627, w_013_1628, w_013_1630, w_013_1631, w_013_1632, w_013_1633, w_013_1634, w_013_1635, w_013_1636, w_013_1637, w_013_1638, w_013_1639, w_013_1640, w_013_1641, w_013_1642, w_013_1643, w_013_1644, w_013_1645, w_013_1646, w_013_1647, w_013_1648, w_013_1649, w_013_1650, w_013_1651, w_013_1652, w_013_1654, w_013_1655, w_013_1656, w_013_1657, w_013_1658, w_013_1659, w_013_1660, w_013_1661, w_013_1662, w_013_1663, w_013_1664, w_013_1665, w_013_1666, w_013_1667, w_013_1668, w_013_1669, w_013_1670, w_013_1671, w_013_1672, w_013_1673, w_013_1676, w_013_1677, w_013_1678, w_013_1679, w_013_1680, w_013_1681, w_013_1682, w_013_1683, w_013_1684, w_013_1685, w_013_1686, w_013_1687, w_013_1688, w_013_1689, w_013_1690, w_013_1691, w_013_1692, w_013_1693, w_013_1694, w_013_1695, w_013_1696, w_013_1697, w_013_1698, w_013_1699, w_013_1700, w_013_1701, w_013_1702, w_013_1703, w_013_1705, w_013_1706, w_013_1707, w_013_1708, w_013_1709, w_013_1710, w_013_1711, w_013_1712, w_013_1713, w_013_1714, w_013_1715, w_013_1716, w_013_1717, w_013_1718, w_013_1719, w_013_1720, w_013_1721, w_013_1722, w_013_1723, w_013_1724, w_013_1725, w_013_1726, w_013_1727, w_013_1728, w_013_1729, w_013_1730, w_013_1731, w_013_1732, w_013_1734, w_013_1735, w_013_1736, w_013_1737, w_013_1738, w_013_1739, w_013_1740, w_013_1741, w_013_1742, w_013_1743, w_013_1744, w_013_1745, w_013_1746, w_013_1747, w_013_1748, w_013_1749, w_013_1750, w_013_1751, w_013_1752, w_013_1753, w_013_1754, w_013_1755, w_013_1756, w_013_1757, w_013_1758, w_013_1759, w_013_1760, w_013_1761, w_013_1762, w_013_1763, w_013_1765, w_013_1767, w_013_1768, w_013_1770, w_013_1771, w_013_1772, w_013_1773, w_013_1775, w_013_1776, w_013_1777, w_013_1778, w_013_1779, w_013_1780, w_013_1781, w_013_1782, w_013_1783, w_013_1784, w_013_1785, w_013_1786, w_013_1788, w_013_1789, w_013_1790, w_013_1791, w_013_1792, w_013_1793, w_013_1795, w_013_1796, w_013_1797, w_013_1798, w_013_1799, w_013_1800, w_013_1801, w_013_1802, w_013_1803, w_013_1804, w_013_1806, w_013_1807, w_013_1808, w_013_1809, w_013_1810, w_013_1812, w_013_1813, w_013_1814, w_013_1815, w_013_1816, w_013_1817, w_013_1818, w_013_1819, w_013_1820, w_013_1821, w_013_1822, w_013_1824, w_013_1825, w_013_1826, w_013_1827, w_013_1828, w_013_1829, w_013_1830, w_013_1831, w_013_1832, w_013_1834, w_013_1835, w_013_1837, w_013_1838, w_013_1839, w_013_1840, w_013_1842, w_013_1843, w_013_1844, w_013_1845, w_013_1846, w_013_1847, w_013_1848, w_013_1849, w_013_1850, w_013_1851, w_013_1852, w_013_1855, w_013_1856, w_013_1857, w_013_1858, w_013_1859, w_013_1860, w_013_1861, w_013_1863, w_013_1864, w_013_1865, w_013_1866, w_013_1867, w_013_1868, w_013_1869, w_013_1870, w_013_1871, w_013_1872, w_013_1873, w_013_1874, w_013_1875, w_013_1876, w_013_1878, w_013_1879, w_013_1880, w_013_1881, w_013_1882, w_013_1883, w_013_1884, w_013_1885, w_013_1886, w_013_1887, w_013_1888, w_013_1889, w_013_1890, w_013_1892, w_013_1893, w_013_1895, w_013_1896, w_013_1897, w_013_1898, w_013_1899, w_013_1900, w_013_1902, w_013_1903, w_013_1904, w_013_1905, w_013_1906, w_013_1907, w_013_1908, w_013_1909, w_013_1910, w_013_1911, w_013_1912, w_013_1913, w_013_1915, w_013_1916, w_013_1917, w_013_1918, w_013_1919, w_013_1920, w_013_1921, w_013_1922, w_013_1923, w_013_1924, w_013_1925, w_013_1926, w_013_1927, w_013_1928, w_013_1929, w_013_1930, w_013_1932, w_013_1933, w_013_1935, w_013_1936, w_013_1937, w_013_1938, w_013_1939, w_013_1940, w_013_1941, w_013_1942, w_013_1943, w_013_1944, w_013_1945, w_013_1946, w_013_1947, w_013_1948, w_013_1949, w_013_1950, w_013_1951, w_013_1953, w_013_1954, w_013_1955, w_013_1956, w_013_1957, w_013_1958, w_013_1959, w_013_1960, w_013_1962, w_013_1963, w_013_1964, w_013_1965, w_013_1966, w_013_1967, w_013_1968, w_013_1969, w_013_1970, w_013_1971, w_013_1972, w_013_1973, w_013_1974, w_013_1975, w_013_1976, w_013_1977, w_013_1978, w_013_1979, w_013_1980, w_013_1981, w_013_1983, w_013_1984, w_013_1985, w_013_1986, w_013_1987, w_013_1988, w_013_1989, w_013_1990, w_013_1991, w_013_1992, w_013_1993, w_013_1994, w_013_1995, w_013_1996, w_013_1997, w_013_1998, w_013_1999, w_013_2000, w_013_2001, w_013_2002, w_013_2003, w_013_2004, w_013_2005, w_013_2006, w_013_2007, w_013_2008, w_013_2009, w_013_2010, w_013_2011, w_013_2012, w_013_2013, w_013_2014, w_013_2015, w_013_2016, w_013_2017, w_013_2018, w_013_2020, w_013_2021, w_013_2022, w_013_2023, w_013_2025, w_013_2026, w_013_2027, w_013_2028, w_013_2029, w_013_2030, w_013_2031, w_013_2032, w_013_2033, w_013_2034, w_013_2035, w_013_2036, w_013_2038, w_013_2039, w_013_2040, w_013_2041, w_013_2042, w_013_2043, w_013_2044, w_013_2045, w_013_2046, w_013_2047, w_013_2048, w_013_2049, w_013_2050, w_013_2051, w_013_2052, w_013_2053, w_013_2055, w_013_2056, w_013_2057, w_013_2058, w_013_2060, w_013_2061, w_013_2062, w_013_2063, w_013_2064, w_013_2065, w_013_2066, w_013_2067, w_013_2069, w_013_2070, w_013_2071, w_013_2072, w_013_2074, w_013_2075, w_013_2076, w_013_2077, w_013_2078, w_013_2079, w_013_2080, w_013_2081, w_013_2084, w_013_2085, w_013_2086, w_013_2087, w_013_2088, w_013_2089, w_013_2090, w_013_2092, w_013_2093, w_013_2094, w_013_2095, w_013_2096, w_013_2097, w_013_2098, w_013_2099, w_013_2100, w_013_2101, w_013_2102, w_013_2104, w_013_2105, w_013_2106, w_013_2107, w_013_2108, w_013_2109, w_013_2110, w_013_2111, w_013_2112, w_013_2114, w_013_2115, w_013_2116, w_013_2117, w_013_2118, w_013_2119, w_013_2120, w_013_2121, w_013_2122, w_013_2125, w_013_2126, w_013_2127, w_013_2128, w_013_2130, w_013_2131, w_013_2132, w_013_2133, w_013_2134, w_013_2135, w_013_2136, w_013_2137, w_013_2138, w_013_2139, w_013_2140, w_013_2141, w_013_2142, w_013_2144, w_013_2145, w_013_2146, w_013_2147, w_013_2148, w_013_2151, w_013_2152, w_013_2153, w_013_2155, w_013_2156, w_013_2157, w_013_2158, w_013_2159, w_013_2160, w_013_2161, w_013_2162, w_013_2163, w_013_2164, w_013_2165, w_013_2166, w_013_2168, w_013_2169, w_013_2170, w_013_2171, w_013_2172, w_013_2173, w_013_2174, w_013_2175, w_013_2177, w_013_2178, w_013_2179, w_013_2180, w_013_2181, w_013_2182, w_013_2183, w_013_2184, w_013_2185, w_013_2186, w_013_2187, w_013_2188, w_013_2190, w_013_2191, w_013_2192, w_013_2193, w_013_2194, w_013_2195, w_013_2196, w_013_2197, w_013_2198, w_013_2201, w_013_2202, w_013_2203, w_013_2204, w_013_2205, w_013_2207, w_013_2208, w_013_2209, w_013_2210, w_013_2211, w_013_2212, w_013_2213, w_013_2214, w_013_2215, w_013_2216, w_013_2217, w_013_2218, w_013_2219, w_013_2220, w_013_2221, w_013_2222, w_013_2223, w_013_2224, w_013_2225, w_013_2226, w_013_2227, w_013_2228, w_013_2229, w_013_2230, w_013_2232, w_013_2233, w_013_2234, w_013_2235, w_013_2236, w_013_2237, w_013_2238, w_013_2239, w_013_2241, w_013_2242, w_013_2243, w_013_2244, w_013_2246, w_013_2247, w_013_2248, w_013_2249, w_013_2250, w_013_2251, w_013_2252, w_013_2253, w_013_2254, w_013_2255, w_013_2256, w_013_2257, w_013_2258, w_013_2259, w_013_2260, w_013_2261, w_013_2262, w_013_2263, w_013_2264, w_013_2265, w_013_2266, w_013_2267, w_013_2268, w_013_2269, w_013_2270, w_013_2271, w_013_2272, w_013_2273, w_013_2274, w_013_2275, w_013_2276, w_013_2277, w_013_2278, w_013_2279, w_013_2280, w_013_2281, w_013_2282, w_013_2283, w_013_2284, w_013_2285, w_013_2286, w_013_2287, w_013_2288, w_013_2289, w_013_2291, w_013_2292, w_013_2293, w_013_2294, w_013_2295, w_013_2297, w_013_2298, w_013_2299, w_013_2300, w_013_2301, w_013_2302, w_013_2303, w_013_2304, w_013_2305, w_013_2307, w_013_2308, w_013_2310, w_013_2311, w_013_2312, w_013_2314, w_013_2315, w_013_2316, w_013_2317, w_013_2318, w_013_2319, w_013_2321, w_013_2323, w_013_2324, w_013_2325, w_013_2326, w_013_2327, w_013_2328, w_013_2329, w_013_2330, w_013_2331, w_013_2332, w_013_2333, w_013_2334, w_013_2335, w_013_2336, w_013_2337, w_013_2338, w_013_2339, w_013_2340, w_013_2341, w_013_2342, w_013_2343, w_013_2344, w_013_2345, w_013_2346, w_013_2349, w_013_2350, w_013_2351, w_013_2352, w_013_2353, w_013_2354, w_013_2355, w_013_2356, w_013_2358, w_013_2359, w_013_2360, w_013_2361, w_013_2362, w_013_2363, w_013_2364, w_013_2366, w_013_2367, w_013_2368, w_013_2369, w_013_2371, w_013_2372, w_013_2373, w_013_2374, w_013_2375, w_013_2376, w_013_2377, w_013_2378, w_013_2379, w_013_2380, w_013_2382, w_013_2383, w_013_2385, w_013_2386, w_013_2387, w_013_2389, w_013_2391, w_013_2392, w_013_2393, w_013_2394, w_013_2395, w_013_2397, w_013_2398, w_013_2399, w_013_2400, w_013_2401, w_013_2402, w_013_2403, w_013_2404, w_013_2405, w_013_2406, w_013_2407, w_013_2408, w_013_2409, w_013_2410, w_013_2411, w_013_2412, w_013_2413, w_013_2414, w_013_2415, w_013_2416, w_013_2417, w_013_2418, w_013_2419, w_013_2420, w_013_2421, w_013_2422, w_013_2423, w_013_2424, w_013_2425, w_013_2427, w_013_2428, w_013_2429, w_013_2430, w_013_2431, w_013_2432, w_013_2433, w_013_2434, w_013_2435, w_013_2436, w_013_2437, w_013_2438, w_013_2439, w_013_2440, w_013_2441, w_013_2443, w_013_2444, w_013_2445, w_013_2446, w_013_2447, w_013_2448, w_013_2449, w_013_2450, w_013_2452, w_013_2453, w_013_2454, w_013_2455, w_013_2456, w_013_2457, w_013_2458, w_013_2459, w_013_2460, w_013_2461, w_013_2462, w_013_2463, w_013_2464, w_013_2465, w_013_2466, w_013_2467, w_013_2468, w_013_2469, w_013_2470, w_013_2471, w_013_2472, w_013_2473, w_013_2474, w_013_2475, w_013_2477, w_013_2478, w_013_2479, w_013_2480, w_013_2481, w_013_2482, w_013_2483, w_013_2484, w_013_2485, w_013_2487, w_013_2488, w_013_2490, w_013_2491, w_013_2492, w_013_2493, w_013_2494, w_013_2495, w_013_2496, w_013_2497, w_013_2498, w_013_2499, w_013_2500, w_013_2501, w_013_2503, w_013_2504, w_013_2505, w_013_2506, w_013_2507, w_013_2508, w_013_2509, w_013_2510, w_013_2511, w_013_2512, w_013_2513, w_013_2514, w_013_2515, w_013_2516, w_013_2517, w_013_2518, w_013_2519, w_013_2522, w_013_2523, w_013_2525, w_013_2527, w_013_2528, w_013_2529, w_013_2530, w_013_2531, w_013_2532, w_013_2533, w_013_2534, w_013_2535, w_013_2536, w_013_2537, w_013_2538, w_013_2539, w_013_2540, w_013_2541, w_013_2542, w_013_2543, w_013_2545, w_013_2546, w_013_2547, w_013_2548, w_013_2549, w_013_2550, w_013_2551, w_013_2552, w_013_2553, w_013_2554, w_013_2555, w_013_2556, w_013_2557, w_013_2558, w_013_2559, w_013_2560, w_013_2561, w_013_2562, w_013_2563, w_013_2564, w_013_2565, w_013_2566, w_013_2567, w_013_2569, w_013_2570, w_013_2571, w_013_2572, w_013_2573, w_013_2574, w_013_2575, w_013_2576, w_013_2577, w_013_2578, w_013_2579, w_013_2580, w_013_2581, w_013_2582, w_013_2583, w_013_2584, w_013_2585, w_013_2586, w_013_2587, w_013_2588, w_013_2589, w_013_2590, w_013_2591, w_013_2592, w_013_2593, w_013_2594, w_013_2595, w_013_2596, w_013_2597, w_013_2598, w_013_2599, w_013_2600, w_013_2601, w_013_2602, w_013_2603, w_013_2604, w_013_2606, w_013_2607, w_013_2609, w_013_2610, w_013_2611, w_013_2612, w_013_2613, w_013_2614, w_013_2615, w_013_2616, w_013_2617, w_013_2618, w_013_2619, w_013_2620, w_013_2621, w_013_2622, w_013_2623, w_013_2624, w_013_2626, w_013_2627, w_013_2629, w_013_2631, w_013_2632, w_013_2633, w_013_2634, w_013_2635, w_013_2636, w_013_2637, w_013_2638, w_013_2639, w_013_2640, w_013_2641, w_013_2642, w_013_2643, w_013_2644, w_013_2645, w_013_2646, w_013_2647, w_013_2648, w_013_2649, w_013_2650, w_013_2651, w_013_2652, w_013_2653, w_013_2654, w_013_2655, w_013_2656, w_013_2657, w_013_2658, w_013_2660, w_013_2661, w_013_2662, w_013_2663, w_013_2664, w_013_2666, w_013_2667, w_013_2668, w_013_2670, w_013_2671, w_013_2674, w_013_2675, w_013_2676, w_013_2677, w_013_2679, w_013_2680, w_013_2681, w_013_2682, w_013_2683, w_013_2684, w_013_2685, w_013_2686, w_013_2687, w_013_2688, w_013_2689, w_013_2690, w_013_2691, w_013_2692, w_013_2693, w_013_2695, w_013_2696, w_013_2697, w_013_2698, w_013_2699, w_013_2700, w_013_2701, w_013_2702, w_013_2703, w_013_2704, w_013_2705, w_013_2706, w_013_2707, w_013_2708, w_013_2709, w_013_2710, w_013_2711, w_013_2712, w_013_2713, w_013_2714, w_013_2715, w_013_2716, w_013_2717, w_013_2718, w_013_2719, w_013_2720, w_013_2721, w_013_2723, w_013_2724, w_013_2725, w_013_2726, w_013_2727, w_013_2728, w_013_2730, w_013_2731, w_013_2732, w_013_2733, w_013_2734, w_013_2735, w_013_2736, w_013_2737, w_013_2738, w_013_2739, w_013_2740, w_013_2741, w_013_2742, w_013_2743, w_013_2744, w_013_2745, w_013_2746, w_013_2747, w_013_2748, w_013_2749, w_013_2750, w_013_2752, w_013_2753, w_013_2754, w_013_2755, w_013_2756, w_013_2757, w_013_2758, w_013_2759, w_013_2760, w_013_2761, w_013_2762, w_013_2763, w_013_2764, w_013_2765, w_013_2766, w_013_2767, w_013_2768, w_013_2769, w_013_2770, w_013_2771, w_013_2772, w_013_2773, w_013_2775, w_013_2776, w_013_2777, w_013_2778, w_013_2779, w_013_2780, w_013_2782, w_013_2783, w_013_2784, w_013_2785, w_013_2786, w_013_2787, w_013_2788, w_013_2789, w_013_2790, w_013_2791, w_013_2792, w_013_2793, w_013_2794, w_013_2795, w_013_2796, w_013_2797, w_013_2798, w_013_2799, w_013_2800, w_013_2801, w_013_2802, w_013_2803, w_013_2804, w_013_2805, w_013_2806, w_013_2807, w_013_2808, w_013_2809, w_013_2810, w_013_2811, w_013_2812, w_013_2814, w_013_2815, w_013_2816, w_013_2817, w_013_2818, w_013_2821, w_013_2822, w_013_2823, w_013_2824, w_013_2825, w_013_2826, w_013_2827, w_013_2828, w_013_2830, w_013_2831, w_013_2832, w_013_2833, w_013_2834, w_013_2835, w_013_2836, w_013_2837, w_013_2838, w_013_2839, w_013_2840, w_013_2841, w_013_2842, w_013_2843, w_013_2844, w_013_2845, w_013_2846, w_013_2847, w_013_2848, w_013_2849, w_013_2850, w_013_2851, w_013_2853, w_013_2855, w_013_2856, w_013_2857, w_013_2858, w_013_2859, w_013_2860, w_013_2861, w_013_2862, w_013_2863, w_013_2864, w_013_2865, w_013_2866, w_013_2867, w_013_2869, w_013_2870, w_013_2871, w_013_2872, w_013_2873, w_013_2874, w_013_2875, w_013_2876, w_013_2877, w_013_2878, w_013_2879, w_013_2880, w_013_2881, w_013_2882, w_013_2883, w_013_2884, w_013_2885, w_013_2886, w_013_2887, w_013_2888, w_013_2889, w_013_2890, w_013_2891, w_013_2892, w_013_2893, w_013_2894, w_013_2895, w_013_2896, w_013_2898, w_013_2899, w_013_2900, w_013_2901, w_013_2902, w_013_2903, w_013_2904, w_013_2906, w_013_2907, w_013_2908, w_013_2909, w_013_2910, w_013_2911, w_013_2912, w_013_2913, w_013_2915, w_013_2916, w_013_2917, w_013_2918, w_013_2919, w_013_2920, w_013_2921, w_013_2922, w_013_2923, w_013_2924, w_013_2925, w_013_2926, w_013_2928, w_013_2929, w_013_2931, w_013_2932, w_013_2933, w_013_2934, w_013_2935, w_013_2936, w_013_2938, w_013_2939, w_013_2940, w_013_2941, w_013_2942, w_013_2944, w_013_2945, w_013_2946, w_013_2947, w_013_2948, w_013_2950, w_013_2951, w_013_2952, w_013_2953, w_013_2954, w_013_2955, w_013_2956, w_013_2958, w_013_2959, w_013_2960, w_013_2961, w_013_2962, w_013_2963, w_013_2964, w_013_2965, w_013_2966, w_013_2967, w_013_2968, w_013_2969, w_013_2971, w_013_2972, w_013_2973, w_013_2974, w_013_2975, w_013_2976, w_013_2977, w_013_2978, w_013_2979, w_013_2980, w_013_2982, w_013_2983, w_013_2984, w_013_2985, w_013_2986, w_013_2987, w_013_2988, w_013_2989, w_013_2990, w_013_2991, w_013_2992, w_013_2993, w_013_2994, w_013_2995, w_013_2996, w_013_2997, w_013_2998, w_013_2999, w_013_3000, w_013_3001, w_013_3002, w_013_3003, w_013_3004, w_013_3005, w_013_3006, w_013_3007, w_013_3008, w_013_3009, w_013_3010, w_013_3011, w_013_3013, w_013_3014, w_013_3015, w_013_3016, w_013_3017, w_013_3018, w_013_3020, w_013_3022, w_013_3024, w_013_3025, w_013_3026, w_013_3027, w_013_3029, w_013_3030, w_013_3032, w_013_3033, w_013_3034, w_013_3035, w_013_3036, w_013_3037, w_013_3038, w_013_3039, w_013_3041, w_013_3042, w_013_3043, w_013_3044, w_013_3045, w_013_3046, w_013_3047, w_013_3048, w_013_3049, w_013_3050, w_013_3051, w_013_3052, w_013_3053, w_013_3054, w_013_3056, w_013_3057, w_013_3059, w_013_3060, w_013_3061, w_013_3062, w_013_3063, w_013_3064, w_013_3065, w_013_3067, w_013_3068, w_013_3069, w_013_3070, w_013_3071, w_013_3072, w_013_3073, w_013_3074, w_013_3075, w_013_3076, w_013_3077, w_013_3078, w_013_3079, w_013_3080, w_013_3081, w_013_3083, w_013_3084, w_013_3085, w_013_3086, w_013_3087, w_013_3088, w_013_3089, w_013_3090, w_013_3091, w_013_3092, w_013_3093, w_013_3094, w_013_3095, w_013_3096, w_013_3097, w_013_3098, w_013_3099, w_013_3100, w_013_3101, w_013_3102, w_013_3103, w_013_3104, w_013_3105, w_013_3106, w_013_3107, w_013_3108, w_013_3109, w_013_3110, w_013_3111, w_013_3112, w_013_3113, w_013_3114, w_013_3115, w_013_3116, w_013_3117, w_013_3118, w_013_3119, w_013_3120, w_013_3121, w_013_3122, w_013_3123, w_013_3124, w_013_3125, w_013_3126, w_013_3128, w_013_3129, w_013_3130, w_013_3131, w_013_3132, w_013_3133, w_013_3134, w_013_3135, w_013_3136, w_013_3137, w_013_3138, w_013_3139, w_013_3140, w_013_3141, w_013_3142, w_013_3143, w_013_3144, w_013_3145, w_013_3146, w_013_3147, w_013_3148, w_013_3150, w_013_3151, w_013_3152, w_013_3153, w_013_3154, w_013_3155, w_013_3156, w_013_3157, w_013_3158, w_013_3160, w_013_3161, w_013_3162, w_013_3163, w_013_3164, w_013_3165, w_013_3166, w_013_3167, w_013_3168, w_013_3171, w_013_3172, w_013_3174, w_013_3175, w_013_3176, w_013_3177, w_013_3178, w_013_3179, w_013_3180, w_013_3181, w_013_3182, w_013_3183, w_013_3184, w_013_3185, w_013_3186, w_013_3187, w_013_3188, w_013_3189, w_013_3190, w_013_3191, w_013_3192, w_013_3193, w_013_3194, w_013_3195, w_013_3196, w_013_3197, w_013_3198, w_013_3201, w_013_3202, w_013_3203, w_013_3204, w_013_3205, w_013_3206, w_013_3207, w_013_3208, w_013_3210, w_013_3211, w_013_3213, w_013_3215, w_013_3216, w_013_3217, w_013_3218, w_013_3219, w_013_3221, w_013_3222, w_013_3223, w_013_3224, w_013_3225, w_013_3226, w_013_3227, w_013_3228, w_013_3229, w_013_3230, w_013_3231, w_013_3232, w_013_3233, w_013_3235, w_013_3236, w_013_3237, w_013_3238, w_013_3239, w_013_3240, w_013_3241, w_013_3243, w_013_3244, w_013_3245, w_013_3246, w_013_3247, w_013_3248, w_013_3249, w_013_3250, w_013_3251, w_013_3252, w_013_3253, w_013_3254, w_013_3255, w_013_3256, w_013_3257, w_013_3258, w_013_3259, w_013_3260, w_013_3261, w_013_3262, w_013_3263, w_013_3264, w_013_3265, w_013_3266, w_013_3267, w_013_3268, w_013_3269, w_013_3271, w_013_3272, w_013_3274, w_013_3275, w_013_3276, w_013_3277, w_013_3279, w_013_3280, w_013_3281, w_013_3282, w_013_3283, w_013_3284, w_013_3286, w_013_3288, w_013_3289, w_013_3290, w_013_3291, w_013_3292, w_013_3293, w_013_3294, w_013_3295, w_013_3297, w_013_3298, w_013_3299, w_013_3300, w_013_3301, w_013_3303, w_013_3304, w_013_3305, w_013_3306, w_013_3307, w_013_3309, w_013_3310, w_013_3311, w_013_3312, w_013_3313, w_013_3315, w_013_3316, w_013_3317, w_013_3318, w_013_3319, w_013_3321, w_013_3323, w_013_3324, w_013_3325, w_013_3326, w_013_3327, w_013_3329, w_013_3330, w_013_3331, w_013_3332, w_013_3333, w_013_3334, w_013_3335, w_013_3336, w_013_3337, w_013_3338, w_013_3339, w_013_3340, w_013_3341, w_013_3342, w_013_3343, w_013_3344, w_013_3345, w_013_3346, w_013_3347, w_013_3348, w_013_3349, w_013_3350, w_013_3351, w_013_3352, w_013_3353, w_013_3354, w_013_3355, w_013_3356, w_013_3359, w_013_3360, w_013_3361, w_013_3362, w_013_3363, w_013_3364, w_013_3366, w_013_3367, w_013_3368, w_013_3369, w_013_3370, w_013_3371, w_013_3372, w_013_3373, w_013_3374, w_013_3376, w_013_3377, w_013_3378, w_013_3379, w_013_3380, w_013_3381, w_013_3382, w_013_3383, w_013_3384, w_013_3385, w_013_3386, w_013_3387, w_013_3388, w_013_3389, w_013_3390, w_013_3391, w_013_3392, w_013_3393, w_013_3394, w_013_3395, w_013_3396, w_013_3397, w_013_3398, w_013_3399, w_013_3400, w_013_3401, w_013_3402, w_013_3404, w_013_3405, w_013_3406, w_013_3407, w_013_3408, w_013_3409, w_013_3410, w_013_3411, w_013_3412, w_013_3413, w_013_3414, w_013_3415, w_013_3417, w_013_3418, w_013_3419, w_013_3420, w_013_3421, w_013_3422, w_013_3423, w_013_3424, w_013_3425, w_013_3426, w_013_3427, w_013_3428, w_013_3429, w_013_3430, w_013_3431, w_013_3432, w_013_3433, w_013_3434, w_013_3435, w_013_3436, w_013_3437, w_013_3438, w_013_3439, w_013_3441, w_013_3443, w_013_3444, w_013_3445, w_013_3447, w_013_3448, w_013_3449, w_013_3450, w_013_3451, w_013_3452, w_013_3453, w_013_3454, w_013_3455, w_013_3456, w_013_3457, w_013_3458, w_013_3459, w_013_3460, w_013_3461, w_013_3462, w_013_3463, w_013_3464, w_013_3465, w_013_3466, w_013_3467, w_013_3468, w_013_3469, w_013_3470, w_013_3471, w_013_3472, w_013_3473, w_013_3475, w_013_3476, w_013_3477, w_013_3478, w_013_3479, w_013_3480, w_013_3481, w_013_3483, w_013_3484, w_013_3485, w_013_3486, w_013_3488, w_013_3491, w_013_3492, w_013_3493, w_013_3494, w_013_3495, w_013_3496, w_013_3497, w_013_3498, w_013_3500, w_013_3501, w_013_3502, w_013_3503, w_013_3504, w_013_3505, w_013_3506, w_013_3507, w_013_3509, w_013_3510, w_013_3511, w_013_3512, w_013_3513, w_013_3514, w_013_3515, w_013_3517, w_013_3518, w_013_3519, w_013_3520, w_013_3521, w_013_3522, w_013_3523, w_013_3524, w_013_3525, w_013_3526, w_013_3527, w_013_3528, w_013_3529, w_013_3530, w_013_3531, w_013_3533, w_013_3534, w_013_3535, w_013_3536, w_013_3537, w_013_3538, w_013_3539, w_013_3540, w_013_3541, w_013_3542, w_013_3544, w_013_3545, w_013_3546, w_013_3547, w_013_3548, w_013_3549, w_013_3550, w_013_3551, w_013_3552, w_013_3553, w_013_3554, w_013_3555, w_013_3556, w_013_3557, w_013_3558, w_013_3559, w_013_3560, w_013_3561, w_013_3562, w_013_3563, w_013_3564, w_013_3565, w_013_3566, w_013_3567, w_013_3568, w_013_3569, w_013_3570, w_013_3571, w_013_3572, w_013_3573, w_013_3574, w_013_3575, w_013_3576, w_013_3577, w_013_3578, w_013_3579, w_013_3581, w_013_3582, w_013_3583, w_013_3585, w_013_3586, w_013_3587, w_013_3588, w_013_3589, w_013_3590, w_013_3591, w_013_3592, w_013_3593, w_013_3594, w_013_3595, w_013_3596, w_013_3597, w_013_3598, w_013_3599, w_013_3600, w_013_3601, w_013_3603, w_013_3605, w_013_3606, w_013_3607, w_013_3608, w_013_3609, w_013_3610, w_013_3611, w_013_3612, w_013_3613, w_013_3614, w_013_3616, w_013_3617, w_013_3618, w_013_3619, w_013_3620, w_013_3621, w_013_3622, w_013_3623, w_013_3624, w_013_3625, w_013_3626, w_013_3627, w_013_3628, w_013_3629, w_013_3630, w_013_3631, w_013_3633, w_013_3634, w_013_3635, w_013_3636, w_013_3637, w_013_3638, w_013_3639, w_013_3640, w_013_3641, w_013_3642, w_013_3644, w_013_3645, w_013_3646, w_013_3648, w_013_3649, w_013_3651, w_013_3653, w_013_3654, w_013_3656, w_013_3657, w_013_3658, w_013_3659, w_013_3660, w_013_3661, w_013_3662, w_013_3663, w_013_3664, w_013_3665, w_013_3667, w_013_3668, w_013_3669, w_013_3670, w_013_3671, w_013_3674, w_013_3675, w_013_3676, w_013_3677, w_013_3678, w_013_3679, w_013_3680, w_013_3681, w_013_3683, w_013_3685, w_013_3686, w_013_3687, w_013_3688, w_013_3689, w_013_3690, w_013_3691, w_013_3692, w_013_3693, w_013_3694, w_013_3695, w_013_3696, w_013_3697, w_013_3698, w_013_3699, w_013_3701, w_013_3702, w_013_3703, w_013_3704, w_013_3705, w_013_3706, w_013_3707, w_013_3709, w_013_3710, w_013_3711, w_013_3712, w_013_3713, w_013_3714, w_013_3715, w_013_3716, w_013_3717, w_013_3718, w_013_3719, w_013_3720, w_013_3721, w_013_3722, w_013_3723, w_013_3724, w_013_3725, w_013_3726, w_013_3727, w_013_3728, w_013_3729, w_013_3730, w_013_3731, w_013_3732, w_013_3733, w_013_3734, w_013_3735, w_013_3736, w_013_3737, w_013_3738, w_013_3739, w_013_3740, w_013_3741, w_013_3742, w_013_3743, w_013_3744, w_013_3745, w_013_3746, w_013_3747, w_013_3748, w_013_3750, w_013_3752, w_013_3753, w_013_3754, w_013_3755, w_013_3756, w_013_3757, w_013_3758, w_013_3760, w_013_3762, w_013_3763, w_013_3764, w_013_3765, w_013_3766, w_013_3767, w_013_3768, w_013_3769, w_013_3770, w_013_3771, w_013_3772, w_013_3773, w_013_3774, w_013_3775, w_013_3776, w_013_3777, w_013_3778, w_013_3779, w_013_3780, w_013_3781, w_013_3782, w_013_3783, w_013_3785, w_013_3786, w_013_3788, w_013_3789, w_013_3791, w_013_3792, w_013_3793, w_013_3794, w_013_3795, w_013_3796, w_013_3797, w_013_3798, w_013_3799, w_013_3800, w_013_3801, w_013_3802, w_013_3803, w_013_3804, w_013_3805, w_013_3806, w_013_3808, w_013_3809, w_013_3810, w_013_3811, w_013_3812, w_013_3813, w_013_3814, w_013_3815, w_013_3817, w_013_3818, w_013_3819, w_013_3820, w_013_3821, w_013_3822, w_013_3823, w_013_3824, w_013_3825, w_013_3826, w_013_3827, w_013_3828, w_013_3829, w_013_3831, w_013_3833, w_013_3834, w_013_3835, w_013_3836, w_013_3837, w_013_3838, w_013_3839, w_013_3840, w_013_3841, w_013_3842, w_013_3843, w_013_3844, w_013_3845, w_013_3847, w_013_3848, w_013_3849, w_013_3850, w_013_3851, w_013_3852, w_013_3853, w_013_3854, w_013_3855, w_013_3856, w_013_3857, w_013_3858, w_013_3861, w_013_3862, w_013_3863, w_013_3864, w_013_3866, w_013_3867, w_013_3868, w_013_3869, w_013_3870, w_013_3872, w_013_3873, w_013_3874, w_013_3875, w_013_3876, w_013_3877, w_013_3878, w_013_3879, w_013_3880, w_013_3881, w_013_3883, w_013_3884, w_013_3885, w_013_3886, w_013_3887, w_013_3888, w_013_3889, w_013_3890, w_013_3891, w_013_3892, w_013_3893, w_013_3894, w_013_3895, w_013_3896, w_013_3897, w_013_3898, w_013_3899, w_013_3900, w_013_3901, w_013_3902, w_013_3903, w_013_3904, w_013_3905, w_013_3908, w_013_3909, w_013_3910, w_013_3911, w_013_3912, w_013_3913, w_013_3914, w_013_3915, w_013_3916, w_013_3917, w_013_3918, w_013_3919, w_013_3920, w_013_3921, w_013_3923, w_013_3925, w_013_3926, w_013_3928, w_013_3929, w_013_3930, w_013_3931, w_013_3932, w_013_3933, w_013_3934, w_013_3935, w_013_3936, w_013_3937, w_013_3938, w_013_3939, w_013_3941, w_013_3942, w_013_3944, w_013_3945, w_013_3946, w_013_3947, w_013_3948, w_013_3949, w_013_3950, w_013_3951, w_013_3952, w_013_3953, w_013_3955, w_013_3956, w_013_3957, w_013_3958, w_013_3959, w_013_3960, w_013_3961, w_013_3962, w_013_3964, w_013_3965, w_013_3966, w_013_3967, w_013_3968, w_013_3969, w_013_3970, w_013_3971, w_013_3972, w_013_3973, w_013_3975, w_013_3976, w_013_3977, w_013_3978, w_013_3979, w_013_3980, w_013_3981, w_013_3982, w_013_3983, w_013_3984, w_013_3985, w_013_3986, w_013_3987, w_013_3988, w_013_3989, w_013_3990, w_013_3991, w_013_3992, w_013_3993, w_013_3994, w_013_3995, w_013_3996, w_013_3997, w_013_3998, w_013_3999, w_013_4000, w_013_4001, w_013_4003, w_013_4004, w_013_4005, w_013_4006, w_013_4007, w_013_4008, w_013_4009, w_013_4010, w_013_4011, w_013_4013, w_013_4014, w_013_4015, w_013_4017, w_013_4018, w_013_4020, w_013_4021, w_013_4022, w_013_4023, w_013_4024, w_013_4025, w_013_4026, w_013_4027, w_013_4028, w_013_4029, w_013_4030, w_013_4031, w_013_4032, w_013_4033, w_013_4034, w_013_4035, w_013_4036, w_013_4038, w_013_4039, w_013_4040, w_013_4041, w_013_4042, w_013_4043, w_013_4044, w_013_4045, w_013_4046, w_013_4047, w_013_4048, w_013_4049, w_013_4050, w_013_4051, w_013_4052, w_013_4053, w_013_4054, w_013_4055, w_013_4056, w_013_4057, w_013_4058, w_013_4060, w_013_4061, w_013_4062, w_013_4063, w_013_4065, w_013_4066, w_013_4067, w_013_4069, w_013_4070, w_013_4071, w_013_4072, w_013_4073, w_013_4074, w_013_4075, w_013_4076, w_013_4077, w_013_4079, w_013_4080, w_013_4081, w_013_4082, w_013_4084, w_013_4085, w_013_4086, w_013_4087, w_013_4088, w_013_4089, w_013_4090, w_013_4091, w_013_4092, w_013_4093, w_013_4094, w_013_4095, w_013_4096, w_013_4097, w_013_4098, w_013_4099, w_013_4100, w_013_4101, w_013_4102, w_013_4104, w_013_4105, w_013_4106, w_013_4107, w_013_4109, w_013_4111, w_013_4112, w_013_4114, w_013_4115, w_013_4116, w_013_4117, w_013_4118, w_013_4119, w_013_4120, w_013_4121, w_013_4122, w_013_4123, w_013_4124, w_013_4125, w_013_4126, w_013_4127, w_013_4128, w_013_4130, w_013_4131, w_013_4132, w_013_4133, w_013_4134, w_013_4135, w_013_4136, w_013_4137, w_013_4138, w_013_4139, w_013_4140, w_013_4141, w_013_4142, w_013_4143, w_013_4144, w_013_4145, w_013_4146, w_013_4147, w_013_4148, w_013_4149, w_013_4150, w_013_4151, w_013_4152, w_013_4153, w_013_4154, w_013_4155, w_013_4156, w_013_4157, w_013_4158, w_013_4159, w_013_4160, w_013_4161, w_013_4162, w_013_4163, w_013_4164, w_013_4165, w_013_4166, w_013_4167, w_013_4168, w_013_4169, w_013_4170, w_013_4171, w_013_4172, w_013_4174, w_013_4175, w_013_4176, w_013_4177, w_013_4178, w_013_4179, w_013_4180, w_013_4181, w_013_4182, w_013_4183, w_013_4184, w_013_4185, w_013_4186, w_013_4187, w_013_4188, w_013_4189, w_013_4190, w_013_4191, w_013_4192, w_013_4193, w_013_4194, w_013_4195, w_013_4196, w_013_4197, w_013_4200, w_013_4201, w_013_4202, w_013_4203, w_013_4205, w_013_4206, w_013_4208, w_013_4209, w_013_4210, w_013_4211, w_013_4212, w_013_4213, w_013_4214, w_013_4215, w_013_4218, w_013_4219, w_013_4221, w_013_4222, w_013_4223, w_013_4224, w_013_4225, w_013_4227, w_013_4230, w_013_4233, w_013_4234, w_013_4238, w_013_4240, w_013_4241, w_013_4242, w_013_4243, w_013_4244, w_013_4247, w_013_4248, w_013_4250, w_013_4252, w_013_4253, w_013_4256, w_013_4257, w_013_4258, w_013_4259, w_013_4260, w_013_4261, w_013_4262, w_013_4264, w_013_4265, w_013_4266, w_013_4267, w_013_4268, w_013_4271, w_013_4272, w_013_4273, w_013_4276, w_013_4278, w_013_4279, w_013_4281, w_013_4282, w_013_4284, w_013_4285, w_013_4286, w_013_4288, w_013_4291, w_013_4294, w_013_4295, w_013_4296, w_013_4297, w_013_4298, w_013_4299, w_013_4300, w_013_4301, w_013_4303, w_013_4304, w_013_4307, w_013_4308, w_013_4309, w_013_4310, w_013_4311, w_013_4312, w_013_4314, w_013_4315, w_013_4316, w_013_4318, w_013_4320, w_013_4322, w_013_4324, w_013_4325, w_013_4326, w_013_4327, w_013_4329, w_013_4330, w_013_4331, w_013_4334, w_013_4335, w_013_4336, w_013_4337, w_013_4338, w_013_4339, w_013_4341, w_013_4344, w_013_4345, w_013_4346, w_013_4348, w_013_4349, w_013_4353, w_013_4356, w_013_4358, w_013_4359, w_013_4360, w_013_4361, w_013_4363, w_013_4366, w_013_4368, w_013_4369, w_013_4370, w_013_4371, w_013_4372, w_013_4373, w_013_4375, w_013_4377, w_013_4378, w_013_4379, w_013_4382, w_013_4383, w_013_4385, w_013_4386, w_013_4387, w_013_4388, w_013_4389, w_013_4390, w_013_4391, w_013_4393, w_013_4395, w_013_4396, w_013_4398, w_013_4399, w_013_4401, w_013_4402, w_013_4403, w_013_4404, w_013_4405, w_013_4406, w_013_4407, w_013_4409, w_013_4412, w_013_4413, w_013_4414, w_013_4416, w_013_4418, w_013_4419, w_013_4421, w_013_4422, w_013_4426, w_013_4429, w_013_4430, w_013_4431, w_013_4432, w_013_4433, w_013_4434, w_013_4436, w_013_4437, w_013_4438, w_013_4439, w_013_4440, w_013_4441, w_013_4442, w_013_4443, w_013_4444, w_013_4445, w_013_4446, w_013_4447, w_013_4448, w_013_4449, w_013_4450, w_013_4452, w_013_4454, w_013_4456, w_013_4458, w_013_4460, w_013_4461, w_013_4463, w_013_4464, w_013_4465, w_013_4466, w_013_4468, w_013_4469, w_013_4470, w_013_4471, w_013_4472, w_013_4473, w_013_4476, w_013_4477, w_013_4478, w_013_4480, w_013_4481, w_013_4482, w_013_4484, w_013_4485, w_013_4487, w_013_4488, w_013_4489, w_013_4491, w_013_4492, w_013_4493, w_013_4494, w_013_4495, w_013_4498, w_013_4501, w_013_4503, w_013_4504, w_013_4506, w_013_4507, w_013_4510, w_013_4513, w_013_4514, w_013_4516, w_013_4520, w_013_4521, w_013_4522, w_013_4523, w_013_4524, w_013_4526, w_013_4528, w_013_4529, w_013_4531, w_013_4532, w_013_4533, w_013_4534, w_013_4539, w_013_4540, w_013_4541, w_013_4543, w_013_4544, w_013_4545, w_013_4546, w_013_4549, w_013_4551, w_013_4552, w_013_4553, w_013_4555, w_013_4557, w_013_4558, w_013_4559, w_013_4560, w_013_4562, w_013_4563, w_013_4564, w_013_4565, w_013_4566, w_013_4567, w_013_4571, w_013_4572, w_013_4573, w_013_4574, w_013_4575, w_013_4576, w_013_4577, w_013_4579, w_013_4581, w_013_4582, w_013_4583, w_013_4588, w_013_4589, w_013_4590, w_013_4591, w_013_4592, w_013_4593, w_013_4594, w_013_4595, w_013_4598, w_013_4599, w_013_4600, w_013_4601, w_013_4603, w_013_4604, w_013_4605, w_013_4606, w_013_4609, w_013_4610, w_013_4615, w_013_4616, w_013_4617, w_013_4618, w_013_4619, w_013_4620, w_013_4621, w_013_4623, w_013_4624, w_013_4625, w_013_4626, w_013_4627, w_013_4628, w_013_4629, w_013_4631, w_013_4632, w_013_4633, w_013_4635, w_013_4636, w_013_4637, w_013_4638, w_013_4639, w_013_4641, w_013_4643, w_013_4644, w_013_4646, w_013_4647, w_013_4648, w_013_4650, w_013_4652, w_013_4653, w_013_4654, w_013_4656, w_013_4657, w_013_4658, w_013_4659, w_013_4660, w_013_4661, w_013_4662, w_013_4664, w_013_4665, w_013_4667, w_013_4668, w_013_4669, w_013_4671, w_013_4679, w_013_4682, w_013_4683, w_013_4684, w_013_4685, w_013_4688, w_013_4690, w_013_4691, w_013_4692, w_013_4693, w_013_4695, w_013_4696, w_013_4697, w_013_4702, w_013_4706, w_013_4709, w_013_4710, w_013_4711, w_013_4712, w_013_4713, w_013_4716, w_013_4717, w_013_4718, w_013_4719, w_013_4721, w_013_4722, w_013_4726, w_013_4727, w_013_4728, w_013_4729, w_013_4730, w_013_4731, w_013_4732, w_013_4734, w_013_4735, w_013_4738, w_013_4739, w_013_4740, w_013_4741, w_013_4742, w_013_4743, w_013_4744, w_013_4745, w_013_4746, w_013_4747, w_013_4750, w_013_4753, w_013_4754, w_013_4756, w_013_4757, w_013_4759, w_013_4761, w_013_4762, w_013_4763, w_013_4764, w_013_4765, w_013_4766, w_013_4768, w_013_4770, w_013_4771, w_013_4772, w_013_4773, w_013_4774, w_013_4776, w_013_4777, w_013_4780, w_013_4781, w_013_4782, w_013_4783, w_013_4785, w_013_4787, w_013_4788, w_013_4790, w_013_4791, w_013_4793, w_013_4796, w_013_4797, w_013_4799, w_013_4800, w_013_4803, w_013_4804, w_013_4805, w_013_4806, w_013_4807, w_013_4810, w_013_4811, w_013_4812, w_013_4814, w_013_4817, w_013_4819, w_013_4820, w_013_4821, w_013_4823, w_013_4824, w_013_4825, w_013_4826, w_013_4828, w_013_4830, w_013_4831, w_013_4832, w_013_4834, w_013_4835, w_013_4836, w_013_4838, w_013_4839, w_013_4840, w_013_4842, w_013_4843, w_013_4845, w_013_4847, w_013_4848, w_013_4849, w_013_4850, w_013_4852, w_013_4853, w_013_4855, w_013_4858, w_013_4859, w_013_4860, w_013_4861, w_013_4862, w_013_4863, w_013_4864, w_013_4866, w_013_4867, w_013_4868, w_013_4869, w_013_4874, w_013_4875, w_013_4878, w_013_4879, w_013_4881, w_013_4882, w_013_4883, w_013_4884, w_013_4886, w_013_4887, w_013_4888, w_013_4889, w_013_4890, w_013_4892, w_013_4894, w_013_4895, w_013_4896, w_013_4897, w_013_4898, w_013_4899, w_013_4900, w_013_4901, w_013_4902, w_013_4904, w_013_4905, w_013_4906, w_013_4908, w_013_4909, w_013_4911, w_013_4912, w_013_4913, w_013_4915, w_013_4916, w_013_4918, w_013_4919, w_013_4920, w_013_4921, w_013_4922, w_013_4923, w_013_4926, w_013_4927, w_013_4928, w_013_4929, w_013_4930, w_013_4932, w_013_4934, w_013_4935, w_013_4937, w_013_4939, w_013_4941, w_013_4942, w_013_4943, w_013_4944, w_013_4945, w_013_4947, w_013_4948, w_013_4949, w_013_4950, w_013_4952, w_013_4953, w_013_4955, w_013_4956, w_013_4957, w_013_4958, w_013_4959, w_013_4960, w_013_4961, w_013_4963, w_013_4964, w_013_4966, w_013_4967, w_013_4969, w_013_4970, w_013_4971, w_013_4972, w_013_4973, w_013_4975, w_013_4976, w_013_4977, w_013_4979, w_013_4981, w_013_4982, w_013_4985, w_013_4987, w_013_4988, w_013_4989, w_013_4993, w_013_4994, w_013_4996, w_013_4999, w_013_5000, w_013_5001, w_013_5002, w_013_5004, w_013_5005, w_013_5006, w_013_5007, w_013_5008, w_013_5009, w_013_5010, w_013_5012, w_013_5013, w_013_5014, w_013_5015, w_013_5016, w_013_5017, w_013_5018, w_013_5019, w_013_5020, w_013_5022, w_013_5023, w_013_5024, w_013_5027, w_013_5028, w_013_5029, w_013_5030, w_013_5031, w_013_5034, w_013_5035, w_013_5036, w_013_5037, w_013_5038, w_013_5039, w_013_5040, w_013_5041, w_013_5043, w_013_5044, w_013_5046, w_013_5047, w_013_5049, w_013_5050, w_013_5051, w_013_5055, w_013_5056, w_013_5058, w_013_5060, w_013_5061, w_013_5062, w_013_5064, w_013_5065, w_013_5067, w_013_5068, w_013_5069, w_013_5071, w_013_5072, w_013_5073, w_013_5074, w_013_5076, w_013_5077, w_013_5078, w_013_5079, w_013_5081, w_013_5082, w_013_5083, w_013_5086, w_013_5087, w_013_5088, w_013_5089, w_013_5091, w_013_5092, w_013_5093, w_013_5094, w_013_5095, w_013_5096, w_013_5097, w_013_5098, w_013_5101, w_013_5102, w_013_5104, w_013_5105, w_013_5109, w_013_5110, w_013_5111, w_013_5112, w_013_5113, w_013_5114, w_013_5117, w_013_5118, w_013_5120, w_013_5125, w_013_5127, w_013_5128, w_013_5130, w_013_5131, w_013_5132, w_013_5133, w_013_5134, w_013_5136, w_013_5137, w_013_5140, w_013_5141, w_013_5144, w_013_5145, w_013_5146, w_013_5148, w_013_5149, w_013_5151, w_013_5152, w_013_5153, w_013_5157, w_013_5158, w_013_5159, w_013_5161, w_013_5163, w_013_5164, w_013_5165, w_013_5167, w_013_5169, w_013_5170, w_013_5171, w_013_5172, w_013_5175, w_013_5176, w_013_5177, w_013_5179, w_013_5180, w_013_5181, w_013_5183, w_013_5184, w_013_5185, w_013_5186, w_013_5187, w_013_5188, w_013_5190, w_013_5191, w_013_5192, w_013_5194, w_013_5195, w_013_5197, w_013_5198, w_013_5199, w_013_5200, w_013_5201, w_013_5203, w_013_5204, w_013_5205, w_013_5207, w_013_5208, w_013_5209, w_013_5211, w_013_5212, w_013_5213, w_013_5215, w_013_5217, w_013_5218, w_013_5219, w_013_5220, w_013_5221, w_013_5222, w_013_5224, w_013_5228, w_013_5229, w_013_5231, w_013_5232, w_013_5233, w_013_5234, w_013_5235, w_013_5236, w_013_5237, w_013_5238, w_013_5239, w_013_5242, w_013_5244, w_013_5247, w_013_5249, w_013_5250, w_013_5251, w_013_5254, w_013_5255, w_013_5258, w_013_5260, w_013_5261, w_013_5263, w_013_5264, w_013_5265, w_013_5266, w_013_5267, w_013_5268, w_013_5270, w_013_5271, w_013_5272, w_013_5274, w_013_5275, w_013_5276, w_013_5278, w_013_5279, w_013_5280, w_013_5281, w_013_5282, w_013_5284, w_013_5285, w_013_5286, w_013_5287, w_013_5289, w_013_5290, w_013_5291, w_013_5292, w_013_5293, w_013_5295, w_013_5296, w_013_5297, w_013_5299, w_013_5300, w_013_5303, w_013_5305, w_013_5306, w_013_5307, w_013_5309, w_013_5312, w_013_5315, w_013_5316, w_013_5317, w_013_5318, w_013_5323, w_013_5324, w_013_5326, w_013_5328, w_013_5329, w_013_5330, w_013_5333, w_013_5334, w_013_5335, w_013_5336, w_013_5339, w_013_5340, w_013_5342, w_013_5345, w_013_5346, w_013_5347, w_013_5348, w_013_5349, w_013_5350, w_013_5351, w_013_5352, w_013_5353, w_013_5354, w_013_5355, w_013_5361, w_013_5363, w_013_5364, w_013_5365, w_013_5366, w_013_5368, w_013_5369, w_013_5370, w_013_5373, w_013_5375, w_013_5376, w_013_5379, w_013_5380, w_013_5381, w_013_5383, w_013_5385, w_013_5386, w_013_5387, w_013_5388, w_013_5389, w_013_5392, w_013_5393, w_013_5395, w_013_5396, w_013_5397, w_013_5398, w_013_5400, w_013_5401, w_013_5402, w_013_5403, w_013_5404, w_013_5405, w_013_5406, w_013_5407, w_013_5408, w_013_5410, w_013_5414, w_013_5416, w_013_5417, w_013_5418, w_013_5419, w_013_5420, w_013_5421, w_013_5422, w_013_5423, w_013_5426, w_013_5427, w_013_5429, w_013_5430, w_013_5432, w_013_5433, w_013_5434, w_013_5435, w_013_5436, w_013_5437, w_013_5438, w_013_5439, w_013_5440, w_013_5441, w_013_5443, w_013_5444, w_013_5446, w_013_5448, w_013_5449, w_013_5450, w_013_5451, w_013_5452, w_013_5453, w_013_5454, w_013_5456, w_013_5457, w_013_5458, w_013_5459, w_013_5460, w_013_5461, w_013_5464, w_013_5465, w_013_5466, w_013_5467, w_013_5468, w_013_5469, w_013_5471, w_013_5472, w_013_5474, w_013_5475, w_013_5476, w_013_5478, w_013_5479, w_013_5480, w_013_5481, w_013_5482, w_013_5483, w_013_5485, w_013_5486, w_013_5487, w_013_5489, w_013_5490, w_013_5491, w_013_5492, w_013_5494, w_013_5496, w_013_5498, w_013_5499, w_013_5500, w_013_5501, w_013_5502, w_013_5503, w_013_5504, w_013_5505, w_013_5507, w_013_5508, w_013_5509, w_013_5510, w_013_5511, w_013_5512, w_013_5514, w_013_5515, w_013_5516, w_013_5517, w_013_5518, w_013_5519, w_013_5520, w_013_5521, w_013_5522, w_013_5523, w_013_5524, w_013_5525, w_013_5526, w_013_5527, w_013_5528, w_013_5529, w_013_5531, w_013_5532, w_013_5534, w_013_5537, w_013_5538, w_013_5539, w_013_5540, w_013_5543, w_013_5544, w_013_5546, w_013_5547, w_013_5549, w_013_5551, w_013_5552, w_013_5553, w_013_5554, w_013_5555, w_013_5556, w_013_5557, w_013_5558, w_013_5559, w_013_5562, w_013_5563, w_013_5566, w_013_5567, w_013_5568, w_013_5569, w_013_5571, w_013_5572, w_013_5575, w_013_5577, w_013_5578, w_013_5580, w_013_5581, w_013_5582, w_013_5583, w_013_5585, w_013_5588, w_013_5589, w_013_5590, w_013_5592, w_013_5593, w_013_5594, w_013_5595, w_013_5596, w_013_5597, w_013_5598, w_013_5599, w_013_5600, w_013_5601, w_013_5602, w_013_5603, w_013_5604, w_013_5606, w_013_5607, w_013_5608, w_013_5609, w_013_5611, w_013_5612, w_013_5613, w_013_5614, w_013_5617, w_013_5619, w_013_5620, w_013_5621, w_013_5622, w_013_5623, w_013_5624, w_013_5626, w_013_5627, w_013_5628, w_013_5629, w_013_5631, w_013_5632, w_013_5634, w_013_5636, w_013_5637, w_013_5638, w_013_5639, w_013_5641, w_013_5644, w_013_5645, w_013_5647, w_013_5648, w_013_5652, w_013_5653, w_013_5654, w_013_5656, w_013_5658, w_013_5659, w_013_5661, w_013_5662, w_013_5664, w_013_5665, w_013_5666, w_013_5667, w_013_5668, w_013_5670, w_013_5671, w_013_5672, w_013_5673, w_013_5674, w_013_5675, w_013_5676, w_013_5677, w_013_5678, w_013_5681, w_013_5682, w_013_5683, w_013_5684, w_013_5685, w_013_5686, w_013_5687, w_013_5688, w_013_5692, w_013_5693, w_013_5694, w_013_5696, w_013_5698, w_013_5700, w_013_5701, w_013_5704, w_013_5705, w_013_5707, w_013_5708, w_013_5709, w_013_5710, w_013_5712, w_013_5713, w_013_5715, w_013_5719, w_013_5722, w_013_5724, w_013_5726, w_013_5727, w_013_5728, w_013_5729, w_013_5731, w_013_5732, w_013_5733, w_013_5735, w_013_5736, w_013_5737, w_013_5739, w_013_5741, w_013_5742, w_013_5743, w_013_5744, w_013_5747, w_013_5748, w_013_5749, w_013_5750, w_013_5752, w_013_5754, w_013_5755, w_013_5756, w_013_5757, w_013_5759, w_013_5760, w_013_5761, w_013_5762, w_013_5763, w_013_5764, w_013_5765, w_013_5767, w_013_5768, w_013_5769, w_013_5772, w_013_5773, w_013_5774, w_013_5775, w_013_5776, w_013_5778, w_013_5779, w_013_5780, w_013_5781, w_013_5783;
  wire w_014_000, w_014_001, w_014_002, w_014_003, w_014_004, w_014_005, w_014_006, w_014_007, w_014_008, w_014_009, w_014_010, w_014_011, w_014_012, w_014_013, w_014_014, w_014_015, w_014_016, w_014_017, w_014_018, w_014_019, w_014_020, w_014_021, w_014_022, w_014_023, w_014_024, w_014_025, w_014_026, w_014_027, w_014_028, w_014_029, w_014_030, w_014_031, w_014_032, w_014_033, w_014_034, w_014_035, w_014_036, w_014_037, w_014_038, w_014_039, w_014_040, w_014_041, w_014_042, w_014_043, w_014_044, w_014_045, w_014_046, w_014_047, w_014_048, w_014_049, w_014_050, w_014_051, w_014_052, w_014_053, w_014_054, w_014_055, w_014_056, w_014_057, w_014_058, w_014_059, w_014_060, w_014_061, w_014_062, w_014_063, w_014_064, w_014_065, w_014_066, w_014_067, w_014_068, w_014_069, w_014_070, w_014_071, w_014_072, w_014_073, w_014_074, w_014_075, w_014_076, w_014_077, w_014_078, w_014_079, w_014_080, w_014_081, w_014_082, w_014_083, w_014_084, w_014_085, w_014_086, w_014_087, w_014_088, w_014_089, w_014_090, w_014_091, w_014_092, w_014_093, w_014_094, w_014_095, w_014_096, w_014_097, w_014_098, w_014_099, w_014_100, w_014_101, w_014_102, w_014_103, w_014_104, w_014_105, w_014_106, w_014_107, w_014_108, w_014_109, w_014_110, w_014_111, w_014_112, w_014_113, w_014_114, w_014_115, w_014_116, w_014_117, w_014_118, w_014_119, w_014_120, w_014_121, w_014_122, w_014_123, w_014_124, w_014_125, w_014_126, w_014_127, w_014_128, w_014_129, w_014_130, w_014_131, w_014_132, w_014_133, w_014_134, w_014_135, w_014_136, w_014_137, w_014_138, w_014_139, w_014_140, w_014_141, w_014_142, w_014_143, w_014_144, w_014_145, w_014_146, w_014_147, w_014_148, w_014_149, w_014_150, w_014_151, w_014_152, w_014_153, w_014_154, w_014_155, w_014_156, w_014_157, w_014_158, w_014_159, w_014_160, w_014_161, w_014_162, w_014_163, w_014_164, w_014_165, w_014_166, w_014_167, w_014_168, w_014_169, w_014_170, w_014_171, w_014_172, w_014_173, w_014_174, w_014_175, w_014_176, w_014_177, w_014_178, w_014_179, w_014_180, w_014_181, w_014_182, w_014_183, w_014_184, w_014_185, w_014_186, w_014_187, w_014_188, w_014_189, w_014_190, w_014_191, w_014_192, w_014_193, w_014_194, w_014_195, w_014_196, w_014_197, w_014_198, w_014_199, w_014_200, w_014_201, w_014_202, w_014_203, w_014_204, w_014_205, w_014_206, w_014_207, w_014_208, w_014_209, w_014_210, w_014_211, w_014_212, w_014_213, w_014_214, w_014_215, w_014_216, w_014_217, w_014_218, w_014_219, w_014_220, w_014_221, w_014_222, w_014_223, w_014_224, w_014_225, w_014_226, w_014_227, w_014_228, w_014_229, w_014_230, w_014_231, w_014_232, w_014_233, w_014_234, w_014_235, w_014_236, w_014_237, w_014_238, w_014_239, w_014_240, w_014_241, w_014_242, w_014_243, w_014_244, w_014_245, w_014_246, w_014_247, w_014_248, w_014_249, w_014_250, w_014_251, w_014_252, w_014_253, w_014_254, w_014_255, w_014_256, w_014_257, w_014_258, w_014_259, w_014_260, w_014_261, w_014_262, w_014_263, w_014_264, w_014_265, w_014_266, w_014_267, w_014_268, w_014_269, w_014_270, w_014_271, w_014_272, w_014_273, w_014_274, w_014_275, w_014_276, w_014_277, w_014_278, w_014_279, w_014_280, w_014_281, w_014_282, w_014_283, w_014_284, w_014_285, w_014_286, w_014_287, w_014_288, w_014_289, w_014_290, w_014_291, w_014_292, w_014_293, w_014_294, w_014_295, w_014_296, w_014_297, w_014_298, w_014_299, w_014_300, w_014_301, w_014_302, w_014_303, w_014_304, w_014_305, w_014_306, w_014_307, w_014_308, w_014_309, w_014_310, w_014_311, w_014_312, w_014_313, w_014_314, w_014_315, w_014_316, w_014_317, w_014_318, w_014_319, w_014_320, w_014_321, w_014_322, w_014_323, w_014_324, w_014_325, w_014_326, w_014_327, w_014_328, w_014_329, w_014_330, w_014_331, w_014_332, w_014_333, w_014_334, w_014_335, w_014_336, w_014_337, w_014_338, w_014_339, w_014_340, w_014_341, w_014_342, w_014_343, w_014_344, w_014_345, w_014_346, w_014_347, w_014_348, w_014_349, w_014_350, w_014_351, w_014_352, w_014_353, w_014_354, w_014_355, w_014_356, w_014_357, w_014_358, w_014_359, w_014_360, w_014_361, w_014_362, w_014_363, w_014_364, w_014_365, w_014_366, w_014_367, w_014_368, w_014_369, w_014_370, w_014_371, w_014_372, w_014_373, w_014_374, w_014_375, w_014_376, w_014_377, w_014_378, w_014_379, w_014_380, w_014_381, w_014_382, w_014_383, w_014_384, w_014_385, w_014_386, w_014_387, w_014_388, w_014_389, w_014_390, w_014_391, w_014_392, w_014_393, w_014_394, w_014_395, w_014_396, w_014_397, w_014_398, w_014_399, w_014_400, w_014_401, w_014_402, w_014_403, w_014_404, w_014_405, w_014_406, w_014_407, w_014_408, w_014_409, w_014_410, w_014_411, w_014_412, w_014_413, w_014_414, w_014_415, w_014_416, w_014_417, w_014_418, w_014_419, w_014_420, w_014_421, w_014_422, w_014_423, w_014_424, w_014_425, w_014_426, w_014_427, w_014_428, w_014_429, w_014_430, w_014_431, w_014_432, w_014_433, w_014_434, w_014_435, w_014_436, w_014_437, w_014_438, w_014_439, w_014_440, w_014_441, w_014_442, w_014_443, w_014_444, w_014_445, w_014_446, w_014_447, w_014_448, w_014_449, w_014_450, w_014_451, w_014_452, w_014_453;
  wire w_015_000, w_015_001, w_015_002, w_015_003, w_015_005, w_015_007, w_015_008, w_015_010, w_015_011, w_015_012, w_015_013, w_015_014, w_015_015, w_015_016, w_015_017, w_015_018, w_015_019, w_015_020, w_015_021, w_015_022, w_015_024, w_015_025, w_015_026, w_015_027, w_015_028, w_015_029, w_015_030, w_015_031, w_015_032, w_015_033, w_015_034, w_015_035, w_015_036, w_015_037, w_015_038, w_015_039, w_015_040, w_015_041, w_015_043, w_015_045, w_015_046, w_015_047, w_015_048, w_015_049, w_015_050, w_015_051, w_015_052, w_015_053, w_015_054, w_015_055, w_015_056, w_015_057, w_015_059, w_015_060, w_015_061, w_015_062, w_015_063, w_015_065, w_015_066, w_015_067, w_015_068, w_015_070, w_015_071, w_015_072, w_015_073, w_015_074, w_015_075, w_015_076, w_015_077, w_015_078, w_015_079, w_015_080, w_015_081, w_015_082, w_015_083, w_015_085, w_015_086, w_015_087, w_015_089, w_015_090, w_015_091, w_015_092, w_015_093, w_015_094, w_015_095, w_015_096, w_015_097, w_015_098, w_015_099, w_015_100, w_015_101, w_015_102, w_015_103, w_015_104, w_015_105, w_015_106, w_015_107, w_015_108, w_015_109, w_015_110, w_015_112, w_015_114, w_015_115, w_015_116, w_015_117, w_015_119, w_015_121, w_015_123, w_015_124, w_015_125, w_015_126, w_015_127, w_015_128, w_015_130, w_015_131, w_015_132, w_015_134, w_015_135, w_015_136, w_015_137, w_015_138, w_015_139, w_015_140, w_015_142, w_015_143, w_015_145, w_015_146, w_015_147, w_015_148, w_015_150, w_015_151, w_015_152, w_015_153, w_015_154, w_015_155, w_015_156, w_015_158, w_015_159, w_015_160, w_015_162, w_015_163, w_015_164, w_015_165, w_015_166, w_015_167, w_015_168, w_015_169, w_015_170, w_015_171, w_015_172, w_015_173, w_015_175, w_015_176, w_015_177, w_015_178, w_015_180, w_015_181, w_015_182, w_015_183, w_015_184, w_015_185, w_015_186, w_015_187, w_015_188, w_015_189, w_015_190, w_015_191, w_015_192, w_015_193, w_015_194, w_015_195, w_015_196, w_015_197, w_015_198, w_015_199, w_015_200, w_015_202, w_015_203, w_015_206, w_015_207, w_015_208, w_015_209, w_015_210, w_015_211, w_015_212, w_015_213, w_015_215, w_015_216, w_015_217, w_015_218, w_015_219, w_015_220, w_015_224, w_015_225, w_015_226, w_015_227, w_015_228, w_015_229, w_015_231, w_015_232, w_015_234, w_015_235, w_015_236, w_015_237, w_015_238, w_015_239, w_015_240, w_015_241, w_015_242, w_015_243, w_015_244, w_015_245, w_015_246, w_015_247, w_015_248, w_015_249, w_015_250, w_015_251, w_015_252, w_015_253, w_015_254, w_015_255, w_015_256, w_015_258, w_015_259, w_015_261, w_015_262, w_015_263, w_015_264, w_015_265, w_015_266, w_015_267, w_015_268, w_015_270, w_015_271, w_015_272, w_015_273, w_015_274, w_015_275, w_015_276, w_015_277, w_015_278, w_015_279, w_015_280, w_015_281, w_015_282, w_015_283, w_015_284, w_015_285, w_015_286, w_015_287, w_015_289, w_015_290, w_015_291, w_015_292, w_015_293, w_015_294, w_015_295, w_015_296, w_015_297, w_015_298, w_015_299, w_015_300, w_015_301, w_015_302, w_015_303, w_015_304, w_015_305, w_015_306, w_015_307, w_015_308, w_015_309, w_015_310, w_015_311, w_015_312, w_015_313, w_015_314, w_015_315, w_015_317, w_015_318, w_015_319, w_015_320, w_015_321, w_015_322, w_015_323, w_015_324, w_015_325, w_015_326, w_015_327, w_015_328, w_015_329, w_015_330, w_015_331, w_015_332, w_015_333, w_015_334, w_015_335, w_015_336, w_015_337, w_015_338, w_015_339, w_015_340, w_015_341, w_015_342, w_015_343, w_015_344, w_015_345, w_015_346, w_015_347, w_015_348, w_015_349, w_015_350, w_015_351, w_015_353, w_015_354, w_015_356, w_015_357, w_015_358, w_015_359, w_015_360, w_015_361, w_015_362, w_015_364, w_015_365, w_015_366, w_015_367, w_015_368, w_015_369, w_015_370, w_015_371, w_015_372, w_015_373, w_015_374, w_015_375, w_015_376, w_015_377, w_015_379, w_015_380, w_015_381, w_015_382, w_015_383, w_015_384, w_015_385, w_015_386, w_015_387, w_015_388, w_015_389, w_015_391, w_015_393, w_015_394, w_015_395, w_015_396, w_015_397, w_015_398, w_015_399, w_015_400, w_015_401, w_015_402, w_015_403, w_015_404, w_015_405, w_015_407, w_015_408, w_015_409, w_015_410, w_015_411, w_015_412, w_015_413, w_015_414, w_015_415, w_015_416, w_015_417, w_015_419, w_015_420, w_015_421, w_015_423, w_015_424, w_015_425, w_015_426, w_015_427, w_015_428, w_015_429, w_015_430, w_015_431, w_015_432, w_015_433, w_015_434, w_015_435, w_015_436, w_015_438, w_015_439, w_015_440, w_015_441, w_015_442, w_015_443, w_015_444, w_015_445, w_015_446, w_015_447, w_015_448, w_015_449, w_015_450, w_015_451, w_015_452, w_015_454, w_015_456, w_015_457, w_015_458, w_015_459, w_015_460, w_015_462, w_015_463, w_015_464, w_015_465, w_015_466, w_015_467, w_015_468, w_015_469, w_015_470, w_015_471, w_015_472, w_015_473, w_015_474, w_015_475, w_015_476, w_015_477, w_015_478, w_015_479, w_015_480, w_015_481, w_015_482, w_015_483, w_015_484, w_015_485, w_015_487, w_015_488, w_015_489, w_015_490, w_015_491, w_015_492, w_015_493, w_015_494, w_015_495, w_015_496, w_015_497, w_015_498, w_015_500, w_015_501, w_015_502, w_015_504, w_015_505, w_015_506, w_015_507, w_015_508, w_015_509, w_015_510, w_015_511, w_015_512, w_015_513, w_015_514, w_015_515, w_015_517, w_015_518, w_015_520, w_015_521, w_015_522, w_015_523, w_015_524, w_015_525, w_015_526, w_015_527, w_015_528, w_015_529, w_015_530, w_015_531, w_015_532, w_015_533, w_015_534, w_015_536, w_015_537, w_015_538, w_015_539, w_015_540, w_015_541, w_015_542, w_015_543, w_015_544, w_015_545, w_015_546, w_015_547, w_015_548, w_015_549, w_015_550, w_015_551, w_015_552, w_015_553, w_015_554, w_015_555, w_015_556, w_015_557, w_015_558, w_015_559, w_015_560, w_015_561, w_015_562, w_015_563, w_015_564, w_015_565, w_015_566, w_015_567, w_015_568, w_015_569, w_015_570, w_015_571, w_015_572, w_015_573, w_015_574, w_015_576, w_015_577, w_015_578, w_015_579, w_015_580, w_015_581, w_015_582, w_015_583, w_015_584, w_015_585, w_015_586, w_015_587, w_015_588, w_015_590, w_015_591, w_015_592, w_015_593, w_015_594, w_015_595, w_015_596, w_015_597, w_015_598, w_015_599, w_015_600, w_015_601, w_015_602, w_015_603, w_015_604, w_015_605, w_015_606, w_015_607, w_015_608, w_015_609, w_015_611, w_015_612, w_015_614, w_015_616, w_015_617, w_015_618, w_015_619, w_015_621, w_015_622, w_015_623, w_015_624, w_015_625, w_015_626, w_015_628, w_015_629, w_015_630, w_015_631, w_015_632, w_015_633, w_015_634, w_015_636, w_015_637, w_015_638, w_015_640, w_015_641, w_015_642, w_015_643, w_015_644, w_015_645, w_015_646, w_015_647, w_015_648, w_015_649, w_015_650, w_015_651, w_015_652, w_015_654, w_015_655, w_015_657, w_015_658, w_015_659, w_015_660, w_015_662, w_015_664, w_015_665, w_015_666, w_015_667, w_015_668, w_015_669, w_015_670, w_015_671, w_015_672, w_015_673, w_015_674, w_015_675, w_015_676, w_015_677, w_015_678, w_015_679, w_015_680, w_015_681, w_015_682, w_015_683, w_015_684, w_015_685, w_015_687, w_015_688, w_015_689, w_015_690, w_015_691, w_015_692, w_015_693, w_015_694, w_015_695, w_015_696, w_015_697, w_015_698, w_015_699, w_015_700, w_015_701, w_015_702, w_015_703, w_015_705, w_015_706, w_015_708, w_015_709, w_015_710, w_015_711, w_015_712, w_015_713, w_015_714, w_015_715, w_015_716, w_015_717, w_015_718, w_015_719, w_015_720, w_015_721, w_015_722, w_015_723, w_015_724, w_015_727, w_015_728, w_015_729, w_015_730, w_015_731, w_015_732, w_015_734, w_015_735, w_015_736, w_015_737, w_015_738, w_015_739, w_015_740, w_015_741, w_015_742, w_015_743, w_015_744, w_015_745, w_015_747, w_015_748, w_015_749, w_015_750, w_015_751, w_015_752, w_015_753, w_015_754, w_015_755, w_015_756, w_015_757, w_015_758, w_015_759, w_015_760, w_015_761, w_015_762, w_015_763, w_015_764, w_015_765, w_015_766, w_015_767, w_015_769, w_015_770, w_015_771, w_015_772, w_015_773, w_015_774, w_015_776, w_015_777, w_015_778, w_015_779, w_015_780, w_015_781, w_015_782, w_015_783, w_015_784, w_015_785, w_015_787, w_015_788, w_015_789, w_015_790, w_015_791, w_015_792, w_015_793, w_015_794, w_015_795, w_015_796, w_015_797, w_015_798, w_015_799, w_015_800, w_015_801, w_015_802, w_015_803, w_015_804, w_015_805, w_015_806, w_015_807, w_015_808, w_015_810, w_015_811, w_015_812, w_015_813, w_015_814, w_015_815, w_015_816, w_015_817, w_015_818, w_015_819, w_015_820, w_015_821, w_015_823, w_015_824, w_015_825, w_015_826, w_015_827, w_015_828, w_015_829, w_015_830, w_015_831, w_015_832, w_015_833, w_015_834, w_015_835, w_015_836, w_015_837, w_015_838, w_015_839, w_015_840, w_015_841, w_015_842, w_015_845, w_015_847, w_015_848, w_015_849, w_015_851, w_015_852, w_015_853, w_015_854, w_015_855, w_015_856, w_015_857, w_015_858, w_015_859, w_015_860, w_015_862, w_015_863, w_015_864, w_015_865, w_015_866, w_015_867, w_015_868, w_015_869, w_015_870, w_015_871, w_015_872, w_015_873, w_015_875, w_015_876, w_015_877, w_015_878, w_015_879, w_015_880, w_015_881, w_015_882, w_015_884, w_015_885, w_015_886, w_015_888, w_015_889, w_015_890, w_015_891, w_015_893, w_015_894, w_015_895, w_015_897, w_015_898, w_015_899, w_015_900, w_015_901, w_015_902, w_015_904, w_015_905, w_015_906, w_015_907, w_015_908, w_015_909, w_015_910, w_015_911, w_015_912, w_015_913, w_015_914, w_015_915, w_015_916, w_015_917, w_015_918, w_015_919, w_015_920, w_015_921, w_015_922, w_015_923, w_015_924, w_015_925, w_015_926, w_015_927, w_015_928, w_015_929, w_015_930, w_015_931, w_015_932, w_015_933, w_015_934, w_015_935, w_015_936, w_015_937, w_015_938, w_015_939, w_015_940, w_015_941, w_015_942, w_015_943, w_015_944, w_015_945, w_015_946, w_015_947, w_015_948, w_015_949, w_015_950, w_015_951, w_015_952, w_015_953, w_015_954, w_015_955, w_015_956, w_015_957, w_015_958, w_015_959, w_015_960, w_015_961, w_015_962, w_015_963, w_015_964, w_015_965, w_015_966, w_015_967, w_015_969, w_015_970, w_015_971, w_015_972, w_015_974, w_015_976, w_015_977, w_015_978, w_015_979, w_015_980, w_015_982, w_015_984, w_015_985, w_015_986, w_015_987, w_015_988, w_015_989, w_015_990, w_015_991, w_015_992, w_015_993, w_015_994, w_015_995, w_015_996, w_015_997, w_015_999, w_015_1000, w_015_1001, w_015_1002, w_015_1003, w_015_1004, w_015_1005, w_015_1006, w_015_1009, w_015_1010, w_015_1011, w_015_1012, w_015_1014, w_015_1015, w_015_1016, w_015_1017, w_015_1018, w_015_1019, w_015_1020, w_015_1021, w_015_1022, w_015_1023, w_015_1024, w_015_1025, w_015_1026, w_015_1028, w_015_1029, w_015_1030, w_015_1032, w_015_1033, w_015_1034, w_015_1035, w_015_1036, w_015_1037, w_015_1038, w_015_1039, w_015_1040, w_015_1042, w_015_1043, w_015_1044, w_015_1045, w_015_1046, w_015_1047, w_015_1048, w_015_1049, w_015_1050, w_015_1051, w_015_1052, w_015_1054, w_015_1055, w_015_1056, w_015_1057, w_015_1058, w_015_1059, w_015_1060, w_015_1061, w_015_1063, w_015_1064, w_015_1065, w_015_1066, w_015_1067, w_015_1068, w_015_1071, w_015_1072, w_015_1073, w_015_1075, w_015_1076, w_015_1077, w_015_1078, w_015_1079, w_015_1080, w_015_1081, w_015_1082, w_015_1084, w_015_1085, w_015_1086, w_015_1087, w_015_1088, w_015_1089, w_015_1090, w_015_1091, w_015_1092, w_015_1093, w_015_1094, w_015_1095, w_015_1096, w_015_1097, w_015_1098, w_015_1099, w_015_1100, w_015_1101, w_015_1102, w_015_1103, w_015_1104, w_015_1105, w_015_1106, w_015_1107, w_015_1108, w_015_1109, w_015_1110, w_015_1111, w_015_1112, w_015_1113, w_015_1114, w_015_1115, w_015_1116, w_015_1118, w_015_1119, w_015_1120, w_015_1121, w_015_1122, w_015_1123, w_015_1124, w_015_1125, w_015_1126, w_015_1127, w_015_1129, w_015_1130, w_015_1131, w_015_1132, w_015_1133, w_015_1134, w_015_1135, w_015_1136, w_015_1137, w_015_1139, w_015_1141, w_015_1142, w_015_1143, w_015_1144, w_015_1145, w_015_1146, w_015_1147, w_015_1148, w_015_1149, w_015_1151, w_015_1152, w_015_1153, w_015_1154, w_015_1157, w_015_1160, w_015_1161, w_015_1162, w_015_1164, w_015_1165, w_015_1166, w_015_1167, w_015_1168, w_015_1169, w_015_1170, w_015_1171, w_015_1172, w_015_1173, w_015_1174, w_015_1175, w_015_1176, w_015_1177, w_015_1178, w_015_1179, w_015_1180, w_015_1181, w_015_1183, w_015_1184, w_015_1185, w_015_1186, w_015_1187, w_015_1188, w_015_1189, w_015_1190, w_015_1191, w_015_1192, w_015_1194, w_015_1195, w_015_1196, w_015_1197, w_015_1198, w_015_1199, w_015_1200, w_015_1201, w_015_1202, w_015_1203, w_015_1204, w_015_1205, w_015_1206, w_015_1207, w_015_1208, w_015_1209, w_015_1210, w_015_1212, w_015_1213, w_015_1214, w_015_1215, w_015_1216, w_015_1217, w_015_1219, w_015_1220, w_015_1221, w_015_1224, w_015_1225, w_015_1227, w_015_1228, w_015_1229, w_015_1230, w_015_1231, w_015_1232, w_015_1233, w_015_1236, w_015_1237, w_015_1238, w_015_1239, w_015_1240, w_015_1241, w_015_1242, w_015_1243, w_015_1244, w_015_1245, w_015_1246, w_015_1247, w_015_1249, w_015_1250, w_015_1251, w_015_1252, w_015_1253, w_015_1254, w_015_1255, w_015_1256, w_015_1257, w_015_1258, w_015_1259, w_015_1261, w_015_1262, w_015_1263, w_015_1264, w_015_1266, w_015_1267, w_015_1268, w_015_1269, w_015_1270, w_015_1271, w_015_1272, w_015_1273, w_015_1274, w_015_1275, w_015_1276, w_015_1277, w_015_1279, w_015_1280, w_015_1281, w_015_1282, w_015_1283, w_015_1284, w_015_1285, w_015_1287, w_015_1288, w_015_1289, w_015_1290, w_015_1291, w_015_1292, w_015_1293, w_015_1294, w_015_1295, w_015_1296, w_015_1297, w_015_1298, w_015_1299, w_015_1300, w_015_1301, w_015_1302, w_015_1303, w_015_1304, w_015_1305, w_015_1306, w_015_1307, w_015_1308, w_015_1309, w_015_1310, w_015_1312, w_015_1313, w_015_1314, w_015_1315, w_015_1316, w_015_1317, w_015_1318, w_015_1319, w_015_1320, w_015_1321, w_015_1322, w_015_1323, w_015_1324, w_015_1325, w_015_1326, w_015_1327, w_015_1328, w_015_1330, w_015_1331, w_015_1332, w_015_1333, w_015_1334, w_015_1335, w_015_1336, w_015_1337, w_015_1338, w_015_1339, w_015_1340, w_015_1341, w_015_1342, w_015_1343, w_015_1344, w_015_1345, w_015_1346, w_015_1348, w_015_1349, w_015_1350, w_015_1352, w_015_1353, w_015_1354, w_015_1355, w_015_1357, w_015_1358, w_015_1359, w_015_1360, w_015_1361, w_015_1362, w_015_1363, w_015_1364, w_015_1366, w_015_1369, w_015_1370, w_015_1371, w_015_1372, w_015_1373, w_015_1375, w_015_1376, w_015_1377, w_015_1379, w_015_1380, w_015_1381, w_015_1382, w_015_1383, w_015_1384, w_015_1385, w_015_1386, w_015_1387, w_015_1388, w_015_1389, w_015_1390, w_015_1391, w_015_1392, w_015_1394, w_015_1395, w_015_1396, w_015_1397, w_015_1398, w_015_1400, w_015_1401, w_015_1402, w_015_1403, w_015_1404, w_015_1406, w_015_1407, w_015_1409, w_015_1410, w_015_1411, w_015_1412, w_015_1413, w_015_1414, w_015_1415, w_015_1416, w_015_1417, w_015_1418, w_015_1419, w_015_1420, w_015_1421, w_015_1422, w_015_1423, w_015_1424, w_015_1425, w_015_1426, w_015_1427, w_015_1428, w_015_1429, w_015_1430, w_015_1431, w_015_1432, w_015_1433, w_015_1434, w_015_1435, w_015_1436, w_015_1437, w_015_1438, w_015_1440, w_015_1441, w_015_1443, w_015_1444, w_015_1445, w_015_1446, w_015_1447, w_015_1448, w_015_1449, w_015_1451, w_015_1452, w_015_1453, w_015_1454, w_015_1455, w_015_1456, w_015_1457, w_015_1458, w_015_1459, w_015_1460, w_015_1461, w_015_1462, w_015_1464, w_015_1465, w_015_1466, w_015_1467, w_015_1468, w_015_1469, w_015_1470, w_015_1471, w_015_1472, w_015_1474, w_015_1476, w_015_1477, w_015_1478, w_015_1479, w_015_1480, w_015_1481, w_015_1482, w_015_1483, w_015_1484, w_015_1485, w_015_1486, w_015_1487, w_015_1488, w_015_1489, w_015_1490, w_015_1491, w_015_1492, w_015_1494, w_015_1496, w_015_1497, w_015_1499, w_015_1501, w_015_1502, w_015_1503, w_015_1504, w_015_1506, w_015_1508, w_015_1509, w_015_1510, w_015_1511, w_015_1512, w_015_1513, w_015_1514, w_015_1515, w_015_1516, w_015_1517, w_015_1518, w_015_1519, w_015_1520, w_015_1521, w_015_1522, w_015_1523, w_015_1524, w_015_1525, w_015_1526, w_015_1527, w_015_1528, w_015_1529, w_015_1530, w_015_1531, w_015_1532, w_015_1533, w_015_1534, w_015_1535, w_015_1536, w_015_1537, w_015_1539, w_015_1540, w_015_1541, w_015_1542, w_015_1543, w_015_1544, w_015_1545, w_015_1546, w_015_1547, w_015_1549, w_015_1550, w_015_1551, w_015_1552, w_015_1553, w_015_1554, w_015_1555, w_015_1556, w_015_1557, w_015_1558, w_015_1559, w_015_1560, w_015_1561, w_015_1563, w_015_1564, w_015_1566, w_015_1567, w_015_1568, w_015_1569, w_015_1570, w_015_1572, w_015_1574, w_015_1575, w_015_1576, w_015_1578, w_015_1579, w_015_1580, w_015_1581, w_015_1582, w_015_1583, w_015_1584, w_015_1585, w_015_1586, w_015_1587, w_015_1588, w_015_1589, w_015_1590, w_015_1591, w_015_1592, w_015_1594, w_015_1595, w_015_1596, w_015_1597, w_015_1598, w_015_1599, w_015_1600, w_015_1602, w_015_1603, w_015_1605, w_015_1606, w_015_1607, w_015_1608, w_015_1609, w_015_1610, w_015_1611, w_015_1612, w_015_1613, w_015_1614, w_015_1615, w_015_1616, w_015_1617, w_015_1618, w_015_1619, w_015_1620, w_015_1621, w_015_1622, w_015_1624, w_015_1625, w_015_1626, w_015_1627, w_015_1628, w_015_1629, w_015_1630, w_015_1632, w_015_1633, w_015_1634, w_015_1635, w_015_1636, w_015_1637, w_015_1638, w_015_1639, w_015_1640, w_015_1641, w_015_1642, w_015_1643, w_015_1644, w_015_1645, w_015_1646, w_015_1647, w_015_1648, w_015_1649, w_015_1650, w_015_1651, w_015_1652, w_015_1653, w_015_1654, w_015_1655, w_015_1656, w_015_1657, w_015_1658, w_015_1659, w_015_1660, w_015_1662, w_015_1663, w_015_1664, w_015_1665, w_015_1666, w_015_1667, w_015_1668, w_015_1669, w_015_1670, w_015_1671, w_015_1672, w_015_1673, w_015_1674, w_015_1675, w_015_1676, w_015_1677, w_015_1678, w_015_1679, w_015_1680, w_015_1682, w_015_1683, w_015_1684, w_015_1685, w_015_1686, w_015_1687, w_015_1688, w_015_1689, w_015_1690, w_015_1692, w_015_1693, w_015_1694, w_015_1695, w_015_1696, w_015_1697, w_015_1698, w_015_1699, w_015_1700, w_015_1701, w_015_1704, w_015_1705, w_015_1706, w_015_1707, w_015_1708, w_015_1709, w_015_1710, w_015_1712, w_015_1713, w_015_1714, w_015_1716, w_015_1717, w_015_1718, w_015_1719, w_015_1720, w_015_1721, w_015_1722, w_015_1723, w_015_1724, w_015_1725, w_015_1726, w_015_1727, w_015_1728, w_015_1729, w_015_1730, w_015_1731, w_015_1732, w_015_1733, w_015_1734, w_015_1735, w_015_1736, w_015_1737, w_015_1740, w_015_1741, w_015_1742, w_015_1743, w_015_1744, w_015_1745, w_015_1747, w_015_1748, w_015_1749, w_015_1750, w_015_1751, w_015_1752, w_015_1753, w_015_1754, w_015_1755, w_015_1757, w_015_1758, w_015_1759, w_015_1760, w_015_1761, w_015_1762, w_015_1764, w_015_1766, w_015_1768, w_015_1769, w_015_1770, w_015_1771, w_015_1772, w_015_1773, w_015_1774, w_015_1775, w_015_1776, w_015_1777, w_015_1778, w_015_1779, w_015_1780, w_015_1781, w_015_1782, w_015_1783, w_015_1784, w_015_1786, w_015_1787, w_015_1788, w_015_1789, w_015_1790, w_015_1791, w_015_1792, w_015_1793, w_015_1794, w_015_1796, w_015_1798, w_015_1799, w_015_1800, w_015_1802, w_015_1803, w_015_1805, w_015_1806, w_015_1807, w_015_1808, w_015_1809, w_015_1810, w_015_1811, w_015_1812, w_015_1813, w_015_1814, w_015_1816, w_015_1817, w_015_1818, w_015_1819, w_015_1820, w_015_1821, w_015_1822, w_015_1823, w_015_1824, w_015_1825, w_015_1826, w_015_1827, w_015_1828, w_015_1829, w_015_1830, w_015_1831, w_015_1832, w_015_1833, w_015_1834, w_015_1835, w_015_1836, w_015_1837, w_015_1838, w_015_1839, w_015_1840, w_015_1841, w_015_1842, w_015_1843, w_015_1844, w_015_1845, w_015_1846, w_015_1847, w_015_1849, w_015_1850, w_015_1851, w_015_1852, w_015_1854, w_015_1855, w_015_1856, w_015_1857, w_015_1858, w_015_1859, w_015_1860, w_015_1861, w_015_1862, w_015_1864, w_015_1865, w_015_1866, w_015_1868, w_015_1869, w_015_1870, w_015_1871, w_015_1873, w_015_1874, w_015_1875, w_015_1876, w_015_1877, w_015_1878, w_015_1879, w_015_1880, w_015_1881, w_015_1882, w_015_1883, w_015_1884, w_015_1885, w_015_1886, w_015_1887, w_015_1888, w_015_1889, w_015_1890, w_015_1891, w_015_1892, w_015_1893, w_015_1894, w_015_1895, w_015_1896, w_015_1897, w_015_1898, w_015_1899, w_015_1900, w_015_1901, w_015_1902, w_015_1903, w_015_1904, w_015_1905, w_015_1906, w_015_1907, w_015_1908, w_015_1909, w_015_1911, w_015_1912, w_015_1913, w_015_1914, w_015_1915, w_015_1916, w_015_1917, w_015_1918, w_015_1919, w_015_1920, w_015_1921, w_015_1922, w_015_1923, w_015_1924, w_015_1925, w_015_1926, w_015_1927, w_015_1930, w_015_1931, w_015_1933, w_015_1934, w_015_1935, w_015_1936, w_015_1938, w_015_1939, w_015_1940, w_015_1941, w_015_1942, w_015_1943, w_015_1944, w_015_1945, w_015_1946, w_015_1948, w_015_1949, w_015_1950, w_015_1951, w_015_1952, w_015_1953, w_015_1954, w_015_1955, w_015_1956, w_015_1957, w_015_1958, w_015_1959, w_015_1960, w_015_1961, w_015_1962, w_015_1963, w_015_1964, w_015_1965, w_015_1966, w_015_1967, w_015_1968, w_015_1969, w_015_1970, w_015_1972, w_015_1973, w_015_1974, w_015_1975, w_015_1976, w_015_1978, w_015_1979, w_015_1980, w_015_1982, w_015_1983, w_015_1985, w_015_1986, w_015_1987, w_015_1988, w_015_1989, w_015_1991, w_015_1992, w_015_1993, w_015_1994, w_015_1995, w_015_1996, w_015_1997, w_015_1998, w_015_1999, w_015_2000, w_015_2001, w_015_2002, w_015_2003, w_015_2004, w_015_2005, w_015_2008, w_015_2009, w_015_2010, w_015_2011, w_015_2012, w_015_2013, w_015_2014, w_015_2015, w_015_2016, w_015_2017, w_015_2018, w_015_2019, w_015_2020, w_015_2021, w_015_2022, w_015_2023, w_015_2024, w_015_2025, w_015_2026, w_015_2027, w_015_2028, w_015_2029, w_015_2030, w_015_2031, w_015_2032, w_015_2033, w_015_2034, w_015_2035, w_015_2036, w_015_2037, w_015_2039, w_015_2040, w_015_2042, w_015_2043, w_015_2044, w_015_2045, w_015_2046, w_015_2047, w_015_2048, w_015_2049, w_015_2050, w_015_2051, w_015_2053, w_015_2054, w_015_2055, w_015_2056, w_015_2057, w_015_2059, w_015_2060, w_015_2061, w_015_2062, w_015_2063, w_015_2064, w_015_2065, w_015_2066, w_015_2067, w_015_2068, w_015_2070, w_015_2071, w_015_2072, w_015_2073, w_015_2075, w_015_2076, w_015_2077, w_015_2079, w_015_2080, w_015_2082, w_015_2083, w_015_2084, w_015_2085, w_015_2086, w_015_2087, w_015_2088, w_015_2089, w_015_2091, w_015_2092, w_015_2093, w_015_2094, w_015_2095, w_015_2096, w_015_2097, w_015_2098, w_015_2099, w_015_2100, w_015_2101, w_015_2102, w_015_2103, w_015_2104, w_015_2105, w_015_2106, w_015_2107, w_015_2108, w_015_2110, w_015_2111, w_015_2112, w_015_2113, w_015_2114, w_015_2115, w_015_2116, w_015_2117, w_015_2118, w_015_2119, w_015_2120, w_015_2121, w_015_2122, w_015_2123, w_015_2126, w_015_2127, w_015_2128, w_015_2129, w_015_2130, w_015_2131, w_015_2132, w_015_2133, w_015_2134, w_015_2135, w_015_2136, w_015_2138, w_015_2139, w_015_2140, w_015_2141, w_015_2142, w_015_2143, w_015_2144, w_015_2145, w_015_2146, w_015_2147, w_015_2148, w_015_2149, w_015_2151, w_015_2152, w_015_2153, w_015_2154, w_015_2155, w_015_2157, w_015_2158, w_015_2159, w_015_2160, w_015_2161, w_015_2162, w_015_2163, w_015_2164, w_015_2165, w_015_2166, w_015_2167, w_015_2168, w_015_2169, w_015_2170, w_015_2171, w_015_2172, w_015_2173, w_015_2174, w_015_2175, w_015_2176, w_015_2177, w_015_2178, w_015_2179, w_015_2180, w_015_2181, w_015_2182, w_015_2183, w_015_2184, w_015_2185, w_015_2186, w_015_2187, w_015_2188, w_015_2190, w_015_2191, w_015_2192, w_015_2193, w_015_2195, w_015_2196, w_015_2197, w_015_2198, w_015_2199, w_015_2200, w_015_2201, w_015_2202, w_015_2203, w_015_2204, w_015_2206, w_015_2207, w_015_2208, w_015_2209, w_015_2210, w_015_2211, w_015_2212, w_015_2213, w_015_2214, w_015_2216, w_015_2217, w_015_2218, w_015_2219, w_015_2220, w_015_2221, w_015_2222, w_015_2223, w_015_2224, w_015_2225, w_015_2226, w_015_2227, w_015_2228, w_015_2229, w_015_2230, w_015_2231, w_015_2233, w_015_2234, w_015_2235, w_015_2236, w_015_2237, w_015_2238, w_015_2239, w_015_2240, w_015_2241, w_015_2244, w_015_2245, w_015_2246, w_015_2247, w_015_2248, w_015_2249, w_015_2250, w_015_2252, w_015_2253, w_015_2255, w_015_2256, w_015_2257, w_015_2258, w_015_2259, w_015_2260, w_015_2261, w_015_2262, w_015_2263, w_015_2264, w_015_2266, w_015_2267, w_015_2268, w_015_2270, w_015_2271, w_015_2272, w_015_2273, w_015_2274, w_015_2275, w_015_2276, w_015_2277, w_015_2278, w_015_2279, w_015_2282, w_015_2283, w_015_2284, w_015_2285, w_015_2286, w_015_2287, w_015_2288, w_015_2289, w_015_2290, w_015_2291, w_015_2292, w_015_2293, w_015_2294, w_015_2295, w_015_2296, w_015_2297, w_015_2299, w_015_2300, w_015_2301, w_015_2303, w_015_2304, w_015_2305, w_015_2306, w_015_2307, w_015_2308, w_015_2310, w_015_2311, w_015_2312, w_015_2313, w_015_2314, w_015_2315, w_015_2316, w_015_2317, w_015_2318, w_015_2321, w_015_2323, w_015_2324, w_015_2325, w_015_2326, w_015_2327, w_015_2328, w_015_2329, w_015_2330, w_015_2331, w_015_2333, w_015_2334, w_015_2335, w_015_2336, w_015_2337, w_015_2338, w_015_2340, w_015_2341, w_015_2342, w_015_2343, w_015_2344, w_015_2345, w_015_2347, w_015_2348, w_015_2349, w_015_2350, w_015_2351, w_015_2352, w_015_2353, w_015_2354, w_015_2355, w_015_2356, w_015_2357, w_015_2358, w_015_2359, w_015_2360, w_015_2361, w_015_2362, w_015_2363, w_015_2364, w_015_2365, w_015_2366, w_015_2367, w_015_2368, w_015_2369, w_015_2370, w_015_2371, w_015_2372, w_015_2375, w_015_2376, w_015_2377, w_015_2378, w_015_2379, w_015_2380, w_015_2382, w_015_2383, w_015_2384, w_015_2385, w_015_2386, w_015_2387, w_015_2388, w_015_2389, w_015_2390, w_015_2391, w_015_2392, w_015_2393, w_015_2394, w_015_2395, w_015_2398, w_015_2399, w_015_2400, w_015_2401, w_015_2402, w_015_2403, w_015_2404, w_015_2405, w_015_2407, w_015_2408, w_015_2409, w_015_2410, w_015_2411, w_015_2413, w_015_2414, w_015_2415, w_015_2416, w_015_2417, w_015_2418, w_015_2419, w_015_2420, w_015_2422, w_015_2423, w_015_2424, w_015_2425, w_015_2426, w_015_2427, w_015_2428, w_015_2429, w_015_2430, w_015_2431, w_015_2432, w_015_2433, w_015_2434, w_015_2435, w_015_2436, w_015_2438, w_015_2439, w_015_2440, w_015_2441, w_015_2442, w_015_2443, w_015_2444, w_015_2445, w_015_2446, w_015_2448, w_015_2449, w_015_2450, w_015_2451, w_015_2452, w_015_2453, w_015_2454, w_015_2455, w_015_2456, w_015_2457, w_015_2458, w_015_2459, w_015_2460, w_015_2461, w_015_2462, w_015_2463, w_015_2464, w_015_2466, w_015_2467, w_015_2469, w_015_2471, w_015_2473, w_015_2474, w_015_2475, w_015_2476, w_015_2477, w_015_2478, w_015_2479, w_015_2480, w_015_2481, w_015_2482, w_015_2484, w_015_2485, w_015_2486, w_015_2487, w_015_2488, w_015_2489, w_015_2490, w_015_2491, w_015_2492, w_015_2493, w_015_2494, w_015_2495, w_015_2496, w_015_2497, w_015_2498, w_015_2499, w_015_2500, w_015_2501, w_015_2502, w_015_2503, w_015_2504, w_015_2505, w_015_2506, w_015_2509, w_015_2510, w_015_2512, w_015_2513, w_015_2514, w_015_2515, w_015_2516, w_015_2517, w_015_2519, w_015_2520, w_015_2521, w_015_2522, w_015_2523, w_015_2525, w_015_2526, w_015_2527, w_015_2528, w_015_2529, w_015_2530, w_015_2531, w_015_2533, w_015_2534, w_015_2535, w_015_2536, w_015_2537, w_015_2538, w_015_2539, w_015_2540, w_015_2541, w_015_2542, w_015_2543, w_015_2544, w_015_2545, w_015_2546, w_015_2547, w_015_2548, w_015_2549, w_015_2550, w_015_2551, w_015_2552, w_015_2553, w_015_2554, w_015_2555, w_015_2556, w_015_2557, w_015_2558, w_015_2559, w_015_2560, w_015_2562, w_015_2563, w_015_2564, w_015_2565, w_015_2566, w_015_2567, w_015_2568, w_015_2569, w_015_2570, w_015_2571, w_015_2572, w_015_2573, w_015_2574, w_015_2575, w_015_2576, w_015_2577, w_015_2578, w_015_2579, w_015_2580, w_015_2581, w_015_2582, w_015_2583, w_015_2584, w_015_2585, w_015_2586, w_015_2587, w_015_2588, w_015_2589, w_015_2590, w_015_2591, w_015_2592, w_015_2593, w_015_2595, w_015_2596, w_015_2597, w_015_2598, w_015_2599, w_015_2600, w_015_2601, w_015_2602, w_015_2603, w_015_2604, w_015_2605, w_015_2606, w_015_2607, w_015_2608, w_015_2609, w_015_2610, w_015_2611, w_015_2612, w_015_2613, w_015_2614, w_015_2615, w_015_2616, w_015_2617, w_015_2619, w_015_2620, w_015_2621, w_015_2622, w_015_2623, w_015_2624, w_015_2625, w_015_2626, w_015_2627, w_015_2629, w_015_2630, w_015_2631, w_015_2632, w_015_2634, w_015_2635, w_015_2636, w_015_2637, w_015_2638, w_015_2639, w_015_2640, w_015_2641, w_015_2642, w_015_2644, w_015_2645, w_015_2646, w_015_2647, w_015_2648, w_015_2649, w_015_2650, w_015_2651, w_015_2652, w_015_2653, w_015_2654, w_015_2655, w_015_2656, w_015_2658, w_015_2659, w_015_2660, w_015_2661, w_015_2662, w_015_2663, w_015_2665, w_015_2666, w_015_2669, w_015_2670, w_015_2671, w_015_2673, w_015_2674, w_015_2675, w_015_2676, w_015_2677, w_015_2679, w_015_2680, w_015_2682, w_015_2683, w_015_2684, w_015_2685, w_015_2686, w_015_2687, w_015_2688, w_015_2689, w_015_2690, w_015_2691, w_015_2692, w_015_2693, w_015_2694, w_015_2695, w_015_2696, w_015_2697, w_015_2698, w_015_2699, w_015_2700, w_015_2701, w_015_2702, w_015_2703, w_015_2704, w_015_2706, w_015_2707, w_015_2708, w_015_2709, w_015_2710, w_015_2711, w_015_2712, w_015_2713, w_015_2714, w_015_2715, w_015_2716, w_015_2717, w_015_2718, w_015_2719, w_015_2720, w_015_2721, w_015_2722, w_015_2723, w_015_2724, w_015_2725, w_015_2726, w_015_2727, w_015_2728, w_015_2729, w_015_2730, w_015_2731, w_015_2732, w_015_2733, w_015_2734, w_015_2736, w_015_2737, w_015_2738, w_015_2739, w_015_2740, w_015_2741, w_015_2743, w_015_2745, w_015_2746, w_015_2747, w_015_2748, w_015_2749, w_015_2751, w_015_2752, w_015_2753, w_015_2754, w_015_2755, w_015_2756, w_015_2757, w_015_2758, w_015_2759, w_015_2760, w_015_2762, w_015_2763, w_015_2765, w_015_2767, w_015_2768, w_015_2769, w_015_2770, w_015_2771, w_015_2772, w_015_2773, w_015_2774, w_015_2775, w_015_2776, w_015_2777, w_015_2778, w_015_2779, w_015_2780, w_015_2781, w_015_2782, w_015_2783, w_015_2786, w_015_2787, w_015_2788, w_015_2789, w_015_2790, w_015_2791, w_015_2792, w_015_2793, w_015_2794, w_015_2795, w_015_2797, w_015_2798, w_015_2799, w_015_2800, w_015_2801, w_015_2804, w_015_2805, w_015_2806, w_015_2807, w_015_2808, w_015_2809, w_015_2810, w_015_2811, w_015_2812, w_015_2813, w_015_2814, w_015_2815, w_015_2816, w_015_2817, w_015_2818, w_015_2819, w_015_2820, w_015_2821, w_015_2822, w_015_2824, w_015_2825, w_015_2826, w_015_2827, w_015_2828, w_015_2829, w_015_2830, w_015_2831, w_015_2832, w_015_2833, w_015_2835, w_015_2836, w_015_2837, w_015_2838, w_015_2839, w_015_2840, w_015_2841, w_015_2842, w_015_2843, w_015_2844, w_015_2845, w_015_2846, w_015_2847, w_015_2848, w_015_2849, w_015_2850, w_015_2851, w_015_2852, w_015_2853, w_015_2854, w_015_2855, w_015_2856, w_015_2857, w_015_2858, w_015_2859, w_015_2860, w_015_2861, w_015_2862, w_015_2863, w_015_2864, w_015_2865, w_015_2866, w_015_2867, w_015_2868, w_015_2869, w_015_2870, w_015_2871, w_015_2872, w_015_2873, w_015_2874, w_015_2875, w_015_2876, w_015_2877, w_015_2878, w_015_2879, w_015_2880, w_015_2881, w_015_2882, w_015_2883, w_015_2884, w_015_2885, w_015_2886, w_015_2887, w_015_2888, w_015_2889, w_015_2891, w_015_2895, w_015_2896, w_015_2897, w_015_2898, w_015_2899, w_015_2900, w_015_2901, w_015_2902, w_015_2904, w_015_2905, w_015_2906, w_015_2907, w_015_2908, w_015_2909, w_015_2911, w_015_2912, w_015_2913, w_015_2914, w_015_2915, w_015_2916, w_015_2918, w_015_2919, w_015_2920, w_015_2921, w_015_2923, w_015_2924, w_015_2925, w_015_2926, w_015_2927, w_015_2928, w_015_2929, w_015_2930, w_015_2931, w_015_2932, w_015_2933, w_015_2935, w_015_2936, w_015_2937, w_015_2938, w_015_2939, w_015_2940, w_015_2941, w_015_2943, w_015_2944, w_015_2945, w_015_2946, w_015_2947, w_015_2949, w_015_2950, w_015_2951, w_015_2952, w_015_2953, w_015_2954, w_015_2955, w_015_2956, w_015_2958, w_015_2959, w_015_2960, w_015_2961, w_015_2962, w_015_2963, w_015_2964, w_015_2965, w_015_2966, w_015_2967, w_015_2968, w_015_2969, w_015_2970, w_015_2971, w_015_2972, w_015_2973, w_015_2974, w_015_2975, w_015_2976, w_015_2977, w_015_2978, w_015_2979, w_015_2981, w_015_2982, w_015_2984, w_015_2985, w_015_2986, w_015_2987, w_015_2988, w_015_2989, w_015_2990, w_015_2991, w_015_2992, w_015_2993, w_015_2994, w_015_2995, w_015_2996, w_015_2997, w_015_2998, w_015_2999, w_015_3000, w_015_3001, w_015_3002, w_015_3003, w_015_3004, w_015_3005, w_015_3006, w_015_3007, w_015_3008, w_015_3009, w_015_3011, w_015_3012, w_015_3013, w_015_3014, w_015_3015, w_015_3016, w_015_3017, w_015_3018, w_015_3019, w_015_3020, w_015_3023, w_015_3025, w_015_3026, w_015_3027, w_015_3028, w_015_3029, w_015_3030, w_015_3031, w_015_3032, w_015_3033, w_015_3034, w_015_3035, w_015_3037, w_015_3038, w_015_3039, w_015_3040, w_015_3042, w_015_3043, w_015_3044, w_015_3045, w_015_3046, w_015_3047, w_015_3048, w_015_3049, w_015_3050, w_015_3051, w_015_3052, w_015_3054, w_015_3055, w_015_3056, w_015_3057, w_015_3058, w_015_3059, w_015_3060, w_015_3061, w_015_3062, w_015_3063, w_015_3064, w_015_3065, w_015_3066, w_015_3067, w_015_3068, w_015_3069, w_015_3070, w_015_3071, w_015_3072, w_015_3073, w_015_3074, w_015_3075, w_015_3076, w_015_3077, w_015_3078, w_015_3079, w_015_3080, w_015_3081, w_015_3082, w_015_3083, w_015_3084, w_015_3085, w_015_3086, w_015_3087, w_015_3089, w_015_3090, w_015_3091, w_015_3092, w_015_3093, w_015_3094, w_015_3095, w_015_3096, w_015_3097, w_015_3098, w_015_3099, w_015_3100, w_015_3101, w_015_3102, w_015_3103, w_015_3104, w_015_3105, w_015_3106, w_015_3108, w_015_3109, w_015_3110, w_015_3111, w_015_3112, w_015_3113, w_015_3115, w_015_3116, w_015_3117, w_015_3118, w_015_3119, w_015_3120, w_015_3122, w_015_3123, w_015_3124, w_015_3125, w_015_3126, w_015_3128, w_015_3130, w_015_3131, w_015_3132, w_015_3133, w_015_3134, w_015_3135, w_015_3136, w_015_3137, w_015_3138, w_015_3139, w_015_3140, w_015_3142, w_015_3145, w_015_3146, w_015_3148, w_015_3149, w_015_3150, w_015_3151, w_015_3155, w_015_3156, w_015_3157, w_015_3158, w_015_3159, w_015_3161, w_015_3163, w_015_3165, w_015_3166, w_015_3167, w_015_3170, w_015_3171, w_015_3172, w_015_3173, w_015_3174, w_015_3177, w_015_3180, w_015_3181, w_015_3182, w_015_3183, w_015_3184, w_015_3185, w_015_3186, w_015_3187, w_015_3188, w_015_3189, w_015_3191, w_015_3192, w_015_3194, w_015_3195, w_015_3197, w_015_3198, w_015_3199, w_015_3200, w_015_3201, w_015_3203, w_015_3204, w_015_3205, w_015_3206, w_015_3207, w_015_3208, w_015_3209, w_015_3210, w_015_3211, w_015_3212, w_015_3215, w_015_3216, w_015_3217, w_015_3218, w_015_3219, w_015_3220, w_015_3221, w_015_3222, w_015_3223, w_015_3224, w_015_3226, w_015_3227, w_015_3228, w_015_3229, w_015_3230, w_015_3231, w_015_3233, w_015_3235, w_015_3238, w_015_3240, w_015_3241, w_015_3245, w_015_3246, w_015_3250, w_015_3253, w_015_3254, w_015_3255, w_015_3256, w_015_3257, w_015_3258, w_015_3259, w_015_3260, w_015_3262, w_015_3264, w_015_3265, w_015_3266, w_015_3267, w_015_3271, w_015_3273, w_015_3275, w_015_3276, w_015_3277, w_015_3278, w_015_3280, w_015_3281, w_015_3282, w_015_3284, w_015_3285, w_015_3286, w_015_3287, w_015_3289, w_015_3290, w_015_3291, w_015_3292, w_015_3293, w_015_3295, w_015_3296, w_015_3298, w_015_3299, w_015_3301, w_015_3304, w_015_3305, w_015_3307, w_015_3308, w_015_3310, w_015_3311, w_015_3313, w_015_3315, w_015_3317, w_015_3318, w_015_3320, w_015_3321, w_015_3322, w_015_3326, w_015_3329, w_015_3330, w_015_3331, w_015_3332, w_015_3333, w_015_3334, w_015_3336, w_015_3337, w_015_3341, w_015_3342, w_015_3343, w_015_3347, w_015_3350, w_015_3351, w_015_3352, w_015_3354, w_015_3357, w_015_3359, w_015_3360, w_015_3361, w_015_3364, w_015_3365, w_015_3366, w_015_3368, w_015_3370, w_015_3372, w_015_3376, w_015_3377, w_015_3379, w_015_3380, w_015_3384, w_015_3387, w_015_3389, w_015_3390, w_015_3391, w_015_3392, w_015_3393, w_015_3395, w_015_3396, w_015_3397, w_015_3398, w_015_3399, w_015_3400, w_015_3401, w_015_3402, w_015_3404, w_015_3410, w_015_3411, w_015_3412, w_015_3413, w_015_3414, w_015_3416, w_015_3417, w_015_3419, w_015_3420, w_015_3422, w_015_3423, w_015_3424, w_015_3425, w_015_3426, w_015_3427, w_015_3428, w_015_3429, w_015_3430, w_015_3432, w_015_3433, w_015_3434, w_015_3435, w_015_3436, w_015_3437, w_015_3438, w_015_3439, w_015_3440, w_015_3441, w_015_3443, w_015_3444, w_015_3446, w_015_3448, w_015_3449, w_015_3450, w_015_3452, w_015_3454, w_015_3456, w_015_3458, w_015_3459, w_015_3461, w_015_3462, w_015_3463, w_015_3464, w_015_3465, w_015_3466, w_015_3468, w_015_3470, w_015_3473, w_015_3474, w_015_3475, w_015_3477, w_015_3479, w_015_3480, w_015_3481, w_015_3482, w_015_3483, w_015_3486, w_015_3488, w_015_3489, w_015_3490, w_015_3491, w_015_3492, w_015_3493, w_015_3494, w_015_3495, w_015_3496, w_015_3497, w_015_3498, w_015_3500, w_015_3502, w_015_3503, w_015_3504, w_015_3505, w_015_3506, w_015_3507, w_015_3508, w_015_3510, w_015_3513, w_015_3514, w_015_3515, w_015_3517, w_015_3518, w_015_3519, w_015_3522, w_015_3523, w_015_3524, w_015_3525, w_015_3526, w_015_3528, w_015_3530, w_015_3531, w_015_3532, w_015_3534, w_015_3535, w_015_3537, w_015_3539, w_015_3540, w_015_3542, w_015_3544, w_015_3545, w_015_3546, w_015_3547, w_015_3549, w_015_3550, w_015_3553, w_015_3554, w_015_3556, w_015_3559, w_015_3560, w_015_3561, w_015_3562, w_015_3563, w_015_3566, w_015_3567, w_015_3568, w_015_3569, w_015_3570, w_015_3571, w_015_3573, w_015_3575, w_015_3576, w_015_3577, w_015_3578, w_015_3579, w_015_3580, w_015_3581, w_015_3586, w_015_3588, w_015_3590, w_015_3591, w_015_3592, w_015_3595, w_015_3596, w_015_3597, w_015_3598, w_015_3599, w_015_3601, w_015_3604, w_015_3605, w_015_3606, w_015_3608, w_015_3609, w_015_3610, w_015_3613, w_015_3615, w_015_3616, w_015_3617, w_015_3618, w_015_3619, w_015_3620, w_015_3621, w_015_3622, w_015_3623, w_015_3625, w_015_3626, w_015_3628, w_015_3629, w_015_3630, w_015_3631, w_015_3632, w_015_3633, w_015_3634, w_015_3636, w_015_3637, w_015_3639, w_015_3640, w_015_3641, w_015_3642, w_015_3645, w_015_3647, w_015_3648, w_015_3649, w_015_3650, w_015_3651, w_015_3652, w_015_3653, w_015_3654, w_015_3656, w_015_3657, w_015_3661, w_015_3662, w_015_3664, w_015_3667, w_015_3668, w_015_3669, w_015_3673, w_015_3675, w_015_3677, w_015_3679, w_015_3683, w_015_3685, w_015_3686, w_015_3687, w_015_3690, w_015_3691, w_015_3693, w_015_3696, w_015_3697, w_015_3698, w_015_3699, w_015_3700, w_015_3701, w_015_3702, w_015_3707, w_015_3709, w_015_3711, w_015_3714, w_015_3715, w_015_3716, w_015_3717, w_015_3718, w_015_3720, w_015_3721, w_015_3722, w_015_3723, w_015_3726, w_015_3727, w_015_3728, w_015_3729, w_015_3730, w_015_3733, w_015_3734, w_015_3735, w_015_3736, w_015_3737, w_015_3739, w_015_3740, w_015_3741, w_015_3743, w_015_3744, w_015_3746, w_015_3747, w_015_3748, w_015_3749, w_015_3753, w_015_3754, w_015_3757, w_015_3759, w_015_3761, w_015_3763, w_015_3764, w_015_3765, w_015_3769, w_015_3770, w_015_3772, w_015_3775, w_015_3776, w_015_3777, w_015_3778, w_015_3780, w_015_3781, w_015_3784, w_015_3785, w_015_3788, w_015_3789, w_015_3792, w_015_3794, w_015_3796, w_015_3797, w_015_3798, w_015_3799, w_015_3800, w_015_3802, w_015_3803, w_015_3807, w_015_3809, w_015_3811, w_015_3812, w_015_3813, w_015_3815, w_015_3816, w_015_3818, w_015_3819, w_015_3820, w_015_3821, w_015_3824, w_015_3825, w_015_3827, w_015_3828, w_015_3829, w_015_3831, w_015_3832, w_015_3834, w_015_3835, w_015_3837, w_015_3839, w_015_3840, w_015_3843, w_015_3846, w_015_3847, w_015_3849, w_015_3850, w_015_3852, w_015_3854, w_015_3856, w_015_3857, w_015_3858, w_015_3859, w_015_3862, w_015_3863, w_015_3864, w_015_3865, w_015_3866, w_015_3867, w_015_3868, w_015_3869, w_015_3870, w_015_3872, w_015_3873, w_015_3874, w_015_3876, w_015_3878, w_015_3879, w_015_3882, w_015_3884, w_015_3885, w_015_3886, w_015_3890, w_015_3892, w_015_3893, w_015_3894, w_015_3895, w_015_3896, w_015_3899, w_015_3900, w_015_3901, w_015_3903, w_015_3904, w_015_3905, w_015_3907, w_015_3908, w_015_3909, w_015_3910, w_015_3911, w_015_3913, w_015_3914, w_015_3915, w_015_3916, w_015_3917, w_015_3918, w_015_3920, w_015_3922, w_015_3923, w_015_3925, w_015_3926, w_015_3927, w_015_3928, w_015_3930, w_015_3931, w_015_3932, w_015_3934, w_015_3935, w_015_3936, w_015_3938, w_015_3939, w_015_3943, w_015_3944, w_015_3945, w_015_3948, w_015_3949, w_015_3952, w_015_3953, w_015_3955, w_015_3956, w_015_3957, w_015_3959, w_015_3962, w_015_3963, w_015_3964, w_015_3965, w_015_3966, w_015_3967, w_015_3968, w_015_3969, w_015_3971, w_015_3973, w_015_3974, w_015_3975, w_015_3976, w_015_3978, w_015_3979, w_015_3983, w_015_3984, w_015_3985, w_015_3986, w_015_3987, w_015_3988, w_015_3989, w_015_3991, w_015_3992, w_015_3994, w_015_3995, w_015_3996, w_015_3997, w_015_3998, w_015_3999, w_015_4000, w_015_4001, w_015_4002, w_015_4004, w_015_4005, w_015_4006, w_015_4007, w_015_4008, w_015_4009, w_015_4011, w_015_4012, w_015_4014, w_015_4020, w_015_4021, w_015_4022, w_015_4023, w_015_4025, w_015_4026, w_015_4027, w_015_4028, w_015_4030, w_015_4031, w_015_4033, w_015_4034, w_015_4036, w_015_4037, w_015_4038, w_015_4040, w_015_4043, w_015_4045, w_015_4046, w_015_4049, w_015_4051, w_015_4055, w_015_4057, w_015_4058, w_015_4059, w_015_4062, w_015_4064, w_015_4065, w_015_4066, w_015_4068, w_015_4070, w_015_4071, w_015_4072, w_015_4073, w_015_4075, w_015_4076, w_015_4077, w_015_4078, w_015_4079, w_015_4080, w_015_4083, w_015_4084, w_015_4085, w_015_4086, w_015_4088, w_015_4089, w_015_4090, w_015_4091, w_015_4092, w_015_4093, w_015_4094, w_015_4095, w_015_4096, w_015_4097, w_015_4100, w_015_4104, w_015_4106, w_015_4108, w_015_4109, w_015_4110, w_015_4111, w_015_4114, w_015_4115, w_015_4118, w_015_4119, w_015_4120, w_015_4121, w_015_4124, w_015_4125, w_015_4126, w_015_4129, w_015_4130, w_015_4132, w_015_4133, w_015_4134, w_015_4137, w_015_4138, w_015_4139, w_015_4140, w_015_4141, w_015_4142, w_015_4143, w_015_4146, w_015_4147, w_015_4149, w_015_4150, w_015_4152, w_015_4154, w_015_4155, w_015_4156, w_015_4157, w_015_4159, w_015_4161, w_015_4164, w_015_4165, w_015_4168, w_015_4169, w_015_4170, w_015_4172, w_015_4173, w_015_4174, w_015_4175, w_015_4177, w_015_4179, w_015_4181, w_015_4182, w_015_4183, w_015_4184, w_015_4186, w_015_4187, w_015_4188, w_015_4190, w_015_4191, w_015_4193, w_015_4197, w_015_4200, w_015_4201, w_015_4204, w_015_4207, w_015_4208, w_015_4212, w_015_4213, w_015_4214, w_015_4215, w_015_4216, w_015_4218, w_015_4219, w_015_4223, w_015_4224, w_015_4225, w_015_4226, w_015_4227, w_015_4228, w_015_4229, w_015_4233, w_015_4235, w_015_4237, w_015_4238, w_015_4239, w_015_4240, w_015_4241, w_015_4242, w_015_4243, w_015_4247, w_015_4248, w_015_4251, w_015_4252, w_015_4253, w_015_4255, w_015_4258, w_015_4259, w_015_4260, w_015_4261, w_015_4263, w_015_4266, w_015_4267, w_015_4269, w_015_4271, w_015_4273, w_015_4274, w_015_4278, w_015_4279, w_015_4280, w_015_4281, w_015_4282, w_015_4283, w_015_4285, w_015_4286, w_015_4288, w_015_4289, w_015_4290, w_015_4291, w_015_4292, w_015_4293, w_015_4295, w_015_4296, w_015_4297, w_015_4299, w_015_4300, w_015_4302, w_015_4303, w_015_4304, w_015_4305, w_015_4307, w_015_4308, w_015_4311, w_015_4314, w_015_4315, w_015_4316, w_015_4318, w_015_4320, w_015_4321, w_015_4322, w_015_4324, w_015_4325, w_015_4326, w_015_4329, w_015_4331, w_015_4333, w_015_4334, w_015_4337, w_015_4338, w_015_4339, w_015_4340, w_015_4341, w_015_4343, w_015_4346, w_015_4348, w_015_4349, w_015_4351, w_015_4352, w_015_4353, w_015_4354, w_015_4358, w_015_4359, w_015_4360, w_015_4362, w_015_4364, w_015_4367, w_015_4368, w_015_4369, w_015_4371, w_015_4373, w_015_4374, w_015_4378, w_015_4379, w_015_4380, w_015_4382, w_015_4384, w_015_4386, w_015_4388, w_015_4394, w_015_4395, w_015_4396, w_015_4397, w_015_4398, w_015_4399, w_015_4400, w_015_4401, w_015_4402, w_015_4403, w_015_4404, w_015_4405, w_015_4407, w_015_4408, w_015_4409, w_015_4410, w_015_4411, w_015_4413, w_015_4415, w_015_4418, w_015_4419, w_015_4420, w_015_4422, w_015_4423, w_015_4424, w_015_4425, w_015_4427, w_015_4431, w_015_4433, w_015_4434, w_015_4436, w_015_4437, w_015_4438, w_015_4439, w_015_4440, w_015_4442, w_015_4443, w_015_4445, w_015_4446, w_015_4447, w_015_4448, w_015_4450, w_015_4451, w_015_4452, w_015_4453, w_015_4454, w_015_4455, w_015_4456, w_015_4457, w_015_4458, w_015_4461, w_015_4462, w_015_4463, w_015_4464, w_015_4465, w_015_4468, w_015_4469, w_015_4470, w_015_4471, w_015_4473, w_015_4475, w_015_4477, w_015_4478, w_015_4479, w_015_4480, w_015_4481, w_015_4483, w_015_4486, w_015_4488, w_015_4489, w_015_4490, w_015_4491, w_015_4492, w_015_4493, w_015_4496, w_015_4498, w_015_4499, w_015_4500, w_015_4501, w_015_4502, w_015_4504, w_015_4505, w_015_4507, w_015_4508, w_015_4510, w_015_4512, w_015_4513, w_015_4514, w_015_4515, w_015_4516, w_015_4518, w_015_4519, w_015_4521, w_015_4524, w_015_4525, w_015_4526, w_015_4527, w_015_4528, w_015_4530, w_015_4531, w_015_4532, w_015_4533, w_015_4534, w_015_4535, w_015_4536, w_015_4537, w_015_4538, w_015_4539, w_015_4540, w_015_4541, w_015_4542, w_015_4544, w_015_4545, w_015_4547, w_015_4548, w_015_4551, w_015_4552, w_015_4553, w_015_4554, w_015_4555, w_015_4556, w_015_4557, w_015_4560, w_015_4561, w_015_4565, w_015_4566, w_015_4568, w_015_4569, w_015_4572, w_015_4574, w_015_4575, w_015_4578, w_015_4579, w_015_4580, w_015_4581, w_015_4583, w_015_4584, w_015_4585, w_015_4586, w_015_4588, w_015_4589, w_015_4592, w_015_4595, w_015_4596, w_015_4597, w_015_4598, w_015_4600, w_015_4601, w_015_4602, w_015_4603, w_015_4604, w_015_4606, w_015_4607, w_015_4609, w_015_4610, w_015_4613, w_015_4614, w_015_4615, w_015_4616, w_015_4617, w_015_4620, w_015_4623, w_015_4624, w_015_4625, w_015_4627, w_015_4628, w_015_4630, w_015_4631, w_015_4635, w_015_4638, w_015_4641, w_015_4642, w_015_4643, w_015_4645, w_015_4647, w_015_4648, w_015_4649, w_015_4651, w_015_4653, w_015_4654, w_015_4656, w_015_4657, w_015_4658, w_015_4659, w_015_4660, w_015_4661, w_015_4663, w_015_4664, w_015_4666, w_015_4667, w_015_4671, w_015_4673, w_015_4675, w_015_4676, w_015_4678, w_015_4679, w_015_4680, w_015_4681, w_015_4682, w_015_4683, w_015_4685, w_015_4686, w_015_4688, w_015_4690, w_015_4692, w_015_4693, w_015_4695, w_015_4696, w_015_4697, w_015_4698, w_015_4699, w_015_4700, w_015_4701, w_015_4702, w_015_4703, w_015_4704, w_015_4705, w_015_4706, w_015_4707, w_015_4709, w_015_4711, w_015_4712, w_015_4713, w_015_4716, w_015_4717, w_015_4718, w_015_4719, w_015_4721, w_015_4722, w_015_4723, w_015_4724, w_015_4725, w_015_4726, w_015_4729, w_015_4732, w_015_4734, w_015_4735, w_015_4736, w_015_4738, w_015_4739, w_015_4740, w_015_4742, w_015_4743, w_015_4744, w_015_4745, w_015_4747, w_015_4749, w_015_4751, w_015_4753, w_015_4754, w_015_4755, w_015_4756, w_015_4757, w_015_4761, w_015_4762, w_015_4763, w_015_4764, w_015_4765, w_015_4766, w_015_4767, w_015_4770, w_015_4771, w_015_4772, w_015_4773, w_015_4774, w_015_4775, w_015_4776, w_015_4777, w_015_4778, w_015_4779, w_015_4780, w_015_4781, w_015_4784, w_015_4785, w_015_4786, w_015_4787, w_015_4788, w_015_4789, w_015_4790, w_015_4791, w_015_4793, w_015_4794, w_015_4795, w_015_4796, w_015_4797, w_015_4800, w_015_4801, w_015_4802, w_015_4803, w_015_4804, w_015_4805, w_015_4810, w_015_4811, w_015_4812, w_015_4813, w_015_4817, w_015_4818, w_015_4820, w_015_4823, w_015_4825, w_015_4826, w_015_4827, w_015_4829, w_015_4830, w_015_4831, w_015_4832, w_015_4834, w_015_4835, w_015_4836, w_015_4840, w_015_4842, w_015_4843, w_015_4844, w_015_4845, w_015_4846, w_015_4848, w_015_4850, w_015_4852, w_015_4854, w_015_4855, w_015_4856, w_015_4862, w_015_4863, w_015_4864, w_015_4865, w_015_4868, w_015_4869, w_015_4870, w_015_4872, w_015_4873, w_015_4875, w_015_4878, w_015_4879, w_015_4881, w_015_4882, w_015_4884, w_015_4885, w_015_4887, w_015_4891, w_015_4892, w_015_4893, w_015_4894, w_015_4895, w_015_4896, w_015_4897, w_015_4899, w_015_4900, w_015_4901, w_015_4902, w_015_4904, w_015_4905, w_015_4906, w_015_4907, w_015_4909, w_015_4910, w_015_4914, w_015_4915, w_015_4917, w_015_4919, w_015_4920, w_015_4921, w_015_4923, w_015_4926, w_015_4929, w_015_4930, w_015_4931, w_015_4932, w_015_4933, w_015_4934, w_015_4937, w_015_4938, w_015_4939, w_015_4940, w_015_4941, w_015_4942, w_015_4944, w_015_4949, w_015_4950, w_015_4952, w_015_4953, w_015_4954, w_015_4955, w_015_4956, w_015_4957, w_015_4959, w_015_4960, w_015_4961, w_015_4963, w_015_4965, w_015_4966, w_015_4969, w_015_4971, w_015_4973, w_015_4974, w_015_4979, w_015_4980, w_015_4982, w_015_4983, w_015_4984, w_015_4987, w_015_4989, w_015_4990, w_015_4991, w_015_4993, w_015_4995, w_015_4996, w_015_4997, w_015_4998, w_015_4999, w_015_5000, w_015_5001, w_015_5003, w_015_5004, w_015_5005, w_015_5006, w_015_5007, w_015_5008, w_015_5009, w_015_5011, w_015_5012, w_015_5013, w_015_5014, w_015_5016, w_015_5018, w_015_5019, w_015_5020, w_015_5023, w_015_5024, w_015_5026, w_015_5028, w_015_5029, w_015_5030, w_015_5031, w_015_5033, w_015_5034, w_015_5035, w_015_5036, w_015_5040, w_015_5041, w_015_5043, w_015_5047, w_015_5048, w_015_5049, w_015_5051, w_015_5052, w_015_5054, w_015_5056, w_015_5058, w_015_5061, w_015_5062, w_015_5063, w_015_5064, w_015_5065, w_015_5067, w_015_5068, w_015_5070, w_015_5072, w_015_5074, w_015_5076, w_015_5077, w_015_5079, w_015_5084, w_015_5085, w_015_5087, w_015_5088, w_015_5090, w_015_5092, w_015_5094, w_015_5095, w_015_5096, w_015_5097, w_015_5098, w_015_5099, w_015_5100, w_015_5101, w_015_5102, w_015_5104, w_015_5107, w_015_5108, w_015_5109, w_015_5110, w_015_5112, w_015_5113, w_015_5114, w_015_5115, w_015_5116, w_015_5118, w_015_5119, w_015_5120, w_015_5122, w_015_5124, w_015_5125, w_015_5128, w_015_5130, w_015_5132, w_015_5133, w_015_5134, w_015_5135, w_015_5136, w_015_5137, w_015_5141, w_015_5143, w_015_5146, w_015_5147, w_015_5148, w_015_5149, w_015_5151, w_015_5153, w_015_5154, w_015_5156, w_015_5158, w_015_5160, w_015_5161, w_015_5163, w_015_5164, w_015_5165, w_015_5167, w_015_5168, w_015_5170, w_015_5172, w_015_5173, w_015_5174, w_015_5175, w_015_5176, w_015_5177, w_015_5179, w_015_5180, w_015_5181, w_015_5183, w_015_5184, w_015_5186, w_015_5187, w_015_5188, w_015_5193, w_015_5194, w_015_5195, w_015_5196, w_015_5197, w_015_5198, w_015_5199, w_015_5200, w_015_5202, w_015_5203, w_015_5205, w_015_5207, w_015_5212, w_015_5214, w_015_5215, w_015_5217, w_015_5218, w_015_5220, w_015_5221, w_015_5222, w_015_5225, w_015_5226, w_015_5227, w_015_5228, w_015_5229, w_015_5230, w_015_5231, w_015_5232, w_015_5233, w_015_5234, w_015_5236, w_015_5238, w_015_5239, w_015_5240, w_015_5241, w_015_5242, w_015_5243, w_015_5244, w_015_5245, w_015_5246, w_015_5247, w_015_5248, w_015_5250, w_015_5251, w_015_5253, w_015_5256, w_015_5257, w_015_5259, w_015_5260, w_015_5261, w_015_5264, w_015_5265, w_015_5266, w_015_5269, w_015_5270, w_015_5271, w_015_5272, w_015_5274, w_015_5275, w_015_5276, w_015_5277, w_015_5278, w_015_5282, w_015_5285, w_015_5286, w_015_5288, w_015_5289, w_015_5290, w_015_5291, w_015_5292, w_015_5294, w_015_5295, w_015_5296, w_015_5298, w_015_5299, w_015_5301, w_015_5305, w_015_5307, w_015_5309, w_015_5310, w_015_5312, w_015_5313, w_015_5314, w_015_5316, w_015_5317, w_015_5319, w_015_5321, w_015_5323, w_015_5324, w_015_5325, w_015_5326, w_015_5327, w_015_5336, w_015_5337, w_015_5338, w_015_5341, w_015_5343, w_015_5344, w_015_5345, w_015_5347, w_015_5349, w_015_5350, w_015_5352, w_015_5353, w_015_5354, w_015_5356, w_015_5357, w_015_5358, w_015_5359, w_015_5362, w_015_5363, w_015_5364, w_015_5367, w_015_5368, w_015_5369, w_015_5371, w_015_5372, w_015_5374, w_015_5376, w_015_5377, w_015_5378, w_015_5379, w_015_5380, w_015_5381, w_015_5382, w_015_5384, w_015_5385, w_015_5386, w_015_5387, w_015_5390, w_015_5391, w_015_5393, w_015_5394, w_015_5395, w_015_5397, w_015_5398, w_015_5399, w_015_5400, w_015_5401, w_015_5403, w_015_5407, w_015_5408, w_015_5409, w_015_5410, w_015_5413, w_015_5414, w_015_5415, w_015_5417, w_015_5419, w_015_5420, w_015_5422, w_015_5423, w_015_5424, w_015_5425, w_015_5428, w_015_5433, w_015_5434, w_015_5435, w_015_5436, w_015_5437, w_015_5438, w_015_5439, w_015_5440, w_015_5441, w_015_5442, w_015_5443, w_015_5444, w_015_5445, w_015_5446, w_015_5448, w_015_5449, w_015_5452, w_015_5453, w_015_5454, w_015_5455, w_015_5456, w_015_5459, w_015_5461, w_015_5464, w_015_5465, w_015_5467, w_015_5468, w_015_5469, w_015_5470, w_015_5471, w_015_5472, w_015_5473, w_015_5474, w_015_5475, w_015_5476, w_015_5477, w_015_5478, w_015_5480, w_015_5481, w_015_5484, w_015_5485, w_015_5486, w_015_5487, w_015_5488, w_015_5490, w_015_5491, w_015_5492, w_015_5493, w_015_5495, w_015_5496, w_015_5497, w_015_5498, w_015_5499, w_015_5500, w_015_5501, w_015_5502, w_015_5504, w_015_5505, w_015_5506, w_015_5507, w_015_5508, w_015_5510, w_015_5511, w_015_5514, w_015_5515, w_015_5516, w_015_5518, w_015_5520, w_015_5521, w_015_5522, w_015_5523, w_015_5524, w_015_5525, w_015_5526, w_015_5527, w_015_5528, w_015_5529, w_015_5530, w_015_5531, w_015_5533, w_015_5534, w_015_5535, w_015_5536, w_015_5537, w_015_5538, w_015_5539, w_015_5543, w_015_5545, w_015_5547, w_015_5548, w_015_5549, w_015_5550, w_015_5551, w_015_5552, w_015_5553, w_015_5554, w_015_5555, w_015_5556, w_015_5557, w_015_5558, w_015_5560, w_015_5561, w_015_5563, w_015_5564, w_015_5565, w_015_5566, w_015_5570, w_015_5572, w_015_5575, w_015_5576, w_015_5577, w_015_5578, w_015_5579, w_015_5580, w_015_5582, w_015_5583, w_015_5585, w_015_5586, w_015_5587, w_015_5588, w_015_5589, w_015_5590, w_015_5592, w_015_5594, w_015_5595, w_015_5596, w_015_5597, w_015_5599, w_015_5600, w_015_5601, w_015_5602, w_015_5603, w_015_5604, w_015_5605, w_015_5607, w_015_5608, w_015_5609, w_015_5610, w_015_5613, w_015_5614, w_015_5615, w_015_5616, w_015_5617, w_015_5618, w_015_5620, w_015_5621, w_015_5622, w_015_5626, w_015_5627, w_015_5629, w_015_5630, w_015_5632, w_015_5633, w_015_5635, w_015_5636, w_015_5638, w_015_5639, w_015_5641, w_015_5642, w_015_5644, w_015_5647, w_015_5648, w_015_5650, w_015_5654, w_015_5656, w_015_5658, w_015_5659, w_015_5662, w_015_5664, w_015_5665, w_015_5666, w_015_5667, w_015_5672, w_015_5674, w_015_5676, w_015_5677, w_015_5679, w_015_5680, w_015_5681, w_015_5682, w_015_5684, w_015_5685, w_015_5686, w_015_5689, w_015_5691, w_015_5692, w_015_5693, w_015_5696, w_015_5697, w_015_5702, w_015_5705, w_015_5707, w_015_5708, w_015_5709, w_015_5711, w_015_5713, w_015_5715, w_015_5716, w_015_5717, w_015_5718, w_015_5719, w_015_5720, w_015_5721, w_015_5723, w_015_5724, w_015_5725, w_015_5727, w_015_5728, w_015_5730, w_015_5733, w_015_5735, w_015_5738, w_015_5739, w_015_5741, w_015_5742, w_015_5743, w_015_5744, w_015_5745, w_015_5748, w_015_5749, w_015_5750, w_015_5753, w_015_5756, w_015_5757, w_015_5758, w_015_5759, w_015_5760, w_015_5761, w_015_5763, w_015_5764, w_015_5765, w_015_5766, w_015_5768, w_015_5769, w_015_5770, w_015_5772, w_015_5774, w_015_5775, w_015_5777, w_015_5778, w_015_5780, w_015_5781, w_015_5782, w_015_5783, w_015_5785, w_015_5786, w_015_5788, w_015_5792, w_015_5793, w_015_5794, w_015_5795, w_015_5796, w_015_5798, w_015_5799, w_015_5800, w_015_5805, w_015_5808, w_015_5810, w_015_5811, w_015_5812, w_015_5813, w_015_5815, w_015_5816, w_015_5817, w_015_5818, w_015_5819, w_015_5820, w_015_5821, w_015_5822, w_015_5826, w_015_5827, w_015_5828, w_015_5829, w_015_5832, w_015_5834, w_015_5835, w_015_5838, w_015_5839, w_015_5840, w_015_5841, w_015_5843, w_015_5844, w_015_5845, w_015_5846, w_015_5849, w_015_5850, w_015_5851, w_015_5852, w_015_5854, w_015_5855, w_015_5856, w_015_5857, w_015_5858, w_015_5859, w_015_5860, w_015_5862, w_015_5863, w_015_5864, w_015_5870, w_015_5871, w_015_5872, w_015_5873, w_015_5874, w_015_5876, w_015_5877, w_015_5878, w_015_5879, w_015_5880, w_015_5882, w_015_5883, w_015_5884, w_015_5885, w_015_5887, w_015_5888, w_015_5890, w_015_5891, w_015_5892, w_015_5893, w_015_5895, w_015_5898, w_015_5900, w_015_5903, w_015_5904, w_015_5906, w_015_5907, w_015_5908, w_015_5909, w_015_5910, w_015_5912, w_015_5913, w_015_5914, w_015_5915, w_015_5916, w_015_5917, w_015_5918, w_015_5920, w_015_5922, w_015_5925, w_015_5928, w_015_5929, w_015_5931, w_015_5932, w_015_5933, w_015_5934, w_015_5938, w_015_5939, w_015_5940, w_015_5943, w_015_5944, w_015_5945, w_015_5946, w_015_5951, w_015_5952, w_015_5953, w_015_5954, w_015_5955, w_015_5956, w_015_5958, w_015_5959, w_015_5960, w_015_5961, w_015_5962, w_015_5963, w_015_5964, w_015_5965, w_015_5966, w_015_5968, w_015_5969, w_015_5972, w_015_5974, w_015_5975, w_015_5977, w_015_5978, w_015_5979, w_015_5980, w_015_5981, w_015_5982, w_015_5983, w_015_5985, w_015_5987, w_015_5988, w_015_5990, w_015_5991, w_015_5992, w_015_5993, w_015_5994, w_015_5996, w_015_5997, w_015_5999, w_015_6000, w_015_6001, w_015_6002, w_015_6004, w_015_6005, w_015_6006, w_015_6007, w_015_6012, w_015_6013, w_015_6015, w_015_6016, w_015_6017, w_015_6018, w_015_6019, w_015_6021, w_015_6022, w_015_6025, w_015_6026, w_015_6027, w_015_6028, w_015_6029, w_015_6030, w_015_6032, w_015_6033, w_015_6034, w_015_6036, w_015_6038, w_015_6039, w_015_6041, w_015_6043, w_015_6044, w_015_6047, w_015_6048, w_015_6049, w_015_6050, w_015_6051, w_015_6052, w_015_6053, w_015_6054, w_015_6055, w_015_6056, w_015_6057, w_015_6059, w_015_6060, w_015_6064, w_015_6065, w_015_6066, w_015_6067, w_015_6069, w_015_6071, w_015_6072, w_015_6073, w_015_6074, w_015_6075, w_015_6077, w_015_6078, w_015_6079, w_015_6080, w_015_6083, w_015_6084, w_015_6086, w_015_6087, w_015_6088, w_015_6089, w_015_6091, w_015_6092, w_015_6093, w_015_6094, w_015_6095, w_015_6096, w_015_6097, w_015_6098, w_015_6100, w_015_6101, w_015_6102, w_015_6104, w_015_6105, w_015_6107, w_015_6108, w_015_6109, w_015_6111, w_015_6112, w_015_6114, w_015_6117, w_015_6118, w_015_6119, w_015_6121, w_015_6122, w_015_6123, w_015_6124, w_015_6125, w_015_6126, w_015_6127, w_015_6128, w_015_6129, w_015_6130, w_015_6131, w_015_6132, w_015_6133, w_015_6134, w_015_6135, w_015_6136, w_015_6137, w_015_6138, w_015_6140, w_015_6141, w_015_6143, w_015_6144, w_015_6145, w_015_6146, w_015_6147, w_015_6148, w_015_6149, w_015_6150, w_015_6151, w_015_6152, w_015_6153, w_015_6154, w_015_6155, w_015_6156, w_015_6157, w_015_6158, w_015_6159, w_015_6161, w_015_6162, w_015_6164, w_015_6166, w_015_6167, w_015_6168, w_015_6169, w_015_6170, w_015_6172, w_015_6173, w_015_6175, w_015_6178, w_015_6181, w_015_6182, w_015_6183, w_015_6184, w_015_6185, w_015_6186, w_015_6187, w_015_6188, w_015_6190, w_015_6192, w_015_6193, w_015_6194, w_015_6197, w_015_6198, w_015_6199, w_015_6200, w_015_6201, w_015_6202, w_015_6204, w_015_6205, w_015_6206, w_015_6207, w_015_6208, w_015_6210, w_015_6211, w_015_6212, w_015_6214, w_015_6215, w_015_6216, w_015_6217, w_015_6219, w_015_6220, w_015_6221, w_015_6222, w_015_6224, w_015_6225, w_015_6226, w_015_6227, w_015_6229, w_015_6233, w_015_6235, w_015_6236, w_015_6237, w_015_6238, w_015_6239, w_015_6242, w_015_6243, w_015_6244, w_015_6245, w_015_6246, w_015_6248, w_015_6250, w_015_6254, w_015_6255, w_015_6256, w_015_6257, w_015_6258, w_015_6260, w_015_6262, w_015_6264, w_015_6266, w_015_6267, w_015_6268, w_015_6269, w_015_6270, w_015_6271, w_015_6273, w_015_6275, w_015_6276, w_015_6277, w_015_6278, w_015_6281, w_015_6282, w_015_6284, w_015_6289, w_015_6290, w_015_6291, w_015_6292, w_015_6297, w_015_6301, w_015_6302, w_015_6304, w_015_6305, w_015_6306, w_015_6307, w_015_6308, w_015_6309, w_015_6310, w_015_6311, w_015_6312, w_015_6314, w_015_6315, w_015_6320, w_015_6321, w_015_6322, w_015_6323, w_015_6324, w_015_6327, w_015_6329, w_015_6330, w_015_6331, w_015_6335, w_015_6336, w_015_6338, w_015_6339, w_015_6340, w_015_6342, w_015_6343, w_015_6344, w_015_6345, w_015_6348, w_015_6349, w_015_6353, w_015_6354, w_015_6356, w_015_6357, w_015_6358, w_015_6359, w_015_6362, w_015_6363, w_015_6365, w_015_6366, w_015_6368, w_015_6369, w_015_6372, w_015_6373, w_015_6374, w_015_6375, w_015_6376, w_015_6380, w_015_6383, w_015_6384, w_015_6385, w_015_6386, w_015_6387, w_015_6388, w_015_6390, w_015_6391, w_015_6392, w_015_6393, w_015_6394, w_015_6395, w_015_6396, w_015_6397, w_015_6398, w_015_6400, w_015_6403, w_015_6404, w_015_6407, w_015_6408, w_015_6409, w_015_6410, w_015_6413, w_015_6414, w_015_6415, w_015_6416, w_015_6418, w_015_6421, w_015_6422, w_015_6423, w_015_6424, w_015_6425, w_015_6426, w_015_6427, w_015_6428, w_015_6430, w_015_6431, w_015_6433, w_015_6435, w_015_6436, w_015_6437, w_015_6438, w_015_6439, w_015_6441, w_015_6442, w_015_6444, w_015_6446, w_015_6447, w_015_6449, w_015_6451, w_015_6452, w_015_6453, w_015_6458, w_015_6459, w_015_6461, w_015_6462, w_015_6463, w_015_6466, w_015_6467, w_015_6469, w_015_6470, w_015_6471, w_015_6472, w_015_6473, w_015_6474, w_015_6475, w_015_6476, w_015_6478, w_015_6479, w_015_6481, w_015_6483, w_015_6484, w_015_6485, w_015_6486, w_015_6487, w_015_6488, w_015_6489, w_015_6490, w_015_6491, w_015_6492, w_015_6493, w_015_6494, w_015_6497, w_015_6498, w_015_6500, w_015_6501, w_015_6502, w_015_6503, w_015_6504, w_015_6505, w_015_6506, w_015_6507, w_015_6509, w_015_6511, w_015_6512, w_015_6514, w_015_6515, w_015_6518, w_015_6521, w_015_6522, w_015_6524, w_015_6525, w_015_6526, w_015_6527, w_015_6528, w_015_6529, w_015_6530, w_015_6531, w_015_6532, w_015_6533, w_015_6534, w_015_6535, w_015_6536, w_015_6537, w_015_6538, w_015_6539, w_015_6540, w_015_6541, w_015_6542, w_015_6543, w_015_6545, w_015_6546, w_015_6548, w_015_6549, w_015_6551, w_015_6553, w_015_6554, w_015_6556, w_015_6557, w_015_6558, w_015_6559, w_015_6560, w_015_6561, w_015_6562, w_015_6563, w_015_6565, w_015_6566, w_015_6569, w_015_6570, w_015_6571, w_015_6572, w_015_6574, w_015_6576, w_015_6578, w_015_6579, w_015_6580, w_015_6581, w_015_6582, w_015_6583, w_015_6584, w_015_6585, w_015_6586, w_015_6587, w_015_6588, w_015_6589, w_015_6593, w_015_6594, w_015_6595, w_015_6596, w_015_6597, w_015_6599, w_015_6601, w_015_6603, w_015_6606, w_015_6609, w_015_6611, w_015_6612, w_015_6616, w_015_6617, w_015_6619, w_015_6620, w_015_6621, w_015_6624, w_015_6626, w_015_6628, w_015_6631, w_015_6633, w_015_6634, w_015_6635, w_015_6636, w_015_6637, w_015_6640, w_015_6641, w_015_6643, w_015_6644, w_015_6647, w_015_6648, w_015_6651, w_015_6656, w_015_6660, w_015_6662, w_015_6663, w_015_6665, w_015_6668, w_015_6669, w_015_6671, w_015_6672, w_015_6676, w_015_6677, w_015_6678, w_015_6679, w_015_6680, w_015_6682, w_015_6684, w_015_6686, w_015_6687, w_015_6688, w_015_6689, w_015_6690, w_015_6691, w_015_6692, w_015_6695, w_015_6696, w_015_6697, w_015_6698, w_015_6699, w_015_6702, w_015_6704, w_015_6705, w_015_6706, w_015_6707, w_015_6708, w_015_6709, w_015_6710, w_015_6711, w_015_6712, w_015_6714, w_015_6716, w_015_6717, w_015_6718, w_015_6719, w_015_6720, w_015_6721, w_015_6722, w_015_6724, w_015_6725, w_015_6726, w_015_6728, w_015_6729, w_015_6731, w_015_6732, w_015_6733, w_015_6734, w_015_6735, w_015_6737, w_015_6738, w_015_6739, w_015_6741, w_015_6743, w_015_6746, w_015_6747, w_015_6748, w_015_6749, w_015_6750, w_015_6752, w_015_6753, w_015_6754, w_015_6755, w_015_6757, w_015_6758, w_015_6759, w_015_6760, w_015_6766, w_015_6767, w_015_6768, w_015_6769, w_015_6770, w_015_6772, w_015_6773, w_015_6774, w_015_6775, w_015_6778, w_015_6779, w_015_6780, w_015_6781, w_015_6782, w_015_6783, w_015_6785, w_015_6786, w_015_6788, w_015_6789, w_015_6790, w_015_6791, w_015_6792, w_015_6793, w_015_6794, w_015_6795, w_015_6799, w_015_6801, w_015_6802, w_015_6804, w_015_6805, w_015_6806, w_015_6807, w_015_6808, w_015_6809, w_015_6810, w_015_6814, w_015_6815, w_015_6816, w_015_6817, w_015_6818, w_015_6820, w_015_6821, w_015_6822, w_015_6823, w_015_6826, w_015_6830, w_015_6831, w_015_6832, w_015_6833, w_015_6834, w_015_6835, w_015_6836, w_015_6838, w_015_6839, w_015_6840, w_015_6843, w_015_6845, w_015_6846, w_015_6847, w_015_6849, w_015_6850, w_015_6853, w_015_6854, w_015_6855, w_015_6857;
  wire w_016_000, w_016_001, w_016_002, w_016_003, w_016_004, w_016_005, w_016_006, w_016_007, w_016_008, w_016_009, w_016_010, w_016_011, w_016_012, w_016_013, w_016_014, w_016_015, w_016_016, w_016_017, w_016_018, w_016_019, w_016_020, w_016_021, w_016_022, w_016_023, w_016_024, w_016_025, w_016_026, w_016_027, w_016_028, w_016_029, w_016_030, w_016_031, w_016_032, w_016_033, w_016_034, w_016_035, w_016_036, w_016_037, w_016_038, w_016_039, w_016_040, w_016_041, w_016_042, w_016_043, w_016_044, w_016_045, w_016_046, w_016_047, w_016_048, w_016_049, w_016_050, w_016_051, w_016_052, w_016_053, w_016_054, w_016_055, w_016_056, w_016_057, w_016_058, w_016_059, w_016_060, w_016_061, w_016_062, w_016_063, w_016_064, w_016_065, w_016_066, w_016_067, w_016_068, w_016_069, w_016_070, w_016_071, w_016_072, w_016_073, w_016_074, w_016_075, w_016_076, w_016_077, w_016_078, w_016_079, w_016_080, w_016_081, w_016_082, w_016_083, w_016_084, w_016_085, w_016_086, w_016_087, w_016_088, w_016_089, w_016_090, w_016_091, w_016_092, w_016_093, w_016_094, w_016_095, w_016_096, w_016_097, w_016_098, w_016_099, w_016_100, w_016_101, w_016_102, w_016_103, w_016_104, w_016_105, w_016_106, w_016_107, w_016_108, w_016_109, w_016_110, w_016_111, w_016_112, w_016_113, w_016_114, w_016_115, w_016_116, w_016_117, w_016_118, w_016_119, w_016_120, w_016_121, w_016_122, w_016_123, w_016_124, w_016_125, w_016_126, w_016_127, w_016_128, w_016_129, w_016_130, w_016_131, w_016_132, w_016_133, w_016_134, w_016_136, w_016_137, w_016_138, w_016_139, w_016_140, w_016_141, w_016_142, w_016_143, w_016_144, w_016_145, w_016_146, w_016_147, w_016_148, w_016_149, w_016_150, w_016_151, w_016_152, w_016_153, w_016_154, w_016_155, w_016_156, w_016_157, w_016_158, w_016_159, w_016_160, w_016_161, w_016_162, w_016_163, w_016_164, w_016_165, w_016_166, w_016_167, w_016_168, w_016_169, w_016_170, w_016_171, w_016_172, w_016_173, w_016_174, w_016_175, w_016_176, w_016_177, w_016_178, w_016_179, w_016_180, w_016_181, w_016_182, w_016_183, w_016_184, w_016_185, w_016_186, w_016_187, w_016_188, w_016_189, w_016_190, w_016_191, w_016_192, w_016_193, w_016_194, w_016_195, w_016_196, w_016_197, w_016_198, w_016_199, w_016_200, w_016_201, w_016_202, w_016_203, w_016_204, w_016_205, w_016_206, w_016_207, w_016_208, w_016_209, w_016_210, w_016_211, w_016_212, w_016_213, w_016_214, w_016_215, w_016_216, w_016_217, w_016_218, w_016_219, w_016_220, w_016_221, w_016_222, w_016_223, w_016_224, w_016_225, w_016_226, w_016_227, w_016_228, w_016_229, w_016_230, w_016_231, w_016_232, w_016_233, w_016_234, w_016_235, w_016_236, w_016_237, w_016_238, w_016_239, w_016_240, w_016_241, w_016_242, w_016_243, w_016_244, w_016_245, w_016_246, w_016_247, w_016_248, w_016_249, w_016_250, w_016_251, w_016_252, w_016_253, w_016_254, w_016_255, w_016_256, w_016_257, w_016_258, w_016_259, w_016_260, w_016_261, w_016_262, w_016_263, w_016_264, w_016_265, w_016_266, w_016_267, w_016_268, w_016_269, w_016_270, w_016_271, w_016_272, w_016_273, w_016_274, w_016_275, w_016_276, w_016_277, w_016_278, w_016_279, w_016_280, w_016_281, w_016_282, w_016_283, w_016_284, w_016_285, w_016_286, w_016_287, w_016_288, w_016_289, w_016_290, w_016_291, w_016_292, w_016_293, w_016_294, w_016_295, w_016_296, w_016_297, w_016_298, w_016_299, w_016_300, w_016_301, w_016_302, w_016_303, w_016_304, w_016_305, w_016_306, w_016_307, w_016_308, w_016_309, w_016_310, w_016_311, w_016_312, w_016_313, w_016_314, w_016_315, w_016_316, w_016_317, w_016_318, w_016_319, w_016_320, w_016_321, w_016_322, w_016_323, w_016_324, w_016_325, w_016_326, w_016_327, w_016_328, w_016_329, w_016_330, w_016_331, w_016_332, w_016_333, w_016_334, w_016_335, w_016_336, w_016_337, w_016_338, w_016_339, w_016_340, w_016_341, w_016_342, w_016_343, w_016_344, w_016_345, w_016_346, w_016_347, w_016_348, w_016_349, w_016_350, w_016_351, w_016_352, w_016_353, w_016_354, w_016_355, w_016_356, w_016_357, w_016_358, w_016_359, w_016_360, w_016_361, w_016_362, w_016_363, w_016_364, w_016_365, w_016_366, w_016_367, w_016_368, w_016_369, w_016_370, w_016_371, w_016_372, w_016_373, w_016_374, w_016_375, w_016_376, w_016_377, w_016_378, w_016_379, w_016_380, w_016_381, w_016_382, w_016_383, w_016_384, w_016_385, w_016_386, w_016_387, w_016_388, w_016_389, w_016_390, w_016_391, w_016_392, w_016_393, w_016_394, w_016_396, w_016_397, w_016_398, w_016_399, w_016_400, w_016_401, w_016_402, w_016_403, w_016_404, w_016_405, w_016_406, w_016_407, w_016_408, w_016_409, w_016_410, w_016_411, w_016_412, w_016_413, w_016_414, w_016_415, w_016_416, w_016_417, w_016_418, w_016_419, w_016_420, w_016_421, w_016_422, w_016_423, w_016_424, w_016_425, w_016_426, w_016_427, w_016_428, w_016_429, w_016_430, w_016_431, w_016_432, w_016_433, w_016_434, w_016_435, w_016_436, w_016_437, w_016_438, w_016_439, w_016_440, w_016_441, w_016_442, w_016_443, w_016_444, w_016_445, w_016_446, w_016_447, w_016_448, w_016_449, w_016_450, w_016_451, w_016_452, w_016_453, w_016_454, w_016_455, w_016_456, w_016_457, w_016_458, w_016_459, w_016_460, w_016_461, w_016_462, w_016_463, w_016_464, w_016_465, w_016_466, w_016_467, w_016_468, w_016_469, w_016_471, w_016_472, w_016_473, w_016_474, w_016_475, w_016_476, w_016_477, w_016_478, w_016_479, w_016_480, w_016_481, w_016_482, w_016_483, w_016_484, w_016_485, w_016_486, w_016_487, w_016_488, w_016_489, w_016_490, w_016_491, w_016_492, w_016_493, w_016_494, w_016_495, w_016_496, w_016_497, w_016_498, w_016_499, w_016_500, w_016_501, w_016_502, w_016_503, w_016_504, w_016_505, w_016_506, w_016_507, w_016_508, w_016_509, w_016_510, w_016_511, w_016_512, w_016_513, w_016_514, w_016_515, w_016_516, w_016_517, w_016_518, w_016_519, w_016_520, w_016_521, w_016_522, w_016_523, w_016_524, w_016_525, w_016_526, w_016_527, w_016_528, w_016_529, w_016_530, w_016_531, w_016_532, w_016_533, w_016_534, w_016_535, w_016_536, w_016_537, w_016_538, w_016_539, w_016_540, w_016_541, w_016_542, w_016_543, w_016_544, w_016_545, w_016_546, w_016_547, w_016_548, w_016_549, w_016_550, w_016_551, w_016_552, w_016_553, w_016_554, w_016_555, w_016_556, w_016_557, w_016_558, w_016_559, w_016_560, w_016_561, w_016_562, w_016_563, w_016_564, w_016_565, w_016_566, w_016_567, w_016_568, w_016_569, w_016_570, w_016_571, w_016_572, w_016_573, w_016_574, w_016_575, w_016_576, w_016_577, w_016_578, w_016_579, w_016_580, w_016_581, w_016_582, w_016_583, w_016_584, w_016_585, w_016_586, w_016_587, w_016_588, w_016_589, w_016_590, w_016_591, w_016_592, w_016_593, w_016_594, w_016_595, w_016_596, w_016_597, w_016_598, w_016_599, w_016_600, w_016_601, w_016_602, w_016_603, w_016_604, w_016_605, w_016_606, w_016_607, w_016_608, w_016_609, w_016_610, w_016_611, w_016_612, w_016_613, w_016_614, w_016_615, w_016_616, w_016_617, w_016_618, w_016_619, w_016_620, w_016_621, w_016_622, w_016_623, w_016_624, w_016_625, w_016_626, w_016_627, w_016_628, w_016_629, w_016_630, w_016_632, w_016_633, w_016_634, w_016_635, w_016_636, w_016_637, w_016_638, w_016_639, w_016_640, w_016_641, w_016_642, w_016_643, w_016_644, w_016_645, w_016_646, w_016_647, w_016_648, w_016_649, w_016_650, w_016_651, w_016_652, w_016_653, w_016_654, w_016_655, w_016_656, w_016_657, w_016_658, w_016_659, w_016_660, w_016_661, w_016_662, w_016_663, w_016_664, w_016_665, w_016_666, w_016_667, w_016_668, w_016_669, w_016_670, w_016_671, w_016_672, w_016_673, w_016_674, w_016_675, w_016_676, w_016_677, w_016_678, w_016_679, w_016_680, w_016_681, w_016_682, w_016_683, w_016_684, w_016_685, w_016_686, w_016_687, w_016_688, w_016_689, w_016_690, w_016_691, w_016_692, w_016_693, w_016_694, w_016_695, w_016_696, w_016_697, w_016_698, w_016_699, w_016_700, w_016_701, w_016_702, w_016_703, w_016_704, w_016_705, w_016_706, w_016_707, w_016_708, w_016_709, w_016_710, w_016_711, w_016_712, w_016_713, w_016_714, w_016_715, w_016_716, w_016_717, w_016_718, w_016_719, w_016_720, w_016_721, w_016_722, w_016_723, w_016_724, w_016_725, w_016_726, w_016_727, w_016_728, w_016_729, w_016_730, w_016_731, w_016_732, w_016_733, w_016_734, w_016_735, w_016_736, w_016_737, w_016_738, w_016_739, w_016_740, w_016_741, w_016_742, w_016_743, w_016_744, w_016_745, w_016_746, w_016_747, w_016_748, w_016_749, w_016_750, w_016_751, w_016_752, w_016_753, w_016_754, w_016_755, w_016_756, w_016_757, w_016_758, w_016_759, w_016_760, w_016_761, w_016_762, w_016_763, w_016_764, w_016_765, w_016_766, w_016_767, w_016_768, w_016_769, w_016_770, w_016_771, w_016_772, w_016_773, w_016_774, w_016_775, w_016_776, w_016_777, w_016_778, w_016_779, w_016_780, w_016_781, w_016_782, w_016_783, w_016_784, w_016_785, w_016_786, w_016_787, w_016_788, w_016_789, w_016_790, w_016_791, w_016_792, w_016_793, w_016_794, w_016_795, w_016_796, w_016_797, w_016_798, w_016_799, w_016_800, w_016_801, w_016_802, w_016_803, w_016_804, w_016_805, w_016_806, w_016_807, w_016_808, w_016_809, w_016_810, w_016_811, w_016_812, w_016_813, w_016_814, w_016_815, w_016_816, w_016_817, w_016_818, w_016_819, w_016_820, w_016_821, w_016_822, w_016_823, w_016_824, w_016_825, w_016_826, w_016_827, w_016_828, w_016_829, w_016_830, w_016_831, w_016_832, w_016_833, w_016_834, w_016_835, w_016_836, w_016_837, w_016_838, w_016_839, w_016_840, w_016_841, w_016_842, w_016_843, w_016_844, w_016_845, w_016_846, w_016_847, w_016_848, w_016_849, w_016_850, w_016_851, w_016_852, w_016_853, w_016_854, w_016_856, w_016_857, w_016_858, w_016_859, w_016_860, w_016_861, w_016_862, w_016_863, w_016_864, w_016_865, w_016_866, w_016_867, w_016_868, w_016_869, w_016_870, w_016_871, w_016_872, w_016_873, w_016_874, w_016_875, w_016_876, w_016_877, w_016_878, w_016_879, w_016_880, w_016_881, w_016_882, w_016_883, w_016_884, w_016_885, w_016_886, w_016_887, w_016_888, w_016_889, w_016_890, w_016_891, w_016_892, w_016_893, w_016_894, w_016_895, w_016_896, w_016_897, w_016_898, w_016_899, w_016_900, w_016_901, w_016_902, w_016_903, w_016_904, w_016_905, w_016_906, w_016_907, w_016_908, w_016_909, w_016_910, w_016_911, w_016_912, w_016_913, w_016_914, w_016_915, w_016_916, w_016_917, w_016_918, w_016_919, w_016_920, w_016_921, w_016_922, w_016_923, w_016_924, w_016_925, w_016_926, w_016_927, w_016_928, w_016_929, w_016_930, w_016_931, w_016_932, w_016_933, w_016_934, w_016_935, w_016_936, w_016_937, w_016_938, w_016_939, w_016_940, w_016_941, w_016_942, w_016_943, w_016_944, w_016_945, w_016_946, w_016_947, w_016_948, w_016_949, w_016_950, w_016_951, w_016_952, w_016_953, w_016_954, w_016_955, w_016_956, w_016_957, w_016_958, w_016_959, w_016_960, w_016_961, w_016_962, w_016_963, w_016_964, w_016_965, w_016_966, w_016_967, w_016_968, w_016_969, w_016_970, w_016_971, w_016_972, w_016_973, w_016_974, w_016_975, w_016_976, w_016_977, w_016_978, w_016_979, w_016_980, w_016_981, w_016_982, w_016_983, w_016_984, w_016_985, w_016_986, w_016_987, w_016_988, w_016_989, w_016_990, w_016_991, w_016_992, w_016_993, w_016_994, w_016_995, w_016_996, w_016_997, w_016_998, w_016_999, w_016_1000, w_016_1001, w_016_1002, w_016_1003, w_016_1004, w_016_1005, w_016_1006, w_016_1007, w_016_1008, w_016_1009, w_016_1010, w_016_1011, w_016_1012, w_016_1013, w_016_1014, w_016_1015, w_016_1016, w_016_1017, w_016_1018, w_016_1019, w_016_1020, w_016_1021, w_016_1022, w_016_1023, w_016_1024, w_016_1025, w_016_1026, w_016_1027, w_016_1028, w_016_1029, w_016_1030, w_016_1031, w_016_1032, w_016_1033, w_016_1034, w_016_1035, w_016_1036, w_016_1037, w_016_1038, w_016_1039, w_016_1040, w_016_1041, w_016_1042, w_016_1043, w_016_1044, w_016_1045, w_016_1046, w_016_1047, w_016_1048, w_016_1049, w_016_1050, w_016_1051, w_016_1052, w_016_1053, w_016_1054, w_016_1055, w_016_1056, w_016_1057, w_016_1058, w_016_1059, w_016_1060, w_016_1061, w_016_1062, w_016_1063, w_016_1064, w_016_1065, w_016_1066, w_016_1067, w_016_1068, w_016_1069, w_016_1070, w_016_1071, w_016_1072, w_016_1073, w_016_1074, w_016_1075, w_016_1076, w_016_1077, w_016_1078, w_016_1079, w_016_1080, w_016_1081, w_016_1082, w_016_1083, w_016_1084, w_016_1085, w_016_1086, w_016_1087, w_016_1088, w_016_1089, w_016_1090, w_016_1091, w_016_1092, w_016_1093, w_016_1094, w_016_1095, w_016_1096, w_016_1097, w_016_1098, w_016_1099, w_016_1100, w_016_1101, w_016_1102, w_016_1103, w_016_1104, w_016_1105, w_016_1106, w_016_1107, w_016_1108, w_016_1109, w_016_1110, w_016_1111, w_016_1112, w_016_1113, w_016_1114, w_016_1115, w_016_1116, w_016_1117, w_016_1118, w_016_1119, w_016_1120, w_016_1121, w_016_1122, w_016_1123, w_016_1124, w_016_1125, w_016_1126, w_016_1127, w_016_1128, w_016_1129, w_016_1130, w_016_1131, w_016_1132, w_016_1133, w_016_1134, w_016_1135, w_016_1136, w_016_1137, w_016_1138, w_016_1139, w_016_1140, w_016_1141, w_016_1142, w_016_1143, w_016_1144, w_016_1145, w_016_1146, w_016_1147, w_016_1148, w_016_1149, w_016_1150, w_016_1151, w_016_1152, w_016_1153, w_016_1154, w_016_1155, w_016_1156, w_016_1157, w_016_1158, w_016_1159, w_016_1160, w_016_1161, w_016_1162, w_016_1163, w_016_1164, w_016_1165, w_016_1166, w_016_1167, w_016_1168, w_016_1169, w_016_1170, w_016_1171, w_016_1172, w_016_1173, w_016_1174, w_016_1175, w_016_1176, w_016_1177, w_016_1178, w_016_1179, w_016_1180, w_016_1181, w_016_1182, w_016_1183, w_016_1184, w_016_1185, w_016_1186, w_016_1187, w_016_1188, w_016_1189, w_016_1190, w_016_1191, w_016_1192, w_016_1193, w_016_1194, w_016_1195, w_016_1196, w_016_1197, w_016_1198, w_016_1199, w_016_1200, w_016_1201, w_016_1202, w_016_1203, w_016_1204, w_016_1205, w_016_1206, w_016_1207, w_016_1208, w_016_1209, w_016_1210, w_016_1211, w_016_1212, w_016_1213, w_016_1214, w_016_1215, w_016_1216, w_016_1217, w_016_1218, w_016_1219, w_016_1220, w_016_1221, w_016_1222, w_016_1223, w_016_1224, w_016_1225, w_016_1226, w_016_1227, w_016_1228, w_016_1229, w_016_1230, w_016_1231, w_016_1232, w_016_1233, w_016_1234, w_016_1235, w_016_1236, w_016_1237, w_016_1238, w_016_1239, w_016_1240, w_016_1241, w_016_1242, w_016_1243, w_016_1244, w_016_1245, w_016_1246, w_016_1247, w_016_1248, w_016_1249, w_016_1250, w_016_1251, w_016_1252, w_016_1253, w_016_1254, w_016_1255, w_016_1256, w_016_1257, w_016_1258, w_016_1259, w_016_1260, w_016_1261, w_016_1262, w_016_1263, w_016_1264, w_016_1265, w_016_1266, w_016_1267, w_016_1268, w_016_1269, w_016_1270, w_016_1271, w_016_1272, w_016_1273, w_016_1274, w_016_1275, w_016_1276, w_016_1277, w_016_1278, w_016_1279, w_016_1280, w_016_1281, w_016_1282, w_016_1283, w_016_1284, w_016_1285, w_016_1286, w_016_1287, w_016_1288, w_016_1289, w_016_1290, w_016_1291, w_016_1292, w_016_1293, w_016_1294, w_016_1295, w_016_1296, w_016_1297, w_016_1298, w_016_1299, w_016_1300, w_016_1301, w_016_1302, w_016_1303, w_016_1304, w_016_1305, w_016_1306, w_016_1307, w_016_1308, w_016_1309, w_016_1310, w_016_1311, w_016_1312, w_016_1313, w_016_1314, w_016_1315, w_016_1316, w_016_1317, w_016_1318, w_016_1319, w_016_1320, w_016_1321, w_016_1322, w_016_1323, w_016_1324, w_016_1325, w_016_1326, w_016_1327, w_016_1328, w_016_1329, w_016_1330, w_016_1331, w_016_1332, w_016_1333, w_016_1334, w_016_1335, w_016_1336, w_016_1337, w_016_1338, w_016_1339, w_016_1340, w_016_1341, w_016_1342, w_016_1343, w_016_1344, w_016_1345, w_016_1346, w_016_1347, w_016_1348, w_016_1349, w_016_1350, w_016_1351, w_016_1352, w_016_1353, w_016_1354, w_016_1355, w_016_1356, w_016_1357, w_016_1358, w_016_1359, w_016_1360, w_016_1361, w_016_1362, w_016_1363, w_016_1364, w_016_1365, w_016_1366, w_016_1367, w_016_1368, w_016_1369, w_016_1370, w_016_1371, w_016_1372, w_016_1373, w_016_1374, w_016_1375, w_016_1376, w_016_1377, w_016_1378, w_016_1379, w_016_1380, w_016_1381, w_016_1382, w_016_1383, w_016_1384, w_016_1385, w_016_1386, w_016_1387, w_016_1388, w_016_1389, w_016_1390, w_016_1391, w_016_1392, w_016_1393, w_016_1394, w_016_1395, w_016_1396, w_016_1397, w_016_1398, w_016_1399, w_016_1400, w_016_1401, w_016_1402, w_016_1403, w_016_1404, w_016_1405, w_016_1406, w_016_1407, w_016_1408, w_016_1409, w_016_1410, w_016_1411, w_016_1412, w_016_1413, w_016_1414, w_016_1415, w_016_1416, w_016_1417, w_016_1418, w_016_1419, w_016_1420, w_016_1421, w_016_1422, w_016_1423, w_016_1424, w_016_1425, w_016_1426, w_016_1427, w_016_1428, w_016_1429, w_016_1430, w_016_1431, w_016_1432, w_016_1433, w_016_1434, w_016_1435, w_016_1436, w_016_1437, w_016_1438, w_016_1439, w_016_1440, w_016_1441, w_016_1442, w_016_1443, w_016_1444, w_016_1445, w_016_1446, w_016_1447, w_016_1448, w_016_1449, w_016_1450, w_016_1451, w_016_1452, w_016_1453, w_016_1454, w_016_1455, w_016_1456, w_016_1457, w_016_1458, w_016_1459, w_016_1460, w_016_1461, w_016_1462, w_016_1463, w_016_1464, w_016_1465, w_016_1466, w_016_1467, w_016_1468, w_016_1469, w_016_1470, w_016_1471, w_016_1472, w_016_1473, w_016_1474, w_016_1475, w_016_1476, w_016_1477, w_016_1478, w_016_1479, w_016_1480, w_016_1481, w_016_1482, w_016_1483, w_016_1484, w_016_1485, w_016_1486, w_016_1487, w_016_1488, w_016_1489, w_016_1490, w_016_1491, w_016_1492, w_016_1493, w_016_1494, w_016_1495, w_016_1496, w_016_1497, w_016_1498, w_016_1499, w_016_1500, w_016_1501, w_016_1502, w_016_1503, w_016_1504, w_016_1505, w_016_1506, w_016_1507, w_016_1508, w_016_1509, w_016_1510, w_016_1511, w_016_1512, w_016_1513, w_016_1514, w_016_1515, w_016_1516, w_016_1517, w_016_1518, w_016_1519, w_016_1520, w_016_1521, w_016_1522, w_016_1523, w_016_1524, w_016_1525, w_016_1526, w_016_1527, w_016_1528, w_016_1529, w_016_1530, w_016_1531, w_016_1532, w_016_1533, w_016_1534, w_016_1535, w_016_1536, w_016_1537, w_016_1538, w_016_1539, w_016_1540, w_016_1541, w_016_1542, w_016_1543, w_016_1544, w_016_1545, w_016_1546, w_016_1547, w_016_1548, w_016_1549, w_016_1550, w_016_1551, w_016_1552, w_016_1553, w_016_1554, w_016_1555, w_016_1556, w_016_1557, w_016_1558, w_016_1559, w_016_1560, w_016_1561, w_016_1562, w_016_1563, w_016_1564, w_016_1565, w_016_1566, w_016_1567, w_016_1568, w_016_1569, w_016_1570, w_016_1571, w_016_1572, w_016_1573, w_016_1574, w_016_1575, w_016_1576, w_016_1577, w_016_1578, w_016_1579, w_016_1580, w_016_1581, w_016_1582, w_016_1583, w_016_1584, w_016_1585, w_016_1586, w_016_1587, w_016_1588, w_016_1589, w_016_1590, w_016_1591, w_016_1592, w_016_1593, w_016_1594, w_016_1595, w_016_1596, w_016_1597, w_016_1598, w_016_1599, w_016_1600, w_016_1601, w_016_1602, w_016_1603, w_016_1604, w_016_1605, w_016_1606, w_016_1607, w_016_1608, w_016_1609, w_016_1610, w_016_1611, w_016_1612, w_016_1613, w_016_1614, w_016_1615, w_016_1616, w_016_1617, w_016_1618, w_016_1619, w_016_1620, w_016_1621, w_016_1622, w_016_1623, w_016_1624, w_016_1625, w_016_1626, w_016_1627, w_016_1628, w_016_1629, w_016_1630, w_016_1631, w_016_1632, w_016_1633, w_016_1634, w_016_1635, w_016_1636, w_016_1637, w_016_1638, w_016_1639, w_016_1640, w_016_1641, w_016_1642, w_016_1643, w_016_1644, w_016_1645, w_016_1646, w_016_1647, w_016_1648, w_016_1649, w_016_1650, w_016_1651, w_016_1652, w_016_1653, w_016_1654, w_016_1655, w_016_1656, w_016_1657, w_016_1658, w_016_1659, w_016_1660, w_016_1661, w_016_1662, w_016_1663, w_016_1664, w_016_1665, w_016_1666, w_016_1667, w_016_1668, w_016_1669, w_016_1670, w_016_1671, w_016_1672, w_016_1673, w_016_1674, w_016_1675, w_016_1676, w_016_1677, w_016_1678, w_016_1679, w_016_1680, w_016_1681, w_016_1682, w_016_1683, w_016_1684, w_016_1685, w_016_1686, w_016_1687, w_016_1688, w_016_1689, w_016_1690, w_016_1691, w_016_1692, w_016_1693, w_016_1694, w_016_1695, w_016_1696, w_016_1697, w_016_1698, w_016_1699, w_016_1700, w_016_1701, w_016_1702, w_016_1703, w_016_1704, w_016_1705, w_016_1706, w_016_1707, w_016_1708, w_016_1709, w_016_1710, w_016_1711, w_016_1712, w_016_1713, w_016_1714, w_016_1715, w_016_1716, w_016_1717, w_016_1718, w_016_1719, w_016_1720, w_016_1721, w_016_1722, w_016_1723, w_016_1724, w_016_1725, w_016_1726, w_016_1727, w_016_1728, w_016_1729, w_016_1730, w_016_1731, w_016_1732, w_016_1733, w_016_1734, w_016_1735, w_016_1736, w_016_1737, w_016_1738, w_016_1739, w_016_1740, w_016_1741, w_016_1742, w_016_1743, w_016_1744, w_016_1745, w_016_1746, w_016_1747, w_016_1748, w_016_1749, w_016_1750, w_016_1751, w_016_1752, w_016_1753, w_016_1754, w_016_1755, w_016_1756, w_016_1757, w_016_1758, w_016_1759, w_016_1760, w_016_1761, w_016_1762, w_016_1763, w_016_1764, w_016_1765, w_016_1766, w_016_1767, w_016_1768, w_016_1769, w_016_1770, w_016_1771, w_016_1772, w_016_1773, w_016_1774, w_016_1775, w_016_1776, w_016_1777, w_016_1778, w_016_1779, w_016_1780, w_016_1781, w_016_1782, w_016_1783, w_016_1784, w_016_1785, w_016_1786, w_016_1787, w_016_1788, w_016_1789, w_016_1790, w_016_1791, w_016_1792, w_016_1793, w_016_1794, w_016_1795, w_016_1796, w_016_1797, w_016_1798, w_016_1799, w_016_1800, w_016_1801, w_016_1802, w_016_1803, w_016_1804, w_016_1805, w_016_1806, w_016_1807, w_016_1808, w_016_1809, w_016_1810, w_016_1811, w_016_1812, w_016_1813, w_016_1814, w_016_1815, w_016_1816, w_016_1817, w_016_1818, w_016_1819, w_016_1820, w_016_1821, w_016_1822, w_016_1823, w_016_1824, w_016_1825, w_016_1826, w_016_1827, w_016_1828, w_016_1829, w_016_1830, w_016_1831, w_016_1832, w_016_1833, w_016_1834, w_016_1835, w_016_1836, w_016_1837, w_016_1838, w_016_1839, w_016_1840, w_016_1841, w_016_1842, w_016_1843, w_016_1844, w_016_1845, w_016_1846, w_016_1847, w_016_1848, w_016_1849, w_016_1850, w_016_1851, w_016_1852, w_016_1853, w_016_1854, w_016_1855, w_016_1856, w_016_1857, w_016_1858, w_016_1859, w_016_1860, w_016_1861, w_016_1862, w_016_1863, w_016_1864, w_016_1865, w_016_1866, w_016_1867, w_016_1868, w_016_1869, w_016_1870, w_016_1871, w_016_1872, w_016_1873, w_016_1874, w_016_1875, w_016_1876, w_016_1877, w_016_1878, w_016_1879, w_016_1880, w_016_1881, w_016_1882, w_016_1883, w_016_1884, w_016_1885, w_016_1886, w_016_1887, w_016_1888, w_016_1889, w_016_1890, w_016_1891, w_016_1892, w_016_1893, w_016_1894, w_016_1895, w_016_1896, w_016_1897, w_016_1898, w_016_1899, w_016_1900, w_016_1901, w_016_1902, w_016_1903, w_016_1904, w_016_1905, w_016_1906, w_016_1907, w_016_1908, w_016_1909, w_016_1910, w_016_1911, w_016_1912, w_016_1913, w_016_1914, w_016_1915, w_016_1916, w_016_1917, w_016_1918, w_016_1919, w_016_1920, w_016_1921, w_016_1922, w_016_1923, w_016_1924, w_016_1925, w_016_1926, w_016_1927, w_016_1928, w_016_1929, w_016_1930, w_016_1931, w_016_1932, w_016_1933, w_016_1934, w_016_1935, w_016_1936, w_016_1937, w_016_1938, w_016_1939, w_016_1940, w_016_1941, w_016_1942, w_016_1943, w_016_1944, w_016_1945, w_016_1946, w_016_1947, w_016_1948, w_016_1949;
  wire w_017_000, w_017_001, w_017_002, w_017_003, w_017_004, w_017_006, w_017_007, w_017_008, w_017_009, w_017_010, w_017_011, w_017_012, w_017_013, w_017_014, w_017_015, w_017_016, w_017_017, w_017_018, w_017_019, w_017_020, w_017_021, w_017_022, w_017_023, w_017_025, w_017_026, w_017_027, w_017_028, w_017_029, w_017_030, w_017_031, w_017_032, w_017_033, w_017_034, w_017_035, w_017_036, w_017_037, w_017_038, w_017_039, w_017_040, w_017_041, w_017_042, w_017_043, w_017_044, w_017_045, w_017_046, w_017_047, w_017_048, w_017_049, w_017_050, w_017_051, w_017_052, w_017_053, w_017_054, w_017_055, w_017_056, w_017_057, w_017_058, w_017_059, w_017_060, w_017_061, w_017_062, w_017_063, w_017_064, w_017_065, w_017_066, w_017_067, w_017_068, w_017_069, w_017_070, w_017_071, w_017_072, w_017_073, w_017_074, w_017_075, w_017_076, w_017_077, w_017_078, w_017_079, w_017_080, w_017_081, w_017_082, w_017_083, w_017_084, w_017_085, w_017_086, w_017_087, w_017_088, w_017_089, w_017_090, w_017_091, w_017_092, w_017_093, w_017_095, w_017_096, w_017_097, w_017_098, w_017_099, w_017_100, w_017_101, w_017_102, w_017_103, w_017_104, w_017_105, w_017_106, w_017_107, w_017_108, w_017_109, w_017_110, w_017_111, w_017_112, w_017_113, w_017_114, w_017_115, w_017_116, w_017_117, w_017_118, w_017_119, w_017_120, w_017_121, w_017_122, w_017_123, w_017_124, w_017_125, w_017_126, w_017_127, w_017_128, w_017_129, w_017_131, w_017_132, w_017_133, w_017_134, w_017_135, w_017_136, w_017_137, w_017_138, w_017_139, w_017_140, w_017_141, w_017_142, w_017_143, w_017_144, w_017_146, w_017_147, w_017_148, w_017_149, w_017_150, w_017_151, w_017_152, w_017_153, w_017_154, w_017_155, w_017_156, w_017_157, w_017_158, w_017_159, w_017_160, w_017_161, w_017_162, w_017_163, w_017_164, w_017_165, w_017_166, w_017_167, w_017_168, w_017_169, w_017_170, w_017_171, w_017_172, w_017_173, w_017_174, w_017_175, w_017_176, w_017_177, w_017_178, w_017_179, w_017_180, w_017_181, w_017_182, w_017_183, w_017_184, w_017_185, w_017_186, w_017_187, w_017_188, w_017_189, w_017_190, w_017_191, w_017_192, w_017_193, w_017_194, w_017_195, w_017_196, w_017_197, w_017_198, w_017_199, w_017_200, w_017_201, w_017_202, w_017_203, w_017_204, w_017_205, w_017_206, w_017_207, w_017_208, w_017_209, w_017_210, w_017_211, w_017_212, w_017_213, w_017_214, w_017_215, w_017_216, w_017_217, w_017_218, w_017_219, w_017_220, w_017_221, w_017_222, w_017_223, w_017_224, w_017_226, w_017_227, w_017_228, w_017_229, w_017_230, w_017_231, w_017_232, w_017_233, w_017_234, w_017_235, w_017_236, w_017_237, w_017_238, w_017_239, w_017_240, w_017_241, w_017_242, w_017_243, w_017_244, w_017_245, w_017_246, w_017_247, w_017_248, w_017_249, w_017_250, w_017_251, w_017_252, w_017_253, w_017_254, w_017_255, w_017_256, w_017_257, w_017_258, w_017_259, w_017_260, w_017_261, w_017_262, w_017_263, w_017_264, w_017_265, w_017_266, w_017_267, w_017_268, w_017_269, w_017_270, w_017_271, w_017_272, w_017_273, w_017_274, w_017_275, w_017_276, w_017_277, w_017_278, w_017_279, w_017_280, w_017_281, w_017_282, w_017_284, w_017_285, w_017_287, w_017_288, w_017_289, w_017_290, w_017_291, w_017_292, w_017_293, w_017_294, w_017_295, w_017_296, w_017_297, w_017_298, w_017_299, w_017_300, w_017_301, w_017_302, w_017_303, w_017_304, w_017_305, w_017_306, w_017_307, w_017_308, w_017_309, w_017_310, w_017_311, w_017_312, w_017_313, w_017_314, w_017_315, w_017_316, w_017_317, w_017_318, w_017_319, w_017_320, w_017_321, w_017_322, w_017_323, w_017_324, w_017_325, w_017_326, w_017_327, w_017_328, w_017_329, w_017_330, w_017_331, w_017_332, w_017_334, w_017_335, w_017_336, w_017_337, w_017_338, w_017_339, w_017_340, w_017_342, w_017_343, w_017_344, w_017_345, w_017_346, w_017_347, w_017_348, w_017_349, w_017_350, w_017_351, w_017_352, w_017_353, w_017_354, w_017_355, w_017_356, w_017_357, w_017_358, w_017_359, w_017_360, w_017_361, w_017_362, w_017_363, w_017_364, w_017_365, w_017_366, w_017_367, w_017_368, w_017_369, w_017_370, w_017_371, w_017_372, w_017_373, w_017_374, w_017_375, w_017_376, w_017_377, w_017_378, w_017_379, w_017_380, w_017_381, w_017_382, w_017_383, w_017_384, w_017_385, w_017_386, w_017_387, w_017_388, w_017_389, w_017_390, w_017_391, w_017_392, w_017_393, w_017_394, w_017_395, w_017_398, w_017_399, w_017_400, w_017_401, w_017_402, w_017_403, w_017_404, w_017_405, w_017_406, w_017_407, w_017_408, w_017_409, w_017_410, w_017_411, w_017_412, w_017_413, w_017_414, w_017_415, w_017_416, w_017_417, w_017_418, w_017_419, w_017_420, w_017_421, w_017_422, w_017_423, w_017_424, w_017_425, w_017_426, w_017_427, w_017_428, w_017_429, w_017_431, w_017_432, w_017_433, w_017_434, w_017_435, w_017_436, w_017_437, w_017_438, w_017_439, w_017_440, w_017_441, w_017_442, w_017_443, w_017_444, w_017_445, w_017_446, w_017_447, w_017_449, w_017_450, w_017_451, w_017_452, w_017_453, w_017_454, w_017_455, w_017_456, w_017_457, w_017_458, w_017_459, w_017_460, w_017_461, w_017_462, w_017_463, w_017_464, w_017_465, w_017_466, w_017_467, w_017_468, w_017_469, w_017_470, w_017_471, w_017_472, w_017_473, w_017_474, w_017_475, w_017_476, w_017_477, w_017_478, w_017_479, w_017_480, w_017_481, w_017_482, w_017_483, w_017_484, w_017_486, w_017_487, w_017_489, w_017_491, w_017_492, w_017_493, w_017_494, w_017_495, w_017_496, w_017_497, w_017_498, w_017_499, w_017_500, w_017_501, w_017_502, w_017_503, w_017_504, w_017_505, w_017_506, w_017_507, w_017_508, w_017_509, w_017_510, w_017_511, w_017_512, w_017_513, w_017_514, w_017_515, w_017_516, w_017_517, w_017_518, w_017_519, w_017_520, w_017_521, w_017_522, w_017_523, w_017_524, w_017_525, w_017_526, w_017_527, w_017_528, w_017_529, w_017_530, w_017_531, w_017_532, w_017_533, w_017_534, w_017_535, w_017_536, w_017_537, w_017_538, w_017_539, w_017_540, w_017_541, w_017_542, w_017_543, w_017_544, w_017_545, w_017_546, w_017_547, w_017_548, w_017_549, w_017_550, w_017_551, w_017_552, w_017_553, w_017_554, w_017_555, w_017_556, w_017_557, w_017_558, w_017_559, w_017_560, w_017_562, w_017_563, w_017_564, w_017_565, w_017_566, w_017_567, w_017_568, w_017_570, w_017_571, w_017_572, w_017_573, w_017_574, w_017_575, w_017_576, w_017_577, w_017_578, w_017_579, w_017_580, w_017_581, w_017_582, w_017_583, w_017_584, w_017_586, w_017_587, w_017_588, w_017_589, w_017_590, w_017_591, w_017_592, w_017_593, w_017_594, w_017_595, w_017_596, w_017_597, w_017_598, w_017_599, w_017_600, w_017_601, w_017_602, w_017_604, w_017_605, w_017_606, w_017_607, w_017_608, w_017_609, w_017_610, w_017_611, w_017_612, w_017_613, w_017_614, w_017_615, w_017_616, w_017_617, w_017_618, w_017_619, w_017_620, w_017_621, w_017_622, w_017_623, w_017_624, w_017_625, w_017_626, w_017_627, w_017_628, w_017_629, w_017_630, w_017_631, w_017_632, w_017_633, w_017_634, w_017_635, w_017_636, w_017_637, w_017_639, w_017_640, w_017_641, w_017_642, w_017_643, w_017_644, w_017_645, w_017_646, w_017_647, w_017_648, w_017_649, w_017_650, w_017_652, w_017_653, w_017_654, w_017_655, w_017_656, w_017_657, w_017_658, w_017_659, w_017_660, w_017_661, w_017_662, w_017_663, w_017_664, w_017_665, w_017_666, w_017_667, w_017_668, w_017_669, w_017_670, w_017_671, w_017_672, w_017_673, w_017_674, w_017_675, w_017_676, w_017_677, w_017_678, w_017_679, w_017_680, w_017_681, w_017_682, w_017_683, w_017_684, w_017_685, w_017_686, w_017_687, w_017_688, w_017_689, w_017_690, w_017_691, w_017_692, w_017_693, w_017_694, w_017_695, w_017_696, w_017_697, w_017_698, w_017_699, w_017_700, w_017_701, w_017_702, w_017_703, w_017_704, w_017_705, w_017_706, w_017_707, w_017_708, w_017_709, w_017_710, w_017_711, w_017_712, w_017_713, w_017_714, w_017_715, w_017_716, w_017_717, w_017_718, w_017_719, w_017_720, w_017_721, w_017_722, w_017_723, w_017_724, w_017_725, w_017_726, w_017_727, w_017_728, w_017_729, w_017_730, w_017_731, w_017_732, w_017_733, w_017_734, w_017_735, w_017_736, w_017_737, w_017_739, w_017_740, w_017_741, w_017_742, w_017_743, w_017_744, w_017_745, w_017_746, w_017_747, w_017_748, w_017_749, w_017_750, w_017_751, w_017_752, w_017_753, w_017_754, w_017_755, w_017_756, w_017_757, w_017_758, w_017_759, w_017_760, w_017_761, w_017_762, w_017_763, w_017_764, w_017_765, w_017_766, w_017_767, w_017_768, w_017_769, w_017_770, w_017_771, w_017_772, w_017_773, w_017_774, w_017_775, w_017_776, w_017_777, w_017_778, w_017_779, w_017_780, w_017_781, w_017_782, w_017_783, w_017_784, w_017_785, w_017_786, w_017_787, w_017_788, w_017_789, w_017_790, w_017_791, w_017_792, w_017_793, w_017_794, w_017_795, w_017_796, w_017_797, w_017_798, w_017_799, w_017_800, w_017_802, w_017_803, w_017_804, w_017_805, w_017_806, w_017_807, w_017_808, w_017_809, w_017_810, w_017_811, w_017_812, w_017_813, w_017_814, w_017_815, w_017_816, w_017_817, w_017_818, w_017_820, w_017_821, w_017_822, w_017_823, w_017_824, w_017_825, w_017_826, w_017_827, w_017_828, w_017_829, w_017_830, w_017_832, w_017_833, w_017_834, w_017_835, w_017_836, w_017_837, w_017_838, w_017_839, w_017_840, w_017_841, w_017_842, w_017_844, w_017_845, w_017_846, w_017_847, w_017_848, w_017_849, w_017_850, w_017_851, w_017_852, w_017_853, w_017_854, w_017_855, w_017_856, w_017_858, w_017_859, w_017_860, w_017_861, w_017_862, w_017_863, w_017_864, w_017_865, w_017_866, w_017_867, w_017_868, w_017_869, w_017_870, w_017_871, w_017_872, w_017_873, w_017_874, w_017_875, w_017_876, w_017_877, w_017_878, w_017_879, w_017_880, w_017_881, w_017_882, w_017_883, w_017_884, w_017_885, w_017_886, w_017_887, w_017_888, w_017_889, w_017_890, w_017_891, w_017_892, w_017_893, w_017_894, w_017_895, w_017_896, w_017_897, w_017_898, w_017_899, w_017_900, w_017_901, w_017_902, w_017_903, w_017_904, w_017_905, w_017_906, w_017_907, w_017_908, w_017_909, w_017_910, w_017_911, w_017_912, w_017_913, w_017_914, w_017_915, w_017_916, w_017_917, w_017_918, w_017_921, w_017_922, w_017_925, w_017_926, w_017_928, w_017_929, w_017_930, w_017_931, w_017_932, w_017_933, w_017_934, w_017_935, w_017_936, w_017_937, w_017_938, w_017_939, w_017_940, w_017_941, w_017_942, w_017_943, w_017_944, w_017_945, w_017_946, w_017_947, w_017_948, w_017_949, w_017_950, w_017_951, w_017_952, w_017_953, w_017_954, w_017_955, w_017_956, w_017_957, w_017_958, w_017_959, w_017_960, w_017_961, w_017_962, w_017_963, w_017_964, w_017_965, w_017_966, w_017_967, w_017_968, w_017_969, w_017_970, w_017_971, w_017_972, w_017_973, w_017_974, w_017_975, w_017_976, w_017_977, w_017_978, w_017_979, w_017_980, w_017_981, w_017_982, w_017_983, w_017_984, w_017_985, w_017_986, w_017_987, w_017_988, w_017_989, w_017_990, w_017_991, w_017_992, w_017_993, w_017_994, w_017_995, w_017_996, w_017_997, w_017_998, w_017_999, w_017_1000, w_017_1001, w_017_1002, w_017_1003, w_017_1004, w_017_1005, w_017_1006, w_017_1007, w_017_1008, w_017_1009, w_017_1010, w_017_1011, w_017_1012, w_017_1013, w_017_1014, w_017_1015, w_017_1016, w_017_1017, w_017_1018, w_017_1019, w_017_1020, w_017_1021, w_017_1022, w_017_1023, w_017_1024, w_017_1025, w_017_1026, w_017_1027, w_017_1028, w_017_1029, w_017_1030, w_017_1031, w_017_1032, w_017_1033, w_017_1034, w_017_1035, w_017_1036, w_017_1037, w_017_1038, w_017_1039, w_017_1040, w_017_1041, w_017_1042, w_017_1043, w_017_1044, w_017_1045, w_017_1046, w_017_1047, w_017_1048, w_017_1049, w_017_1050, w_017_1051, w_017_1052, w_017_1053, w_017_1054, w_017_1055, w_017_1056, w_017_1057, w_017_1058, w_017_1059, w_017_1060, w_017_1061, w_017_1062, w_017_1063, w_017_1064, w_017_1065, w_017_1066, w_017_1067, w_017_1069, w_017_1070, w_017_1071, w_017_1072, w_017_1073, w_017_1074, w_017_1075, w_017_1076, w_017_1077, w_017_1078, w_017_1079, w_017_1080, w_017_1081, w_017_1082, w_017_1083, w_017_1084, w_017_1085, w_017_1086, w_017_1088, w_017_1089, w_017_1090, w_017_1091, w_017_1092, w_017_1093, w_017_1094, w_017_1095, w_017_1096, w_017_1097, w_017_1098, w_017_1099, w_017_1100, w_017_1101, w_017_1102, w_017_1103, w_017_1104, w_017_1105, w_017_1106, w_017_1107, w_017_1108, w_017_1109, w_017_1110, w_017_1111, w_017_1112, w_017_1113, w_017_1114, w_017_1115, w_017_1116, w_017_1117, w_017_1118, w_017_1119, w_017_1120, w_017_1121, w_017_1122, w_017_1123, w_017_1124, w_017_1125, w_017_1126, w_017_1127, w_017_1128, w_017_1129, w_017_1130, w_017_1131, w_017_1132, w_017_1133, w_017_1134, w_017_1135, w_017_1136, w_017_1137, w_017_1138, w_017_1139, w_017_1140, w_017_1141, w_017_1142, w_017_1145, w_017_1146, w_017_1147, w_017_1148, w_017_1149, w_017_1150, w_017_1151, w_017_1152, w_017_1153, w_017_1154, w_017_1155, w_017_1156, w_017_1157, w_017_1158, w_017_1159, w_017_1160, w_017_1161, w_017_1162, w_017_1163, w_017_1164, w_017_1165, w_017_1166, w_017_1167, w_017_1168, w_017_1169, w_017_1170, w_017_1171, w_017_1172, w_017_1173, w_017_1174, w_017_1175, w_017_1176, w_017_1177, w_017_1178, w_017_1179, w_017_1180, w_017_1181, w_017_1182, w_017_1183, w_017_1184, w_017_1185, w_017_1186, w_017_1187, w_017_1188, w_017_1189, w_017_1190, w_017_1191, w_017_1192, w_017_1193, w_017_1194, w_017_1195, w_017_1196, w_017_1197, w_017_1198, w_017_1199, w_017_1200, w_017_1201, w_017_1202, w_017_1203, w_017_1204, w_017_1205, w_017_1206, w_017_1207, w_017_1208, w_017_1209, w_017_1210, w_017_1211, w_017_1212, w_017_1213, w_017_1214, w_017_1215, w_017_1216, w_017_1217, w_017_1218, w_017_1219, w_017_1220, w_017_1221, w_017_1222, w_017_1223, w_017_1224, w_017_1225, w_017_1226, w_017_1227, w_017_1228, w_017_1229, w_017_1230, w_017_1231, w_017_1232, w_017_1233, w_017_1234, w_017_1235, w_017_1236, w_017_1237, w_017_1238, w_017_1239, w_017_1240, w_017_1241, w_017_1242, w_017_1243, w_017_1244, w_017_1245, w_017_1246, w_017_1247, w_017_1248, w_017_1249, w_017_1250, w_017_1251, w_017_1253, w_017_1254, w_017_1255, w_017_1256, w_017_1257, w_017_1258, w_017_1259, w_017_1260, w_017_1261, w_017_1262, w_017_1263, w_017_1264, w_017_1265, w_017_1266, w_017_1267, w_017_1268, w_017_1269, w_017_1270, w_017_1271, w_017_1272, w_017_1273, w_017_1274, w_017_1275, w_017_1276, w_017_1277, w_017_1278, w_017_1279, w_017_1281, w_017_1282, w_017_1283, w_017_1284, w_017_1285, w_017_1286, w_017_1287, w_017_1288, w_017_1289, w_017_1290, w_017_1291, w_017_1292, w_017_1293, w_017_1294, w_017_1295, w_017_1296, w_017_1297, w_017_1298, w_017_1299, w_017_1300, w_017_1301, w_017_1302, w_017_1303, w_017_1304, w_017_1305, w_017_1306, w_017_1307, w_017_1308, w_017_1310, w_017_1311, w_017_1312, w_017_1313, w_017_1314, w_017_1315, w_017_1316, w_017_1317, w_017_1318, w_017_1319, w_017_1320, w_017_1321, w_017_1322, w_017_1323, w_017_1324, w_017_1325, w_017_1326, w_017_1327, w_017_1329, w_017_1330, w_017_1331, w_017_1332, w_017_1333, w_017_1334, w_017_1335, w_017_1336, w_017_1337, w_017_1338, w_017_1339, w_017_1340, w_017_1341, w_017_1342, w_017_1344, w_017_1345, w_017_1346, w_017_1347, w_017_1349, w_017_1350, w_017_1351, w_017_1352, w_017_1353, w_017_1354, w_017_1355, w_017_1356, w_017_1357, w_017_1358, w_017_1359, w_017_1360, w_017_1361, w_017_1362, w_017_1363, w_017_1364, w_017_1365, w_017_1366, w_017_1367, w_017_1368, w_017_1369, w_017_1370, w_017_1371, w_017_1372, w_017_1373, w_017_1374, w_017_1375, w_017_1376, w_017_1377, w_017_1378, w_017_1379, w_017_1380, w_017_1381, w_017_1383, w_017_1384, w_017_1385, w_017_1386, w_017_1387, w_017_1388, w_017_1389, w_017_1390, w_017_1391, w_017_1392, w_017_1393, w_017_1394, w_017_1395, w_017_1396, w_017_1397, w_017_1398, w_017_1399, w_017_1400, w_017_1403, w_017_1404, w_017_1405, w_017_1406, w_017_1407, w_017_1408, w_017_1409, w_017_1410, w_017_1411, w_017_1412, w_017_1413, w_017_1414, w_017_1415, w_017_1416, w_017_1417, w_017_1418, w_017_1419, w_017_1420, w_017_1421, w_017_1422, w_017_1423, w_017_1425, w_017_1426, w_017_1427, w_017_1428, w_017_1429, w_017_1430, w_017_1431, w_017_1432, w_017_1433, w_017_1434, w_017_1435, w_017_1436, w_017_1437, w_017_1438, w_017_1439, w_017_1440, w_017_1441, w_017_1442, w_017_1443, w_017_1444, w_017_1445, w_017_1446, w_017_1447, w_017_1448, w_017_1450, w_017_1451, w_017_1452, w_017_1453, w_017_1454, w_017_1455, w_017_1456, w_017_1457, w_017_1458, w_017_1459, w_017_1460, w_017_1461, w_017_1462, w_017_1463, w_017_1464, w_017_1465, w_017_1466, w_017_1467, w_017_1468, w_017_1469, w_017_1470, w_017_1471, w_017_1472, w_017_1473, w_017_1474, w_017_1475, w_017_1476, w_017_1477, w_017_1478, w_017_1479, w_017_1480, w_017_1481, w_017_1482, w_017_1483, w_017_1484, w_017_1485, w_017_1486, w_017_1487, w_017_1488, w_017_1490, w_017_1491, w_017_1492, w_017_1493, w_017_1494, w_017_1495, w_017_1496, w_017_1497, w_017_1498, w_017_1499, w_017_1500, w_017_1501, w_017_1502, w_017_1503, w_017_1504, w_017_1505, w_017_1506, w_017_1508, w_017_1509, w_017_1510, w_017_1511, w_017_1512, w_017_1513, w_017_1514, w_017_1515, w_017_1516, w_017_1517, w_017_1519, w_017_1520, w_017_1521, w_017_1522, w_017_1523, w_017_1524, w_017_1525, w_017_1526, w_017_1527, w_017_1528, w_017_1529, w_017_1530, w_017_1531, w_017_1532, w_017_1533, w_017_1534, w_017_1535, w_017_1536, w_017_1537, w_017_1538, w_017_1539, w_017_1540, w_017_1541, w_017_1542, w_017_1543, w_017_1544, w_017_1545, w_017_1546, w_017_1548, w_017_1549, w_017_1550, w_017_1551, w_017_1552, w_017_1553, w_017_1554, w_017_1555, w_017_1556, w_017_1557, w_017_1558, w_017_1559, w_017_1560, w_017_1561, w_017_1562, w_017_1563, w_017_1564, w_017_1565, w_017_1566, w_017_1567, w_017_1568, w_017_1569, w_017_1570, w_017_1571, w_017_1572, w_017_1573, w_017_1574, w_017_1575, w_017_1576, w_017_1577, w_017_1578, w_017_1580, w_017_1581, w_017_1582, w_017_1583, w_017_1584, w_017_1585, w_017_1586, w_017_1587, w_017_1588, w_017_1589, w_017_1590, w_017_1591, w_017_1592, w_017_1593, w_017_1594, w_017_1595, w_017_1596, w_017_1597, w_017_1598, w_017_1599, w_017_1600, w_017_1601, w_017_1602, w_017_1604, w_017_1605, w_017_1606, w_017_1607, w_017_1608, w_017_1609, w_017_1610, w_017_1611, w_017_1612, w_017_1613, w_017_1614, w_017_1615, w_017_1616, w_017_1617, w_017_1618, w_017_1619, w_017_1620, w_017_1621, w_017_1622, w_017_1623, w_017_1624, w_017_1625, w_017_1626, w_017_1627, w_017_1628, w_017_1629, w_017_1633, w_017_1634, w_017_1635, w_017_1636, w_017_1637, w_017_1638, w_017_1639, w_017_1640, w_017_1642, w_017_1643, w_017_1644, w_017_1645, w_017_1646, w_017_1647, w_017_1648, w_017_1649, w_017_1650, w_017_1651, w_017_1652, w_017_1653, w_017_1654, w_017_1655, w_017_1656, w_017_1657, w_017_1658, w_017_1659, w_017_1661, w_017_1662, w_017_1663, w_017_1664, w_017_1665, w_017_1666, w_017_1667, w_017_1668, w_017_1669, w_017_1670, w_017_1671, w_017_1672, w_017_1673, w_017_1674, w_017_1675, w_017_1676, w_017_1677, w_017_1678, w_017_1679, w_017_1680, w_017_1681, w_017_1682, w_017_1683, w_017_1684, w_017_1685, w_017_1686, w_017_1687, w_017_1688, w_017_1689, w_017_1690, w_017_1691, w_017_1692, w_017_1693, w_017_1694, w_017_1695, w_017_1696, w_017_1697, w_017_1698, w_017_1699, w_017_1700, w_017_1701, w_017_1702, w_017_1703, w_017_1704, w_017_1705, w_017_1706, w_017_1707, w_017_1708, w_017_1709, w_017_1710, w_017_1711, w_017_1712, w_017_1713, w_017_1714, w_017_1715, w_017_1716, w_017_1717, w_017_1718, w_017_1719, w_017_1720, w_017_1721, w_017_1722, w_017_1724, w_017_1725, w_017_1726, w_017_1727, w_017_1728, w_017_1729, w_017_1730, w_017_1731, w_017_1732, w_017_1733, w_017_1734, w_017_1735, w_017_1736, w_017_1737, w_017_1738, w_017_1739, w_017_1741, w_017_1742, w_017_1743, w_017_1744, w_017_1745, w_017_1746, w_017_1747, w_017_1748, w_017_1749, w_017_1750, w_017_1751, w_017_1752, w_017_1753, w_017_1754, w_017_1755, w_017_1756, w_017_1757, w_017_1758, w_017_1759, w_017_1760, w_017_1761, w_017_1762, w_017_1763, w_017_1764, w_017_1765, w_017_1766, w_017_1767, w_017_1768, w_017_1769, w_017_1770, w_017_1771, w_017_1772, w_017_1773, w_017_1775, w_017_1776, w_017_1777, w_017_1778, w_017_1779, w_017_1780, w_017_1781, w_017_1782, w_017_1783, w_017_1784, w_017_1786, w_017_1787, w_017_1788, w_017_1789, w_017_1790, w_017_1791, w_017_1792, w_017_1793, w_017_1794, w_017_1795, w_017_1796, w_017_1797, w_017_1798, w_017_1799, w_017_1800, w_017_1801, w_017_1802, w_017_1803, w_017_1804, w_017_1805, w_017_1806, w_017_1807, w_017_1808, w_017_1809, w_017_1810, w_017_1811, w_017_1812, w_017_1813, w_017_1814, w_017_1815, w_017_1816, w_017_1817, w_017_1818, w_017_1819, w_017_1820, w_017_1821, w_017_1822, w_017_1823, w_017_1824, w_017_1825, w_017_1826, w_017_1827, w_017_1828, w_017_1829, w_017_1830, w_017_1831, w_017_1832, w_017_1833, w_017_1834, w_017_1835, w_017_1837, w_017_1838, w_017_1839, w_017_1840, w_017_1841, w_017_1842, w_017_1843, w_017_1844, w_017_1845, w_017_1846, w_017_1847, w_017_1848, w_017_1849, w_017_1850, w_017_1851, w_017_1852, w_017_1853, w_017_1854, w_017_1855, w_017_1856, w_017_1857, w_017_1858, w_017_1861, w_017_1862, w_017_1863, w_017_1864, w_017_1865, w_017_1866, w_017_1867, w_017_1868, w_017_1869, w_017_1870, w_017_1871, w_017_1872, w_017_1874, w_017_1875, w_017_1876, w_017_1877, w_017_1878, w_017_1880, w_017_1881, w_017_1882, w_017_1883, w_017_1884, w_017_1885, w_017_1886, w_017_1887, w_017_1888, w_017_1889, w_017_1890, w_017_1891, w_017_1892, w_017_1893, w_017_1894, w_017_1895, w_017_1896, w_017_1897, w_017_1898, w_017_1899, w_017_1900, w_017_1901, w_017_1902, w_017_1903, w_017_1904, w_017_1905, w_017_1906, w_017_1907, w_017_1908, w_017_1909, w_017_1910, w_017_1911, w_017_1912, w_017_1913, w_017_1914, w_017_1915, w_017_1916, w_017_1918, w_017_1919, w_017_1920, w_017_1921, w_017_1922, w_017_1923, w_017_1924, w_017_1925, w_017_1926, w_017_1927, w_017_1928, w_017_1929, w_017_1930, w_017_1931, w_017_1932, w_017_1933, w_017_1934, w_017_1935, w_017_1936, w_017_1937, w_017_1939, w_017_1940, w_017_1941, w_017_1943, w_017_1944, w_017_1945, w_017_1946, w_017_1947, w_017_1948, w_017_1949, w_017_1950, w_017_1951, w_017_1952, w_017_1953, w_017_1954, w_017_1955, w_017_1956, w_017_1957, w_017_1958, w_017_1959, w_017_1960, w_017_1961, w_017_1962, w_017_1963, w_017_1964, w_017_1965, w_017_1966, w_017_1967, w_017_1968, w_017_1969, w_017_1970, w_017_1971, w_017_1972, w_017_1973, w_017_1974, w_017_1975, w_017_1976, w_017_1977, w_017_1978, w_017_1979, w_017_1980, w_017_1981, w_017_1982, w_017_1983, w_017_1984, w_017_1985, w_017_1987, w_017_1988, w_017_1989, w_017_1990, w_017_1991, w_017_1992, w_017_1993, w_017_1994, w_017_1995, w_017_1996, w_017_1997, w_017_1998, w_017_1999, w_017_2000, w_017_2001, w_017_2002, w_017_2003, w_017_2004, w_017_2005, w_017_2006, w_017_2007, w_017_2008, w_017_2009, w_017_2010, w_017_2011, w_017_2012, w_017_2013, w_017_2014, w_017_2015, w_017_2016, w_017_2017, w_017_2018, w_017_2019, w_017_2020, w_017_2021, w_017_2022, w_017_2023, w_017_2024, w_017_2025, w_017_2026, w_017_2027, w_017_2028, w_017_2029, w_017_2030, w_017_2031, w_017_2032, w_017_2033, w_017_2034, w_017_2035, w_017_2036, w_017_2037, w_017_2038, w_017_2039, w_017_2040, w_017_2041, w_017_2042, w_017_2043, w_017_2044, w_017_2045, w_017_2046, w_017_2047, w_017_2048, w_017_2049, w_017_2050, w_017_2052, w_017_2053, w_017_2054, w_017_2055, w_017_2056, w_017_2057, w_017_2058, w_017_2059, w_017_2060, w_017_2061, w_017_2062, w_017_2063, w_017_2064, w_017_2065, w_017_2066, w_017_2067, w_017_2068, w_017_2069, w_017_2070, w_017_2071, w_017_2072, w_017_2073, w_017_2074, w_017_2075, w_017_2076, w_017_2077, w_017_2078, w_017_2079, w_017_2080, w_017_2081, w_017_2083, w_017_2084, w_017_2085, w_017_2086, w_017_2087, w_017_2088, w_017_2089, w_017_2090, w_017_2091, w_017_2092, w_017_2093, w_017_2094, w_017_2095, w_017_2096, w_017_2097, w_017_2098, w_017_2099, w_017_2100, w_017_2101, w_017_2102, w_017_2103, w_017_2104, w_017_2105, w_017_2106, w_017_2107, w_017_2108, w_017_2109, w_017_2110, w_017_2111, w_017_2112, w_017_2113, w_017_2115, w_017_2116, w_017_2117, w_017_2118, w_017_2119, w_017_2120, w_017_2121, w_017_2122, w_017_2123, w_017_2124, w_017_2125, w_017_2126, w_017_2127, w_017_2128, w_017_2129, w_017_2130, w_017_2131, w_017_2132, w_017_2133, w_017_2134, w_017_2135, w_017_2136, w_017_2137, w_017_2138, w_017_2139, w_017_2140, w_017_2141, w_017_2142, w_017_2143, w_017_2144, w_017_2145, w_017_2146, w_017_2147, w_017_2148, w_017_2149, w_017_2150, w_017_2151, w_017_2152, w_017_2153, w_017_2154, w_017_2155, w_017_2156, w_017_2157, w_017_2158, w_017_2159, w_017_2160, w_017_2161, w_017_2163, w_017_2164, w_017_2165, w_017_2166, w_017_2167, w_017_2168, w_017_2169, w_017_2170, w_017_2171, w_017_2172, w_017_2173, w_017_2174, w_017_2175, w_017_2176, w_017_2177, w_017_2178, w_017_2179, w_017_2181, w_017_2182, w_017_2183, w_017_2184, w_017_2185, w_017_2187, w_017_2188, w_017_2189, w_017_2190, w_017_2191, w_017_2192, w_017_2193, w_017_2194, w_017_2195, w_017_2196, w_017_2197, w_017_2198, w_017_2199, w_017_2200, w_017_2201, w_017_2202, w_017_2203, w_017_2204, w_017_2205, w_017_2206, w_017_2207, w_017_2209, w_017_2210, w_017_2211, w_017_2212, w_017_2213, w_017_2214, w_017_2215, w_017_2216, w_017_2217, w_017_2218, w_017_2219, w_017_2220, w_017_2221, w_017_2222, w_017_2223, w_017_2224, w_017_2225, w_017_2226, w_017_2227, w_017_2228, w_017_2229, w_017_2230, w_017_2231, w_017_2232, w_017_2233, w_017_2234, w_017_2235, w_017_2236, w_017_2237, w_017_2238, w_017_2239, w_017_2240, w_017_2241, w_017_2242, w_017_2243, w_017_2244, w_017_2245, w_017_2246, w_017_2247, w_017_2248, w_017_2249, w_017_2250, w_017_2251, w_017_2252, w_017_2253, w_017_2254, w_017_2255, w_017_2256, w_017_2257, w_017_2258, w_017_2259, w_017_2260, w_017_2261, w_017_2262, w_017_2263, w_017_2264, w_017_2265, w_017_2266, w_017_2267, w_017_2268, w_017_2269, w_017_2270, w_017_2271, w_017_2272, w_017_2273, w_017_2274, w_017_2275, w_017_2276, w_017_2277, w_017_2278, w_017_2279, w_017_2280, w_017_2281, w_017_2282, w_017_2283, w_017_2284, w_017_2285, w_017_2286, w_017_2288, w_017_2289, w_017_2290, w_017_2291, w_017_2292, w_017_2293, w_017_2294, w_017_2295, w_017_2296, w_017_2297, w_017_2298, w_017_2299, w_017_2300, w_017_2301, w_017_2302, w_017_2303, w_017_2304, w_017_2306, w_017_2307, w_017_2308, w_017_2309, w_017_2310, w_017_2311, w_017_2312, w_017_2313, w_017_2314, w_017_2315, w_017_2316, w_017_2317, w_017_2318, w_017_2319, w_017_2320, w_017_2321, w_017_2322, w_017_2323, w_017_2324, w_017_2325, w_017_2326, w_017_2327, w_017_2328, w_017_2329, w_017_2331, w_017_2332, w_017_2334, w_017_2335, w_017_2336, w_017_2337, w_017_2338, w_017_2339, w_017_2340, w_017_2341, w_017_2342, w_017_2343, w_017_2344, w_017_2345, w_017_2346, w_017_2347, w_017_2348, w_017_2349, w_017_2350, w_017_2351, w_017_2352, w_017_2353, w_017_2354, w_017_2355, w_017_2356, w_017_2357, w_017_2358, w_017_2359, w_017_2360, w_017_2361, w_017_2362, w_017_2363, w_017_2364, w_017_2365, w_017_2366, w_017_2367, w_017_2368, w_017_2369, w_017_2370, w_017_2371, w_017_2372, w_017_2373, w_017_2374, w_017_2375, w_017_2376, w_017_2377, w_017_2378, w_017_2379, w_017_2381, w_017_2382, w_017_2383, w_017_2384, w_017_2385, w_017_2386, w_017_2387, w_017_2388, w_017_2389, w_017_2390, w_017_2391, w_017_2392, w_017_2393, w_017_2394, w_017_2395, w_017_2396, w_017_2397, w_017_2398, w_017_2399, w_017_2400, w_017_2401, w_017_2402, w_017_2403, w_017_2404, w_017_2405, w_017_2406, w_017_2407, w_017_2408, w_017_2409, w_017_2410, w_017_2412, w_017_2413, w_017_2414, w_017_2415, w_017_2416, w_017_2417, w_017_2418, w_017_2419, w_017_2421, w_017_2422, w_017_2423, w_017_2424, w_017_2425, w_017_2426, w_017_2427, w_017_2428, w_017_2429, w_017_2430, w_017_2431, w_017_2432, w_017_2433, w_017_2434, w_017_2435, w_017_2436, w_017_2437, w_017_2438, w_017_2439, w_017_2440, w_017_2441, w_017_2442, w_017_2443, w_017_2444, w_017_2446, w_017_2447, w_017_2448, w_017_2449, w_017_2450, w_017_2451, w_017_2452, w_017_2454, w_017_2455, w_017_2456, w_017_2457, w_017_2458, w_017_2459, w_017_2460, w_017_2461, w_017_2462, w_017_2463, w_017_2464, w_017_2465, w_017_2466, w_017_2467, w_017_2469, w_017_2470, w_017_2471, w_017_2472, w_017_2473, w_017_2474, w_017_2475, w_017_2476, w_017_2477, w_017_2479, w_017_2480, w_017_2481, w_017_2482, w_017_2483, w_017_2484, w_017_2485, w_017_2486, w_017_2487, w_017_2488, w_017_2489, w_017_2490, w_017_2491, w_017_2492, w_017_2493, w_017_2494, w_017_2495, w_017_2496, w_017_2497, w_017_2498, w_017_2499, w_017_2500, w_017_2501, w_017_2502, w_017_2503, w_017_2504, w_017_2505, w_017_2506, w_017_2507, w_017_2508, w_017_2509, w_017_2510, w_017_2511, w_017_2512, w_017_2513, w_017_2514, w_017_2515, w_017_2516, w_017_2517, w_017_2518, w_017_2519, w_017_2520, w_017_2521, w_017_2522, w_017_2523, w_017_2524, w_017_2526, w_017_2527, w_017_2528, w_017_2529, w_017_2530, w_017_2531, w_017_2532, w_017_2533, w_017_2534, w_017_2535, w_017_2536, w_017_2537, w_017_2538, w_017_2539, w_017_2540, w_017_2541, w_017_2542, w_017_2543, w_017_2544, w_017_2545, w_017_2546, w_017_2547, w_017_2548, w_017_2549, w_017_2550, w_017_2551, w_017_2552, w_017_2553, w_017_2554, w_017_2555, w_017_2556, w_017_2557, w_017_2558, w_017_2559, w_017_2560, w_017_2561, w_017_2562, w_017_2563, w_017_2564, w_017_2565, w_017_2566, w_017_2567, w_017_2568, w_017_2569, w_017_2570, w_017_2571, w_017_2572, w_017_2573, w_017_2574, w_017_2576, w_017_2577, w_017_2578, w_017_2580, w_017_2581, w_017_2582, w_017_2583, w_017_2584, w_017_2585, w_017_2586, w_017_2588, w_017_2589, w_017_2590, w_017_2591, w_017_2592, w_017_2593, w_017_2594, w_017_2595, w_017_2596, w_017_2597, w_017_2598, w_017_2599, w_017_2600, w_017_2601, w_017_2602, w_017_2603, w_017_2604, w_017_2605, w_017_2606, w_017_2607, w_017_2608, w_017_2609, w_017_2610, w_017_2611, w_017_2612, w_017_2613, w_017_2614, w_017_2615, w_017_2616, w_017_2617, w_017_2618, w_017_2619, w_017_2620, w_017_2621, w_017_2622, w_017_2623, w_017_2624, w_017_2625, w_017_2626, w_017_2627, w_017_2628, w_017_2629, w_017_2630, w_017_2631, w_017_2632, w_017_2633, w_017_2634, w_017_2635, w_017_2636, w_017_2637, w_017_2639, w_017_2640, w_017_2641, w_017_2642, w_017_2643, w_017_2644, w_017_2645, w_017_2646, w_017_2647, w_017_2648, w_017_2649, w_017_2650, w_017_2651, w_017_2652, w_017_2654, w_017_2655, w_017_2656, w_017_2657, w_017_2658, w_017_2659, w_017_2660, w_017_2661, w_017_2662, w_017_2663, w_017_2664, w_017_2666, w_017_2667, w_017_2668, w_017_2669, w_017_2670, w_017_2671, w_017_2672, w_017_2673, w_017_2674, w_017_2675, w_017_2676, w_017_2677, w_017_2678, w_017_2679, w_017_2680, w_017_2681, w_017_2683, w_017_2684, w_017_2685, w_017_2686, w_017_2687, w_017_2688, w_017_2689, w_017_2690, w_017_2691, w_017_2692, w_017_2693, w_017_2694, w_017_2695, w_017_2696, w_017_2697, w_017_2698, w_017_2699, w_017_2700, w_017_2701, w_017_2702, w_017_2703, w_017_2704, w_017_2705, w_017_2706, w_017_2707, w_017_2708, w_017_2709, w_017_2710, w_017_2711, w_017_2712, w_017_2714, w_017_2715, w_017_2716, w_017_2717, w_017_2718, w_017_2719, w_017_2720, w_017_2721, w_017_2722, w_017_2723, w_017_2724, w_017_2725, w_017_2726, w_017_2727, w_017_2728, w_017_2729, w_017_2731, w_017_2732, w_017_2734, w_017_2735, w_017_2736, w_017_2737, w_017_2738, w_017_2739, w_017_2740, w_017_2741, w_017_2742, w_017_2743, w_017_2744, w_017_2745, w_017_2746, w_017_2747, w_017_2748, w_017_2749, w_017_2750, w_017_2751, w_017_2753, w_017_2754, w_017_2755, w_017_2756, w_017_2757, w_017_2758, w_017_2759, w_017_2760, w_017_2761, w_017_2762, w_017_2763, w_017_2764, w_017_2765, w_017_2766, w_017_2767, w_017_2768, w_017_2769, w_017_2770, w_017_2771, w_017_2772, w_017_2773, w_017_2774, w_017_2775, w_017_2776, w_017_2777, w_017_2778, w_017_2779, w_017_2780, w_017_2781, w_017_2782, w_017_2783, w_017_2784, w_017_2785, w_017_2786, w_017_2788, w_017_2789, w_017_2790, w_017_2791, w_017_2792, w_017_2793, w_017_2794, w_017_2795, w_017_2796, w_017_2797, w_017_2798, w_017_2799, w_017_2801, w_017_2802, w_017_2803, w_017_2804, w_017_2805, w_017_2806, w_017_2807, w_017_2808, w_017_2809, w_017_2810, w_017_2811, w_017_2812, w_017_2813, w_017_2814, w_017_2815, w_017_2816, w_017_2817, w_017_2818, w_017_2819, w_017_2820, w_017_2821, w_017_2822, w_017_2823, w_017_2824, w_017_2825, w_017_2826, w_017_2827, w_017_2828, w_017_2829, w_017_2830, w_017_2831, w_017_2832, w_017_2833, w_017_2834, w_017_2835, w_017_2836, w_017_2837, w_017_2838, w_017_2839, w_017_2840, w_017_2841, w_017_2842, w_017_2843, w_017_2844, w_017_2845, w_017_2846, w_017_2847, w_017_2848, w_017_2849, w_017_2850, w_017_2851, w_017_2852, w_017_2853, w_017_2854, w_017_2855, w_017_2856, w_017_2857, w_017_2858, w_017_2859, w_017_2860, w_017_2861, w_017_2862, w_017_2863, w_017_2865, w_017_2866, w_017_2867, w_017_2868, w_017_2869, w_017_2870, w_017_2871, w_017_2872, w_017_2873, w_017_2874, w_017_2875, w_017_2876, w_017_2877, w_017_2878, w_017_2879, w_017_2880, w_017_2881, w_017_2882, w_017_2883, w_017_2884, w_017_2885, w_017_2886, w_017_2887, w_017_2888, w_017_2889, w_017_2890, w_017_2891, w_017_2892, w_017_2893, w_017_2894, w_017_2895, w_017_2896, w_017_2897, w_017_2898, w_017_2899, w_017_2900, w_017_2901, w_017_2902, w_017_2903, w_017_2904, w_017_2905, w_017_2906, w_017_2907, w_017_2908, w_017_2909, w_017_2910, w_017_2911, w_017_2912, w_017_2913, w_017_2914, w_017_2915, w_017_2916, w_017_2917, w_017_2918, w_017_2919, w_017_2920, w_017_2921, w_017_2922, w_017_2923, w_017_2924, w_017_2925, w_017_2926, w_017_2927, w_017_2928, w_017_2929, w_017_2930, w_017_2931, w_017_2932, w_017_2933, w_017_2934, w_017_2935, w_017_2936, w_017_2937, w_017_2938, w_017_2939, w_017_2940, w_017_2941, w_017_2942, w_017_2943, w_017_2944, w_017_2945, w_017_2946, w_017_2947, w_017_2948, w_017_2949, w_017_2950, w_017_2951, w_017_2952, w_017_2953, w_017_2954, w_017_2955, w_017_2956, w_017_2957, w_017_2958, w_017_2959, w_017_2961, w_017_2962, w_017_2963, w_017_2965, w_017_2966, w_017_2967, w_017_2968, w_017_2969, w_017_2970, w_017_2971, w_017_2972, w_017_2973, w_017_2974, w_017_2975, w_017_2976, w_017_2977, w_017_2978, w_017_2979, w_017_2980, w_017_2981, w_017_2982, w_017_2983, w_017_2984, w_017_2985, w_017_2986, w_017_2987, w_017_2988, w_017_2989, w_017_2990, w_017_2991, w_017_2992, w_017_2993, w_017_2994, w_017_2995, w_017_2996, w_017_2997, w_017_2998, w_017_2999, w_017_3000, w_017_3001, w_017_3002, w_017_3003, w_017_3004, w_017_3005, w_017_3006, w_017_3007, w_017_3008, w_017_3009, w_017_3010, w_017_3011, w_017_3012, w_017_3013, w_017_3014, w_017_3016, w_017_3017, w_017_3018, w_017_3019, w_017_3020, w_017_3021, w_017_3022, w_017_3023, w_017_3024, w_017_3025, w_017_3026, w_017_3027, w_017_3028, w_017_3029, w_017_3030, w_017_3031, w_017_3032, w_017_3033, w_017_3034, w_017_3035, w_017_3036, w_017_3037, w_017_3038, w_017_3039, w_017_3040, w_017_3041, w_017_3042, w_017_3043, w_017_3044, w_017_3045, w_017_3046, w_017_3047, w_017_3048, w_017_3049, w_017_3050, w_017_3051, w_017_3052, w_017_3053, w_017_3054, w_017_3055, w_017_3056, w_017_3057, w_017_3058, w_017_3059, w_017_3060, w_017_3061, w_017_3062, w_017_3063, w_017_3064, w_017_3065, w_017_3066, w_017_3067, w_017_3068, w_017_3069, w_017_3070, w_017_3072, w_017_3073, w_017_3074, w_017_3075, w_017_3076, w_017_3077, w_017_3078, w_017_3079, w_017_3080, w_017_3081, w_017_3082, w_017_3083, w_017_3084, w_017_3085, w_017_3086, w_017_3087, w_017_3088, w_017_3089, w_017_3090, w_017_3091, w_017_3092, w_017_3093, w_017_3094, w_017_3095, w_017_3096, w_017_3097, w_017_3098, w_017_3099, w_017_3100, w_017_3101, w_017_3102, w_017_3103, w_017_3104, w_017_3105, w_017_3106, w_017_3107, w_017_3108, w_017_3109, w_017_3110, w_017_3111, w_017_3112, w_017_3113, w_017_3114, w_017_3115, w_017_3116, w_017_3117, w_017_3118, w_017_3119, w_017_3120, w_017_3121, w_017_3122, w_017_3123, w_017_3124, w_017_3125, w_017_3126, w_017_3127, w_017_3129, w_017_3130, w_017_3131, w_017_3132, w_017_3134, w_017_3135, w_017_3136, w_017_3137, w_017_3138, w_017_3139, w_017_3140, w_017_3141, w_017_3142, w_017_3143, w_017_3144, w_017_3145, w_017_3146, w_017_3147, w_017_3148, w_017_3149, w_017_3150, w_017_3151, w_017_3152, w_017_3153, w_017_3154, w_017_3155, w_017_3157, w_017_3158, w_017_3159, w_017_3160, w_017_3161, w_017_3162, w_017_3163, w_017_3164, w_017_3165, w_017_3166, w_017_3168, w_017_3169, w_017_3171, w_017_3172, w_017_3173, w_017_3174, w_017_3175, w_017_3176, w_017_3177, w_017_3178, w_017_3179, w_017_3180, w_017_3181, w_017_3182, w_017_3183, w_017_3184, w_017_3185, w_017_3186, w_017_3187, w_017_3188, w_017_3189, w_017_3190, w_017_3191, w_017_3192, w_017_3193, w_017_3194, w_017_3195, w_017_3196, w_017_3197, w_017_3198, w_017_3199, w_017_3200, w_017_3201, w_017_3202, w_017_3203, w_017_3204, w_017_3205, w_017_3206, w_017_3207, w_017_3208, w_017_3209, w_017_3210, w_017_3211, w_017_3212, w_017_3213, w_017_3214, w_017_3215, w_017_3216, w_017_3217, w_017_3218, w_017_3219, w_017_3220, w_017_3221, w_017_3222, w_017_3223, w_017_3224, w_017_3225, w_017_3226, w_017_3227, w_017_3228, w_017_3229, w_017_3230, w_017_3231, w_017_3232, w_017_3233, w_017_3234, w_017_3235, w_017_3236, w_017_3238, w_017_3239, w_017_3240, w_017_3241, w_017_3242, w_017_3243, w_017_3244, w_017_3245, w_017_3246, w_017_3247, w_017_3248, w_017_3249, w_017_3250, w_017_3251, w_017_3252, w_017_3254, w_017_3255, w_017_3256, w_017_3257, w_017_3258, w_017_3259, w_017_3260, w_017_3261, w_017_3262, w_017_3263, w_017_3264, w_017_3265, w_017_3266, w_017_3267, w_017_3268, w_017_3269;
  wire w_018_000, w_018_001, w_018_002, w_018_003, w_018_004, w_018_005, w_018_006, w_018_007, w_018_008, w_018_009, w_018_010, w_018_011, w_018_012, w_018_013, w_018_014, w_018_015, w_018_016, w_018_017, w_018_019, w_018_020, w_018_021, w_018_022, w_018_023, w_018_024, w_018_025, w_018_026, w_018_027, w_018_028, w_018_029, w_018_030, w_018_031, w_018_032, w_018_033, w_018_034, w_018_035, w_018_036, w_018_037, w_018_038, w_018_039, w_018_040, w_018_041, w_018_043, w_018_044, w_018_045, w_018_046, w_018_047, w_018_048, w_018_049, w_018_050, w_018_051, w_018_052, w_018_053, w_018_054, w_018_055, w_018_056, w_018_057, w_018_058, w_018_059, w_018_060, w_018_061, w_018_062, w_018_063, w_018_064, w_018_065, w_018_066, w_018_067, w_018_068, w_018_069, w_018_070, w_018_071, w_018_072, w_018_073, w_018_074, w_018_075, w_018_076, w_018_077, w_018_078, w_018_079, w_018_080, w_018_081, w_018_082, w_018_083, w_018_084, w_018_085, w_018_086, w_018_087, w_018_088, w_018_089, w_018_090, w_018_091, w_018_092, w_018_093, w_018_094, w_018_095, w_018_096, w_018_097, w_018_098, w_018_099, w_018_100, w_018_101, w_018_102, w_018_103, w_018_104, w_018_105, w_018_106, w_018_107, w_018_108, w_018_109, w_018_110, w_018_111, w_018_112, w_018_113, w_018_114, w_018_115, w_018_116, w_018_117, w_018_118, w_018_119, w_018_120, w_018_121, w_018_122, w_018_123, w_018_124, w_018_125, w_018_126, w_018_127, w_018_128, w_018_129, w_018_130, w_018_131, w_018_132, w_018_133, w_018_134, w_018_135, w_018_136, w_018_137, w_018_138, w_018_139, w_018_140, w_018_141, w_018_142, w_018_143, w_018_144, w_018_145, w_018_146, w_018_147, w_018_148, w_018_149, w_018_150, w_018_151, w_018_152, w_018_153, w_018_154, w_018_155, w_018_156, w_018_157, w_018_158, w_018_159, w_018_160, w_018_161, w_018_162, w_018_163, w_018_164, w_018_165, w_018_166, w_018_167, w_018_168, w_018_169, w_018_170, w_018_171, w_018_172, w_018_173, w_018_174, w_018_175, w_018_176, w_018_177, w_018_178, w_018_179, w_018_180, w_018_181, w_018_182, w_018_183, w_018_184, w_018_185, w_018_186, w_018_187, w_018_188, w_018_189, w_018_190, w_018_191, w_018_192, w_018_193, w_018_194, w_018_195, w_018_196, w_018_197, w_018_198, w_018_199, w_018_200, w_018_201, w_018_202, w_018_203, w_018_204, w_018_205, w_018_206, w_018_207, w_018_208, w_018_209, w_018_210, w_018_211, w_018_212, w_018_213, w_018_214, w_018_215, w_018_216, w_018_217, w_018_218, w_018_219, w_018_220, w_018_221, w_018_222, w_018_223, w_018_224, w_018_225, w_018_226, w_018_227, w_018_228, w_018_229, w_018_230, w_018_231, w_018_232, w_018_233, w_018_234, w_018_235, w_018_236, w_018_238, w_018_239, w_018_240, w_018_241, w_018_242, w_018_243, w_018_244, w_018_245, w_018_246, w_018_247, w_018_248, w_018_249, w_018_250, w_018_251, w_018_252, w_018_253, w_018_254, w_018_255, w_018_256, w_018_257, w_018_258, w_018_259, w_018_260, w_018_261, w_018_262, w_018_263, w_018_264, w_018_265, w_018_266, w_018_267, w_018_268, w_018_269, w_018_270, w_018_271, w_018_272, w_018_273, w_018_274, w_018_275, w_018_276, w_018_277, w_018_278, w_018_279, w_018_280, w_018_281, w_018_282, w_018_283, w_018_284, w_018_285, w_018_286, w_018_287, w_018_288, w_018_289, w_018_290, w_018_291, w_018_292, w_018_293, w_018_294, w_018_295, w_018_296, w_018_297, w_018_298, w_018_299, w_018_300, w_018_301, w_018_302, w_018_303, w_018_304, w_018_305, w_018_306, w_018_307, w_018_308, w_018_309, w_018_310, w_018_312, w_018_313, w_018_314, w_018_315, w_018_316, w_018_317, w_018_318, w_018_319, w_018_320, w_018_321, w_018_322, w_018_323, w_018_324, w_018_325, w_018_326, w_018_327, w_018_328, w_018_329, w_018_330, w_018_331, w_018_332, w_018_333, w_018_334, w_018_335, w_018_336, w_018_337, w_018_338, w_018_339, w_018_340, w_018_341, w_018_342, w_018_343, w_018_344, w_018_345, w_018_346, w_018_347, w_018_348, w_018_349, w_018_350, w_018_351, w_018_352, w_018_353, w_018_355, w_018_356, w_018_357, w_018_358, w_018_359, w_018_360, w_018_361, w_018_362, w_018_363, w_018_364, w_018_365, w_018_366, w_018_367, w_018_368, w_018_370, w_018_371, w_018_372, w_018_373, w_018_374, w_018_375, w_018_376, w_018_377, w_018_378, w_018_379, w_018_380, w_018_381, w_018_382, w_018_383, w_018_384, w_018_385, w_018_386, w_018_387, w_018_388, w_018_389, w_018_390, w_018_391, w_018_392, w_018_393, w_018_394, w_018_395, w_018_396, w_018_397, w_018_398, w_018_399, w_018_400, w_018_401, w_018_402, w_018_403, w_018_404, w_018_405, w_018_406, w_018_407, w_018_408, w_018_409, w_018_410, w_018_411, w_018_412, w_018_413, w_018_414, w_018_415, w_018_416, w_018_417, w_018_418, w_018_419, w_018_420, w_018_421, w_018_422, w_018_423, w_018_424, w_018_425, w_018_426, w_018_427, w_018_428, w_018_429, w_018_430, w_018_431, w_018_432, w_018_433, w_018_435, w_018_436, w_018_437, w_018_438, w_018_440, w_018_441, w_018_442, w_018_443, w_018_444, w_018_445, w_018_446, w_018_447, w_018_448, w_018_449, w_018_450, w_018_451, w_018_452, w_018_453, w_018_454, w_018_455, w_018_456, w_018_457, w_018_458, w_018_459, w_018_460, w_018_461, w_018_462, w_018_463, w_018_464, w_018_465, w_018_466, w_018_468, w_018_469, w_018_470, w_018_471, w_018_472, w_018_473, w_018_474, w_018_475, w_018_476, w_018_477, w_018_478, w_018_479, w_018_480, w_018_481, w_018_482, w_018_483, w_018_484, w_018_485, w_018_486, w_018_487, w_018_488, w_018_489, w_018_490, w_018_491, w_018_492, w_018_493, w_018_494, w_018_495, w_018_496, w_018_497, w_018_498, w_018_499, w_018_500, w_018_501, w_018_502, w_018_503, w_018_504, w_018_505, w_018_506, w_018_507, w_018_508, w_018_509, w_018_510, w_018_511, w_018_512, w_018_513, w_018_514, w_018_515, w_018_516, w_018_517, w_018_518, w_018_519, w_018_520, w_018_521, w_018_522, w_018_523, w_018_524, w_018_525, w_018_526, w_018_527, w_018_528, w_018_529, w_018_530, w_018_531, w_018_532, w_018_533, w_018_534, w_018_535, w_018_536, w_018_537, w_018_538, w_018_539, w_018_540, w_018_541, w_018_542, w_018_543, w_018_544, w_018_545, w_018_546, w_018_547, w_018_548, w_018_549, w_018_550, w_018_551, w_018_552, w_018_553, w_018_554, w_018_555, w_018_556, w_018_557, w_018_558, w_018_559, w_018_560, w_018_561, w_018_562, w_018_563, w_018_565, w_018_566, w_018_567, w_018_568, w_018_569, w_018_571, w_018_572, w_018_573, w_018_574, w_018_575, w_018_576, w_018_577, w_018_578, w_018_579, w_018_580, w_018_581, w_018_582, w_018_583, w_018_584, w_018_585, w_018_586, w_018_587, w_018_588, w_018_589, w_018_590, w_018_591, w_018_592, w_018_593, w_018_594, w_018_595, w_018_596, w_018_597, w_018_599, w_018_600, w_018_601, w_018_602, w_018_603, w_018_604, w_018_605, w_018_606, w_018_607, w_018_608, w_018_609, w_018_610, w_018_611, w_018_612, w_018_613, w_018_614, w_018_615, w_018_616, w_018_617, w_018_618, w_018_619, w_018_620, w_018_621, w_018_622, w_018_623, w_018_624, w_018_625, w_018_626, w_018_627, w_018_628, w_018_629, w_018_630, w_018_631, w_018_632, w_018_633, w_018_634, w_018_635, w_018_636, w_018_637, w_018_638, w_018_639, w_018_640, w_018_641, w_018_642, w_018_643, w_018_644, w_018_645, w_018_646, w_018_647, w_018_648, w_018_649, w_018_650, w_018_652, w_018_653, w_018_654, w_018_655, w_018_656, w_018_657, w_018_658, w_018_659, w_018_660, w_018_661, w_018_662, w_018_663, w_018_664, w_018_665, w_018_666, w_018_667, w_018_668, w_018_669, w_018_670, w_018_671, w_018_672, w_018_673, w_018_674, w_018_675, w_018_676, w_018_677, w_018_678, w_018_679, w_018_680, w_018_681, w_018_682, w_018_683, w_018_684, w_018_685, w_018_686, w_018_687, w_018_688, w_018_689, w_018_690, w_018_691, w_018_692, w_018_693, w_018_694, w_018_695, w_018_696, w_018_697, w_018_698, w_018_699, w_018_700, w_018_701, w_018_703, w_018_704, w_018_706, w_018_708, w_018_709, w_018_710, w_018_711, w_018_712, w_018_713, w_018_714, w_018_715, w_018_716, w_018_717, w_018_718, w_018_719, w_018_720, w_018_721, w_018_722, w_018_723, w_018_724, w_018_726, w_018_727, w_018_728, w_018_729, w_018_730, w_018_731, w_018_733, w_018_734, w_018_735, w_018_736, w_018_737, w_018_738, w_018_739, w_018_740, w_018_741, w_018_742, w_018_743, w_018_744, w_018_745, w_018_746, w_018_747, w_018_748, w_018_750, w_018_751, w_018_752, w_018_753, w_018_754, w_018_755, w_018_756, w_018_757, w_018_758, w_018_759, w_018_760, w_018_762, w_018_763, w_018_764, w_018_765, w_018_766, w_018_767, w_018_769, w_018_771, w_018_772, w_018_773, w_018_774, w_018_775, w_018_776, w_018_777, w_018_778, w_018_779, w_018_781, w_018_782, w_018_783, w_018_784, w_018_785, w_018_786, w_018_787, w_018_788, w_018_789, w_018_790, w_018_791, w_018_792, w_018_793, w_018_794, w_018_796, w_018_797, w_018_798, w_018_799, w_018_800, w_018_801, w_018_802, w_018_803, w_018_804, w_018_805, w_018_806, w_018_807, w_018_808, w_018_809, w_018_810, w_018_811, w_018_812, w_018_813, w_018_814, w_018_815, w_018_816, w_018_817, w_018_818, w_018_819, w_018_820, w_018_821, w_018_823, w_018_824, w_018_825, w_018_826, w_018_827, w_018_828, w_018_830, w_018_831, w_018_832, w_018_833, w_018_834, w_018_835, w_018_836, w_018_837, w_018_838, w_018_840, w_018_841, w_018_842, w_018_844, w_018_845, w_018_846, w_018_847, w_018_848, w_018_849, w_018_850, w_018_851, w_018_852, w_018_853, w_018_854, w_018_855, w_018_856, w_018_857, w_018_858, w_018_859, w_018_860, w_018_861, w_018_862, w_018_863, w_018_864, w_018_865, w_018_866, w_018_867, w_018_868, w_018_869, w_018_870, w_018_871, w_018_872, w_018_873, w_018_874, w_018_875, w_018_876, w_018_877, w_018_878, w_018_879, w_018_880, w_018_881, w_018_883, w_018_884, w_018_885, w_018_886, w_018_887, w_018_888, w_018_889, w_018_890, w_018_891, w_018_892, w_018_893, w_018_894, w_018_895, w_018_896, w_018_897, w_018_898, w_018_899, w_018_900, w_018_901, w_018_902, w_018_903, w_018_904, w_018_905, w_018_907, w_018_908, w_018_909, w_018_910, w_018_911, w_018_912, w_018_913, w_018_914, w_018_915, w_018_916, w_018_917, w_018_918, w_018_919, w_018_920, w_018_921, w_018_922, w_018_923, w_018_924, w_018_925, w_018_926, w_018_927, w_018_928, w_018_929, w_018_930, w_018_932, w_018_933, w_018_935, w_018_936, w_018_937, w_018_938, w_018_939, w_018_940, w_018_941, w_018_942, w_018_943, w_018_944, w_018_945, w_018_946, w_018_947, w_018_948, w_018_949, w_018_951, w_018_952, w_018_953, w_018_954, w_018_955, w_018_956, w_018_957, w_018_958, w_018_959, w_018_960, w_018_961, w_018_962, w_018_963, w_018_964, w_018_965, w_018_966, w_018_967, w_018_968, w_018_969, w_018_970, w_018_971, w_018_972, w_018_973, w_018_974, w_018_975, w_018_976, w_018_977, w_018_978, w_018_979, w_018_980, w_018_981, w_018_982, w_018_983, w_018_984, w_018_985, w_018_986, w_018_987, w_018_988, w_018_989, w_018_990, w_018_991, w_018_992, w_018_993, w_018_994, w_018_995, w_018_996, w_018_997, w_018_998, w_018_999, w_018_1000, w_018_1001, w_018_1002, w_018_1003, w_018_1004, w_018_1005, w_018_1006, w_018_1007, w_018_1008, w_018_1009, w_018_1010, w_018_1011, w_018_1012, w_018_1013, w_018_1014, w_018_1015, w_018_1016, w_018_1018, w_018_1019, w_018_1020, w_018_1021, w_018_1022, w_018_1023, w_018_1024, w_018_1025, w_018_1026, w_018_1027, w_018_1028, w_018_1029, w_018_1030, w_018_1031, w_018_1032, w_018_1033, w_018_1034, w_018_1036, w_018_1037, w_018_1038, w_018_1039, w_018_1040, w_018_1041, w_018_1042, w_018_1043, w_018_1044, w_018_1045, w_018_1046, w_018_1047, w_018_1048, w_018_1049, w_018_1050, w_018_1051, w_018_1052, w_018_1053, w_018_1054, w_018_1055, w_018_1056, w_018_1057, w_018_1058, w_018_1061, w_018_1063, w_018_1064, w_018_1065, w_018_1066, w_018_1067, w_018_1068, w_018_1069, w_018_1070, w_018_1071, w_018_1072, w_018_1073, w_018_1074, w_018_1075, w_018_1076, w_018_1077, w_018_1078, w_018_1080, w_018_1081, w_018_1082, w_018_1083, w_018_1084, w_018_1085, w_018_1086, w_018_1087, w_018_1088, w_018_1089, w_018_1091, w_018_1092, w_018_1093, w_018_1094, w_018_1096, w_018_1097, w_018_1098, w_018_1099, w_018_1100, w_018_1101, w_018_1103, w_018_1104, w_018_1105, w_018_1107, w_018_1108, w_018_1109, w_018_1110, w_018_1111, w_018_1112, w_018_1113, w_018_1114, w_018_1115, w_018_1116, w_018_1117, w_018_1118, w_018_1119, w_018_1120, w_018_1121, w_018_1122, w_018_1123, w_018_1124, w_018_1125, w_018_1126, w_018_1127, w_018_1128, w_018_1129, w_018_1130, w_018_1131, w_018_1132, w_018_1134, w_018_1135, w_018_1136, w_018_1137, w_018_1138, w_018_1139, w_018_1140, w_018_1141, w_018_1142, w_018_1143, w_018_1144, w_018_1145, w_018_1146, w_018_1147, w_018_1148, w_018_1149, w_018_1150, w_018_1151, w_018_1152, w_018_1153, w_018_1154, w_018_1156, w_018_1157, w_018_1158, w_018_1159, w_018_1160, w_018_1161, w_018_1162, w_018_1163, w_018_1164, w_018_1165, w_018_1166, w_018_1167, w_018_1168, w_018_1169, w_018_1170, w_018_1171, w_018_1173, w_018_1174, w_018_1176, w_018_1177, w_018_1178, w_018_1179, w_018_1180, w_018_1181, w_018_1182, w_018_1183, w_018_1184, w_018_1185, w_018_1186, w_018_1187, w_018_1188, w_018_1189, w_018_1190, w_018_1191, w_018_1192, w_018_1193, w_018_1194, w_018_1195, w_018_1196, w_018_1197, w_018_1198, w_018_1199, w_018_1200, w_018_1201, w_018_1202, w_018_1203, w_018_1204, w_018_1205, w_018_1206, w_018_1207, w_018_1208, w_018_1209, w_018_1210, w_018_1211, w_018_1212, w_018_1213, w_018_1214, w_018_1215, w_018_1216, w_018_1217, w_018_1218, w_018_1219, w_018_1220, w_018_1221, w_018_1222, w_018_1223, w_018_1224, w_018_1225, w_018_1226, w_018_1227, w_018_1228, w_018_1229, w_018_1230, w_018_1231, w_018_1232, w_018_1233, w_018_1234, w_018_1235, w_018_1237, w_018_1238, w_018_1239, w_018_1240, w_018_1241, w_018_1242, w_018_1243, w_018_1244, w_018_1245, w_018_1246, w_018_1247, w_018_1248, w_018_1249, w_018_1250, w_018_1251, w_018_1252, w_018_1253, w_018_1254, w_018_1255, w_018_1256, w_018_1257, w_018_1258, w_018_1259, w_018_1260, w_018_1262, w_018_1263, w_018_1264, w_018_1265, w_018_1266, w_018_1267, w_018_1268, w_018_1269, w_018_1270, w_018_1271, w_018_1272, w_018_1273, w_018_1274, w_018_1275, w_018_1276, w_018_1277, w_018_1278, w_018_1280, w_018_1281, w_018_1282, w_018_1283, w_018_1284, w_018_1285, w_018_1286, w_018_1287, w_018_1288, w_018_1290, w_018_1291, w_018_1292, w_018_1293, w_018_1294, w_018_1295, w_018_1296, w_018_1297, w_018_1298, w_018_1299, w_018_1300, w_018_1301, w_018_1302, w_018_1303, w_018_1304, w_018_1305, w_018_1306, w_018_1307, w_018_1308, w_018_1309, w_018_1310, w_018_1311, w_018_1312, w_018_1313, w_018_1314, w_018_1315, w_018_1316, w_018_1317, w_018_1318, w_018_1319, w_018_1320, w_018_1321, w_018_1322, w_018_1323, w_018_1324, w_018_1325, w_018_1326, w_018_1327, w_018_1328, w_018_1329, w_018_1330, w_018_1331, w_018_1332, w_018_1333, w_018_1334, w_018_1335, w_018_1336, w_018_1337, w_018_1338, w_018_1339, w_018_1340, w_018_1341, w_018_1342, w_018_1343, w_018_1344, w_018_1345, w_018_1346, w_018_1347, w_018_1348, w_018_1349, w_018_1350, w_018_1351, w_018_1352, w_018_1353, w_018_1354, w_018_1355, w_018_1356, w_018_1357, w_018_1358, w_018_1359, w_018_1360, w_018_1361, w_018_1362, w_018_1363, w_018_1364, w_018_1366, w_018_1367, w_018_1368, w_018_1369, w_018_1370, w_018_1371, w_018_1372, w_018_1373, w_018_1374, w_018_1375, w_018_1376, w_018_1377, w_018_1378, w_018_1379, w_018_1380, w_018_1381, w_018_1382, w_018_1383, w_018_1384, w_018_1385, w_018_1386, w_018_1387, w_018_1388, w_018_1389, w_018_1390, w_018_1391, w_018_1392, w_018_1393, w_018_1394, w_018_1395, w_018_1396, w_018_1397, w_018_1398, w_018_1399, w_018_1400, w_018_1401, w_018_1402, w_018_1403, w_018_1404, w_018_1405, w_018_1406, w_018_1407, w_018_1408, w_018_1409, w_018_1410, w_018_1411, w_018_1412, w_018_1413, w_018_1414, w_018_1415, w_018_1416, w_018_1417, w_018_1418, w_018_1419, w_018_1420, w_018_1421, w_018_1422, w_018_1423, w_018_1424, w_018_1425, w_018_1427, w_018_1429, w_018_1430, w_018_1431, w_018_1432, w_018_1433, w_018_1434, w_018_1435, w_018_1436, w_018_1437, w_018_1439, w_018_1440, w_018_1441, w_018_1442, w_018_1443, w_018_1444, w_018_1445, w_018_1446, w_018_1447, w_018_1448, w_018_1449, w_018_1450, w_018_1451, w_018_1452, w_018_1453, w_018_1454, w_018_1455, w_018_1456, w_018_1457, w_018_1458, w_018_1459, w_018_1460, w_018_1461, w_018_1462, w_018_1463, w_018_1464, w_018_1465, w_018_1466, w_018_1467, w_018_1468, w_018_1469, w_018_1470, w_018_1471, w_018_1472, w_018_1473, w_018_1474, w_018_1475, w_018_1476, w_018_1477, w_018_1478, w_018_1479, w_018_1480, w_018_1481, w_018_1482, w_018_1483, w_018_1484, w_018_1485, w_018_1486, w_018_1488, w_018_1489, w_018_1490, w_018_1491, w_018_1492, w_018_1493, w_018_1494, w_018_1495, w_018_1496, w_018_1497, w_018_1498, w_018_1499, w_018_1500, w_018_1501, w_018_1502, w_018_1504, w_018_1505, w_018_1506, w_018_1507, w_018_1508, w_018_1509, w_018_1510, w_018_1511, w_018_1512, w_018_1513, w_018_1514, w_018_1515, w_018_1516, w_018_1517, w_018_1518, w_018_1519, w_018_1520, w_018_1521, w_018_1522, w_018_1523, w_018_1524, w_018_1525, w_018_1526, w_018_1527, w_018_1528, w_018_1529, w_018_1530, w_018_1531, w_018_1532, w_018_1533, w_018_1534, w_018_1535, w_018_1536, w_018_1537, w_018_1538, w_018_1539, w_018_1540, w_018_1542, w_018_1543, w_018_1544, w_018_1545, w_018_1546, w_018_1547, w_018_1548, w_018_1549, w_018_1550, w_018_1551, w_018_1552, w_018_1553, w_018_1554, w_018_1555, w_018_1556, w_018_1557, w_018_1558, w_018_1559, w_018_1560, w_018_1561, w_018_1562, w_018_1563, w_018_1564, w_018_1565, w_018_1566, w_018_1567, w_018_1568, w_018_1569, w_018_1570, w_018_1571, w_018_1572, w_018_1573, w_018_1574, w_018_1575, w_018_1576, w_018_1577, w_018_1578, w_018_1580, w_018_1581, w_018_1582, w_018_1583, w_018_1584, w_018_1585, w_018_1586, w_018_1587, w_018_1588, w_018_1589, w_018_1590, w_018_1591, w_018_1592, w_018_1593, w_018_1594, w_018_1595, w_018_1596, w_018_1597, w_018_1599, w_018_1600, w_018_1601, w_018_1602, w_018_1603, w_018_1605, w_018_1606, w_018_1607, w_018_1608, w_018_1609, w_018_1610, w_018_1611, w_018_1612, w_018_1613, w_018_1614, w_018_1615, w_018_1616, w_018_1618, w_018_1619, w_018_1621, w_018_1622, w_018_1623, w_018_1624, w_018_1625, w_018_1626, w_018_1627, w_018_1628, w_018_1629, w_018_1631, w_018_1632, w_018_1633, w_018_1634, w_018_1635, w_018_1636, w_018_1637, w_018_1638, w_018_1639, w_018_1640, w_018_1641, w_018_1642, w_018_1643, w_018_1644, w_018_1647, w_018_1649, w_018_1650, w_018_1651, w_018_1652, w_018_1653, w_018_1655, w_018_1656, w_018_1657, w_018_1658, w_018_1659, w_018_1660, w_018_1661, w_018_1662, w_018_1663, w_018_1664, w_018_1665, w_018_1666, w_018_1667, w_018_1668, w_018_1669, w_018_1670, w_018_1671, w_018_1672, w_018_1673, w_018_1674, w_018_1675, w_018_1676, w_018_1677, w_018_1678, w_018_1679, w_018_1680, w_018_1681, w_018_1682, w_018_1683, w_018_1684, w_018_1685, w_018_1686, w_018_1687, w_018_1688, w_018_1690, w_018_1691, w_018_1693, w_018_1694, w_018_1695, w_018_1696, w_018_1697, w_018_1698, w_018_1700, w_018_1701, w_018_1702, w_018_1703, w_018_1704, w_018_1705, w_018_1706, w_018_1707, w_018_1708, w_018_1709, w_018_1710, w_018_1711, w_018_1712, w_018_1713, w_018_1714, w_018_1715, w_018_1716, w_018_1717, w_018_1718, w_018_1719, w_018_1720, w_018_1721, w_018_1722, w_018_1723, w_018_1724, w_018_1725, w_018_1726, w_018_1727, w_018_1728, w_018_1729, w_018_1730, w_018_1731, w_018_1732, w_018_1733, w_018_1734, w_018_1735, w_018_1736, w_018_1737, w_018_1738, w_018_1739, w_018_1740, w_018_1741, w_018_1742, w_018_1743, w_018_1744, w_018_1745, w_018_1746, w_018_1747, w_018_1748, w_018_1749, w_018_1750, w_018_1751, w_018_1752, w_018_1754, w_018_1755, w_018_1756, w_018_1757, w_018_1758, w_018_1759, w_018_1760, w_018_1761, w_018_1762, w_018_1763, w_018_1764, w_018_1765, w_018_1766, w_018_1767, w_018_1768, w_018_1769, w_018_1770, w_018_1771, w_018_1773, w_018_1774, w_018_1776, w_018_1777, w_018_1778, w_018_1779, w_018_1780, w_018_1781, w_018_1782, w_018_1783, w_018_1784, w_018_1785, w_018_1786, w_018_1787, w_018_1788, w_018_1789, w_018_1790, w_018_1791, w_018_1792, w_018_1793, w_018_1794, w_018_1795, w_018_1796, w_018_1797, w_018_1798, w_018_1799, w_018_1800, w_018_1801, w_018_1802, w_018_1803, w_018_1804, w_018_1805, w_018_1806, w_018_1807, w_018_1808, w_018_1809, w_018_1810, w_018_1811, w_018_1812, w_018_1813, w_018_1814, w_018_1815, w_018_1816, w_018_1817, w_018_1818, w_018_1819, w_018_1820, w_018_1821, w_018_1822, w_018_1823, w_018_1825, w_018_1826, w_018_1827, w_018_1828, w_018_1829, w_018_1830, w_018_1831, w_018_1832, w_018_1833, w_018_1834, w_018_1835, w_018_1836, w_018_1837, w_018_1838, w_018_1839, w_018_1840, w_018_1841, w_018_1842, w_018_1843, w_018_1844, w_018_1845, w_018_1847, w_018_1848, w_018_1849, w_018_1850, w_018_1851, w_018_1853, w_018_1854, w_018_1855, w_018_1856, w_018_1857, w_018_1858, w_018_1859, w_018_1860, w_018_1861, w_018_1862, w_018_1863, w_018_1864, w_018_1865, w_018_1866, w_018_1867, w_018_1868, w_018_1869, w_018_1870, w_018_1871, w_018_1873, w_018_1874, w_018_1875, w_018_1876, w_018_1877, w_018_1878, w_018_1879, w_018_1880, w_018_1881, w_018_1882, w_018_1883, w_018_1884, w_018_1885, w_018_1886, w_018_1887, w_018_1888, w_018_1889, w_018_1890, w_018_1891, w_018_1892, w_018_1893, w_018_1894, w_018_1895, w_018_1896, w_018_1897, w_018_1898, w_018_1899, w_018_1900, w_018_1901, w_018_1902, w_018_1903, w_018_1904, w_018_1905, w_018_1906, w_018_1907, w_018_1908, w_018_1909, w_018_1910, w_018_1911, w_018_1912, w_018_1913, w_018_1914, w_018_1915, w_018_1916, w_018_1917, w_018_1918, w_018_1919, w_018_1920, w_018_1921, w_018_1922, w_018_1923, w_018_1924, w_018_1925, w_018_1927, w_018_1928, w_018_1929, w_018_1930, w_018_1932, w_018_1933, w_018_1934, w_018_1935, w_018_1936, w_018_1937, w_018_1938, w_018_1939, w_018_1940, w_018_1941, w_018_1942, w_018_1943, w_018_1945, w_018_1946, w_018_1947, w_018_1948, w_018_1949, w_018_1950, w_018_1951, w_018_1952, w_018_1953, w_018_1954, w_018_1955, w_018_1956, w_018_1957, w_018_1958, w_018_1959, w_018_1960, w_018_1961, w_018_1962, w_018_1963, w_018_1964, w_018_1965, w_018_1966, w_018_1967, w_018_1968, w_018_1969, w_018_1970, w_018_1971, w_018_1972, w_018_1973, w_018_1974, w_018_1975, w_018_1976, w_018_1977, w_018_1978, w_018_1979, w_018_1980, w_018_1981, w_018_1982, w_018_1984, w_018_1985, w_018_1986, w_018_1987, w_018_1988, w_018_1989, w_018_1990, w_018_1991, w_018_1992, w_018_1993, w_018_1994, w_018_1995, w_018_1996, w_018_1997, w_018_1998, w_018_1999, w_018_2000, w_018_2001, w_018_2002, w_018_2003, w_018_2004, w_018_2005, w_018_2006, w_018_2007, w_018_2008, w_018_2009, w_018_2010, w_018_2011, w_018_2012, w_018_2013, w_018_2014, w_018_2015, w_018_2016, w_018_2017, w_018_2018, w_018_2019, w_018_2020, w_018_2021, w_018_2022, w_018_2023, w_018_2024, w_018_2025, w_018_2026, w_018_2027, w_018_2028, w_018_2029, w_018_2030, w_018_2032, w_018_2033, w_018_2034, w_018_2035, w_018_2036, w_018_2037, w_018_2038, w_018_2039, w_018_2040, w_018_2041, w_018_2042, w_018_2043, w_018_2044, w_018_2045, w_018_2046, w_018_2047, w_018_2048, w_018_2049, w_018_2050, w_018_2051, w_018_2052, w_018_2053, w_018_2054, w_018_2055, w_018_2056, w_018_2057, w_018_2058, w_018_2059, w_018_2060, w_018_2061, w_018_2062, w_018_2064, w_018_2065, w_018_2066, w_018_2067, w_018_2068, w_018_2069, w_018_2070, w_018_2071, w_018_2072, w_018_2073, w_018_2074, w_018_2075, w_018_2076, w_018_2077, w_018_2078, w_018_2079, w_018_2080, w_018_2081, w_018_2082, w_018_2083, w_018_2084, w_018_2085, w_018_2086, w_018_2087, w_018_2088, w_018_2089, w_018_2090, w_018_2091, w_018_2092, w_018_2094, w_018_2095, w_018_2097, w_018_2098, w_018_2099, w_018_2100, w_018_2101, w_018_2102, w_018_2103, w_018_2104, w_018_2105, w_018_2106, w_018_2107, w_018_2108, w_018_2109, w_018_2111, w_018_2112, w_018_2113, w_018_2114, w_018_2115, w_018_2116, w_018_2117, w_018_2118, w_018_2119, w_018_2120, w_018_2121, w_018_2122, w_018_2123, w_018_2124, w_018_2125, w_018_2126, w_018_2127, w_018_2128, w_018_2129, w_018_2130, w_018_2131, w_018_2132, w_018_2133, w_018_2134, w_018_2135, w_018_2136, w_018_2137, w_018_2138, w_018_2139, w_018_2140, w_018_2141, w_018_2142, w_018_2143, w_018_2144, w_018_2145, w_018_2146, w_018_2147, w_018_2148, w_018_2149, w_018_2150, w_018_2151, w_018_2152, w_018_2153, w_018_2154, w_018_2155, w_018_2156, w_018_2157, w_018_2158, w_018_2159, w_018_2160, w_018_2161, w_018_2162, w_018_2163, w_018_2164, w_018_2165, w_018_2166, w_018_2167, w_018_2168, w_018_2169, w_018_2170, w_018_2172, w_018_2173, w_018_2174, w_018_2175, w_018_2176, w_018_2178, w_018_2179, w_018_2180, w_018_2181, w_018_2182, w_018_2183, w_018_2184, w_018_2185, w_018_2186, w_018_2187, w_018_2188, w_018_2189, w_018_2190, w_018_2191, w_018_2192, w_018_2193, w_018_2194, w_018_2195, w_018_2196, w_018_2197, w_018_2198, w_018_2199, w_018_2200, w_018_2201, w_018_2202, w_018_2203, w_018_2204, w_018_2205, w_018_2206, w_018_2207, w_018_2208, w_018_2209, w_018_2210, w_018_2211, w_018_2212, w_018_2213, w_018_2214, w_018_2215, w_018_2216, w_018_2217, w_018_2218, w_018_2219, w_018_2220, w_018_2221, w_018_2222, w_018_2223, w_018_2224, w_018_2225, w_018_2226, w_018_2227, w_018_2228, w_018_2229, w_018_2230, w_018_2231, w_018_2232, w_018_2233, w_018_2234, w_018_2235, w_018_2236, w_018_2237, w_018_2238, w_018_2239, w_018_2240, w_018_2241, w_018_2242, w_018_2243, w_018_2244, w_018_2246, w_018_2247, w_018_2249, w_018_2250, w_018_2251, w_018_2253, w_018_2254, w_018_2255, w_018_2256, w_018_2257, w_018_2258, w_018_2259, w_018_2260, w_018_2261, w_018_2262, w_018_2263, w_018_2265, w_018_2266, w_018_2267, w_018_2268, w_018_2269, w_018_2270, w_018_2271, w_018_2272, w_018_2273, w_018_2274, w_018_2275, w_018_2276, w_018_2277, w_018_2278, w_018_2279, w_018_2280, w_018_2281, w_018_2282, w_018_2283, w_018_2285, w_018_2287, w_018_2288, w_018_2289, w_018_2290, w_018_2291, w_018_2292, w_018_2293, w_018_2294, w_018_2295, w_018_2296, w_018_2297, w_018_2299, w_018_2300, w_018_2301, w_018_2302, w_018_2303, w_018_2304, w_018_2305, w_018_2306, w_018_2307, w_018_2308, w_018_2309, w_018_2310, w_018_2311, w_018_2312, w_018_2313, w_018_2314, w_018_2315, w_018_2316, w_018_2317, w_018_2318, w_018_2319, w_018_2321, w_018_2322, w_018_2323, w_018_2324, w_018_2325, w_018_2326, w_018_2327, w_018_2328, w_018_2329, w_018_2330, w_018_2331, w_018_2332, w_018_2333, w_018_2334, w_018_2335, w_018_2336, w_018_2337, w_018_2338, w_018_2340, w_018_2341, w_018_2342, w_018_2343, w_018_2344, w_018_2345, w_018_2346, w_018_2347, w_018_2348, w_018_2349, w_018_2350, w_018_2351, w_018_2352, w_018_2353, w_018_2354, w_018_2355, w_018_2356, w_018_2357, w_018_2358, w_018_2359, w_018_2361, w_018_2362, w_018_2363, w_018_2364, w_018_2366, w_018_2367, w_018_2368, w_018_2369, w_018_2370, w_018_2371, w_018_2373, w_018_2374, w_018_2375, w_018_2376, w_018_2377, w_018_2378, w_018_2379, w_018_2380, w_018_2381, w_018_2382, w_018_2383, w_018_2384, w_018_2385, w_018_2386, w_018_2387, w_018_2388, w_018_2389, w_018_2390, w_018_2391, w_018_2392, w_018_2393, w_018_2394, w_018_2395, w_018_2396, w_018_2397, w_018_2398, w_018_2399, w_018_2400, w_018_2401, w_018_2402, w_018_2403, w_018_2404, w_018_2405, w_018_2406, w_018_2407, w_018_2408, w_018_2409, w_018_2410, w_018_2411, w_018_2412, w_018_2413, w_018_2414, w_018_2416, w_018_2417, w_018_2418, w_018_2419, w_018_2420, w_018_2421, w_018_2422, w_018_2423, w_018_2424, w_018_2425, w_018_2426, w_018_2427, w_018_2428, w_018_2429, w_018_2430, w_018_2431, w_018_2432, w_018_2433, w_018_2434, w_018_2435, w_018_2436, w_018_2437, w_018_2438, w_018_2439, w_018_2440, w_018_2441, w_018_2442, w_018_2443, w_018_2444, w_018_2446, w_018_2447, w_018_2448, w_018_2449, w_018_2450, w_018_2451, w_018_2452, w_018_2453, w_018_2454, w_018_2455, w_018_2456, w_018_2457, w_018_2458, w_018_2459, w_018_2460, w_018_2461, w_018_2462, w_018_2463, w_018_2464, w_018_2465, w_018_2466, w_018_2467, w_018_2468, w_018_2469, w_018_2470, w_018_2471, w_018_2472, w_018_2473, w_018_2474, w_018_2475, w_018_2476, w_018_2477, w_018_2478, w_018_2479, w_018_2480, w_018_2481, w_018_2482, w_018_2484, w_018_2485, w_018_2486, w_018_2487, w_018_2488, w_018_2489, w_018_2490, w_018_2491, w_018_2492, w_018_2493, w_018_2494, w_018_2495, w_018_2497, w_018_2498, w_018_2499, w_018_2500, w_018_2501, w_018_2502, w_018_2503, w_018_2504, w_018_2505, w_018_2506, w_018_2507, w_018_2508, w_018_2509, w_018_2510, w_018_2511, w_018_2512, w_018_2513, w_018_2514, w_018_2515, w_018_2516, w_018_2517, w_018_2518, w_018_2519, w_018_2520, w_018_2521, w_018_2522, w_018_2523, w_018_2524, w_018_2525, w_018_2526, w_018_2527, w_018_2528, w_018_2529, w_018_2530, w_018_2531, w_018_2532, w_018_2533, w_018_2534, w_018_2535, w_018_2536, w_018_2537, w_018_2538, w_018_2539, w_018_2540, w_018_2541, w_018_2542, w_018_2543, w_018_2544, w_018_2545, w_018_2546, w_018_2547, w_018_2548, w_018_2549, w_018_2550, w_018_2551, w_018_2552, w_018_2554, w_018_2555, w_018_2556, w_018_2557, w_018_2558, w_018_2559, w_018_2560, w_018_2561, w_018_2562, w_018_2563, w_018_2564, w_018_2565, w_018_2566, w_018_2567, w_018_2568, w_018_2569, w_018_2570, w_018_2571, w_018_2572, w_018_2573, w_018_2574, w_018_2575, w_018_2576, w_018_2577, w_018_2578, w_018_2580, w_018_2581, w_018_2582, w_018_2583, w_018_2584, w_018_2585, w_018_2586, w_018_2587, w_018_2588, w_018_2589, w_018_2590, w_018_2591, w_018_2592, w_018_2593, w_018_2594, w_018_2595, w_018_2596, w_018_2597, w_018_2598, w_018_2599, w_018_2600, w_018_2601, w_018_2602, w_018_2604, w_018_2605, w_018_2606, w_018_2607, w_018_2608, w_018_2609, w_018_2610, w_018_2611, w_018_2612, w_018_2613, w_018_2614, w_018_2615, w_018_2616, w_018_2617, w_018_2618, w_018_2619, w_018_2620, w_018_2621, w_018_2622, w_018_2623, w_018_2624, w_018_2625, w_018_2626, w_018_2627, w_018_2628, w_018_2629, w_018_2630, w_018_2631, w_018_2632, w_018_2633, w_018_2634, w_018_2635, w_018_2636, w_018_2637, w_018_2639, w_018_2640, w_018_2641, w_018_2642, w_018_2643, w_018_2645, w_018_2647, w_018_2648, w_018_2649, w_018_2650, w_018_2651, w_018_2652, w_018_2653, w_018_2654, w_018_2655, w_018_2656, w_018_2657, w_018_2658, w_018_2659, w_018_2660, w_018_2661, w_018_2662, w_018_2663, w_018_2664, w_018_2665, w_018_2666, w_018_2667, w_018_2668, w_018_2669, w_018_2670, w_018_2671, w_018_2672, w_018_2673, w_018_2675, w_018_2676, w_018_2677, w_018_2678, w_018_2679, w_018_2680, w_018_2681, w_018_2682, w_018_2683, w_018_2684, w_018_2685, w_018_2686, w_018_2687, w_018_2688, w_018_2690, w_018_2691, w_018_2692, w_018_2693, w_018_2694, w_018_2695, w_018_2696, w_018_2697, w_018_2698, w_018_2699, w_018_2700, w_018_2701, w_018_2702, w_018_2705, w_018_2706, w_018_2707, w_018_2708, w_018_2709, w_018_2711, w_018_2712, w_018_2713, w_018_2715, w_018_2716, w_018_2717, w_018_2718, w_018_2719, w_018_2720, w_018_2721, w_018_2722, w_018_2723, w_018_2724, w_018_2725, w_018_2726, w_018_2727, w_018_2728, w_018_2729, w_018_2730, w_018_2731, w_018_2732, w_018_2733, w_018_2734, w_018_2735, w_018_2736, w_018_2737, w_018_2738, w_018_2739, w_018_2740, w_018_2741, w_018_2742, w_018_2743, w_018_2744, w_018_2745, w_018_2746, w_018_2747, w_018_2748, w_018_2749, w_018_2750, w_018_2751, w_018_2752, w_018_2753, w_018_2754, w_018_2755, w_018_2756, w_018_2757, w_018_2758, w_018_2759, w_018_2760, w_018_2761, w_018_2762, w_018_2764, w_018_2765, w_018_2766, w_018_2768, w_018_2769, w_018_2770, w_018_2771, w_018_2772, w_018_2773, w_018_2774, w_018_2776, w_018_2777, w_018_2778, w_018_2779, w_018_2780, w_018_2781, w_018_2782, w_018_2783, w_018_2784, w_018_2785, w_018_2786, w_018_2787, w_018_2788, w_018_2789, w_018_2790, w_018_2791, w_018_2792, w_018_2793, w_018_2794, w_018_2795, w_018_2796, w_018_2797, w_018_2798, w_018_2799, w_018_2800, w_018_2801, w_018_2802, w_018_2803, w_018_2804, w_018_2805, w_018_2806, w_018_2807, w_018_2808, w_018_2809, w_018_2810, w_018_2811, w_018_2812, w_018_2813, w_018_2814, w_018_2815, w_018_2816, w_018_2817, w_018_2818, w_018_2819, w_018_2820, w_018_2821, w_018_2822, w_018_2823, w_018_2824, w_018_2825, w_018_2826, w_018_2827, w_018_2828, w_018_2829, w_018_2830, w_018_2831, w_018_2832, w_018_2833, w_018_2834, w_018_2835, w_018_2836, w_018_2837, w_018_2838, w_018_2839, w_018_2840, w_018_2841, w_018_2842, w_018_2843, w_018_2844, w_018_2845, w_018_2846, w_018_2847, w_018_2848, w_018_2849, w_018_2850, w_018_2851, w_018_2852, w_018_2853, w_018_2854, w_018_2855, w_018_2856, w_018_2857, w_018_2858, w_018_2859, w_018_2860, w_018_2861, w_018_2862, w_018_2863, w_018_2864, w_018_2865, w_018_2866, w_018_2867, w_018_2869, w_018_2870, w_018_2871, w_018_2872, w_018_2873, w_018_2874, w_018_2875, w_018_2876, w_018_2877, w_018_2878, w_018_2879, w_018_2880, w_018_2881, w_018_2882, w_018_2883, w_018_2884, w_018_2885, w_018_2886, w_018_2887, w_018_2889, w_018_2890, w_018_2891, w_018_2893, w_018_2894, w_018_2895, w_018_2897, w_018_2898, w_018_2899, w_018_2900, w_018_2901, w_018_2902, w_018_2903, w_018_2904, w_018_2905, w_018_2906, w_018_2907, w_018_2908, w_018_2909, w_018_2910, w_018_2911, w_018_2912, w_018_2913, w_018_2914, w_018_2915, w_018_2916, w_018_2917, w_018_2918, w_018_2919, w_018_2920, w_018_2921, w_018_2922, w_018_2923, w_018_2924, w_018_2925, w_018_2926, w_018_2927, w_018_2928, w_018_2929, w_018_2930, w_018_2931, w_018_2932, w_018_2933, w_018_2934, w_018_2935, w_018_2936, w_018_2937, w_018_2938, w_018_2939, w_018_2941, w_018_2942, w_018_2944, w_018_2945, w_018_2947, w_018_2948, w_018_2949, w_018_2950, w_018_2951, w_018_2952, w_018_2953, w_018_2954, w_018_2955, w_018_2956, w_018_2957, w_018_2958, w_018_2959, w_018_2960, w_018_2961, w_018_2962, w_018_2963, w_018_2964, w_018_2965, w_018_2966, w_018_2967, w_018_2968, w_018_2969, w_018_2970, w_018_2971, w_018_2972, w_018_2973, w_018_2974, w_018_2975, w_018_2976, w_018_2977, w_018_2978, w_018_2979, w_018_2980, w_018_2981, w_018_2982, w_018_2983, w_018_2984, w_018_2985, w_018_2986, w_018_2987, w_018_2988, w_018_2989, w_018_2990, w_018_2991, w_018_2992, w_018_2993, w_018_2994, w_018_2996, w_018_2997, w_018_2998, w_018_2999, w_018_3000, w_018_3001, w_018_3003, w_018_3004, w_018_3005, w_018_3006, w_018_3007, w_018_3008, w_018_3009, w_018_3010, w_018_3011, w_018_3012, w_018_3013, w_018_3014, w_018_3015, w_018_3016, w_018_3017, w_018_3018, w_018_3019, w_018_3020, w_018_3021, w_018_3022, w_018_3023, w_018_3024, w_018_3025, w_018_3026, w_018_3027, w_018_3028, w_018_3029, w_018_3030, w_018_3031, w_018_3032, w_018_3033, w_018_3034, w_018_3035, w_018_3036, w_018_3037, w_018_3038, w_018_3039, w_018_3040, w_018_3041, w_018_3042, w_018_3043, w_018_3044, w_018_3045, w_018_3047, w_018_3048, w_018_3049, w_018_3050, w_018_3051, w_018_3052, w_018_3053, w_018_3054, w_018_3055, w_018_3056, w_018_3057, w_018_3058, w_018_3059, w_018_3060, w_018_3061, w_018_3062, w_018_3063, w_018_3065, w_018_3066, w_018_3067, w_018_3068, w_018_3069, w_018_3070, w_018_3071, w_018_3072, w_018_3073, w_018_3074, w_018_3075, w_018_3076, w_018_3077, w_018_3078, w_018_3079, w_018_3080, w_018_3081, w_018_3082, w_018_3083, w_018_3084, w_018_3085, w_018_3086, w_018_3087, w_018_3088, w_018_3089, w_018_3090, w_018_3091, w_018_3092, w_018_3093, w_018_3094, w_018_3095, w_018_3097, w_018_3098, w_018_3099, w_018_3100, w_018_3101, w_018_3102, w_018_3103, w_018_3105, w_018_3106, w_018_3107, w_018_3108, w_018_3109;
  wire w_019_000, w_019_001, w_019_002, w_019_003, w_019_004, w_019_005, w_019_006, w_019_007, w_019_008, w_019_009, w_019_010, w_019_011, w_019_012, w_019_013, w_019_014, w_019_015, w_019_016, w_019_017, w_019_018, w_019_019, w_019_020, w_019_021, w_019_022, w_019_023, w_019_024, w_019_025, w_019_026, w_019_027, w_019_028, w_019_029, w_019_030, w_019_031, w_019_032, w_019_033, w_019_034, w_019_035, w_019_036, w_019_037, w_019_038, w_019_039, w_019_040, w_019_041, w_019_042, w_019_043, w_019_044, w_019_045, w_019_046, w_019_047, w_019_048, w_019_049, w_019_050, w_019_051, w_019_052, w_019_053, w_019_054, w_019_055, w_019_056, w_019_057, w_019_058, w_019_059, w_019_060, w_019_061, w_019_062, w_019_063, w_019_064, w_019_065, w_019_066, w_019_067, w_019_068, w_019_069, w_019_070, w_019_071, w_019_072, w_019_073, w_019_074, w_019_075, w_019_076, w_019_077, w_019_078, w_019_079, w_019_080, w_019_081, w_019_082, w_019_083, w_019_084, w_019_085, w_019_086, w_019_087, w_019_088, w_019_089, w_019_090, w_019_091, w_019_092, w_019_093, w_019_094, w_019_095, w_019_096, w_019_097, w_019_098, w_019_099, w_019_100, w_019_101, w_019_102, w_019_103, w_019_104, w_019_105, w_019_106, w_019_107, w_019_108, w_019_109, w_019_110, w_019_111, w_019_112, w_019_113, w_019_114, w_019_115, w_019_116, w_019_117, w_019_118, w_019_119, w_019_120, w_019_121, w_019_122, w_019_123, w_019_124, w_019_125, w_019_126, w_019_127, w_019_128, w_019_129, w_019_130, w_019_131, w_019_132, w_019_133, w_019_134, w_019_135, w_019_136, w_019_137, w_019_138, w_019_139, w_019_140, w_019_141, w_019_142, w_019_143, w_019_144, w_019_145, w_019_146, w_019_147, w_019_148, w_019_149, w_019_150, w_019_151, w_019_152, w_019_153, w_019_154, w_019_155, w_019_156, w_019_157, w_019_158, w_019_159, w_019_160, w_019_161, w_019_162, w_019_163, w_019_164, w_019_165, w_019_166, w_019_167, w_019_168, w_019_169, w_019_170, w_019_171, w_019_172, w_019_173, w_019_174, w_019_175, w_019_176, w_019_177, w_019_178, w_019_179, w_019_180, w_019_181, w_019_182, w_019_183, w_019_184, w_019_185, w_019_186, w_019_187, w_019_188, w_019_189, w_019_190, w_019_191, w_019_192, w_019_193, w_019_194, w_019_195, w_019_196, w_019_197, w_019_198, w_019_199, w_019_200, w_019_201, w_019_202, w_019_203, w_019_204, w_019_205, w_019_206, w_019_207, w_019_208, w_019_209, w_019_210, w_019_211, w_019_212, w_019_213, w_019_214, w_019_215, w_019_216, w_019_217, w_019_218, w_019_219, w_019_220, w_019_221, w_019_222, w_019_223, w_019_224, w_019_225, w_019_226, w_019_227, w_019_228, w_019_229, w_019_230, w_019_231, w_019_232, w_019_233, w_019_234, w_019_235, w_019_236, w_019_237, w_019_238, w_019_239, w_019_240, w_019_241, w_019_242, w_019_243, w_019_244, w_019_245, w_019_246, w_019_247, w_019_248, w_019_249, w_019_250, w_019_251, w_019_252, w_019_253, w_019_254, w_019_255, w_019_256, w_019_257, w_019_258, w_019_259, w_019_260, w_019_261, w_019_262, w_019_263, w_019_264, w_019_265, w_019_266, w_019_267, w_019_268, w_019_269, w_019_270, w_019_271, w_019_272, w_019_273, w_019_274, w_019_275, w_019_276, w_019_277, w_019_278, w_019_279, w_019_280, w_019_281, w_019_282, w_019_283, w_019_284, w_019_285, w_019_286, w_019_287, w_019_288, w_019_289, w_019_290, w_019_291, w_019_292, w_019_293, w_019_294, w_019_295, w_019_296, w_019_297, w_019_298, w_019_299, w_019_300, w_019_301, w_019_302, w_019_303, w_019_304, w_019_305, w_019_306, w_019_307, w_019_308, w_019_309, w_019_310, w_019_311, w_019_312, w_019_313, w_019_314, w_019_315, w_019_316, w_019_317, w_019_318, w_019_319, w_019_320, w_019_321, w_019_322, w_019_323, w_019_324, w_019_325, w_019_326, w_019_327, w_019_328, w_019_329, w_019_330, w_019_331, w_019_332, w_019_333, w_019_334, w_019_335, w_019_336, w_019_337, w_019_338, w_019_339, w_019_340, w_019_341, w_019_342, w_019_343, w_019_344, w_019_345, w_019_346, w_019_347, w_019_348, w_019_349, w_019_350, w_019_351, w_019_352, w_019_353, w_019_354, w_019_355, w_019_356, w_019_357, w_019_358, w_019_359, w_019_360, w_019_361, w_019_362, w_019_363, w_019_364, w_019_365, w_019_366, w_019_367, w_019_368, w_019_369, w_019_370, w_019_371, w_019_372, w_019_373, w_019_374, w_019_375, w_019_376, w_019_377, w_019_378, w_019_379, w_019_380, w_019_381, w_019_382, w_019_383, w_019_384, w_019_385, w_019_386, w_019_387, w_019_388, w_019_389, w_019_390, w_019_391, w_019_392, w_019_393, w_019_394, w_019_395, w_019_396, w_019_397, w_019_398, w_019_399, w_019_400, w_019_401, w_019_402, w_019_403, w_019_404, w_019_405, w_019_406, w_019_407, w_019_408, w_019_409, w_019_410, w_019_411, w_019_412, w_019_413, w_019_414, w_019_415, w_019_416, w_019_417, w_019_418, w_019_419, w_019_420, w_019_421, w_019_422, w_019_423, w_019_424, w_019_425, w_019_426, w_019_427, w_019_428, w_019_429, w_019_430, w_019_431, w_019_432, w_019_433, w_019_434, w_019_435, w_019_436, w_019_437, w_019_438, w_019_439, w_019_440, w_019_441, w_019_442, w_019_443, w_019_444, w_019_445, w_019_446, w_019_447, w_019_448, w_019_449, w_019_450, w_019_451, w_019_452, w_019_453, w_019_454, w_019_455, w_019_456, w_019_457, w_019_458, w_019_459, w_019_460, w_019_461, w_019_462, w_019_463, w_019_464, w_019_465, w_019_466, w_019_467, w_019_468, w_019_469, w_019_470, w_019_471, w_019_472, w_019_473, w_019_474, w_019_475, w_019_476, w_019_477, w_019_478, w_019_479, w_019_480, w_019_481, w_019_482, w_019_483, w_019_484, w_019_485, w_019_486, w_019_487, w_019_488, w_019_489, w_019_490, w_019_491, w_019_492, w_019_493, w_019_494, w_019_495, w_019_496, w_019_497, w_019_498, w_019_499, w_019_500, w_019_501, w_019_502, w_019_503, w_019_504, w_019_505, w_019_506, w_019_507, w_019_508, w_019_509, w_019_510, w_019_511, w_019_512, w_019_513, w_019_514, w_019_515, w_019_516, w_019_517, w_019_518, w_019_519, w_019_520, w_019_521, w_019_522, w_019_523, w_019_524, w_019_525, w_019_526, w_019_527, w_019_528, w_019_529, w_019_530, w_019_531, w_019_532, w_019_533, w_019_534, w_019_535, w_019_536, w_019_537, w_019_538, w_019_539, w_019_540, w_019_541, w_019_542, w_019_543, w_019_544, w_019_545, w_019_546, w_019_547, w_019_548, w_019_549, w_019_550, w_019_551, w_019_552, w_019_553, w_019_554, w_019_555, w_019_556, w_019_557, w_019_558, w_019_559, w_019_560, w_019_561, w_019_562, w_019_563, w_019_564, w_019_565, w_019_566, w_019_567, w_019_568, w_019_569, w_019_570, w_019_571, w_019_572, w_019_573, w_019_574, w_019_575, w_019_576, w_019_577, w_019_578, w_019_579, w_019_580, w_019_581, w_019_582, w_019_583, w_019_584, w_019_585, w_019_586, w_019_587, w_019_588, w_019_589, w_019_590, w_019_591, w_019_592, w_019_593, w_019_594, w_019_595, w_019_596, w_019_597, w_019_598, w_019_599, w_019_600, w_019_601, w_019_602, w_019_603, w_019_604, w_019_605, w_019_606, w_019_607, w_019_608, w_019_609, w_019_610, w_019_611, w_019_612, w_019_613, w_019_614, w_019_615, w_019_616, w_019_617, w_019_618, w_019_619, w_019_620, w_019_621, w_019_622, w_019_623, w_019_624, w_019_625, w_019_626, w_019_627, w_019_628, w_019_629, w_019_630, w_019_631, w_019_632, w_019_633, w_019_634, w_019_635, w_019_636, w_019_637, w_019_638, w_019_639, w_019_640, w_019_641, w_019_642, w_019_643, w_019_644, w_019_645, w_019_646, w_019_647, w_019_648, w_019_649, w_019_650, w_019_651, w_019_652, w_019_653, w_019_654, w_019_655, w_019_656, w_019_657, w_019_658, w_019_659, w_019_660, w_019_661, w_019_662, w_019_663, w_019_664, w_019_665, w_019_666, w_019_667, w_019_668, w_019_669, w_019_670, w_019_671, w_019_672, w_019_673, w_019_674, w_019_675, w_019_676, w_019_677, w_019_678, w_019_679, w_019_680, w_019_681, w_019_682, w_019_683, w_019_684, w_019_685, w_019_686, w_019_687, w_019_688, w_019_689, w_019_690, w_019_691, w_019_692, w_019_693, w_019_694, w_019_695, w_019_696, w_019_697, w_019_698, w_019_699, w_019_700, w_019_701, w_019_702, w_019_703, w_019_704, w_019_705, w_019_706, w_019_707, w_019_708, w_019_709, w_019_710, w_019_711, w_019_712, w_019_713, w_019_714, w_019_715, w_019_716, w_019_717, w_019_718, w_019_719, w_019_720, w_019_721, w_019_722, w_019_723, w_019_724, w_019_725, w_019_726, w_019_727, w_019_728, w_019_729, w_019_730, w_019_731, w_019_732, w_019_733, w_019_734, w_019_735, w_019_736, w_019_737, w_019_738, w_019_739, w_019_740, w_019_741, w_019_742, w_019_743, w_019_744, w_019_745, w_019_746, w_019_747, w_019_748, w_019_749, w_019_750, w_019_751, w_019_752, w_019_753, w_019_754, w_019_755, w_019_756, w_019_757, w_019_758, w_019_759, w_019_760, w_019_761, w_019_762, w_019_763, w_019_764, w_019_765, w_019_766, w_019_767, w_019_768, w_019_769, w_019_770, w_019_771, w_019_772, w_019_773, w_019_774, w_019_775, w_019_776, w_019_777, w_019_778, w_019_779, w_019_780, w_019_781, w_019_782, w_019_783, w_019_784, w_019_785, w_019_786, w_019_787, w_019_788, w_019_789, w_019_790, w_019_791, w_019_792, w_019_793, w_019_794, w_019_795, w_019_796, w_019_797, w_019_798, w_019_799, w_019_800, w_019_801, w_019_802, w_019_803, w_019_804, w_019_805, w_019_806, w_019_807, w_019_808, w_019_809, w_019_810, w_019_811, w_019_812, w_019_813, w_019_814, w_019_815, w_019_816, w_019_817, w_019_818, w_019_819, w_019_820, w_019_821, w_019_822, w_019_823, w_019_824, w_019_825, w_019_826, w_019_827, w_019_828, w_019_829, w_019_830, w_019_831, w_019_832, w_019_833, w_019_834, w_019_835, w_019_836, w_019_837, w_019_838, w_019_839, w_019_840, w_019_841, w_019_842, w_019_843, w_019_844, w_019_845, w_019_846, w_019_847, w_019_848, w_019_849, w_019_850, w_019_851, w_019_852, w_019_853, w_019_854, w_019_855, w_019_856, w_019_857, w_019_858, w_019_859, w_019_860, w_019_861, w_019_862, w_019_863, w_019_864, w_019_865, w_019_866, w_019_867, w_019_868, w_019_869, w_019_870, w_019_871, w_019_872, w_019_873, w_019_874, w_019_875, w_019_876, w_019_877, w_019_878, w_019_879, w_019_880, w_019_881, w_019_882, w_019_883, w_019_884, w_019_885, w_019_886, w_019_887, w_019_888, w_019_889, w_019_890, w_019_891, w_019_892, w_019_893, w_019_894, w_019_895, w_019_896, w_019_897, w_019_898, w_019_899, w_019_900, w_019_901, w_019_902, w_019_903, w_019_904, w_019_905, w_019_906, w_019_907, w_019_908, w_019_909, w_019_910, w_019_911, w_019_912, w_019_913, w_019_914, w_019_915, w_019_916, w_019_917, w_019_918, w_019_919, w_019_920, w_019_921, w_019_922, w_019_923, w_019_924;
  wire w_020_000, w_020_001, w_020_002, w_020_003, w_020_005, w_020_006, w_020_007, w_020_008, w_020_009, w_020_010, w_020_011, w_020_012, w_020_013, w_020_014, w_020_016, w_020_017, w_020_018, w_020_019, w_020_021, w_020_022, w_020_023, w_020_024, w_020_025, w_020_026, w_020_028, w_020_029, w_020_030, w_020_031, w_020_032, w_020_033, w_020_034, w_020_035, w_020_036, w_020_037, w_020_038, w_020_039, w_020_040, w_020_041, w_020_042, w_020_044, w_020_045, w_020_047, w_020_048, w_020_049, w_020_050, w_020_051, w_020_052, w_020_053, w_020_054, w_020_055, w_020_056, w_020_057, w_020_058, w_020_059, w_020_060, w_020_061, w_020_062, w_020_064, w_020_065, w_020_066, w_020_067, w_020_068, w_020_070, w_020_071, w_020_072, w_020_073, w_020_074, w_020_075, w_020_076, w_020_077, w_020_078, w_020_079, w_020_081, w_020_082, w_020_084, w_020_085, w_020_086, w_020_087, w_020_088, w_020_089, w_020_090, w_020_091, w_020_092, w_020_093, w_020_094, w_020_095, w_020_096, w_020_097, w_020_098, w_020_099, w_020_100, w_020_101, w_020_102, w_020_103, w_020_104, w_020_105, w_020_107, w_020_108, w_020_109, w_020_110, w_020_111, w_020_112, w_020_113, w_020_114, w_020_115, w_020_117, w_020_118, w_020_119, w_020_120, w_020_121, w_020_122, w_020_123, w_020_124, w_020_127, w_020_128, w_020_129, w_020_130, w_020_131, w_020_133, w_020_134, w_020_135, w_020_136, w_020_137, w_020_138, w_020_140, w_020_141, w_020_142, w_020_143, w_020_144, w_020_145, w_020_146, w_020_147, w_020_148, w_020_149, w_020_150, w_020_151, w_020_152, w_020_153, w_020_155, w_020_156, w_020_157, w_020_158, w_020_159, w_020_160, w_020_161, w_020_162, w_020_163, w_020_164, w_020_166, w_020_167, w_020_168, w_020_169, w_020_170, w_020_171, w_020_172, w_020_173, w_020_175, w_020_176, w_020_177, w_020_178, w_020_179, w_020_180, w_020_181, w_020_182, w_020_183, w_020_184, w_020_185, w_020_186, w_020_187, w_020_189, w_020_190, w_020_191, w_020_192, w_020_193, w_020_194, w_020_195, w_020_196, w_020_197, w_020_198, w_020_200, w_020_201, w_020_202, w_020_203, w_020_204, w_020_205, w_020_206, w_020_207, w_020_208, w_020_209, w_020_210, w_020_211, w_020_212, w_020_213, w_020_214, w_020_215, w_020_216, w_020_217, w_020_218, w_020_219, w_020_220, w_020_221, w_020_223, w_020_224, w_020_225, w_020_227, w_020_228, w_020_229, w_020_230, w_020_231, w_020_232, w_020_233, w_020_234, w_020_235, w_020_236, w_020_237, w_020_238, w_020_239, w_020_240, w_020_242, w_020_243, w_020_244, w_020_245, w_020_247, w_020_248, w_020_250, w_020_251, w_020_252, w_020_253, w_020_255, w_020_256, w_020_257, w_020_258, w_020_259, w_020_261, w_020_263, w_020_265, w_020_266, w_020_267, w_020_268, w_020_269, w_020_270, w_020_271, w_020_272, w_020_273, w_020_274, w_020_275, w_020_276, w_020_277, w_020_278, w_020_279, w_020_283, w_020_284, w_020_285, w_020_286, w_020_287, w_020_288, w_020_289, w_020_290, w_020_291, w_020_293, w_020_294, w_020_295, w_020_296, w_020_297, w_020_298, w_020_299, w_020_300, w_020_301, w_020_302, w_020_303, w_020_306, w_020_307, w_020_308, w_020_309, w_020_310, w_020_311, w_020_312, w_020_313, w_020_314, w_020_315, w_020_316, w_020_317, w_020_318, w_020_319, w_020_320, w_020_321, w_020_322, w_020_323, w_020_324, w_020_326, w_020_327, w_020_328, w_020_329, w_020_330, w_020_331, w_020_332, w_020_334, w_020_335, w_020_336, w_020_337, w_020_338, w_020_339, w_020_340, w_020_341, w_020_342, w_020_343, w_020_344, w_020_345, w_020_346, w_020_348, w_020_349, w_020_350, w_020_351, w_020_352, w_020_353, w_020_354, w_020_355, w_020_356, w_020_357, w_020_358, w_020_359, w_020_360, w_020_361, w_020_362, w_020_363, w_020_364, w_020_365, w_020_366, w_020_367, w_020_368, w_020_369, w_020_370, w_020_371, w_020_372, w_020_373, w_020_374, w_020_375, w_020_376, w_020_377, w_020_378, w_020_379, w_020_380, w_020_381, w_020_382, w_020_383, w_020_384, w_020_386, w_020_387, w_020_388, w_020_389, w_020_390, w_020_391, w_020_392, w_020_393, w_020_394, w_020_395, w_020_396, w_020_397, w_020_398, w_020_399, w_020_400, w_020_401, w_020_403, w_020_404, w_020_405, w_020_406, w_020_407, w_020_408, w_020_409, w_020_410, w_020_411, w_020_412, w_020_413, w_020_414, w_020_415, w_020_416, w_020_417, w_020_418, w_020_420, w_020_421, w_020_422, w_020_423, w_020_424, w_020_425, w_020_426, w_020_427, w_020_429, w_020_430, w_020_431, w_020_432, w_020_433, w_020_434, w_020_435, w_020_436, w_020_437, w_020_439, w_020_440, w_020_441, w_020_442, w_020_443, w_020_444, w_020_445, w_020_446, w_020_447, w_020_448, w_020_449, w_020_450, w_020_451, w_020_453, w_020_454, w_020_456, w_020_458, w_020_461, w_020_464, w_020_465, w_020_466, w_020_467, w_020_468, w_020_469, w_020_471, w_020_473, w_020_474, w_020_475, w_020_476, w_020_477, w_020_478, w_020_479, w_020_480, w_020_481, w_020_483, w_020_484, w_020_485, w_020_486, w_020_487, w_020_488, w_020_489, w_020_490, w_020_491, w_020_493, w_020_494, w_020_495, w_020_496, w_020_497, w_020_498, w_020_499, w_020_500, w_020_501, w_020_502, w_020_503, w_020_504, w_020_506, w_020_507, w_020_508, w_020_509, w_020_510, w_020_511, w_020_512, w_020_513, w_020_514, w_020_515, w_020_517, w_020_519, w_020_520, w_020_521, w_020_522, w_020_524, w_020_525, w_020_526, w_020_527, w_020_528, w_020_529, w_020_530, w_020_533, w_020_534, w_020_535, w_020_536, w_020_537, w_020_538, w_020_539, w_020_540, w_020_541, w_020_542, w_020_543, w_020_544, w_020_545, w_020_546, w_020_547, w_020_548, w_020_549, w_020_551, w_020_552, w_020_553, w_020_554, w_020_555, w_020_556, w_020_557, w_020_559, w_020_560, w_020_561, w_020_562, w_020_563, w_020_564, w_020_565, w_020_566, w_020_567, w_020_569, w_020_570, w_020_572, w_020_573, w_020_574, w_020_575, w_020_576, w_020_577, w_020_578, w_020_579, w_020_580, w_020_581, w_020_582, w_020_583, w_020_584, w_020_585, w_020_586, w_020_587, w_020_588, w_020_590, w_020_591, w_020_592, w_020_593, w_020_595, w_020_596, w_020_597, w_020_598, w_020_599, w_020_600, w_020_601, w_020_602, w_020_603, w_020_605, w_020_606, w_020_607, w_020_609, w_020_610, w_020_611, w_020_612, w_020_614, w_020_615, w_020_616, w_020_617, w_020_618, w_020_619, w_020_620, w_020_621, w_020_622, w_020_624, w_020_626, w_020_627, w_020_628, w_020_629, w_020_630, w_020_632, w_020_633, w_020_634, w_020_635, w_020_636, w_020_637, w_020_638, w_020_639, w_020_641, w_020_642, w_020_643, w_020_644, w_020_645, w_020_646, w_020_647, w_020_650, w_020_651, w_020_652, w_020_653, w_020_654, w_020_655, w_020_656, w_020_657, w_020_658, w_020_660, w_020_662, w_020_666, w_020_667, w_020_670, w_020_671, w_020_672, w_020_673, w_020_674, w_020_675, w_020_676, w_020_677, w_020_678, w_020_679, w_020_680, w_020_681, w_020_682, w_020_684, w_020_689, w_020_690, w_020_691, w_020_692, w_020_693, w_020_695, w_020_697, w_020_698, w_020_699, w_020_700, w_020_701, w_020_702, w_020_704, w_020_705, w_020_706, w_020_707, w_020_708, w_020_709, w_020_710, w_020_711, w_020_712, w_020_713, w_020_714, w_020_715, w_020_716, w_020_717, w_020_718, w_020_719, w_020_720, w_020_721, w_020_722, w_020_723, w_020_724, w_020_725, w_020_726, w_020_727, w_020_728, w_020_729, w_020_730, w_020_731, w_020_732, w_020_733, w_020_734, w_020_735, w_020_736, w_020_738, w_020_739, w_020_740, w_020_741, w_020_742, w_020_743, w_020_744, w_020_745, w_020_746, w_020_747, w_020_748, w_020_749, w_020_750, w_020_752, w_020_753, w_020_754, w_020_755, w_020_756, w_020_757, w_020_758, w_020_759, w_020_760, w_020_761, w_020_762, w_020_763, w_020_764, w_020_765, w_020_766, w_020_767, w_020_768, w_020_769, w_020_771, w_020_772, w_020_773, w_020_774, w_020_775, w_020_776, w_020_777, w_020_780, w_020_781, w_020_782, w_020_784, w_020_785, w_020_787, w_020_788, w_020_789, w_020_790, w_020_791, w_020_792, w_020_793, w_020_794, w_020_795, w_020_796, w_020_797, w_020_798, w_020_799, w_020_801, w_020_802, w_020_803, w_020_804, w_020_805, w_020_806, w_020_807, w_020_808, w_020_809, w_020_811, w_020_812, w_020_813, w_020_814, w_020_815, w_020_816, w_020_817, w_020_818, w_020_819, w_020_820, w_020_821, w_020_822, w_020_824, w_020_826, w_020_827, w_020_829, w_020_830, w_020_831, w_020_832, w_020_833, w_020_834, w_020_835, w_020_836, w_020_837, w_020_838, w_020_839, w_020_840, w_020_841, w_020_842, w_020_843, w_020_845, w_020_846, w_020_847, w_020_848, w_020_849, w_020_850, w_020_851, w_020_852, w_020_853, w_020_854, w_020_855, w_020_856, w_020_857, w_020_858, w_020_862, w_020_863, w_020_864, w_020_865, w_020_866, w_020_867, w_020_868, w_020_869, w_020_871, w_020_872, w_020_873, w_020_874, w_020_875, w_020_876, w_020_877, w_020_878, w_020_879, w_020_880, w_020_881, w_020_882, w_020_883, w_020_884, w_020_885, w_020_886, w_020_887, w_020_888, w_020_889, w_020_890, w_020_892, w_020_893, w_020_894, w_020_895, w_020_896, w_020_897, w_020_898, w_020_901, w_020_903, w_020_904, w_020_905, w_020_906, w_020_907, w_020_908, w_020_909, w_020_910, w_020_911, w_020_913, w_020_914, w_020_915, w_020_917, w_020_918, w_020_919, w_020_920, w_020_921, w_020_922, w_020_923, w_020_924, w_020_925, w_020_926, w_020_927, w_020_928, w_020_929, w_020_930, w_020_931, w_020_932, w_020_933, w_020_934, w_020_935, w_020_936, w_020_937, w_020_938, w_020_939, w_020_940, w_020_941, w_020_942, w_020_943, w_020_944, w_020_948, w_020_950, w_020_951, w_020_952, w_020_953, w_020_954, w_020_955, w_020_956, w_020_957, w_020_959, w_020_960, w_020_961, w_020_962, w_020_963, w_020_964, w_020_966, w_020_967, w_020_969, w_020_970, w_020_971, w_020_972, w_020_973, w_020_974, w_020_976, w_020_977, w_020_978, w_020_979, w_020_980, w_020_981, w_020_982, w_020_984, w_020_985, w_020_986, w_020_989, w_020_991, w_020_992, w_020_993, w_020_994, w_020_995, w_020_996, w_020_997, w_020_998, w_020_1000, w_020_1001, w_020_1002, w_020_1003, w_020_1005, w_020_1006, w_020_1007, w_020_1008, w_020_1010, w_020_1011, w_020_1012, w_020_1013, w_020_1014, w_020_1016, w_020_1017, w_020_1018, w_020_1019, w_020_1020, w_020_1021, w_020_1022, w_020_1023, w_020_1024, w_020_1025, w_020_1026, w_020_1028, w_020_1029, w_020_1030, w_020_1031, w_020_1032, w_020_1033, w_020_1034, w_020_1035, w_020_1036, w_020_1037, w_020_1038, w_020_1039, w_020_1040, w_020_1041, w_020_1042, w_020_1043, w_020_1044, w_020_1045, w_020_1046, w_020_1047, w_020_1048, w_020_1049, w_020_1050, w_020_1051, w_020_1052, w_020_1053, w_020_1054, w_020_1055, w_020_1056, w_020_1057, w_020_1058, w_020_1059, w_020_1060, w_020_1062, w_020_1063, w_020_1064, w_020_1065, w_020_1066, w_020_1067, w_020_1068, w_020_1069, w_020_1070, w_020_1071, w_020_1072, w_020_1073, w_020_1074, w_020_1076, w_020_1077, w_020_1078, w_020_1079, w_020_1080, w_020_1083, w_020_1084, w_020_1085, w_020_1086, w_020_1087, w_020_1089, w_020_1090, w_020_1091, w_020_1092, w_020_1093, w_020_1094, w_020_1095, w_020_1096, w_020_1097, w_020_1099, w_020_1100, w_020_1101, w_020_1102, w_020_1103, w_020_1105, w_020_1106, w_020_1107, w_020_1108, w_020_1109, w_020_1110, w_020_1111, w_020_1112, w_020_1113, w_020_1115, w_020_1118, w_020_1119, w_020_1120, w_020_1121, w_020_1122, w_020_1123, w_020_1124, w_020_1125, w_020_1126, w_020_1127, w_020_1128, w_020_1129, w_020_1130, w_020_1131, w_020_1132, w_020_1133, w_020_1134, w_020_1135, w_020_1136, w_020_1137, w_020_1139, w_020_1140, w_020_1141, w_020_1142, w_020_1143, w_020_1144, w_020_1145, w_020_1146, w_020_1147, w_020_1148, w_020_1149, w_020_1150, w_020_1151, w_020_1153, w_020_1154, w_020_1155, w_020_1156, w_020_1157, w_020_1158, w_020_1159, w_020_1160, w_020_1161, w_020_1162, w_020_1163, w_020_1164, w_020_1165, w_020_1166, w_020_1167, w_020_1168, w_020_1169, w_020_1170, w_020_1171, w_020_1172, w_020_1173, w_020_1174, w_020_1175, w_020_1176, w_020_1177, w_020_1178, w_020_1179, w_020_1180, w_020_1182, w_020_1183, w_020_1184, w_020_1185, w_020_1186, w_020_1187, w_020_1188, w_020_1189, w_020_1190, w_020_1191, w_020_1192, w_020_1193, w_020_1195, w_020_1196, w_020_1197, w_020_1199, w_020_1200, w_020_1201, w_020_1202, w_020_1204, w_020_1205, w_020_1206, w_020_1207, w_020_1208, w_020_1209, w_020_1210, w_020_1211, w_020_1212, w_020_1213, w_020_1214, w_020_1215, w_020_1216, w_020_1217, w_020_1218, w_020_1219, w_020_1220, w_020_1221, w_020_1224, w_020_1225, w_020_1226, w_020_1227, w_020_1228, w_020_1229, w_020_1230, w_020_1231, w_020_1232, w_020_1233, w_020_1235, w_020_1236, w_020_1237, w_020_1239, w_020_1240, w_020_1242, w_020_1243, w_020_1244, w_020_1245, w_020_1246, w_020_1247, w_020_1248, w_020_1249, w_020_1250, w_020_1251, w_020_1252, w_020_1253, w_020_1255, w_020_1256, w_020_1258, w_020_1259, w_020_1260, w_020_1261, w_020_1262, w_020_1263, w_020_1264, w_020_1265, w_020_1266, w_020_1267, w_020_1268, w_020_1269, w_020_1270, w_020_1271, w_020_1272, w_020_1273, w_020_1274, w_020_1275, w_020_1276, w_020_1277, w_020_1278, w_020_1279, w_020_1282, w_020_1283, w_020_1284, w_020_1286, w_020_1288, w_020_1289, w_020_1290, w_020_1291, w_020_1292, w_020_1294, w_020_1295, w_020_1296, w_020_1297, w_020_1298, w_020_1299, w_020_1300, w_020_1302, w_020_1304, w_020_1305, w_020_1306, w_020_1307, w_020_1308, w_020_1309, w_020_1310, w_020_1312, w_020_1313, w_020_1314, w_020_1315, w_020_1316, w_020_1317, w_020_1318, w_020_1320, w_020_1321, w_020_1322, w_020_1323, w_020_1324, w_020_1325, w_020_1326, w_020_1327, w_020_1328, w_020_1329, w_020_1330, w_020_1331, w_020_1332, w_020_1333, w_020_1334, w_020_1335, w_020_1336, w_020_1337, w_020_1338, w_020_1339, w_020_1340, w_020_1341, w_020_1342, w_020_1343, w_020_1344, w_020_1345, w_020_1347, w_020_1348, w_020_1349, w_020_1350, w_020_1352, w_020_1353, w_020_1354, w_020_1355, w_020_1356, w_020_1357, w_020_1358, w_020_1359, w_020_1360, w_020_1361, w_020_1362, w_020_1364, w_020_1365, w_020_1366, w_020_1367, w_020_1370, w_020_1371, w_020_1372, w_020_1373, w_020_1374, w_020_1376, w_020_1377, w_020_1379, w_020_1380, w_020_1381, w_020_1382, w_020_1384, w_020_1385, w_020_1386, w_020_1387, w_020_1388, w_020_1389, w_020_1390, w_020_1391, w_020_1392, w_020_1393, w_020_1394, w_020_1395, w_020_1396, w_020_1397, w_020_1398, w_020_1399, w_020_1400, w_020_1401, w_020_1402, w_020_1403, w_020_1404, w_020_1405, w_020_1406, w_020_1407, w_020_1408, w_020_1409, w_020_1411, w_020_1412, w_020_1413, w_020_1414, w_020_1415, w_020_1416, w_020_1417, w_020_1418, w_020_1419, w_020_1422, w_020_1423, w_020_1425, w_020_1426, w_020_1427, w_020_1428, w_020_1429, w_020_1430, w_020_1431, w_020_1432, w_020_1433, w_020_1434, w_020_1435, w_020_1436, w_020_1437, w_020_1438, w_020_1439, w_020_1440, w_020_1441, w_020_1442, w_020_1443, w_020_1444, w_020_1445, w_020_1446, w_020_1447, w_020_1449, w_020_1450, w_020_1451, w_020_1452, w_020_1453, w_020_1454, w_020_1455, w_020_1456, w_020_1457, w_020_1458, w_020_1459, w_020_1460, w_020_1461, w_020_1463, w_020_1464, w_020_1465, w_020_1466, w_020_1467, w_020_1470, w_020_1471, w_020_1472, w_020_1473, w_020_1475, w_020_1476, w_020_1477, w_020_1478, w_020_1479, w_020_1480, w_020_1481, w_020_1482, w_020_1483, w_020_1484, w_020_1485, w_020_1486, w_020_1488, w_020_1489, w_020_1491, w_020_1493, w_020_1494, w_020_1495, w_020_1496, w_020_1497, w_020_1498, w_020_1499, w_020_1500, w_020_1501, w_020_1502, w_020_1503, w_020_1504, w_020_1505, w_020_1506, w_020_1507, w_020_1508, w_020_1509, w_020_1510, w_020_1511, w_020_1512, w_020_1513, w_020_1514, w_020_1516, w_020_1517, w_020_1518, w_020_1519, w_020_1520, w_020_1521, w_020_1522, w_020_1523, w_020_1524, w_020_1527, w_020_1528, w_020_1529, w_020_1530, w_020_1532, w_020_1533, w_020_1535, w_020_1537, w_020_1538, w_020_1539, w_020_1540, w_020_1541, w_020_1542, w_020_1543, w_020_1544, w_020_1545, w_020_1546, w_020_1547, w_020_1548, w_020_1549, w_020_1550, w_020_1552, w_020_1553, w_020_1554, w_020_1555, w_020_1556, w_020_1557, w_020_1558, w_020_1559, w_020_1560, w_020_1561, w_020_1562, w_020_1563, w_020_1564, w_020_1565, w_020_1566, w_020_1567, w_020_1568, w_020_1569, w_020_1571, w_020_1572, w_020_1573, w_020_1574, w_020_1575, w_020_1576, w_020_1577, w_020_1578, w_020_1579, w_020_1580, w_020_1581, w_020_1582, w_020_1583, w_020_1584, w_020_1585, w_020_1586, w_020_1587, w_020_1588, w_020_1589, w_020_1590, w_020_1591, w_020_1592, w_020_1593, w_020_1594, w_020_1595, w_020_1596, w_020_1597, w_020_1598, w_020_1599, w_020_1600, w_020_1601, w_020_1602, w_020_1604, w_020_1605, w_020_1606, w_020_1607, w_020_1608, w_020_1610, w_020_1611, w_020_1612, w_020_1613, w_020_1614, w_020_1615, w_020_1616, w_020_1617, w_020_1618, w_020_1620, w_020_1621, w_020_1622, w_020_1623, w_020_1624, w_020_1626, w_020_1629, w_020_1631, w_020_1632, w_020_1633, w_020_1634, w_020_1635, w_020_1636, w_020_1637, w_020_1638, w_020_1639, w_020_1640, w_020_1641, w_020_1643, w_020_1645, w_020_1646, w_020_1647, w_020_1648, w_020_1649, w_020_1651, w_020_1652, w_020_1654, w_020_1655, w_020_1657, w_020_1658, w_020_1659, w_020_1660, w_020_1661, w_020_1662, w_020_1663, w_020_1664, w_020_1665, w_020_1666, w_020_1667, w_020_1668, w_020_1669, w_020_1670, w_020_1671, w_020_1672, w_020_1673, w_020_1674, w_020_1675, w_020_1677, w_020_1678, w_020_1679, w_020_1680, w_020_1681, w_020_1682, w_020_1683, w_020_1684, w_020_1685, w_020_1686, w_020_1687, w_020_1688, w_020_1689, w_020_1690, w_020_1691, w_020_1692, w_020_1695, w_020_1696, w_020_1697, w_020_1699, w_020_1700, w_020_1701, w_020_1702, w_020_1703, w_020_1704, w_020_1705, w_020_1706, w_020_1707, w_020_1710, w_020_1711, w_020_1712, w_020_1713, w_020_1714, w_020_1715, w_020_1716, w_020_1717, w_020_1721, w_020_1722, w_020_1723, w_020_1725, w_020_1726, w_020_1727, w_020_1728, w_020_1731, w_020_1732, w_020_1733, w_020_1734, w_020_1735, w_020_1736, w_020_1738, w_020_1739, w_020_1740, w_020_1741, w_020_1742, w_020_1743, w_020_1744, w_020_1745, w_020_1746, w_020_1747, w_020_1748, w_020_1749, w_020_1750, w_020_1751, w_020_1752, w_020_1754, w_020_1755, w_020_1756, w_020_1757, w_020_1758, w_020_1759, w_020_1760, w_020_1761, w_020_1762, w_020_1763, w_020_1764, w_020_1765, w_020_1766, w_020_1767, w_020_1768, w_020_1769, w_020_1770, w_020_1772, w_020_1774, w_020_1775, w_020_1777, w_020_1778, w_020_1779, w_020_1780, w_020_1781, w_020_1782, w_020_1783, w_020_1784, w_020_1785, w_020_1786, w_020_1787, w_020_1788, w_020_1789, w_020_1790, w_020_1791, w_020_1793, w_020_1794, w_020_1795, w_020_1796, w_020_1799, w_020_1800, w_020_1802, w_020_1803, w_020_1804, w_020_1805, w_020_1806, w_020_1807, w_020_1808, w_020_1809, w_020_1811, w_020_1812, w_020_1813, w_020_1814, w_020_1815, w_020_1816, w_020_1817, w_020_1819, w_020_1820, w_020_1821, w_020_1822, w_020_1823, w_020_1824, w_020_1825, w_020_1827, w_020_1828, w_020_1829, w_020_1830, w_020_1831, w_020_1832, w_020_1833, w_020_1834, w_020_1835, w_020_1836, w_020_1839, w_020_1840, w_020_1841, w_020_1842, w_020_1843, w_020_1844, w_020_1845, w_020_1846, w_020_1848, w_020_1849, w_020_1851, w_020_1852, w_020_1853, w_020_1854, w_020_1855, w_020_1856, w_020_1858, w_020_1859, w_020_1860, w_020_1862, w_020_1863, w_020_1865, w_020_1866, w_020_1867, w_020_1868, w_020_1869, w_020_1870, w_020_1871, w_020_1873, w_020_1874, w_020_1875, w_020_1876, w_020_1877, w_020_1879, w_020_1880, w_020_1881, w_020_1882, w_020_1883, w_020_1884, w_020_1885, w_020_1887, w_020_1888, w_020_1889, w_020_1890, w_020_1891, w_020_1892, w_020_1893, w_020_1894, w_020_1895, w_020_1896, w_020_1897, w_020_1898, w_020_1899, w_020_1900, w_020_1901, w_020_1902, w_020_1903, w_020_1904, w_020_1906, w_020_1907, w_020_1908, w_020_1909, w_020_1910, w_020_1911, w_020_1912, w_020_1913, w_020_1914, w_020_1916, w_020_1917, w_020_1918, w_020_1919, w_020_1920, w_020_1921, w_020_1922, w_020_1924, w_020_1925, w_020_1926, w_020_1927, w_020_1928, w_020_1930, w_020_1931, w_020_1934, w_020_1936, w_020_1938, w_020_1939, w_020_1940, w_020_1941, w_020_1942, w_020_1943, w_020_1944, w_020_1945, w_020_1946, w_020_1947, w_020_1949, w_020_1950, w_020_1951, w_020_1952, w_020_1953, w_020_1954, w_020_1955, w_020_1956, w_020_1957, w_020_1958, w_020_1959, w_020_1960, w_020_1961, w_020_1962, w_020_1963, w_020_1964, w_020_1965, w_020_1968, w_020_1970, w_020_1971, w_020_1972, w_020_1974, w_020_1976, w_020_1977, w_020_1978, w_020_1979, w_020_1980, w_020_1981, w_020_1983, w_020_1984, w_020_1986, w_020_1987, w_020_1988, w_020_1990, w_020_1991, w_020_1992, w_020_1993, w_020_1994, w_020_1996, w_020_1997, w_020_1998, w_020_1999, w_020_2000, w_020_2001, w_020_2002, w_020_2003, w_020_2004, w_020_2005, w_020_2006, w_020_2007, w_020_2008, w_020_2009, w_020_2010, w_020_2011, w_020_2012, w_020_2014, w_020_2015, w_020_2017, w_020_2018, w_020_2019, w_020_2021, w_020_2022, w_020_2023, w_020_2024, w_020_2025, w_020_2027, w_020_2029, w_020_2030, w_020_2031, w_020_2032, w_020_2033, w_020_2034, w_020_2035, w_020_2036, w_020_2037, w_020_2038, w_020_2040, w_020_2042, w_020_2044, w_020_2045, w_020_2046, w_020_2047, w_020_2048, w_020_2049, w_020_2050, w_020_2052, w_020_2053, w_020_2054, w_020_2055, w_020_2056, w_020_2057, w_020_2058, w_020_2059, w_020_2060, w_020_2061, w_020_2062, w_020_2063, w_020_2065, w_020_2066, w_020_2067, w_020_2068, w_020_2069, w_020_2070, w_020_2071, w_020_2072, w_020_2073, w_020_2075, w_020_2076, w_020_2077, w_020_2078, w_020_2079, w_020_2080, w_020_2081, w_020_2082, w_020_2083, w_020_2084, w_020_2085, w_020_2086, w_020_2088, w_020_2089, w_020_2090, w_020_2092, w_020_2093, w_020_2094, w_020_2095, w_020_2096, w_020_2097, w_020_2098, w_020_2100, w_020_2101, w_020_2102, w_020_2103, w_020_2104, w_020_2105, w_020_2108, w_020_2110, w_020_2111, w_020_2112, w_020_2113, w_020_2114, w_020_2115, w_020_2117, w_020_2118, w_020_2119, w_020_2121, w_020_2122, w_020_2123, w_020_2124, w_020_2125, w_020_2126, w_020_2127, w_020_2128, w_020_2130, w_020_2131, w_020_2132, w_020_2133, w_020_2134, w_020_2135, w_020_2137, w_020_2138, w_020_2141, w_020_2142, w_020_2143, w_020_2144, w_020_2145, w_020_2146, w_020_2147, w_020_2149, w_020_2150, w_020_2153, w_020_2154, w_020_2155, w_020_2156, w_020_2157, w_020_2158, w_020_2159, w_020_2160, w_020_2161, w_020_2162, w_020_2163, w_020_2165, w_020_2167, w_020_2168, w_020_2169, w_020_2170, w_020_2171, w_020_2172, w_020_2173, w_020_2174, w_020_2175, w_020_2178, w_020_2179, w_020_2180, w_020_2181, w_020_2182, w_020_2183, w_020_2184, w_020_2186, w_020_2187, w_020_2188, w_020_2189, w_020_2190, w_020_2193, w_020_2194, w_020_2195, w_020_2196, w_020_2197, w_020_2198, w_020_2199, w_020_2200, w_020_2201, w_020_2203, w_020_2204, w_020_2205, w_020_2206, w_020_2207, w_020_2208, w_020_2209, w_020_2210, w_020_2211, w_020_2212, w_020_2213, w_020_2214, w_020_2215, w_020_2216, w_020_2217, w_020_2218, w_020_2219, w_020_2220, w_020_2222, w_020_2223, w_020_2224, w_020_2225, w_020_2226, w_020_2227, w_020_2228, w_020_2229, w_020_2230, w_020_2231, w_020_2232, w_020_2236, w_020_2239, w_020_2241, w_020_2243, w_020_2245, w_020_2246, w_020_2247, w_020_2248, w_020_2250, w_020_2253, w_020_2254, w_020_2255, w_020_2256, w_020_2257, w_020_2259, w_020_2260, w_020_2261, w_020_2264, w_020_2265, w_020_2266, w_020_2267, w_020_2271, w_020_2274, w_020_2275, w_020_2276, w_020_2277, w_020_2278, w_020_2279, w_020_2280, w_020_2281, w_020_2282, w_020_2283, w_020_2285, w_020_2288, w_020_2289, w_020_2291, w_020_2292, w_020_2294, w_020_2296, w_020_2298, w_020_2299, w_020_2300, w_020_2303, w_020_2305, w_020_2306, w_020_2307, w_020_2309, w_020_2310, w_020_2313, w_020_2314, w_020_2317, w_020_2318, w_020_2319, w_020_2320, w_020_2321, w_020_2323, w_020_2324, w_020_2325, w_020_2326, w_020_2327, w_020_2328, w_020_2329, w_020_2331, w_020_2332, w_020_2333, w_020_2334, w_020_2335, w_020_2336, w_020_2338, w_020_2339, w_020_2340, w_020_2343, w_020_2344, w_020_2345, w_020_2346, w_020_2348, w_020_2350, w_020_2351, w_020_2353, w_020_2356, w_020_2357, w_020_2360, w_020_2361, w_020_2364, w_020_2366, w_020_2369, w_020_2370, w_020_2371, w_020_2372, w_020_2373, w_020_2374, w_020_2375, w_020_2376, w_020_2377, w_020_2378, w_020_2379, w_020_2383, w_020_2384, w_020_2385, w_020_2386, w_020_2387, w_020_2389, w_020_2390, w_020_2393, w_020_2394, w_020_2395, w_020_2397, w_020_2398, w_020_2399, w_020_2400, w_020_2402, w_020_2404, w_020_2405, w_020_2406, w_020_2407, w_020_2409, w_020_2411, w_020_2414, w_020_2415, w_020_2416, w_020_2417, w_020_2418, w_020_2422, w_020_2423, w_020_2426, w_020_2428, w_020_2429, w_020_2432, w_020_2433, w_020_2435, w_020_2436, w_020_2439, w_020_2440, w_020_2441, w_020_2442, w_020_2444, w_020_2445, w_020_2446, w_020_2447, w_020_2449, w_020_2450, w_020_2451, w_020_2452, w_020_2454, w_020_2456, w_020_2457, w_020_2459, w_020_2460, w_020_2461, w_020_2462, w_020_2464, w_020_2466, w_020_2468, w_020_2470, w_020_2473, w_020_2476, w_020_2477, w_020_2479, w_020_2480, w_020_2485, w_020_2486, w_020_2487, w_020_2489, w_020_2490, w_020_2491, w_020_2492, w_020_2496, w_020_2499, w_020_2500, w_020_2501, w_020_2502, w_020_2505, w_020_2506, w_020_2507, w_020_2509, w_020_2510, w_020_2512, w_020_2514, w_020_2515, w_020_2516, w_020_2517, w_020_2519, w_020_2520, w_020_2521, w_020_2524, w_020_2525, w_020_2527, w_020_2528, w_020_2529, w_020_2530, w_020_2531, w_020_2532, w_020_2533, w_020_2535, w_020_2539, w_020_2540, w_020_2541, w_020_2549, w_020_2550, w_020_2551, w_020_2552, w_020_2553, w_020_2554, w_020_2557, w_020_2558, w_020_2560, w_020_2561, w_020_2562, w_020_2564, w_020_2565, w_020_2566, w_020_2567, w_020_2569, w_020_2573, w_020_2574, w_020_2575, w_020_2576, w_020_2577, w_020_2578, w_020_2579, w_020_2580, w_020_2581, w_020_2582, w_020_2583, w_020_2584, w_020_2585, w_020_2586, w_020_2587, w_020_2588, w_020_2589, w_020_2590, w_020_2591, w_020_2592, w_020_2594, w_020_2596, w_020_2597, w_020_2598, w_020_2599, w_020_2601, w_020_2602, w_020_2603, w_020_2604, w_020_2605, w_020_2608, w_020_2612, w_020_2614, w_020_2616, w_020_2618, w_020_2619, w_020_2620, w_020_2621, w_020_2622, w_020_2623, w_020_2624, w_020_2627, w_020_2628, w_020_2629, w_020_2630, w_020_2632, w_020_2633, w_020_2634, w_020_2635, w_020_2636, w_020_2637, w_020_2639, w_020_2644, w_020_2645, w_020_2646, w_020_2650, w_020_2652, w_020_2653, w_020_2654, w_020_2655, w_020_2657, w_020_2658, w_020_2660, w_020_2662, w_020_2663, w_020_2664, w_020_2665, w_020_2666, w_020_2668, w_020_2670, w_020_2677, w_020_2679, w_020_2680, w_020_2681, w_020_2682, w_020_2683, w_020_2685, w_020_2686, w_020_2689, w_020_2691, w_020_2693, w_020_2694, w_020_2696, w_020_2698, w_020_2699, w_020_2700, w_020_2702, w_020_2703, w_020_2705, w_020_2708, w_020_2709, w_020_2710, w_020_2713, w_020_2714, w_020_2718, w_020_2719, w_020_2720, w_020_2721, w_020_2723, w_020_2725, w_020_2726, w_020_2729, w_020_2730, w_020_2731, w_020_2732, w_020_2733, w_020_2734, w_020_2735, w_020_2736, w_020_2737, w_020_2738, w_020_2740, w_020_2741, w_020_2744, w_020_2745, w_020_2747, w_020_2750, w_020_2751, w_020_2752, w_020_2753, w_020_2754, w_020_2755, w_020_2758, w_020_2759, w_020_2761, w_020_2762, w_020_2763, w_020_2764, w_020_2767, w_020_2768, w_020_2771, w_020_2772, w_020_2774, w_020_2775, w_020_2776, w_020_2779, w_020_2781, w_020_2782, w_020_2783, w_020_2785, w_020_2786, w_020_2788, w_020_2789, w_020_2792, w_020_2795, w_020_2796, w_020_2797, w_020_2798, w_020_2799, w_020_2800, w_020_2801, w_020_2802, w_020_2803, w_020_2804, w_020_2807, w_020_2808, w_020_2813, w_020_2814, w_020_2815, w_020_2816, w_020_2817, w_020_2818, w_020_2820, w_020_2821, w_020_2822, w_020_2823, w_020_2824, w_020_2827, w_020_2829, w_020_2830, w_020_2832, w_020_2833, w_020_2834, w_020_2835, w_020_2836, w_020_2839, w_020_2840, w_020_2841, w_020_2842, w_020_2844, w_020_2845, w_020_2846, w_020_2847, w_020_2848, w_020_2849, w_020_2850, w_020_2853, w_020_2854, w_020_2860, w_020_2861, w_020_2862, w_020_2864, w_020_2867, w_020_2868, w_020_2869, w_020_2873, w_020_2875, w_020_2876, w_020_2880, w_020_2881, w_020_2883, w_020_2884, w_020_2886, w_020_2887, w_020_2888, w_020_2889, w_020_2891, w_020_2893, w_020_2894, w_020_2896, w_020_2899, w_020_2900, w_020_2901, w_020_2902, w_020_2905, w_020_2906, w_020_2908, w_020_2911, w_020_2915, w_020_2918, w_020_2919, w_020_2920, w_020_2921, w_020_2923, w_020_2924, w_020_2927, w_020_2929, w_020_2931, w_020_2934, w_020_2935, w_020_2937, w_020_2938, w_020_2940, w_020_2942, w_020_2944, w_020_2945, w_020_2946, w_020_2947, w_020_2948, w_020_2949, w_020_2950, w_020_2951, w_020_2952, w_020_2954, w_020_2956, w_020_2957, w_020_2958, w_020_2959, w_020_2962, w_020_2963, w_020_2964, w_020_2967, w_020_2968, w_020_2969, w_020_2971, w_020_2975, w_020_2976, w_020_2977, w_020_2978, w_020_2980, w_020_2981, w_020_2982, w_020_2983, w_020_2986, w_020_2987, w_020_2988, w_020_2991, w_020_2992, w_020_2994, w_020_2997, w_020_2998, w_020_2999, w_020_3000, w_020_3002, w_020_3003, w_020_3004, w_020_3005, w_020_3007, w_020_3009, w_020_3011, w_020_3012, w_020_3016, w_020_3019, w_020_3020, w_020_3022, w_020_3023, w_020_3024, w_020_3025, w_020_3029, w_020_3030, w_020_3032, w_020_3036, w_020_3037, w_020_3038, w_020_3042, w_020_3044, w_020_3045, w_020_3047, w_020_3048, w_020_3050, w_020_3051, w_020_3052, w_020_3053, w_020_3054, w_020_3055, w_020_3056, w_020_3058, w_020_3059, w_020_3060, w_020_3061, w_020_3064, w_020_3065, w_020_3066, w_020_3067, w_020_3071, w_020_3072, w_020_3074, w_020_3075, w_020_3076, w_020_3078, w_020_3081, w_020_3084, w_020_3087, w_020_3088, w_020_3089, w_020_3090, w_020_3092, w_020_3094, w_020_3095, w_020_3096, w_020_3097, w_020_3098, w_020_3099, w_020_3101, w_020_3103, w_020_3105, w_020_3106, w_020_3109, w_020_3110, w_020_3111, w_020_3112, w_020_3113, w_020_3114, w_020_3115, w_020_3116, w_020_3119, w_020_3121, w_020_3122, w_020_3123, w_020_3124, w_020_3125, w_020_3127, w_020_3130, w_020_3131, w_020_3133, w_020_3135, w_020_3136, w_020_3139, w_020_3143, w_020_3145, w_020_3146, w_020_3147, w_020_3148, w_020_3149, w_020_3150, w_020_3151, w_020_3152, w_020_3153, w_020_3154, w_020_3155, w_020_3156, w_020_3157, w_020_3158, w_020_3161, w_020_3162, w_020_3163, w_020_3165, w_020_3166, w_020_3168, w_020_3170, w_020_3171, w_020_3176, w_020_3177, w_020_3178, w_020_3179, w_020_3181, w_020_3182, w_020_3183, w_020_3185, w_020_3188, w_020_3190, w_020_3192, w_020_3194, w_020_3195, w_020_3196, w_020_3197, w_020_3198, w_020_3199, w_020_3200, w_020_3201, w_020_3202, w_020_3203, w_020_3205, w_020_3206, w_020_3208, w_020_3210, w_020_3212, w_020_3214, w_020_3216, w_020_3218, w_020_3220, w_020_3222, w_020_3223, w_020_3224, w_020_3225, w_020_3227, w_020_3228, w_020_3229, w_020_3230, w_020_3231, w_020_3232, w_020_3233, w_020_3235, w_020_3236, w_020_3237, w_020_3238, w_020_3240, w_020_3244, w_020_3245, w_020_3249, w_020_3251, w_020_3252, w_020_3253, w_020_3256, w_020_3257, w_020_3258, w_020_3259, w_020_3260, w_020_3262, w_020_3263, w_020_3264, w_020_3265, w_020_3269, w_020_3270, w_020_3272, w_020_3274, w_020_3275, w_020_3277, w_020_3278, w_020_3279, w_020_3280, w_020_3282, w_020_3283, w_020_3284, w_020_3285, w_020_3286, w_020_3287, w_020_3289, w_020_3290, w_020_3292, w_020_3294, w_020_3296, w_020_3297, w_020_3302, w_020_3303, w_020_3304, w_020_3305, w_020_3308, w_020_3310, w_020_3313, w_020_3314, w_020_3316, w_020_3317, w_020_3319, w_020_3320, w_020_3324, w_020_3326, w_020_3327, w_020_3330, w_020_3331, w_020_3332, w_020_3333, w_020_3334, w_020_3335, w_020_3336, w_020_3338, w_020_3341, w_020_3343, w_020_3346, w_020_3347, w_020_3349, w_020_3351, w_020_3353, w_020_3356, w_020_3357, w_020_3359, w_020_3360, w_020_3361, w_020_3364, w_020_3366, w_020_3368, w_020_3369, w_020_3370, w_020_3371, w_020_3372, w_020_3375, w_020_3377, w_020_3382, w_020_3383, w_020_3384, w_020_3386, w_020_3388, w_020_3389, w_020_3390, w_020_3391, w_020_3392, w_020_3393, w_020_3395, w_020_3396, w_020_3397, w_020_3398, w_020_3399, w_020_3400, w_020_3403, w_020_3405, w_020_3407, w_020_3410, w_020_3411, w_020_3412, w_020_3413, w_020_3414, w_020_3418, w_020_3419, w_020_3420, w_020_3421, w_020_3422, w_020_3430, w_020_3431, w_020_3437, w_020_3439, w_020_3441, w_020_3443, w_020_3444, w_020_3446, w_020_3449, w_020_3450, w_020_3451, w_020_3452, w_020_3453, w_020_3455, w_020_3456, w_020_3457, w_020_3459, w_020_3460, w_020_3461, w_020_3462, w_020_3464, w_020_3465, w_020_3466, w_020_3470, w_020_3472, w_020_3473, w_020_3477, w_020_3478, w_020_3481, w_020_3482, w_020_3483, w_020_3484, w_020_3485, w_020_3486, w_020_3487, w_020_3488, w_020_3489, w_020_3492, w_020_3494, w_020_3496, w_020_3498, w_020_3499, w_020_3500, w_020_3502, w_020_3505, w_020_3508, w_020_3509, w_020_3510, w_020_3511, w_020_3512, w_020_3513, w_020_3514, w_020_3515, w_020_3517, w_020_3518, w_020_3520, w_020_3522, w_020_3523, w_020_3525, w_020_3529, w_020_3532, w_020_3533, w_020_3535, w_020_3536, w_020_3539, w_020_3540, w_020_3541, w_020_3544, w_020_3545, w_020_3546, w_020_3548, w_020_3550, w_020_3551, w_020_3555, w_020_3556, w_020_3557, w_020_3558, w_020_3560, w_020_3561, w_020_3563, w_020_3564, w_020_3566, w_020_3567, w_020_3568, w_020_3570, w_020_3572, w_020_3575, w_020_3576, w_020_3578, w_020_3580, w_020_3581, w_020_3583, w_020_3584, w_020_3587, w_020_3589, w_020_3592, w_020_3593, w_020_3595, w_020_3596, w_020_3598, w_020_3599, w_020_3600, w_020_3602, w_020_3605, w_020_3606, w_020_3607, w_020_3608, w_020_3610, w_020_3611, w_020_3612, w_020_3613, w_020_3614, w_020_3616, w_020_3617, w_020_3618, w_020_3620, w_020_3622, w_020_3623, w_020_3625, w_020_3626, w_020_3627, w_020_3628, w_020_3629, w_020_3630, w_020_3631, w_020_3633, w_020_3635, w_020_3636, w_020_3637, w_020_3639, w_020_3640, w_020_3641, w_020_3642, w_020_3643, w_020_3644, w_020_3645, w_020_3647, w_020_3648, w_020_3650, w_020_3654, w_020_3656, w_020_3657, w_020_3659, w_020_3662, w_020_3664, w_020_3665, w_020_3666, w_020_3668, w_020_3671, w_020_3672, w_020_3674, w_020_3675, w_020_3676, w_020_3677, w_020_3679, w_020_3681, w_020_3682, w_020_3683, w_020_3684, w_020_3685, w_020_3688, w_020_3690, w_020_3692, w_020_3693, w_020_3697, w_020_3698, w_020_3699, w_020_3700, w_020_3701, w_020_3705, w_020_3706, w_020_3707, w_020_3708, w_020_3709, w_020_3710, w_020_3711, w_020_3712, w_020_3713, w_020_3715, w_020_3716, w_020_3717, w_020_3719, w_020_3720, w_020_3722, w_020_3723, w_020_3724, w_020_3725, w_020_3727, w_020_3728, w_020_3729, w_020_3730, w_020_3734, w_020_3735, w_020_3738, w_020_3741, w_020_3742, w_020_3744, w_020_3745, w_020_3747, w_020_3748, w_020_3749, w_020_3750, w_020_3751, w_020_3752, w_020_3753, w_020_3754, w_020_3756, w_020_3757, w_020_3758, w_020_3759, w_020_3761, w_020_3765, w_020_3767, w_020_3771, w_020_3773, w_020_3774, w_020_3775, w_020_3777, w_020_3778, w_020_3781, w_020_3782, w_020_3783, w_020_3784, w_020_3785, w_020_3786, w_020_3787, w_020_3788, w_020_3791, w_020_3792, w_020_3794, w_020_3795, w_020_3797, w_020_3798, w_020_3799, w_020_3801, w_020_3802, w_020_3803, w_020_3804, w_020_3806, w_020_3807, w_020_3808, w_020_3809, w_020_3811, w_020_3813, w_020_3814, w_020_3815, w_020_3817, w_020_3819, w_020_3821, w_020_3822, w_020_3823, w_020_3825, w_020_3826, w_020_3832, w_020_3834, w_020_3835, w_020_3836, w_020_3837, w_020_3839, w_020_3840, w_020_3841, w_020_3842, w_020_3843, w_020_3845, w_020_3848, w_020_3849, w_020_3851, w_020_3853, w_020_3854, w_020_3856, w_020_3861, w_020_3862, w_020_3863, w_020_3865, w_020_3867, w_020_3872, w_020_3874, w_020_3875, w_020_3876, w_020_3877, w_020_3878, w_020_3880, w_020_3881, w_020_3882, w_020_3884, w_020_3885, w_020_3886, w_020_3888, w_020_3889, w_020_3890, w_020_3891, w_020_3893, w_020_3894, w_020_3895, w_020_3896, w_020_3898, w_020_3899, w_020_3900, w_020_3901, w_020_3904, w_020_3905, w_020_3906, w_020_3907, w_020_3908, w_020_3909, w_020_3910, w_020_3911, w_020_3914, w_020_3915, w_020_3916, w_020_3917, w_020_3919, w_020_3920, w_020_3921, w_020_3923, w_020_3924, w_020_3925, w_020_3926, w_020_3927, w_020_3928, w_020_3930, w_020_3936, w_020_3937, w_020_3938, w_020_3940, w_020_3941, w_020_3943, w_020_3945, w_020_3949, w_020_3950, w_020_3951, w_020_3952, w_020_3953, w_020_3954, w_020_3957, w_020_3958, w_020_3959, w_020_3960, w_020_3961, w_020_3962, w_020_3963, w_020_3966, w_020_3967, w_020_3968, w_020_3970, w_020_3971, w_020_3972, w_020_3973, w_020_3974, w_020_3975, w_020_3976, w_020_3978, w_020_3979, w_020_3980, w_020_3981, w_020_3982, w_020_3983, w_020_3984, w_020_3985, w_020_3986, w_020_3989, w_020_3990, w_020_3991, w_020_3992, w_020_3993, w_020_3995, w_020_3996, w_020_3997, w_020_3998, w_020_4000, w_020_4001, w_020_4003, w_020_4005, w_020_4007, w_020_4010, w_020_4013, w_020_4016, w_020_4017, w_020_4019, w_020_4020, w_020_4022, w_020_4023, w_020_4024, w_020_4025, w_020_4026, w_020_4027, w_020_4028, w_020_4029, w_020_4031, w_020_4032, w_020_4034, w_020_4035, w_020_4037, w_020_4039, w_020_4040, w_020_4041, w_020_4042, w_020_4043, w_020_4044, w_020_4046, w_020_4047, w_020_4049, w_020_4050, w_020_4051, w_020_4052, w_020_4054, w_020_4056, w_020_4057, w_020_4064, w_020_4065, w_020_4066, w_020_4069, w_020_4070, w_020_4071, w_020_4072, w_020_4076, w_020_4077, w_020_4078, w_020_4080, w_020_4084, w_020_4086, w_020_4091, w_020_4096, w_020_4097, w_020_4098, w_020_4100, w_020_4101, w_020_4104, w_020_4105, w_020_4106, w_020_4110, w_020_4111, w_020_4113, w_020_4114, w_020_4115, w_020_4116, w_020_4117, w_020_4119, w_020_4120, w_020_4121, w_020_4122, w_020_4123, w_020_4124, w_020_4126, w_020_4127, w_020_4128, w_020_4131, w_020_4133, w_020_4134, w_020_4135, w_020_4136, w_020_4138, w_020_4139, w_020_4140, w_020_4142, w_020_4144, w_020_4145, w_020_4147, w_020_4148, w_020_4149, w_020_4150, w_020_4151, w_020_4152, w_020_4156, w_020_4157, w_020_4160, w_020_4161, w_020_4162, w_020_4163, w_020_4164, w_020_4165, w_020_4166, w_020_4167, w_020_4170, w_020_4171, w_020_4174, w_020_4175, w_020_4176, w_020_4177, w_020_4179, w_020_4181, w_020_4182, w_020_4184, w_020_4187, w_020_4188, w_020_4190, w_020_4191, w_020_4193, w_020_4196, w_020_4199, w_020_4200, w_020_4205, w_020_4210, w_020_4211, w_020_4212, w_020_4214, w_020_4215, w_020_4216, w_020_4217, w_020_4220, w_020_4222, w_020_4223, w_020_4224, w_020_4225, w_020_4227, w_020_4228, w_020_4229, w_020_4230, w_020_4231, w_020_4234, w_020_4236, w_020_4237, w_020_4238, w_020_4239, w_020_4240, w_020_4242, w_020_4243, w_020_4246, w_020_4247, w_020_4250, w_020_4255, w_020_4256, w_020_4260, w_020_4261, w_020_4264, w_020_4265, w_020_4266, w_020_4267, w_020_4268, w_020_4271, w_020_4272, w_020_4274, w_020_4276, w_020_4277, w_020_4279, w_020_4280, w_020_4281, w_020_4282, w_020_4283, w_020_4284, w_020_4285, w_020_4286, w_020_4287, w_020_4288, w_020_4289, w_020_4293, w_020_4294, w_020_4297, w_020_4299, w_020_4301, w_020_4304, w_020_4305, w_020_4306, w_020_4308, w_020_4310, w_020_4313, w_020_4314, w_020_4315, w_020_4318, w_020_4319, w_020_4320, w_020_4324, w_020_4325, w_020_4328, w_020_4329, w_020_4330, w_020_4332, w_020_4334, w_020_4335, w_020_4336, w_020_4337, w_020_4339, w_020_4340, w_020_4342, w_020_4346, w_020_4349, w_020_4356, w_020_4357, w_020_4359, w_020_4361, w_020_4362, w_020_4363, w_020_4364, w_020_4365, w_020_4367, w_020_4369, w_020_4370, w_020_4372, w_020_4374, w_020_4375, w_020_4379, w_020_4380, w_020_4381, w_020_4383, w_020_4384, w_020_4385, w_020_4386, w_020_4387, w_020_4390, w_020_4391, w_020_4393, w_020_4398, w_020_4399, w_020_4401, w_020_4404, w_020_4406, w_020_4408, w_020_4410, w_020_4411, w_020_4413, w_020_4415, w_020_4416, w_020_4417, w_020_4418, w_020_4420, w_020_4422, w_020_4424, w_020_4425, w_020_4427, w_020_4428, w_020_4429, w_020_4430, w_020_4433, w_020_4436, w_020_4437, w_020_4439, w_020_4440, w_020_4442, w_020_4443, w_020_4444, w_020_4445, w_020_4446, w_020_4447, w_020_4448, w_020_4451, w_020_4453, w_020_4455, w_020_4457, w_020_4458, w_020_4459, w_020_4460, w_020_4461, w_020_4462, w_020_4465, w_020_4466, w_020_4467, w_020_4468, w_020_4469, w_020_4470, w_020_4472, w_020_4473, w_020_4475, w_020_4476, w_020_4477, w_020_4478, w_020_4480, w_020_4481, w_020_4482, w_020_4483, w_020_4484, w_020_4486, w_020_4487, w_020_4488, w_020_4490, w_020_4493, w_020_4496, w_020_4498, w_020_4500, w_020_4501, w_020_4502, w_020_4503, w_020_4505, w_020_4506, w_020_4507, w_020_4510, w_020_4511, w_020_4512, w_020_4515, w_020_4517, w_020_4518, w_020_4520, w_020_4523, w_020_4526, w_020_4527, w_020_4528, w_020_4529, w_020_4530, w_020_4532, w_020_4534, w_020_4535, w_020_4536, w_020_4540, w_020_4543, w_020_4544, w_020_4545, w_020_4546, w_020_4547, w_020_4549, w_020_4550, w_020_4551, w_020_4552, w_020_4553, w_020_4554, w_020_4555, w_020_4556, w_020_4557, w_020_4558, w_020_4559, w_020_4560, w_020_4561, w_020_4562, w_020_4563, w_020_4564, w_020_4567, w_020_4569, w_020_4572, w_020_4574, w_020_4575, w_020_4576, w_020_4581, w_020_4582, w_020_4583, w_020_4586, w_020_4587, w_020_4588, w_020_4589, w_020_4590, w_020_4593, w_020_4595, w_020_4596, w_020_4597, w_020_4599, w_020_4600, w_020_4603, w_020_4604, w_020_4605, w_020_4606, w_020_4607, w_020_4608, w_020_4609, w_020_4610, w_020_4613, w_020_4614, w_020_4615, w_020_4619, w_020_4620, w_020_4622, w_020_4623, w_020_4624, w_020_4627, w_020_4629, w_020_4630, w_020_4631, w_020_4636, w_020_4637, w_020_4640, w_020_4641, w_020_4643, w_020_4644, w_020_4646, w_020_4648, w_020_4649, w_020_4650, w_020_4651, w_020_4652, w_020_4653, w_020_4655, w_020_4656, w_020_4657, w_020_4658, w_020_4659, w_020_4660, w_020_4661, w_020_4662, w_020_4664, w_020_4666, w_020_4667, w_020_4668, w_020_4669, w_020_4670, w_020_4671, w_020_4673, w_020_4675, w_020_4676, w_020_4680, w_020_4681, w_020_4682, w_020_4684, w_020_4685, w_020_4686, w_020_4687, w_020_4688, w_020_4689, w_020_4690, w_020_4691, w_020_4692, w_020_4695, w_020_4696, w_020_4697, w_020_4698, w_020_4700, w_020_4702, w_020_4703, w_020_4704, w_020_4706, w_020_4707, w_020_4708, w_020_4709, w_020_4710, w_020_4711, w_020_4712, w_020_4715, w_020_4717, w_020_4718, w_020_4720, w_020_4722, w_020_4723, w_020_4724, w_020_4726, w_020_4727, w_020_4728, w_020_4729, w_020_4730, w_020_4731, w_020_4732, w_020_4735, w_020_4736, w_020_4737, w_020_4738, w_020_4739, w_020_4740, w_020_4742, w_020_4743, w_020_4745, w_020_4746, w_020_4747, w_020_4748, w_020_4749, w_020_4750, w_020_4751, w_020_4752, w_020_4753, w_020_4754, w_020_4755, w_020_4757, w_020_4761, w_020_4764, w_020_4765, w_020_4766, w_020_4767, w_020_4768, w_020_4769, w_020_4772, w_020_4773, w_020_4774, w_020_4775, w_020_4776, w_020_4777, w_020_4778, w_020_4779, w_020_4780, w_020_4781, w_020_4782, w_020_4783, w_020_4785, w_020_4786, w_020_4788, w_020_4789, w_020_4790, w_020_4791, w_020_4792, w_020_4794, w_020_4795, w_020_4796, w_020_4797, w_020_4799, w_020_4801, w_020_4804, w_020_4806, w_020_4807, w_020_4809, w_020_4810, w_020_4811, w_020_4814, w_020_4818, w_020_4820, w_020_4822, w_020_4823, w_020_4824, w_020_4825, w_020_4826, w_020_4828, w_020_4829, w_020_4831, w_020_4832, w_020_4833, w_020_4835, w_020_4836, w_020_4839, w_020_4841, w_020_4842, w_020_4843, w_020_4844, w_020_4845, w_020_4846, w_020_4847, w_020_4848, w_020_4849, w_020_4850, w_020_4851, w_020_4852, w_020_4854, w_020_4855, w_020_4856, w_020_4857, w_020_4859, w_020_4860, w_020_4862, w_020_4863, w_020_4865, w_020_4866, w_020_4867, w_020_4869, w_020_4870, w_020_4872, w_020_4874, w_020_4875, w_020_4877, w_020_4879, w_020_4881, w_020_4882, w_020_4883, w_020_4885, w_020_4886, w_020_4888, w_020_4889, w_020_4890, w_020_4892, w_020_4893, w_020_4894, w_020_4896, w_020_4897, w_020_4898, w_020_4901, w_020_4902, w_020_4903, w_020_4904, w_020_4909, w_020_4910, w_020_4912, w_020_4913, w_020_4915, w_020_4916, w_020_4917, w_020_4918, w_020_4919, w_020_4920, w_020_4923, w_020_4925, w_020_4927, w_020_4928, w_020_4929, w_020_4930, w_020_4931, w_020_4932, w_020_4936, w_020_4937, w_020_4938, w_020_4939, w_020_4940, w_020_4941, w_020_4942, w_020_4943, w_020_4947, w_020_4949, w_020_4950, w_020_4951, w_020_4952, w_020_4954, w_020_4957, w_020_4958, w_020_4959, w_020_4961, w_020_4963, w_020_4965, w_020_4967, w_020_4969, w_020_4970, w_020_4972, w_020_4973, w_020_4975, w_020_4977, w_020_4979, w_020_4983, w_020_4984, w_020_4985, w_020_4986, w_020_4987, w_020_4988, w_020_4989, w_020_4991, w_020_4992, w_020_4994, w_020_4997, w_020_4998, w_020_4999, w_020_5001, w_020_5003, w_020_5005, w_020_5006, w_020_5007, w_020_5008, w_020_5009, w_020_5016, w_020_5017, w_020_5018, w_020_5021, w_020_5022, w_020_5023, w_020_5026, w_020_5027, w_020_5028, w_020_5029, w_020_5030, w_020_5033, w_020_5037, w_020_5040, w_020_5041, w_020_5042, w_020_5043, w_020_5044, w_020_5045, w_020_5046, w_020_5047, w_020_5048, w_020_5049, w_020_5050, w_020_5051, w_020_5052, w_020_5054, w_020_5056, w_020_5058, w_020_5059, w_020_5060, w_020_5061, w_020_5062, w_020_5063, w_020_5064, w_020_5066, w_020_5069, w_020_5070, w_020_5072, w_020_5074, w_020_5076, w_020_5077, w_020_5078, w_020_5079, w_020_5080, w_020_5081, w_020_5082, w_020_5086, w_020_5087, w_020_5088, w_020_5090, w_020_5092, w_020_5093, w_020_5095, w_020_5097, w_020_5098, w_020_5100, w_020_5101, w_020_5102, w_020_5103, w_020_5104, w_020_5106, w_020_5110, w_020_5111, w_020_5112, w_020_5114, w_020_5115, w_020_5116, w_020_5117, w_020_5118, w_020_5119, w_020_5120, w_020_5121, w_020_5122, w_020_5123, w_020_5124, w_020_5125, w_020_5126, w_020_5127, w_020_5129, w_020_5130, w_020_5131, w_020_5132, w_020_5135, w_020_5136, w_020_5138, w_020_5140, w_020_5143, w_020_5144, w_020_5147, w_020_5149, w_020_5150, w_020_5153, w_020_5154, w_020_5155, w_020_5156, w_020_5158, w_020_5161, w_020_5163, w_020_5164, w_020_5166, w_020_5167, w_020_5172, w_020_5173, w_020_5174, w_020_5176, w_020_5177, w_020_5178, w_020_5179, w_020_5181, w_020_5182, w_020_5184, w_020_5185, w_020_5186, w_020_5187, w_020_5190, w_020_5191, w_020_5194, w_020_5195, w_020_5196, w_020_5197, w_020_5198, w_020_5199, w_020_5201, w_020_5202, w_020_5205, w_020_5207, w_020_5210, w_020_5212, w_020_5213, w_020_5217, w_020_5218, w_020_5220, w_020_5221, w_020_5222, w_020_5223, w_020_5224, w_020_5225, w_020_5226, w_020_5230, w_020_5231, w_020_5232, w_020_5233, w_020_5236, w_020_5238, w_020_5240, w_020_5241, w_020_5242, w_020_5243, w_020_5244, w_020_5247, w_020_5248, w_020_5249, w_020_5250, w_020_5253, w_020_5254, w_020_5256, w_020_5259, w_020_5260, w_020_5261, w_020_5263, w_020_5264, w_020_5266, w_020_5267, w_020_5268, w_020_5269, w_020_5273, w_020_5274, w_020_5275, w_020_5276, w_020_5277, w_020_5278, w_020_5280, w_020_5283, w_020_5284, w_020_5286, w_020_5288, w_020_5296, w_020_5297, w_020_5298, w_020_5300, w_020_5301, w_020_5304, w_020_5305, w_020_5306, w_020_5309, w_020_5310, w_020_5313, w_020_5316, w_020_5317, w_020_5318, w_020_5321, w_020_5322, w_020_5323, w_020_5325, w_020_5330, w_020_5331, w_020_5332, w_020_5334, w_020_5335, w_020_5336, w_020_5338, w_020_5341, w_020_5343, w_020_5344, w_020_5345, w_020_5347, w_020_5348, w_020_5349, w_020_5350, w_020_5351, w_020_5353, w_020_5354, w_020_5356, w_020_5357, w_020_5358, w_020_5359, w_020_5361, w_020_5362, w_020_5363, w_020_5364, w_020_5365, w_020_5367, w_020_5370, w_020_5371, w_020_5373, w_020_5376, w_020_5379, w_020_5381, w_020_5382, w_020_5387, w_020_5389, w_020_5390, w_020_5391, w_020_5392, w_020_5394, w_020_5396, w_020_5397, w_020_5398, w_020_5400, w_020_5402, w_020_5406, w_020_5407, w_020_5409, w_020_5410, w_020_5411, w_020_5412, w_020_5415, w_020_5418, w_020_5420, w_020_5421, w_020_5425, w_020_5426, w_020_5429, w_020_5431, w_020_5432, w_020_5435, w_020_5436, w_020_5437, w_020_5438, w_020_5440, w_020_5442, w_020_5445, w_020_5446, w_020_5447, w_020_5450, w_020_5451, w_020_5452, w_020_5457, w_020_5458, w_020_5459, w_020_5461, w_020_5462, w_020_5463, w_020_5464, w_020_5465, w_020_5467, w_020_5471, w_020_5474, w_020_5476, w_020_5477, w_020_5478, w_020_5480, w_020_5481, w_020_5482, w_020_5483, w_020_5485, w_020_5486, w_020_5487, w_020_5488, w_020_5489, w_020_5490, w_020_5491, w_020_5492, w_020_5494, w_020_5496, w_020_5497, w_020_5500, w_020_5501, w_020_5502, w_020_5503, w_020_5505, w_020_5506, w_020_5508, w_020_5511, w_020_5512, w_020_5514, w_020_5516, w_020_5517, w_020_5519, w_020_5521, w_020_5526, w_020_5529, w_020_5530, w_020_5531, w_020_5532, w_020_5535, w_020_5537, w_020_5540, w_020_5544, w_020_5546, w_020_5548, w_020_5549, w_020_5551, w_020_5552, w_020_5554, w_020_5556, w_020_5557, w_020_5559, w_020_5562, w_020_5563, w_020_5568, w_020_5569, w_020_5570, w_020_5571, w_020_5572, w_020_5573, w_020_5575, w_020_5576, w_020_5578, w_020_5582, w_020_5584, w_020_5585, w_020_5586, w_020_5587, w_020_5588, w_020_5589, w_020_5590, w_020_5591, w_020_5593, w_020_5594, w_020_5595, w_020_5598, w_020_5599, w_020_5603, w_020_5604, w_020_5606, w_020_5607, w_020_5608, w_020_5609, w_020_5611, w_020_5613, w_020_5614, w_020_5615, w_020_5617, w_020_5618, w_020_5620, w_020_5623, w_020_5628, w_020_5633, w_020_5635, w_020_5636, w_020_5637, w_020_5638, w_020_5641, w_020_5644, w_020_5645, w_020_5647, w_020_5648, w_020_5650, w_020_5652, w_020_5654, w_020_5656, w_020_5660, w_020_5661, w_020_5662, w_020_5664, w_020_5665, w_020_5666, w_020_5668, w_020_5670, w_020_5671, w_020_5672, w_020_5673, w_020_5674, w_020_5675, w_020_5677, w_020_5681, w_020_5686, w_020_5687, w_020_5688, w_020_5691, w_020_5692, w_020_5693, w_020_5696, w_020_5697, w_020_5699, w_020_5700, w_020_5701, w_020_5702, w_020_5703, w_020_5704, w_020_5705, w_020_5706, w_020_5707, w_020_5708, w_020_5710, w_020_5711, w_020_5713, w_020_5714, w_020_5715, w_020_5716, w_020_5718, w_020_5720, w_020_5724, w_020_5725, w_020_5726, w_020_5727, w_020_5728, w_020_5729, w_020_5732, w_020_5735, w_020_5738, w_020_5739, w_020_5741, w_020_5742, w_020_5744, w_020_5745, w_020_5746, w_020_5751, w_020_5753, w_020_5755, w_020_5757, w_020_5758, w_020_5759, w_020_5760, w_020_5761, w_020_5765, w_020_5767, w_020_5771, w_020_5773, w_020_5774, w_020_5775, w_020_5776, w_020_5778, w_020_5779, w_020_5782, w_020_5784, w_020_5785, w_020_5786, w_020_5787, w_020_5788, w_020_5790, w_020_5792, w_020_5793, w_020_5794, w_020_5795, w_020_5797, w_020_5798, w_020_5801, w_020_5802, w_020_5803, w_020_5804, w_020_5807, w_020_5810, w_020_5811, w_020_5813, w_020_5814, w_020_5815, w_020_5816, w_020_5817, w_020_5818, w_020_5819, w_020_5822, w_020_5823, w_020_5824, w_020_5827, w_020_5828, w_020_5830, w_020_5831, w_020_5832, w_020_5833, w_020_5835, w_020_5837, w_020_5839, w_020_5840, w_020_5853, w_020_5855, w_020_5856, w_020_5862, w_020_5863, w_020_5864, w_020_5866, w_020_5867, w_020_5868, w_020_5869, w_020_5870, w_020_5871, w_020_5873, w_020_5874, w_020_5877, w_020_5881, w_020_5882, w_020_5883, w_020_5884, w_020_5885, w_020_5886, w_020_5889, w_020_5890, w_020_5891, w_020_5892, w_020_5894, w_020_5896, w_020_5898, w_020_5899, w_020_5901, w_020_5902, w_020_5903, w_020_5905, w_020_5906, w_020_5907, w_020_5908, w_020_5910, w_020_5911, w_020_5912, w_020_5914, w_020_5915, w_020_5916, w_020_5918, w_020_5921, w_020_5922, w_020_5923, w_020_5924, w_020_5925, w_020_5926, w_020_5927, w_020_5929, w_020_5930, w_020_5933, w_020_5934, w_020_5935, w_020_5936, w_020_5938, w_020_5939, w_020_5940, w_020_5941, w_020_5942, w_020_5943, w_020_5945, w_020_5946, w_020_5948, w_020_5949, w_020_5952, w_020_5953, w_020_5955, w_020_5956, w_020_5957, w_020_5958, w_020_5959, w_020_5961, w_020_5962, w_020_5963, w_020_5964, w_020_5965, w_020_5966, w_020_5967, w_020_5968, w_020_5969, w_020_5970, w_020_5971, w_020_5972, w_020_5973, w_020_5976, w_020_5977, w_020_5978, w_020_5980, w_020_5981, w_020_5982, w_020_5983, w_020_5986, w_020_5987, w_020_5988, w_020_5989, w_020_5991, w_020_5992, w_020_5993, w_020_5994, w_020_5996, w_020_5997, w_020_5998, w_020_6000, w_020_6001, w_020_6002, w_020_6003, w_020_6007, w_020_6008, w_020_6009, w_020_6010, w_020_6011, w_020_6012, w_020_6014, w_020_6017, w_020_6018, w_020_6020, w_020_6022, w_020_6023, w_020_6024, w_020_6027, w_020_6029, w_020_6030, w_020_6031, w_020_6032, w_020_6033, w_020_6036, w_020_6038, w_020_6039, w_020_6041, w_020_6042, w_020_6043, w_020_6044, w_020_6045, w_020_6046, w_020_6047, w_020_6048, w_020_6050, w_020_6051, w_020_6055, w_020_6057, w_020_6058, w_020_6060, w_020_6061, w_020_6063, w_020_6064, w_020_6065, w_020_6066, w_020_6067, w_020_6068, w_020_6069, w_020_6070, w_020_6071, w_020_6072, w_020_6073, w_020_6074, w_020_6075, w_020_6076, w_020_6077, w_020_6078, w_020_6079, w_020_6080, w_020_6083, w_020_6085, w_020_6087, w_020_6088, w_020_6089, w_020_6092, w_020_6093, w_020_6094, w_020_6095, w_020_6096, w_020_6098, w_020_6099, w_020_6101, w_020_6103, w_020_6104, w_020_6108, w_020_6109, w_020_6110, w_020_6112, w_020_6114, w_020_6116, w_020_6117, w_020_6119, w_020_6120, w_020_6121, w_020_6122, w_020_6123, w_020_6125, w_020_6126, w_020_6128, w_020_6129, w_020_6132, w_020_6135, w_020_6136, w_020_6137, w_020_6138, w_020_6139, w_020_6140, w_020_6141, w_020_6142, w_020_6143, w_020_6144, w_020_6145, w_020_6146, w_020_6147, w_020_6148, w_020_6150, w_020_6152, w_020_6153, w_020_6154, w_020_6155, w_020_6163, w_020_6164, w_020_6166, w_020_6167, w_020_6170, w_020_6171, w_020_6172, w_020_6175, w_020_6177, w_020_6178, w_020_6179, w_020_6182, w_020_6184, w_020_6186, w_020_6187, w_020_6188, w_020_6189, w_020_6190, w_020_6191, w_020_6192, w_020_6193, w_020_6194, w_020_6195, w_020_6196, w_020_6197, w_020_6198, w_020_6199, w_020_6203, w_020_6204, w_020_6205, w_020_6206, w_020_6207, w_020_6208, w_020_6209, w_020_6211, w_020_6212, w_020_6213, w_020_6214, w_020_6215, w_020_6216, w_020_6219, w_020_6220, w_020_6224, w_020_6225, w_020_6228, w_020_6229, w_020_6230, w_020_6231, w_020_6232, w_020_6234, w_020_6236, w_020_6237, w_020_6238, w_020_6239, w_020_6241, w_020_6245, w_020_6246, w_020_6249, w_020_6251, w_020_6252, w_020_6257, w_020_6260, w_020_6261, w_020_6262, w_020_6263, w_020_6264, w_020_6266, w_020_6267, w_020_6269, w_020_6270, w_020_6271, w_020_6272, w_020_6274, w_020_6276, w_020_6277, w_020_6280, w_020_6281, w_020_6282, w_020_6283, w_020_6284, w_020_6286, w_020_6289, w_020_6290, w_020_6292, w_020_6293, w_020_6294, w_020_6295, w_020_6296, w_020_6298, w_020_6299, w_020_6300, w_020_6304, w_020_6308, w_020_6310, w_020_6311, w_020_6313, w_020_6316, w_020_6317, w_020_6318, w_020_6319, w_020_6320, w_020_6322, w_020_6325, w_020_6327, w_020_6328, w_020_6331, w_020_6334, w_020_6335, w_020_6336, w_020_6337, w_020_6338, w_020_6339, w_020_6343, w_020_6344, w_020_6345, w_020_6346, w_020_6347, w_020_6348, w_020_6349, w_020_6351, w_020_6354, w_020_6356, w_020_6357, w_020_6359, w_020_6361, w_020_6362, w_020_6363, w_020_6366, w_020_6367, w_020_6368, w_020_6369, w_020_6370, w_020_6372, w_020_6373, w_020_6374, w_020_6375, w_020_6377, w_020_6380, w_020_6381, w_020_6385, w_020_6388, w_020_6389, w_020_6390, w_020_6391, w_020_6392, w_020_6393, w_020_6394, w_020_6395, w_020_6396, w_020_6397, w_020_6399, w_020_6400, w_020_6402, w_020_6403, w_020_6404, w_020_6405, w_020_6406, w_020_6407, w_020_6412, w_020_6416, w_020_6417, w_020_6420, w_020_6422, w_020_6424, w_020_6426, w_020_6427, w_020_6429, w_020_6430, w_020_6431, w_020_6434, w_020_6435, w_020_6437, w_020_6438, w_020_6439, w_020_6440, w_020_6441, w_020_6442, w_020_6444, w_020_6447, w_020_6448, w_020_6449, w_020_6450, w_020_6451, w_020_6452, w_020_6453, w_020_6456, w_020_6457, w_020_6458, w_020_6461, w_020_6462, w_020_6466, w_020_6470, w_020_6472, w_020_6473, w_020_6474, w_020_6476, w_020_6478, w_020_6479, w_020_6481, w_020_6484, w_020_6486, w_020_6488, w_020_6489, w_020_6490, w_020_6491, w_020_6492, w_020_6493, w_020_6494, w_020_6496, w_020_6497, w_020_6498, w_020_6499, w_020_6500, w_020_6502, w_020_6506, w_020_6507, w_020_6508, w_020_6509, w_020_6510, w_020_6512, w_020_6513, w_020_6515, w_020_6516, w_020_6518, w_020_6520, w_020_6521, w_020_6523, w_020_6525, w_020_6527, w_020_6529, w_020_6530, w_020_6531, w_020_6532, w_020_6533, w_020_6534, w_020_6536, w_020_6537, w_020_6538, w_020_6539, w_020_6540, w_020_6542, w_020_6543, w_020_6544, w_020_6545, w_020_6547, w_020_6548, w_020_6550, w_020_6551, w_020_6552, w_020_6553, w_020_6555, w_020_6560, w_020_6561, w_020_6564, w_020_6566, w_020_6570, w_020_6573, w_020_6576, w_020_6577, w_020_6578, w_020_6581, w_020_6584, w_020_6585, w_020_6586, w_020_6587, w_020_6589, w_020_6591, w_020_6592, w_020_6595, w_020_6596, w_020_6597, w_020_6598, w_020_6602, w_020_6603, w_020_6604, w_020_6605, w_020_6607, w_020_6608, w_020_6612, w_020_6615, w_020_6617, w_020_6620, w_020_6621, w_020_6622, w_020_6623, w_020_6627, w_020_6629, w_020_6631, w_020_6633, w_020_6635, w_020_6640, w_020_6643, w_020_6645, w_020_6646, w_020_6647, w_020_6648, w_020_6649, w_020_6650, w_020_6651, w_020_6652, w_020_6653, w_020_6654, w_020_6658, w_020_6661, w_020_6665, w_020_6666, w_020_6667, w_020_6668, w_020_6670, w_020_6671, w_020_6672, w_020_6673, w_020_6674, w_020_6675, w_020_6676, w_020_6677, w_020_6679, w_020_6680, w_020_6681, w_020_6682, w_020_6683, w_020_6684, w_020_6685, w_020_6686, w_020_6690, w_020_6691, w_020_6692, w_020_6693, w_020_6695, w_020_6696, w_020_6697, w_020_6698, w_020_6702, w_020_6703, w_020_6704, w_020_6705, w_020_6706, w_020_6707, w_020_6708, w_020_6710, w_020_6711, w_020_6712, w_020_6713, w_020_6714, w_020_6718, w_020_6720, w_020_6725, w_020_6726, w_020_6731, w_020_6732, w_020_6734, w_020_6735, w_020_6737, w_020_6738, w_020_6739, w_020_6740, w_020_6743, w_020_6745, w_020_6746, w_020_6747, w_020_6749, w_020_6751, w_020_6752, w_020_6754, w_020_6755, w_020_6756, w_020_6757, w_020_6758, w_020_6763, w_020_6764, w_020_6766, w_020_6767, w_020_6768, w_020_6769, w_020_6770, w_020_6771, w_020_6772, w_020_6775, w_020_6777, w_020_6779, w_020_6780, w_020_6781, w_020_6783, w_020_6785, w_020_6786, w_020_6787, w_020_6788, w_020_6791, w_020_6793, w_020_6794, w_020_6795, w_020_6797, w_020_6800, w_020_6803, w_020_6804, w_020_6805, w_020_6807, w_020_6809, w_020_6815, w_020_6816, w_020_6817, w_020_6819, w_020_6821, w_020_6822, w_020_6823, w_020_6824, w_020_6825, w_020_6826, w_020_6827, w_020_6830, w_020_6831, w_020_6833, w_020_6834, w_020_6835, w_020_6836, w_020_6838, w_020_6839, w_020_6842, w_020_6843, w_020_6844, w_020_6847, w_020_6848, w_020_6849, w_020_6850, w_020_6854, w_020_6855, w_020_6856, w_020_6857, w_020_6858, w_020_6859, w_020_6860, w_020_6861, w_020_6863, w_020_6864, w_020_6867, w_020_6868, w_020_6869, w_020_6870, w_020_6871, w_020_6872, w_020_6873, w_020_6874, w_020_6877, w_020_6881, w_020_6882, w_020_6883, w_020_6884, w_020_6886, w_020_6887, w_020_6888, w_020_6894, w_020_6895, w_020_6898, w_020_6901, w_020_6903, w_020_6904, w_020_6906, w_020_6907, w_020_6908, w_020_6909, w_020_6910, w_020_6911, w_020_6913, w_020_6914, w_020_6917, w_020_6918, w_020_6919, w_020_6921, w_020_6922, w_020_6924, w_020_6925, w_020_6926, w_020_6927, w_020_6928, w_020_6930, w_020_6931, w_020_6934, w_020_6935, w_020_6938, w_020_6939, w_020_6943, w_020_6945, w_020_6948, w_020_6949, w_020_6950, w_020_6951, w_020_6952, w_020_6953, w_020_6954, w_020_6956, w_020_6959, w_020_6964, w_020_6966, w_020_6967, w_020_6968, w_020_6969, w_020_6970, w_020_6971, w_020_6976, w_020_6977, w_020_6979, w_020_6981, w_020_6982, w_020_6984, w_020_6986, w_020_6987, w_020_6990, w_020_6993, w_020_6994, w_020_6995, w_020_6996, w_020_6999, w_020_7000, w_020_7001, w_020_7002, w_020_7005, w_020_7007, w_020_7008, w_020_7009, w_020_7010, w_020_7011, w_020_7013, w_020_7014, w_020_7015, w_020_7016, w_020_7019, w_020_7021, w_020_7022, w_020_7023, w_020_7025, w_020_7026, w_020_7027, w_020_7028, w_020_7030, w_020_7032, w_020_7033, w_020_7035, w_020_7036, w_020_7037, w_020_7038, w_020_7039, w_020_7040, w_020_7042, w_020_7043, w_020_7045, w_020_7046, w_020_7047, w_020_7048, w_020_7049, w_020_7051, w_020_7055, w_020_7058, w_020_7059, w_020_7060, w_020_7061, w_020_7062, w_020_7065, w_020_7066, w_020_7069, w_020_7070, w_020_7072, w_020_7073, w_020_7074, w_020_7075, w_020_7076, w_020_7078, w_020_7079, w_020_7080, w_020_7081, w_020_7084, w_020_7085, w_020_7086, w_020_7087, w_020_7089, w_020_7090, w_020_7091, w_020_7092, w_020_7093, w_020_7094, w_020_7096, w_020_7098, w_020_7099, w_020_7100, w_020_7101, w_020_7102, w_020_7106, w_020_7108, w_020_7109, w_020_7110, w_020_7111, w_020_7112, w_020_7113, w_020_7117, w_020_7118, w_020_7119, w_020_7123, w_020_7124, w_020_7126, w_020_7127, w_020_7128, w_020_7129, w_020_7130, w_020_7135, w_020_7136, w_020_7137, w_020_7142, w_020_7143, w_020_7144, w_020_7145, w_020_7146, w_020_7147, w_020_7149, w_020_7150, w_020_7151, w_020_7152, w_020_7153, w_020_7154, w_020_7155, w_020_7157, w_020_7158, w_020_7160, w_020_7163, w_020_7164, w_020_7165, w_020_7166, w_020_7168, w_020_7171, w_020_7174, w_020_7176, w_020_7177, w_020_7179, w_020_7180, w_020_7181, w_020_7182, w_020_7184, w_020_7185, w_020_7186, w_020_7189, w_020_7190, w_020_7191, w_020_7192, w_020_7193, w_020_7194, w_020_7197, w_020_7198, w_020_7199, w_020_7200, w_020_7201, w_020_7205, w_020_7207, w_020_7208, w_020_7209, w_020_7210, w_020_7211, w_020_7212, w_020_7213, w_020_7214, w_020_7215, w_020_7216, w_020_7217, w_020_7218, w_020_7223, w_020_7225, w_020_7231, w_020_7237, w_020_7238, w_020_7239, w_020_7241, w_020_7243, w_020_7248, w_020_7249, w_020_7251, w_020_7253, w_020_7256, w_020_7258, w_020_7260, w_020_7261, w_020_7262, w_020_7263, w_020_7264, w_020_7267, w_020_7268, w_020_7269, w_020_7271, w_020_7272, w_020_7273, w_020_7275, w_020_7278, w_020_7279, w_020_7280, w_020_7282, w_020_7285, w_020_7287, w_020_7288, w_020_7289, w_020_7290, w_020_7293, w_020_7295, w_020_7296, w_020_7297, w_020_7298, w_020_7300, w_020_7301, w_020_7302, w_020_7303, w_020_7307, w_020_7309, w_020_7310, w_020_7311, w_020_7312, w_020_7314, w_020_7315, w_020_7316, w_020_7317, w_020_7321, w_020_7331, w_020_7332, w_020_7335, w_020_7336, w_020_7337, w_020_7338, w_020_7340, w_020_7342, w_020_7345, w_020_7346, w_020_7348, w_020_7349, w_020_7351, w_020_7352, w_020_7353, w_020_7356, w_020_7357, w_020_7358, w_020_7359, w_020_7360, w_020_7361, w_020_7362, w_020_7364, w_020_7365, w_020_7369, w_020_7370, w_020_7371, w_020_7372, w_020_7376, w_020_7377, w_020_7379, w_020_7382, w_020_7386, w_020_7389, w_020_7390, w_020_7391, w_020_7392, w_020_7393, w_020_7395, w_020_7399, w_020_7401, w_020_7403, w_020_7406, w_020_7407, w_020_7408, w_020_7409, w_020_7410, w_020_7415, w_020_7416, w_020_7417, w_020_7420, w_020_7421, w_020_7422, w_020_7423, w_020_7424, w_020_7426, w_020_7428, w_020_7430, w_020_7431, w_020_7433, w_020_7436, w_020_7438, w_020_7439, w_020_7441, w_020_7443, w_020_7445, w_020_7448, w_020_7449, w_020_7451, w_020_7453, w_020_7454, w_020_7456, w_020_7459, w_020_7461, w_020_7462, w_020_7463, w_020_7464, w_020_7465, w_020_7466, w_020_7467, w_020_7468, w_020_7469, w_020_7470, w_020_7471, w_020_7472, w_020_7473, w_020_7474, w_020_7479, w_020_7480, w_020_7481, w_020_7484, w_020_7487, w_020_7490, w_020_7494, w_020_7495, w_020_7496, w_020_7497, w_020_7498, w_020_7500, w_020_7501, w_020_7503, w_020_7504, w_020_7505, w_020_7507, w_020_7508, w_020_7509, w_020_7513, w_020_7515, w_020_7516, w_020_7517, w_020_7518, w_020_7519, w_020_7520, w_020_7524, w_020_7525, w_020_7527, w_020_7528, w_020_7529, w_020_7530, w_020_7531, w_020_7532, w_020_7535, w_020_7537, w_020_7538, w_020_7539, w_020_7540, w_020_7543, w_020_7544, w_020_7546, w_020_7547, w_020_7548, w_020_7549, w_020_7550, w_020_7551, w_020_7552, w_020_7554, w_020_7555, w_020_7557, w_020_7558, w_020_7559, w_020_7564, w_020_7565, w_020_7568, w_020_7569, w_020_7571, w_020_7574, w_020_7577, w_020_7578, w_020_7579, w_020_7580, w_020_7581, w_020_7586, w_020_7588, w_020_7589, w_020_7591, w_020_7592, w_020_7593, w_020_7594, w_020_7595, w_020_7596, w_020_7597, w_020_7598, w_020_7599, w_020_7600, w_020_7604, w_020_7605, w_020_7606, w_020_7609, w_020_7610, w_020_7611, w_020_7612, w_020_7613, w_020_7614, w_020_7615, w_020_7616, w_020_7617, w_020_7618, w_020_7620, w_020_7623, w_020_7624, w_020_7625, w_020_7626, w_020_7628, w_020_7629, w_020_7633, w_020_7636, w_020_7638, w_020_7641, w_020_7642, w_020_7643, w_020_7646, w_020_7647, w_020_7648, w_020_7649, w_020_7650, w_020_7651, w_020_7652, w_020_7655, w_020_7657, w_020_7658, w_020_7659, w_020_7663, w_020_7664, w_020_7665, w_020_7666, w_020_7669, w_020_7670, w_020_7672, w_020_7674, w_020_7676, w_020_7678, w_020_7680, w_020_7685, w_020_7687, w_020_7688, w_020_7689, w_020_7690, w_020_7692, w_020_7694, w_020_7696, w_020_7697, w_020_7698, w_020_7700, w_020_7704, w_020_7710, w_020_7712, w_020_7714, w_020_7715, w_020_7716, w_020_7718, w_020_7719, w_020_7720, w_020_7721, w_020_7723, w_020_7724, w_020_7725, w_020_7727, w_020_7728, w_020_7729, w_020_7730, w_020_7734, w_020_7736, w_020_7739, w_020_7740, w_020_7742, w_020_7743, w_020_7745, w_020_7746, w_020_7749, w_020_7752, w_020_7753, w_020_7754, w_020_7756, w_020_7757, w_020_7759, w_020_7760, w_020_7761, w_020_7762, w_020_7763;
  wire w_021_000, w_021_001, w_021_002, w_021_003, w_021_004, w_021_005, w_021_006, w_021_007, w_021_008, w_021_009, w_021_010, w_021_011, w_021_012, w_021_013, w_021_014, w_021_015, w_021_016, w_021_017, w_021_018, w_021_019, w_021_020, w_021_021, w_021_022, w_021_023, w_021_024, w_021_025, w_021_026, w_021_027, w_021_028, w_021_029, w_021_030, w_021_031, w_021_032, w_021_033, w_021_034, w_021_035, w_021_036, w_021_037, w_021_038, w_021_039, w_021_040, w_021_041, w_021_042, w_021_043, w_021_044, w_021_045, w_021_046, w_021_047, w_021_048, w_021_049, w_021_050, w_021_051, w_021_052, w_021_053, w_021_054, w_021_055, w_021_056, w_021_057, w_021_058, w_021_059, w_021_060, w_021_061, w_021_062, w_021_063, w_021_064, w_021_065, w_021_066, w_021_067, w_021_068, w_021_069, w_021_070, w_021_071, w_021_072, w_021_073, w_021_074, w_021_075, w_021_076, w_021_077, w_021_078, w_021_079, w_021_080, w_021_081, w_021_082, w_021_083, w_021_084, w_021_085, w_021_086, w_021_087, w_021_088, w_021_089, w_021_090, w_021_091, w_021_092, w_021_093, w_021_094, w_021_095, w_021_096, w_021_097, w_021_098, w_021_099, w_021_100, w_021_101, w_021_102, w_021_103, w_021_104, w_021_105, w_021_106, w_021_107, w_021_108, w_021_109, w_021_110, w_021_111, w_021_112, w_021_113, w_021_114, w_021_115, w_021_116, w_021_117, w_021_118, w_021_119, w_021_120, w_021_121, w_021_122, w_021_123, w_021_124, w_021_125, w_021_126, w_021_127, w_021_128, w_021_129, w_021_130, w_021_131, w_021_132, w_021_133, w_021_134, w_021_135, w_021_136, w_021_137, w_021_138, w_021_139, w_021_140, w_021_141, w_021_142, w_021_143, w_021_144, w_021_145, w_021_146, w_021_147, w_021_148, w_021_149, w_021_150, w_021_151, w_021_152, w_021_153, w_021_154, w_021_155, w_021_156, w_021_157, w_021_158, w_021_159, w_021_160, w_021_161, w_021_162, w_021_163, w_021_164, w_021_165, w_021_166, w_021_167, w_021_168, w_021_169, w_021_170, w_021_171, w_021_172, w_021_173, w_021_174, w_021_175, w_021_176, w_021_177, w_021_178, w_021_179, w_021_180, w_021_181, w_021_182, w_021_183, w_021_184, w_021_185, w_021_186, w_021_187, w_021_188, w_021_189, w_021_190, w_021_191, w_021_192, w_021_193, w_021_194, w_021_195, w_021_196, w_021_197, w_021_198, w_021_199, w_021_200, w_021_201, w_021_202, w_021_203, w_021_204, w_021_205, w_021_206, w_021_207, w_021_208, w_021_209, w_021_210, w_021_211, w_021_212, w_021_213, w_021_214, w_021_215, w_021_216, w_021_217, w_021_218, w_021_219, w_021_220, w_021_221, w_021_222, w_021_223, w_021_224, w_021_225, w_021_226, w_021_227, w_021_228, w_021_229, w_021_230, w_021_231, w_021_232, w_021_233, w_021_234, w_021_235, w_021_236, w_021_237, w_021_238, w_021_239, w_021_240, w_021_241, w_021_242, w_021_243, w_021_244, w_021_245, w_021_246, w_021_247, w_021_248, w_021_249, w_021_250, w_021_251, w_021_252, w_021_253, w_021_254, w_021_255, w_021_256, w_021_257, w_021_258, w_021_259, w_021_260, w_021_261, w_021_262, w_021_263, w_021_264, w_021_265, w_021_266, w_021_267, w_021_268, w_021_269, w_021_270, w_021_271, w_021_272, w_021_273, w_021_274, w_021_275, w_021_276, w_021_277, w_021_278, w_021_279, w_021_280, w_021_281, w_021_282, w_021_283, w_021_284, w_021_285, w_021_286, w_021_287, w_021_288, w_021_289, w_021_290, w_021_291, w_021_292, w_021_293, w_021_294, w_021_295, w_021_296, w_021_297, w_021_298, w_021_299, w_021_300, w_021_301, w_021_302, w_021_303, w_021_304, w_021_305, w_021_306, w_021_307, w_021_308, w_021_309, w_021_310, w_021_311, w_021_312, w_021_313, w_021_314, w_021_315, w_021_316, w_021_317, w_021_318, w_021_319, w_021_320, w_021_321, w_021_322, w_021_323, w_021_324, w_021_325, w_021_326, w_021_327, w_021_328, w_021_329, w_021_330, w_021_331, w_021_332, w_021_333, w_021_334, w_021_335, w_021_336, w_021_337, w_021_338, w_021_339, w_021_340, w_021_341, w_021_342, w_021_343, w_021_344, w_021_345, w_021_346, w_021_347, w_021_348, w_021_349, w_021_350, w_021_351, w_021_352, w_021_353, w_021_354, w_021_355, w_021_356, w_021_357, w_021_358, w_021_359, w_021_360, w_021_361, w_021_362, w_021_363, w_021_364, w_021_365, w_021_366, w_021_367, w_021_368, w_021_369, w_021_370, w_021_371, w_021_372, w_021_373, w_021_374, w_021_375, w_021_376, w_021_377, w_021_378, w_021_379, w_021_380, w_021_381, w_021_382, w_021_383, w_021_384, w_021_385, w_021_386, w_021_387, w_021_388, w_021_389, w_021_390, w_021_391, w_021_392, w_021_393, w_021_394, w_021_395, w_021_396, w_021_397, w_021_398, w_021_399, w_021_400, w_021_401, w_021_402, w_021_403, w_021_404, w_021_405, w_021_406, w_021_407, w_021_408, w_021_409, w_021_410, w_021_411, w_021_412, w_021_413, w_021_414, w_021_415, w_021_416, w_021_417, w_021_418, w_021_419, w_021_420, w_021_421, w_021_422, w_021_423, w_021_424, w_021_425, w_021_426, w_021_427, w_021_428, w_021_429, w_021_430, w_021_431, w_021_432, w_021_433, w_021_434, w_021_435, w_021_436, w_021_437, w_021_438, w_021_439, w_021_440, w_021_441, w_021_442, w_021_443, w_021_444, w_021_445, w_021_446, w_021_447, w_021_448, w_021_449, w_021_450, w_021_451, w_021_452, w_021_453, w_021_454, w_021_455, w_021_456, w_021_457, w_021_458, w_021_459, w_021_460, w_021_461, w_021_462, w_021_463, w_021_464, w_021_465, w_021_466, w_021_467, w_021_468, w_021_469, w_021_470, w_021_471, w_021_472, w_021_473, w_021_474, w_021_475, w_021_476, w_021_477, w_021_478, w_021_479, w_021_480, w_021_481, w_021_482, w_021_483, w_021_484, w_021_485, w_021_486, w_021_487, w_021_488, w_021_489, w_021_490, w_021_491, w_021_492, w_021_493, w_021_494, w_021_495, w_021_496, w_021_497, w_021_498, w_021_499, w_021_500, w_021_501, w_021_502, w_021_503, w_021_504, w_021_505, w_021_506, w_021_507, w_021_508, w_021_509, w_021_510, w_021_511, w_021_512, w_021_513, w_021_514, w_021_515, w_021_516, w_021_517, w_021_518, w_021_519, w_021_520, w_021_521, w_021_522, w_021_523, w_021_524, w_021_525, w_021_526, w_021_527, w_021_528, w_021_529, w_021_530, w_021_531, w_021_532, w_021_533, w_021_534, w_021_535, w_021_536, w_021_537, w_021_538, w_021_539, w_021_540, w_021_541, w_021_542, w_021_543, w_021_544, w_021_545, w_021_546, w_021_547, w_021_548, w_021_549, w_021_550, w_021_551, w_021_552, w_021_553, w_021_554, w_021_555, w_021_556, w_021_557, w_021_558, w_021_559, w_021_560, w_021_561, w_021_562, w_021_563, w_021_564, w_021_565, w_021_566, w_021_567, w_021_568, w_021_569, w_021_570, w_021_571, w_021_572, w_021_573, w_021_574, w_021_575, w_021_576, w_021_577, w_021_578, w_021_579, w_021_580, w_021_581, w_021_582, w_021_583, w_021_584, w_021_585, w_021_586, w_021_587, w_021_588, w_021_589, w_021_590, w_021_591, w_021_592, w_021_593, w_021_594, w_021_595, w_021_596, w_021_597, w_021_598, w_021_599, w_021_600, w_021_601, w_021_602, w_021_603, w_021_604, w_021_605, w_021_606, w_021_607, w_021_608, w_021_609, w_021_610, w_021_611, w_021_612, w_021_613, w_021_614, w_021_615, w_021_616, w_021_617, w_021_618, w_021_619, w_021_620, w_021_621, w_021_622, w_021_623, w_021_624, w_021_625, w_021_626, w_021_627, w_021_628, w_021_629, w_021_630, w_021_631, w_021_632, w_021_633, w_021_634, w_021_635, w_021_636, w_021_637, w_021_638, w_021_639, w_021_640, w_021_641, w_021_642, w_021_643, w_021_644, w_021_645, w_021_646, w_021_647, w_021_648, w_021_649, w_021_650, w_021_651, w_021_652, w_021_653, w_021_654, w_021_655, w_021_656, w_021_657, w_021_658, w_021_659, w_021_660, w_021_661, w_021_662, w_021_663, w_021_664, w_021_665, w_021_666, w_021_667, w_021_668, w_021_669, w_021_670, w_021_671, w_021_672, w_021_673, w_021_674, w_021_675, w_021_676, w_021_677, w_021_678, w_021_679, w_021_680, w_021_681, w_021_682, w_021_683, w_021_684, w_021_685, w_021_686, w_021_687, w_021_688, w_021_689, w_021_690, w_021_691, w_021_692, w_021_693, w_021_694, w_021_695, w_021_696, w_021_697, w_021_698, w_021_699, w_021_700, w_021_701, w_021_702, w_021_703, w_021_704, w_021_705, w_021_706, w_021_707, w_021_708, w_021_709, w_021_710, w_021_711, w_021_712, w_021_713, w_021_714, w_021_715, w_021_716, w_021_717, w_021_718, w_021_719, w_021_720, w_021_721, w_021_722, w_021_723, w_021_724, w_021_725, w_021_726, w_021_727, w_021_728, w_021_729, w_021_730, w_021_731, w_021_732, w_021_733, w_021_734, w_021_735, w_021_736, w_021_737, w_021_738, w_021_739, w_021_740, w_021_741, w_021_742, w_021_743, w_021_744, w_021_745, w_021_746, w_021_747, w_021_748, w_021_749, w_021_750, w_021_751, w_021_752, w_021_753, w_021_754, w_021_755, w_021_756, w_021_757, w_021_758, w_021_759, w_021_760, w_021_761, w_021_762, w_021_763, w_021_764, w_021_765, w_021_766, w_021_767, w_021_768, w_021_769, w_021_770, w_021_771, w_021_772, w_021_773, w_021_774, w_021_775, w_021_776, w_021_777, w_021_778, w_021_779, w_021_780, w_021_781, w_021_782, w_021_783, w_021_784, w_021_785, w_021_786, w_021_787, w_021_788, w_021_789, w_021_790, w_021_791, w_021_792, w_021_793, w_021_794, w_021_795, w_021_796, w_021_797, w_021_798, w_021_799, w_021_800, w_021_801, w_021_802, w_021_803, w_021_804, w_021_805, w_021_806, w_021_807, w_021_808, w_021_809, w_021_810, w_021_811, w_021_812, w_021_813, w_021_814, w_021_815, w_021_816, w_021_817, w_021_818, w_021_819, w_021_820, w_021_821, w_021_822, w_021_823, w_021_824, w_021_825, w_021_826, w_021_827, w_021_828, w_021_829, w_021_830, w_021_831, w_021_832, w_021_833, w_021_834, w_021_835, w_021_836, w_021_837, w_021_838, w_021_839, w_021_840, w_021_841, w_021_842, w_021_843, w_021_844, w_021_845, w_021_846, w_021_847, w_021_848, w_021_849, w_021_850, w_021_851;
  wire w_022_000, w_022_001, w_022_002, w_022_003, w_022_004, w_022_005, w_022_006, w_022_008, w_022_010, w_022_011, w_022_012, w_022_013, w_022_016, w_022_018, w_022_019, w_022_020, w_022_022, w_022_023, w_022_025, w_022_026, w_022_027, w_022_028, w_022_029, w_022_030, w_022_031, w_022_032, w_022_033, w_022_035, w_022_036, w_022_037, w_022_038, w_022_039, w_022_040, w_022_041, w_022_042, w_022_043, w_022_044, w_022_045, w_022_047, w_022_048, w_022_050, w_022_051, w_022_055, w_022_058, w_022_060, w_022_061, w_022_065, w_022_067, w_022_070, w_022_072, w_022_073, w_022_074, w_022_076, w_022_080, w_022_083, w_022_084, w_022_086, w_022_087, w_022_088, w_022_092, w_022_093, w_022_094, w_022_099, w_022_100, w_022_101, w_022_105, w_022_106, w_022_107, w_022_108, w_022_115, w_022_116, w_022_118, w_022_121, w_022_122, w_022_123, w_022_124, w_022_126, w_022_130, w_022_131, w_022_133, w_022_134, w_022_135, w_022_136, w_022_137, w_022_138, w_022_140, w_022_142, w_022_144, w_022_146, w_022_147, w_022_148, w_022_149, w_022_152, w_022_153, w_022_154, w_022_155, w_022_157, w_022_158, w_022_159, w_022_160, w_022_161, w_022_163, w_022_164, w_022_165, w_022_169, w_022_172, w_022_174, w_022_175, w_022_178, w_022_179, w_022_180, w_022_182, w_022_184, w_022_185, w_022_189, w_022_191, w_022_192, w_022_193, w_022_197, w_022_199, w_022_201, w_022_202, w_022_205, w_022_206, w_022_208, w_022_210, w_022_213, w_022_214, w_022_215, w_022_216, w_022_218, w_022_219, w_022_220, w_022_221, w_022_222, w_022_223, w_022_224, w_022_225, w_022_227, w_022_230, w_022_232, w_022_233, w_022_236, w_022_237, w_022_238, w_022_239, w_022_240, w_022_241, w_022_242, w_022_243, w_022_244, w_022_246, w_022_248, w_022_250, w_022_251, w_022_252, w_022_254, w_022_255, w_022_257, w_022_258, w_022_259, w_022_260, w_022_263, w_022_265, w_022_266, w_022_267, w_022_268, w_022_269, w_022_270, w_022_274, w_022_276, w_022_277, w_022_280, w_022_282, w_022_283, w_022_284, w_022_286, w_022_289, w_022_291, w_022_292, w_022_294, w_022_295, w_022_297, w_022_298, w_022_300, w_022_302, w_022_303, w_022_304, w_022_305, w_022_306, w_022_308, w_022_310, w_022_312, w_022_316, w_022_317, w_022_319, w_022_320, w_022_322, w_022_323, w_022_324, w_022_325, w_022_326, w_022_327, w_022_330, w_022_331, w_022_333, w_022_334, w_022_336, w_022_337, w_022_339, w_022_340, w_022_341, w_022_344, w_022_345, w_022_350, w_022_351, w_022_352, w_022_353, w_022_355, w_022_356, w_022_357, w_022_358, w_022_359, w_022_360, w_022_361, w_022_362, w_022_365, w_022_367, w_022_368, w_022_371, w_022_373, w_022_374, w_022_377, w_022_380, w_022_381, w_022_382, w_022_383, w_022_385, w_022_387, w_022_388, w_022_391, w_022_395, w_022_397, w_022_398, w_022_399, w_022_400, w_022_402, w_022_403, w_022_405, w_022_406, w_022_407, w_022_408, w_022_410, w_022_411, w_022_413, w_022_414, w_022_415, w_022_417, w_022_418, w_022_419, w_022_420, w_022_422, w_022_424, w_022_425, w_022_427, w_022_428, w_022_429, w_022_430, w_022_432, w_022_433, w_022_434, w_022_435, w_022_436, w_022_438, w_022_439, w_022_440, w_022_441, w_022_443, w_022_445, w_022_446, w_022_447, w_022_448, w_022_451, w_022_452, w_022_453, w_022_454, w_022_458, w_022_459, w_022_460, w_022_461, w_022_462, w_022_464, w_022_465, w_022_467, w_022_468, w_022_469, w_022_470, w_022_473, w_022_474, w_022_475, w_022_476, w_022_477, w_022_480, w_022_482, w_022_484, w_022_485, w_022_486, w_022_487, w_022_489, w_022_490, w_022_491, w_022_492, w_022_495, w_022_498, w_022_499, w_022_500, w_022_501, w_022_502, w_022_503, w_022_504, w_022_506, w_022_508, w_022_509, w_022_510, w_022_512, w_022_513, w_022_515, w_022_517, w_022_519, w_022_520, w_022_521, w_022_522, w_022_523, w_022_524, w_022_525, w_022_529, w_022_530, w_022_532, w_022_533, w_022_534, w_022_535, w_022_536, w_022_537, w_022_538, w_022_539, w_022_541, w_022_542, w_022_543, w_022_544, w_022_545, w_022_548, w_022_549, w_022_550, w_022_551, w_022_552, w_022_553, w_022_556, w_022_557, w_022_558, w_022_560, w_022_565, w_022_570, w_022_571, w_022_572, w_022_575, w_022_576, w_022_580, w_022_581, w_022_584, w_022_585, w_022_586, w_022_587, w_022_588, w_022_590, w_022_591, w_022_592, w_022_594, w_022_597, w_022_600, w_022_601, w_022_602, w_022_603, w_022_604, w_022_605, w_022_609, w_022_611, w_022_612, w_022_614, w_022_615, w_022_620, w_022_621, w_022_622, w_022_623, w_022_624, w_022_626, w_022_627, w_022_629, w_022_631, w_022_632, w_022_633, w_022_634, w_022_636, w_022_639, w_022_640, w_022_641, w_022_642, w_022_643, w_022_644, w_022_646, w_022_647, w_022_648, w_022_649, w_022_650, w_022_652, w_022_653, w_022_654, w_022_655, w_022_660, w_022_661, w_022_663, w_022_664, w_022_666, w_022_668, w_022_669, w_022_672, w_022_673, w_022_674, w_022_676, w_022_677, w_022_678, w_022_679, w_022_680, w_022_681, w_022_682, w_022_684, w_022_686, w_022_687, w_022_688, w_022_690, w_022_691, w_022_693, w_022_694, w_022_697, w_022_700, w_022_702, w_022_704, w_022_706, w_022_707, w_022_708, w_022_709, w_022_710, w_022_713, w_022_715, w_022_717, w_022_721, w_022_723, w_022_724, w_022_725, w_022_727, w_022_730, w_022_731, w_022_732, w_022_733, w_022_734, w_022_735, w_022_736, w_022_739, w_022_740, w_022_741, w_022_742, w_022_745, w_022_746, w_022_747, w_022_751, w_022_753, w_022_755, w_022_756, w_022_758, w_022_759, w_022_762, w_022_763, w_022_764, w_022_766, w_022_768, w_022_769, w_022_770, w_022_771, w_022_772, w_022_774, w_022_775, w_022_776, w_022_778, w_022_782, w_022_783, w_022_786, w_022_787, w_022_788, w_022_793, w_022_795, w_022_796, w_022_797, w_022_798, w_022_799, w_022_801, w_022_802, w_022_803, w_022_804, w_022_805, w_022_808, w_022_811, w_022_812, w_022_813, w_022_814, w_022_817, w_022_818, w_022_819, w_022_821, w_022_822, w_022_825, w_022_826, w_022_827, w_022_829, w_022_833, w_022_835, w_022_836, w_022_837, w_022_847, w_022_848, w_022_849, w_022_850, w_022_851, w_022_852, w_022_853, w_022_854, w_022_855, w_022_856, w_022_857, w_022_858, w_022_860, w_022_862, w_022_866, w_022_867, w_022_868, w_022_869, w_022_870, w_022_873, w_022_874, w_022_876, w_022_878, w_022_879, w_022_880, w_022_882, w_022_888, w_022_889, w_022_890, w_022_892, w_022_893, w_022_896, w_022_897, w_022_898, w_022_899, w_022_902, w_022_903, w_022_904, w_022_905, w_022_908, w_022_909, w_022_910, w_022_911, w_022_913, w_022_914, w_022_915, w_022_916, w_022_917, w_022_921, w_022_922, w_022_923, w_022_924, w_022_925, w_022_926, w_022_927, w_022_930, w_022_931, w_022_934, w_022_935, w_022_937, w_022_941, w_022_942, w_022_944, w_022_945, w_022_947, w_022_948, w_022_952, w_022_953, w_022_954, w_022_955, w_022_956, w_022_957, w_022_958, w_022_959, w_022_960, w_022_961, w_022_965, w_022_967, w_022_969, w_022_971, w_022_972, w_022_975, w_022_978, w_022_980, w_022_981, w_022_983, w_022_985, w_022_986, w_022_987, w_022_989, w_022_990, w_022_992, w_022_994, w_022_995, w_022_1001, w_022_1002, w_022_1003, w_022_1004, w_022_1005, w_022_1010, w_022_1011, w_022_1012, w_022_1013, w_022_1015, w_022_1016, w_022_1017, w_022_1018, w_022_1019, w_022_1021, w_022_1023, w_022_1024, w_022_1025, w_022_1027, w_022_1029, w_022_1033, w_022_1035, w_022_1036, w_022_1038, w_022_1039, w_022_1040, w_022_1041, w_022_1043, w_022_1044, w_022_1047, w_022_1048, w_022_1049, w_022_1052, w_022_1053, w_022_1054, w_022_1055, w_022_1056, w_022_1057, w_022_1058, w_022_1061, w_022_1065, w_022_1068, w_022_1069, w_022_1070, w_022_1072, w_022_1073, w_022_1074, w_022_1075, w_022_1076, w_022_1078, w_022_1079, w_022_1080, w_022_1083, w_022_1084, w_022_1085, w_022_1087, w_022_1090, w_022_1091, w_022_1093, w_022_1094, w_022_1098, w_022_1102, w_022_1113, w_022_1114, w_022_1116, w_022_1118, w_022_1119, w_022_1121, w_022_1122, w_022_1123, w_022_1124, w_022_1126, w_022_1129, w_022_1130, w_022_1132, w_022_1133, w_022_1135, w_022_1138, w_022_1141, w_022_1144, w_022_1147, w_022_1148, w_022_1149, w_022_1150, w_022_1152, w_022_1154, w_022_1157, w_022_1159, w_022_1162, w_022_1165, w_022_1166, w_022_1167, w_022_1168, w_022_1169, w_022_1170, w_022_1172, w_022_1173, w_022_1175, w_022_1176, w_022_1178, w_022_1179, w_022_1180, w_022_1183, w_022_1185, w_022_1187, w_022_1189, w_022_1190, w_022_1191, w_022_1192, w_022_1193, w_022_1194, w_022_1195, w_022_1198, w_022_1199, w_022_1200, w_022_1201, w_022_1202, w_022_1203, w_022_1205, w_022_1207, w_022_1208, w_022_1209, w_022_1212, w_022_1213, w_022_1214, w_022_1215, w_022_1216, w_022_1217, w_022_1220, w_022_1221, w_022_1222, w_022_1224, w_022_1226, w_022_1231, w_022_1232, w_022_1233, w_022_1234, w_022_1235, w_022_1236, w_022_1238, w_022_1243, w_022_1244, w_022_1248, w_022_1251, w_022_1253, w_022_1254, w_022_1255, w_022_1257, w_022_1258, w_022_1259, w_022_1260, w_022_1266, w_022_1268, w_022_1269, w_022_1271, w_022_1273, w_022_1274, w_022_1276, w_022_1279, w_022_1280, w_022_1281, w_022_1282, w_022_1283, w_022_1284, w_022_1286, w_022_1290, w_022_1292, w_022_1293, w_022_1296, w_022_1297, w_022_1298, w_022_1299, w_022_1301, w_022_1305, w_022_1306, w_022_1309, w_022_1310, w_022_1311, w_022_1314, w_022_1315, w_022_1316, w_022_1318, w_022_1319, w_022_1320, w_022_1322, w_022_1323, w_022_1324, w_022_1325, w_022_1326, w_022_1328, w_022_1329, w_022_1330, w_022_1332, w_022_1333, w_022_1339, w_022_1342, w_022_1343, w_022_1344, w_022_1348, w_022_1351, w_022_1352, w_022_1353, w_022_1357, w_022_1358, w_022_1361, w_022_1362, w_022_1363, w_022_1364, w_022_1365, w_022_1366, w_022_1369, w_022_1370, w_022_1373, w_022_1376, w_022_1378, w_022_1379, w_022_1380, w_022_1382, w_022_1383, w_022_1384, w_022_1385, w_022_1386, w_022_1387, w_022_1389, w_022_1392, w_022_1393, w_022_1395, w_022_1396, w_022_1397, w_022_1398, w_022_1400, w_022_1401, w_022_1402, w_022_1403, w_022_1405, w_022_1406, w_022_1407, w_022_1408, w_022_1409, w_022_1411, w_022_1412, w_022_1413, w_022_1415, w_022_1416, w_022_1417, w_022_1418, w_022_1419, w_022_1421, w_022_1422, w_022_1423, w_022_1424, w_022_1425, w_022_1427, w_022_1428, w_022_1429, w_022_1430, w_022_1431, w_022_1433, w_022_1434, w_022_1435, w_022_1441, w_022_1442, w_022_1443, w_022_1444, w_022_1446, w_022_1447, w_022_1451, w_022_1453, w_022_1455, w_022_1459, w_022_1460, w_022_1461, w_022_1462, w_022_1463, w_022_1464, w_022_1465, w_022_1466, w_022_1468, w_022_1473, w_022_1478, w_022_1479, w_022_1480, w_022_1481, w_022_1483, w_022_1486, w_022_1487, w_022_1488, w_022_1490, w_022_1491, w_022_1492, w_022_1493, w_022_1494, w_022_1495, w_022_1496, w_022_1497, w_022_1501, w_022_1504, w_022_1505, w_022_1506, w_022_1507, w_022_1508, w_022_1512, w_022_1513, w_022_1516, w_022_1517, w_022_1521, w_022_1523, w_022_1525, w_022_1526, w_022_1528, w_022_1529, w_022_1530, w_022_1533, w_022_1534, w_022_1536, w_022_1539, w_022_1540, w_022_1542, w_022_1543, w_022_1545, w_022_1547, w_022_1549, w_022_1550, w_022_1551, w_022_1554, w_022_1556, w_022_1559, w_022_1560, w_022_1561, w_022_1563, w_022_1567, w_022_1568, w_022_1569, w_022_1570, w_022_1571, w_022_1573, w_022_1574, w_022_1577, w_022_1578, w_022_1580, w_022_1581, w_022_1583, w_022_1588, w_022_1590, w_022_1591, w_022_1592, w_022_1593, w_022_1595, w_022_1597, w_022_1598, w_022_1599, w_022_1601, w_022_1602, w_022_1603, w_022_1606, w_022_1607, w_022_1609, w_022_1610, w_022_1611, w_022_1612, w_022_1614, w_022_1615, w_022_1616, w_022_1620, w_022_1622, w_022_1623, w_022_1625, w_022_1626, w_022_1627, w_022_1628, w_022_1630, w_022_1631, w_022_1634, w_022_1636, w_022_1637, w_022_1638, w_022_1639, w_022_1640, w_022_1645, w_022_1646, w_022_1649, w_022_1650, w_022_1652, w_022_1653, w_022_1654, w_022_1655, w_022_1656, w_022_1657, w_022_1658, w_022_1661, w_022_1662, w_022_1663, w_022_1665, w_022_1669, w_022_1670, w_022_1671, w_022_1672, w_022_1674, w_022_1676, w_022_1677, w_022_1681, w_022_1683, w_022_1685, w_022_1687, w_022_1690, w_022_1691, w_022_1692, w_022_1695, w_022_1696, w_022_1698, w_022_1701, w_022_1702, w_022_1703, w_022_1704, w_022_1705, w_022_1706, w_022_1707, w_022_1710, w_022_1714, w_022_1715, w_022_1716, w_022_1717, w_022_1719, w_022_1720, w_022_1721, w_022_1722, w_022_1724, w_022_1725, w_022_1727, w_022_1730, w_022_1731, w_022_1732, w_022_1736, w_022_1737, w_022_1741, w_022_1742, w_022_1744, w_022_1745, w_022_1746, w_022_1748, w_022_1749, w_022_1753, w_022_1754, w_022_1756, w_022_1757, w_022_1758, w_022_1759, w_022_1762, w_022_1763, w_022_1764, w_022_1766, w_022_1767, w_022_1768, w_022_1769, w_022_1770, w_022_1773, w_022_1774, w_022_1775, w_022_1776, w_022_1777, w_022_1778, w_022_1781, w_022_1782, w_022_1783, w_022_1785, w_022_1786, w_022_1789, w_022_1791, w_022_1792, w_022_1794, w_022_1798, w_022_1801, w_022_1803, w_022_1804, w_022_1805, w_022_1808, w_022_1810, w_022_1811, w_022_1812, w_022_1814, w_022_1816, w_022_1819, w_022_1820, w_022_1821, w_022_1824, w_022_1826, w_022_1827, w_022_1830, w_022_1831, w_022_1832, w_022_1833, w_022_1834, w_022_1835, w_022_1837, w_022_1838, w_022_1839, w_022_1840, w_022_1844, w_022_1845, w_022_1849, w_022_1850, w_022_1851, w_022_1853, w_022_1854, w_022_1857, w_022_1858, w_022_1859, w_022_1860, w_022_1863, w_022_1864, w_022_1865, w_022_1868, w_022_1870, w_022_1873, w_022_1874, w_022_1876, w_022_1879, w_022_1880, w_022_1881, w_022_1884, w_022_1888, w_022_1890, w_022_1892, w_022_1896, w_022_1898, w_022_1901, w_022_1904, w_022_1905, w_022_1907, w_022_1908, w_022_1909, w_022_1910, w_022_1911, w_022_1913, w_022_1914, w_022_1915, w_022_1918, w_022_1919, w_022_1922, w_022_1923, w_022_1924, w_022_1926, w_022_1927, w_022_1928, w_022_1931, w_022_1932, w_022_1933, w_022_1934, w_022_1938, w_022_1942, w_022_1945, w_022_1946, w_022_1947, w_022_1948, w_022_1949, w_022_1950, w_022_1951, w_022_1952, w_022_1953, w_022_1954, w_022_1956, w_022_1957, w_022_1963, w_022_1964, w_022_1965, w_022_1969, w_022_1971, w_022_1974, w_022_1978, w_022_1982, w_022_1983, w_022_1984, w_022_1986, w_022_1989, w_022_1990, w_022_1993, w_022_1994, w_022_1995, w_022_1996, w_022_1997, w_022_1998, w_022_2001, w_022_2003, w_022_2005, w_022_2007, w_022_2009, w_022_2012, w_022_2013, w_022_2018, w_022_2020, w_022_2021, w_022_2022, w_022_2023, w_022_2026, w_022_2027, w_022_2028, w_022_2029, w_022_2030, w_022_2031, w_022_2032, w_022_2034, w_022_2037, w_022_2041, w_022_2042, w_022_2043, w_022_2044, w_022_2046, w_022_2049, w_022_2050, w_022_2051, w_022_2052, w_022_2054, w_022_2057, w_022_2058, w_022_2061, w_022_2062, w_022_2063, w_022_2064, w_022_2066, w_022_2067, w_022_2070, w_022_2072, w_022_2073, w_022_2075, w_022_2076, w_022_2078, w_022_2080, w_022_2081, w_022_2082, w_022_2083, w_022_2085, w_022_2086, w_022_2087, w_022_2088, w_022_2090, w_022_2093, w_022_2098, w_022_2101, w_022_2104, w_022_2105, w_022_2106, w_022_2107, w_022_2108, w_022_2109, w_022_2110, w_022_2111, w_022_2112, w_022_2114, w_022_2117, w_022_2120, w_022_2121, w_022_2122, w_022_2123, w_022_2124, w_022_2125, w_022_2127, w_022_2128, w_022_2130, w_022_2131, w_022_2132, w_022_2133, w_022_2135, w_022_2136, w_022_2137, w_022_2138, w_022_2140, w_022_2141, w_022_2142, w_022_2143, w_022_2144, w_022_2145, w_022_2147, w_022_2149, w_022_2151, w_022_2154, w_022_2157, w_022_2158, w_022_2159, w_022_2163, w_022_2164, w_022_2166, w_022_2171, w_022_2172, w_022_2174, w_022_2176, w_022_2179, w_022_2182, w_022_2183, w_022_2185, w_022_2188, w_022_2189, w_022_2190, w_022_2192, w_022_2194, w_022_2195, w_022_2196, w_022_2197, w_022_2198, w_022_2199, w_022_2200, w_022_2202, w_022_2203, w_022_2204, w_022_2205, w_022_2206, w_022_2207, w_022_2208, w_022_2210, w_022_2211, w_022_2212, w_022_2215, w_022_2216, w_022_2218, w_022_2220, w_022_2221, w_022_2224, w_022_2225, w_022_2229, w_022_2233, w_022_2235, w_022_2237, w_022_2238, w_022_2239, w_022_2240, w_022_2241, w_022_2242, w_022_2243, w_022_2244, w_022_2248, w_022_2251, w_022_2252, w_022_2255, w_022_2257, w_022_2258, w_022_2260, w_022_2261, w_022_2265, w_022_2268, w_022_2271, w_022_2272, w_022_2279, w_022_2281, w_022_2282, w_022_2285, w_022_2286, w_022_2295, w_022_2297, w_022_2298, w_022_2299, w_022_2301, w_022_2302, w_022_2304, w_022_2305, w_022_2307, w_022_2308, w_022_2309, w_022_2310, w_022_2311, w_022_2312, w_022_2314, w_022_2315, w_022_2318, w_022_2319, w_022_2321, w_022_2322, w_022_2323, w_022_2324, w_022_2325, w_022_2326, w_022_2327, w_022_2332, w_022_2333, w_022_2334, w_022_2335, w_022_2336, w_022_2337, w_022_2340, w_022_2341, w_022_2342, w_022_2344, w_022_2346, w_022_2347, w_022_2348, w_022_2350, w_022_2351, w_022_2354, w_022_2355, w_022_2356, w_022_2358, w_022_2360, w_022_2361, w_022_2363, w_022_2364, w_022_2365, w_022_2366, w_022_2367, w_022_2368, w_022_2371, w_022_2372, w_022_2373, w_022_2377, w_022_2378, w_022_2381, w_022_2382, w_022_2383, w_022_2384, w_022_2385, w_022_2387, w_022_2388, w_022_2389, w_022_2390, w_022_2391, w_022_2396, w_022_2398, w_022_2399, w_022_2401, w_022_2402, w_022_2403, w_022_2404, w_022_2406, w_022_2407, w_022_2408, w_022_2409, w_022_2412, w_022_2414, w_022_2415, w_022_2416, w_022_2418, w_022_2419, w_022_2422, w_022_2428, w_022_2429, w_022_2431, w_022_2432, w_022_2434, w_022_2435, w_022_2436, w_022_2437, w_022_2438, w_022_2439, w_022_2440, w_022_2443, w_022_2448, w_022_2449, w_022_2451, w_022_2453, w_022_2455, w_022_2456, w_022_2457, w_022_2458, w_022_2460, w_022_2462, w_022_2465, w_022_2468, w_022_2471, w_022_2474, w_022_2475, w_022_2476, w_022_2477, w_022_2478, w_022_2480, w_022_2481, w_022_2484, w_022_2486, w_022_2488, w_022_2489, w_022_2490, w_022_2491, w_022_2494, w_022_2495, w_022_2497, w_022_2498, w_022_2500, w_022_2501, w_022_2502, w_022_2503, w_022_2504, w_022_2505, w_022_2506, w_022_2507, w_022_2509, w_022_2510, w_022_2511, w_022_2512, w_022_2514, w_022_2515, w_022_2517, w_022_2518, w_022_2519, w_022_2521, w_022_2526, w_022_2527, w_022_2528, w_022_2530, w_022_2536, w_022_2538, w_022_2539, w_022_2541, w_022_2543, w_022_2545, w_022_2548, w_022_2550, w_022_2551, w_022_2553, w_022_2555, w_022_2556, w_022_2557, w_022_2558, w_022_2559, w_022_2560, w_022_2561, w_022_2562, w_022_2564, w_022_2566, w_022_2568, w_022_2569, w_022_2571, w_022_2572, w_022_2574, w_022_2575, w_022_2576, w_022_2577, w_022_2578, w_022_2580, w_022_2583, w_022_2585, w_022_2586, w_022_2589, w_022_2590, w_022_2591, w_022_2594, w_022_2595, w_022_2597, w_022_2598, w_022_2602, w_022_2603, w_022_2604, w_022_2605, w_022_2606, w_022_2607, w_022_2608, w_022_2610, w_022_2611, w_022_2613, w_022_2614, w_022_2615, w_022_2616, w_022_2617, w_022_2618, w_022_2619, w_022_2621, w_022_2622, w_022_2623, w_022_2624, w_022_2625, w_022_2626, w_022_2628, w_022_2629, w_022_2630, w_022_2632, w_022_2633, w_022_2635, w_022_2636, w_022_2640, w_022_2642, w_022_2643, w_022_2645, w_022_2646, w_022_2647, w_022_2649, w_022_2650, w_022_2651, w_022_2652, w_022_2653, w_022_2654, w_022_2656, w_022_2657, w_022_2658, w_022_2660, w_022_2661, w_022_2662, w_022_2663, w_022_2665, w_022_2667, w_022_2668, w_022_2670, w_022_2671, w_022_2673, w_022_2674, w_022_2675, w_022_2677, w_022_2679, w_022_2680, w_022_2686, w_022_2687, w_022_2688, w_022_2689, w_022_2690, w_022_2691, w_022_2694, w_022_2695, w_022_2698, w_022_2700, w_022_2701, w_022_2704, w_022_2705, w_022_2708, w_022_2710, w_022_2711, w_022_2712, w_022_2714, w_022_2716, w_022_2718, w_022_2719, w_022_2720, w_022_2722, w_022_2723, w_022_2724, w_022_2725, w_022_2726, w_022_2728, w_022_2729, w_022_2730, w_022_2734, w_022_2735, w_022_2737, w_022_2738, w_022_2740, w_022_2742, w_022_2743, w_022_2746, w_022_2747, w_022_2754, w_022_2757, w_022_2758, w_022_2761, w_022_2764, w_022_2765, w_022_2766, w_022_2769, w_022_2771, w_022_2772, w_022_2775, w_022_2776, w_022_2778, w_022_2780, w_022_2781, w_022_2782, w_022_2785, w_022_2786, w_022_2787, w_022_2794, w_022_2795, w_022_2797, w_022_2798, w_022_2799, w_022_2801, w_022_2802, w_022_2803, w_022_2804, w_022_2805, w_022_2807, w_022_2808, w_022_2811, w_022_2812, w_022_2813, w_022_2814, w_022_2815, w_022_2816, w_022_2819, w_022_2820, w_022_2821, w_022_2823, w_022_2824, w_022_2827, w_022_2828, w_022_2829, w_022_2831, w_022_2832, w_022_2834, w_022_2835, w_022_2838, w_022_2841, w_022_2842, w_022_2843, w_022_2844, w_022_2845, w_022_2846, w_022_2847, w_022_2850, w_022_2853, w_022_2855, w_022_2856, w_022_2857, w_022_2858, w_022_2861, w_022_2862, w_022_2863, w_022_2865, w_022_2867, w_022_2868, w_022_2869, w_022_2872, w_022_2873, w_022_2875, w_022_2878, w_022_2879, w_022_2880, w_022_2881, w_022_2882, w_022_2883, w_022_2885, w_022_2887, w_022_2888, w_022_2891, w_022_2893, w_022_2896, w_022_2897, w_022_2898, w_022_2899, w_022_2900, w_022_2901, w_022_2902, w_022_2903, w_022_2906, w_022_2908, w_022_2909, w_022_2910, w_022_2911, w_022_2912, w_022_2914, w_022_2915, w_022_2918, w_022_2919, w_022_2920, w_022_2921, w_022_2922, w_022_2923, w_022_2926, w_022_2928, w_022_2930, w_022_2931, w_022_2932, w_022_2933, w_022_2936, w_022_2937, w_022_2941, w_022_2943, w_022_2944, w_022_2945, w_022_2947, w_022_2948, w_022_2949, w_022_2951, w_022_2952, w_022_2953, w_022_2954, w_022_2955, w_022_2957, w_022_2958, w_022_2959, w_022_2961, w_022_2962, w_022_2963, w_022_2968, w_022_2969, w_022_2972, w_022_2973, w_022_2974, w_022_2976, w_022_2977, w_022_2978, w_022_2979, w_022_2980, w_022_2981, w_022_2982, w_022_2983, w_022_2984, w_022_2986, w_022_2988, w_022_2989, w_022_2992, w_022_2996, w_022_2999, w_022_3000, w_022_3001, w_022_3002, w_022_3003, w_022_3004, w_022_3005, w_022_3007, w_022_3008, w_022_3009, w_022_3010, w_022_3012, w_022_3013, w_022_3014, w_022_3016, w_022_3018, w_022_3020, w_022_3021, w_022_3024, w_022_3025, w_022_3026, w_022_3027, w_022_3028, w_022_3031, w_022_3032, w_022_3034, w_022_3035, w_022_3038, w_022_3039, w_022_3042, w_022_3043, w_022_3044, w_022_3045, w_022_3046, w_022_3050, w_022_3051, w_022_3052, w_022_3054, w_022_3055, w_022_3056, w_022_3058, w_022_3060, w_022_3062, w_022_3063, w_022_3065, w_022_3066, w_022_3067, w_022_3069, w_022_3070, w_022_3071, w_022_3073, w_022_3074, w_022_3075, w_022_3077, w_022_3079, w_022_3080, w_022_3081, w_022_3083, w_022_3084, w_022_3085, w_022_3088, w_022_3090, w_022_3091, w_022_3092, w_022_3093, w_022_3095, w_022_3096, w_022_3097, w_022_3098, w_022_3102, w_022_3103, w_022_3104, w_022_3106, w_022_3107, w_022_3111, w_022_3113, w_022_3115, w_022_3116, w_022_3117, w_022_3118, w_022_3121, w_022_3126, w_022_3128, w_022_3131, w_022_3132, w_022_3134, w_022_3136, w_022_3137, w_022_3139, w_022_3140, w_022_3141, w_022_3142, w_022_3143, w_022_3144, w_022_3146, w_022_3149, w_022_3150, w_022_3151, w_022_3154, w_022_3155, w_022_3159, w_022_3160, w_022_3162, w_022_3163, w_022_3165, w_022_3166, w_022_3167, w_022_3168, w_022_3170, w_022_3171, w_022_3172, w_022_3173, w_022_3176, w_022_3177, w_022_3178, w_022_3179, w_022_3180, w_022_3182, w_022_3185, w_022_3186, w_022_3188, w_022_3189, w_022_3190, w_022_3195, w_022_3196, w_022_3198, w_022_3199, w_022_3201, w_022_3202, w_022_3203, w_022_3204, w_022_3205, w_022_3207, w_022_3209, w_022_3211, w_022_3214, w_022_3215, w_022_3216, w_022_3219, w_022_3220, w_022_3222, w_022_3224, w_022_3227, w_022_3229, w_022_3230, w_022_3231, w_022_3232, w_022_3233, w_022_3235, w_022_3236, w_022_3237, w_022_3238, w_022_3239, w_022_3241, w_022_3243, w_022_3246, w_022_3247, w_022_3248, w_022_3254, w_022_3256, w_022_3257, w_022_3259, w_022_3260, w_022_3264, w_022_3267, w_022_3268, w_022_3270, w_022_3273, w_022_3274, w_022_3275, w_022_3277, w_022_3279, w_022_3280, w_022_3281, w_022_3282, w_022_3283, w_022_3286, w_022_3287, w_022_3288, w_022_3289, w_022_3290, w_022_3291, w_022_3292, w_022_3293, w_022_3294, w_022_3295, w_022_3296, w_022_3297, w_022_3298, w_022_3301, w_022_3302, w_022_3303, w_022_3304, w_022_3305, w_022_3306, w_022_3307, w_022_3311, w_022_3312, w_022_3314, w_022_3315, w_022_3317, w_022_3319, w_022_3320, w_022_3321, w_022_3324, w_022_3325, w_022_3327, w_022_3328, w_022_3330, w_022_3332, w_022_3334, w_022_3335, w_022_3336, w_022_3337, w_022_3338, w_022_3340, w_022_3343, w_022_3344, w_022_3346, w_022_3347, w_022_3351, w_022_3353, w_022_3354, w_022_3355, w_022_3356, w_022_3357, w_022_3358, w_022_3359, w_022_3360, w_022_3361, w_022_3364, w_022_3365, w_022_3366, w_022_3368, w_022_3369, w_022_3370, w_022_3372, w_022_3373, w_022_3376, w_022_3378, w_022_3380, w_022_3381, w_022_3382, w_022_3383, w_022_3384, w_022_3385, w_022_3389, w_022_3391, w_022_3392, w_022_3393, w_022_3394, w_022_3396, w_022_3397, w_022_3398, w_022_3399, w_022_3402, w_022_3403, w_022_3404, w_022_3406, w_022_3407, w_022_3408, w_022_3409, w_022_3410, w_022_3411, w_022_3412, w_022_3413, w_022_3415, w_022_3416, w_022_3418, w_022_3420, w_022_3421, w_022_3423, w_022_3424, w_022_3425, w_022_3429, w_022_3431, w_022_3433, w_022_3434, w_022_3435, w_022_3437, w_022_3439, w_022_3440, w_022_3441, w_022_3442, w_022_3443, w_022_3444, w_022_3445, w_022_3446, w_022_3447, w_022_3448, w_022_3451, w_022_3454, w_022_3456, w_022_3457, w_022_3458, w_022_3465, w_022_3468, w_022_3469, w_022_3470, w_022_3471, w_022_3474, w_022_3475, w_022_3476, w_022_3477, w_022_3478, w_022_3479, w_022_3480, w_022_3481, w_022_3482, w_022_3484, w_022_3485, w_022_3488, w_022_3490, w_022_3491, w_022_3492, w_022_3493, w_022_3495, w_022_3496, w_022_3497, w_022_3498, w_022_3499, w_022_3501, w_022_3502, w_022_3504, w_022_3505, w_022_3509, w_022_3510, w_022_3513, w_022_3514, w_022_3517, w_022_3518, w_022_3519, w_022_3520, w_022_3521, w_022_3522, w_022_3524, w_022_3525, w_022_3526, w_022_3527, w_022_3529, w_022_3531, w_022_3532, w_022_3534, w_022_3536, w_022_3537, w_022_3539, w_022_3540, w_022_3542, w_022_3544, w_022_3546, w_022_3547, w_022_3549, w_022_3551, w_022_3552, w_022_3553, w_022_3554, w_022_3555, w_022_3556, w_022_3557, w_022_3559, w_022_3560, w_022_3561, w_022_3562, w_022_3563, w_022_3565, w_022_3566, w_022_3568, w_022_3569, w_022_3570, w_022_3572, w_022_3575, w_022_3576, w_022_3578, w_022_3581, w_022_3583, w_022_3585, w_022_3587, w_022_3589, w_022_3590, w_022_3591, w_022_3594, w_022_3596, w_022_3598, w_022_3599, w_022_3600, w_022_3601, w_022_3603, w_022_3606, w_022_3610, w_022_3612, w_022_3613, w_022_3614, w_022_3616, w_022_3617, w_022_3619, w_022_3620, w_022_3622, w_022_3623, w_022_3624, w_022_3625, w_022_3628, w_022_3631, w_022_3634, w_022_3635, w_022_3637, w_022_3639, w_022_3641, w_022_3642, w_022_3643, w_022_3645, w_022_3646, w_022_3648, w_022_3649, w_022_3650, w_022_3651, w_022_3652, w_022_3653, w_022_3655, w_022_3656, w_022_3657, w_022_3658, w_022_3659, w_022_3661, w_022_3663, w_022_3664, w_022_3666, w_022_3669, w_022_3670, w_022_3676, w_022_3677, w_022_3678, w_022_3679, w_022_3680, w_022_3681, w_022_3682, w_022_3683, w_022_3684, w_022_3685, w_022_3689, w_022_3690, w_022_3691, w_022_3693, w_022_3695, w_022_3697, w_022_3698, w_022_3699, w_022_3700, w_022_3701, w_022_3702, w_022_3704, w_022_3707, w_022_3711, w_022_3713, w_022_3714, w_022_3715, w_022_3716, w_022_3717, w_022_3719, w_022_3722, w_022_3723, w_022_3724, w_022_3725, w_022_3726, w_022_3730, w_022_3731, w_022_3732, w_022_3734, w_022_3735, w_022_3736, w_022_3737, w_022_3738, w_022_3740, w_022_3743, w_022_3744, w_022_3745, w_022_3746, w_022_3747, w_022_3749, w_022_3750, w_022_3751, w_022_3754, w_022_3756, w_022_3758, w_022_3759, w_022_3760, w_022_3761, w_022_3762, w_022_3766, w_022_3767, w_022_3768, w_022_3771, w_022_3773, w_022_3777, w_022_3778, w_022_3779, w_022_3780, w_022_3781, w_022_3782, w_022_3783, w_022_3784, w_022_3785, w_022_3786, w_022_3787, w_022_3788, w_022_3789, w_022_3790, w_022_3791, w_022_3794, w_022_3797, w_022_3800, w_022_3801, w_022_3802, w_022_3804, w_022_3805, w_022_3806, w_022_3807, w_022_3809, w_022_3810, w_022_3812, w_022_3813, w_022_3815, w_022_3816, w_022_3818, w_022_3819, w_022_3821, w_022_3822, w_022_3824, w_022_3825, w_022_3826, w_022_3830, w_022_3834, w_022_3835, w_022_3836, w_022_3837, w_022_3838, w_022_3841, w_022_3843, w_022_3844, w_022_3845, w_022_3846, w_022_3850, w_022_3851, w_022_3852, w_022_3853, w_022_3855, w_022_3856, w_022_3857, w_022_3860, w_022_3861, w_022_3866, w_022_3868, w_022_3869, w_022_3870, w_022_3871, w_022_3872, w_022_3873, w_022_3876, w_022_3878, w_022_3882, w_022_3883, w_022_3885, w_022_3886, w_022_3888, w_022_3890, w_022_3891, w_022_3892, w_022_3894, w_022_3898, w_022_3902, w_022_3903, w_022_3905, w_022_3907, w_022_3910, w_022_3911, w_022_3915, w_022_3919, w_022_3920, w_022_3921, w_022_3922, w_022_3924, w_022_3927, w_022_3928, w_022_3931, w_022_3932, w_022_3933, w_022_3935, w_022_3937, w_022_3938, w_022_3939, w_022_3940, w_022_3942, w_022_3943, w_022_3944, w_022_3945, w_022_3946, w_022_3947, w_022_3948, w_022_3949, w_022_3950, w_022_3951, w_022_3952, w_022_3953, w_022_3954, w_022_3955, w_022_3957, w_022_3958, w_022_3959, w_022_3960, w_022_3961, w_022_3962, w_022_3963, w_022_3964, w_022_3965, w_022_3966, w_022_3967, w_022_3968, w_022_3969, w_022_3971, w_022_3973, w_022_3974, w_022_3976, w_022_3977, w_022_3978, w_022_3979, w_022_3982, w_022_3983, w_022_3984, w_022_3985, w_022_3986, w_022_3988, w_022_3990, w_022_3991, w_022_3992, w_022_3993, w_022_3994, w_022_3995, w_022_3996, w_022_3998, w_022_4000, w_022_4002, w_022_4003, w_022_4004, w_022_4005, w_022_4007, w_022_4010, w_022_4013, w_022_4015, w_022_4017, w_022_4019, w_022_4020, w_022_4021, w_022_4022, w_022_4025, w_022_4026, w_022_4029, w_022_4030, w_022_4031, w_022_4032, w_022_4033, w_022_4035, w_022_4038, w_022_4040, w_022_4041, w_022_4044, w_022_4045, w_022_4046, w_022_4047, w_022_4049, w_022_4050, w_022_4051, w_022_4053, w_022_4056, w_022_4057, w_022_4058, w_022_4059, w_022_4061, w_022_4064, w_022_4066, w_022_4068, w_022_4069, w_022_4070, w_022_4071, w_022_4072, w_022_4076, w_022_4077, w_022_4078, w_022_4079, w_022_4081, w_022_4082, w_022_4083, w_022_4086, w_022_4088, w_022_4089, w_022_4090, w_022_4093, w_022_4094, w_022_4095, w_022_4097, w_022_4099, w_022_4100, w_022_4101, w_022_4102, w_022_4107, w_022_4109, w_022_4111, w_022_4113, w_022_4114, w_022_4116, w_022_4118, w_022_4120, w_022_4121, w_022_4122, w_022_4123, w_022_4124, w_022_4125, w_022_4126, w_022_4128, w_022_4131, w_022_4132, w_022_4134, w_022_4135, w_022_4136, w_022_4137, w_022_4140, w_022_4141, w_022_4146, w_022_4147, w_022_4150, w_022_4151, w_022_4152, w_022_4153, w_022_4155, w_022_4156, w_022_4158, w_022_4159, w_022_4160, w_022_4161, w_022_4162, w_022_4163, w_022_4164, w_022_4165, w_022_4166, w_022_4167, w_022_4170, w_022_4171, w_022_4172, w_022_4173, w_022_4174, w_022_4177, w_022_4178, w_022_4179, w_022_4183, w_022_4184, w_022_4187, w_022_4188, w_022_4190, w_022_4192, w_022_4194, w_022_4195, w_022_4196, w_022_4198, w_022_4199, w_022_4202, w_022_4203, w_022_4207, w_022_4210, w_022_4211, w_022_4212, w_022_4216, w_022_4217, w_022_4221, w_022_4222, w_022_4223, w_022_4224, w_022_4225, w_022_4229, w_022_4230, w_022_4233, w_022_4234, w_022_4235, w_022_4236, w_022_4237, w_022_4238, w_022_4239, w_022_4240, w_022_4241, w_022_4244, w_022_4245, w_022_4247, w_022_4249, w_022_4254, w_022_4257, w_022_4258, w_022_4260, w_022_4261, w_022_4262, w_022_4264, w_022_4266, w_022_4267, w_022_4270, w_022_4271, w_022_4272, w_022_4273, w_022_4275, w_022_4276, w_022_4278, w_022_4279, w_022_4280, w_022_4281, w_022_4282, w_022_4283, w_022_4284, w_022_4286, w_022_4287, w_022_4288, w_022_4289, w_022_4290, w_022_4291, w_022_4293, w_022_4295, w_022_4296, w_022_4297, w_022_4299, w_022_4300, w_022_4301, w_022_4302, w_022_4303, w_022_4304, w_022_4305, w_022_4307, w_022_4308, w_022_4310, w_022_4311, w_022_4312, w_022_4313, w_022_4314, w_022_4315, w_022_4316, w_022_4317, w_022_4318, w_022_4320, w_022_4323, w_022_4324, w_022_4325, w_022_4326, w_022_4327, w_022_4329, w_022_4330, w_022_4333, w_022_4334, w_022_4335, w_022_4336, w_022_4337, w_022_4338, w_022_4339, w_022_4340, w_022_4341, w_022_4347, w_022_4351, w_022_4354, w_022_4355, w_022_4357, w_022_4358, w_022_4359, w_022_4361, w_022_4362, w_022_4363, w_022_4366, w_022_4367, w_022_4370, w_022_4371, w_022_4373, w_022_4376, w_022_4377, w_022_4378, w_022_4379, w_022_4381, w_022_4382, w_022_4385, w_022_4386, w_022_4388, w_022_4390, w_022_4391, w_022_4393, w_022_4397, w_022_4399, w_022_4401, w_022_4402, w_022_4404, w_022_4409, w_022_4410, w_022_4411, w_022_4412, w_022_4413, w_022_4414, w_022_4415, w_022_4417, w_022_4420, w_022_4423, w_022_4425, w_022_4426, w_022_4427, w_022_4428, w_022_4430, w_022_4431, w_022_4434, w_022_4435, w_022_4436, w_022_4437, w_022_4438, w_022_4440, w_022_4442, w_022_4444, w_022_4450, w_022_4451, w_022_4452, w_022_4453, w_022_4454, w_022_4456, w_022_4457, w_022_4460, w_022_4461, w_022_4462, w_022_4463, w_022_4464, w_022_4465, w_022_4466, w_022_4467, w_022_4468, w_022_4469, w_022_4475, w_022_4477, w_022_4478, w_022_4479, w_022_4480, w_022_4481, w_022_4482, w_022_4484, w_022_4485, w_022_4486, w_022_4488, w_022_4490, w_022_4491, w_022_4493, w_022_4497, w_022_4499, w_022_4500, w_022_4501, w_022_4502, w_022_4503, w_022_4505, w_022_4507, w_022_4511, w_022_4512, w_022_4513, w_022_4515, w_022_4516, w_022_4518, w_022_4520, w_022_4522, w_022_4523, w_022_4524, w_022_4527, w_022_4530, w_022_4533, w_022_4535, w_022_4538, w_022_4539, w_022_4540, w_022_4542, w_022_4543, w_022_4544, w_022_4547, w_022_4548, w_022_4549, w_022_4551, w_022_4552, w_022_4555, w_022_4557, w_022_4560, w_022_4561, w_022_4562, w_022_4563, w_022_4565, w_022_4566, w_022_4569, w_022_4570, w_022_4571, w_022_4572, w_022_4573, w_022_4574, w_022_4575, w_022_4577, w_022_4578, w_022_4579, w_022_4582, w_022_4583, w_022_4584, w_022_4585, w_022_4586, w_022_4591, w_022_4592, w_022_4593, w_022_4594, w_022_4595, w_022_4598, w_022_4600, w_022_4602, w_022_4603, w_022_4604, w_022_4605, w_022_4607, w_022_4612, w_022_4613, w_022_4616, w_022_4617, w_022_4619, w_022_4621, w_022_4623, w_022_4624, w_022_4625, w_022_4627, w_022_4628, w_022_4629, w_022_4630, w_022_4631, w_022_4634, w_022_4635, w_022_4639, w_022_4640, w_022_4642, w_022_4643, w_022_4645, w_022_4648, w_022_4649, w_022_4651, w_022_4652, w_022_4653, w_022_4654, w_022_4655, w_022_4656, w_022_4657, w_022_4658, w_022_4661, w_022_4662, w_022_4666, w_022_4667, w_022_4668, w_022_4670, w_022_4671, w_022_4672, w_022_4673, w_022_4674, w_022_4675, w_022_4677, w_022_4678, w_022_4679, w_022_4682, w_022_4683, w_022_4684, w_022_4685, w_022_4686, w_022_4687, w_022_4688, w_022_4690, w_022_4691, w_022_4692, w_022_4693, w_022_4695, w_022_4696, w_022_4697, w_022_4698, w_022_4700, w_022_4702, w_022_4704, w_022_4705, w_022_4706, w_022_4707, w_022_4708, w_022_4712, w_022_4713, w_022_4715, w_022_4716, w_022_4717, w_022_4719, w_022_4721, w_022_4722, w_022_4723, w_022_4724, w_022_4725, w_022_4727, w_022_4728, w_022_4729, w_022_4730, w_022_4732, w_022_4733, w_022_4734, w_022_4736, w_022_4738, w_022_4739, w_022_4746, w_022_4747, w_022_4750, w_022_4752, w_022_4754, w_022_4755, w_022_4756, w_022_4758, w_022_4760, w_022_4762, w_022_4763, w_022_4764, w_022_4765, w_022_4767, w_022_4768, w_022_4769, w_022_4773, w_022_4774, w_022_4775, w_022_4776, w_022_4777, w_022_4778, w_022_4779, w_022_4781, w_022_4782, w_022_4786, w_022_4787, w_022_4789, w_022_4790, w_022_4794, w_022_4795, w_022_4797, w_022_4798, w_022_4799, w_022_4801, w_022_4802, w_022_4805, w_022_4806, w_022_4807, w_022_4808, w_022_4810, w_022_4811, w_022_4812, w_022_4814, w_022_4815, w_022_4816, w_022_4817, w_022_4819, w_022_4820, w_022_4821, w_022_4822, w_022_4824, w_022_4825, w_022_4826, w_022_4827, w_022_4828, w_022_4830, w_022_4831, w_022_4832, w_022_4834, w_022_4835, w_022_4837, w_022_4839, w_022_4840, w_022_4842, w_022_4843, w_022_4846, w_022_4848, w_022_4849, w_022_4850, w_022_4852, w_022_4853, w_022_4854, w_022_4855, w_022_4856, w_022_4860, w_022_4863, w_022_4865, w_022_4867, w_022_4869, w_022_4872, w_022_4873, w_022_4875, w_022_4876, w_022_4877, w_022_4879, w_022_4882, w_022_4883, w_022_4885, w_022_4887, w_022_4889, w_022_4891, w_022_4895, w_022_4898, w_022_4900, w_022_4901, w_022_4902, w_022_4904, w_022_4905, w_022_4906, w_022_4907, w_022_4909, w_022_4910, w_022_4913, w_022_4914, w_022_4916, w_022_4917, w_022_4919, w_022_4920, w_022_4921, w_022_4923, w_022_4924, w_022_4925, w_022_4930, w_022_4932, w_022_4934, w_022_4936, w_022_4938, w_022_4946, w_022_4947, w_022_4948, w_022_4949, w_022_4950, w_022_4951, w_022_4952, w_022_4953, w_022_4959, w_022_4960, w_022_4961, w_022_4964, w_022_4965, w_022_4967, w_022_4968, w_022_4972, w_022_4976, w_022_4978, w_022_4979, w_022_4980, w_022_4981, w_022_4982, w_022_4984, w_022_4985, w_022_4986, w_022_4988, w_022_4990, w_022_4994, w_022_4997, w_022_4998, w_022_4999, w_022_5000, w_022_5001, w_022_5004, w_022_5005, w_022_5007, w_022_5008, w_022_5009, w_022_5010, w_022_5013, w_022_5018, w_022_5020, w_022_5022, w_022_5023, w_022_5024, w_022_5025, w_022_5026, w_022_5027, w_022_5032, w_022_5033, w_022_5034, w_022_5035, w_022_5043, w_022_5044, w_022_5045, w_022_5046, w_022_5047, w_022_5050, w_022_5051, w_022_5055, w_022_5056, w_022_5057, w_022_5058, w_022_5060, w_022_5061, w_022_5062, w_022_5064, w_022_5066, w_022_5067, w_022_5069, w_022_5071, w_022_5072, w_022_5076, w_022_5080, w_022_5082, w_022_5083, w_022_5085, w_022_5086, w_022_5087, w_022_5090, w_022_5094, w_022_5095, w_022_5098, w_022_5099, w_022_5101, w_022_5102, w_022_5103, w_022_5104, w_022_5105, w_022_5108, w_022_5109, w_022_5110, w_022_5113, w_022_5117, w_022_5120, w_022_5121, w_022_5123, w_022_5125, w_022_5127, w_022_5128, w_022_5129, w_022_5130, w_022_5131, w_022_5134, w_022_5135, w_022_5136, w_022_5138, w_022_5139, w_022_5142, w_022_5146, w_022_5147, w_022_5148, w_022_5149, w_022_5151, w_022_5153, w_022_5158, w_022_5161, w_022_5162, w_022_5163, w_022_5165, w_022_5167, w_022_5169, w_022_5170, w_022_5171, w_022_5172, w_022_5173, w_022_5174, w_022_5175, w_022_5178, w_022_5179, w_022_5180, w_022_5181, w_022_5182, w_022_5183, w_022_5184, w_022_5185, w_022_5186, w_022_5187, w_022_5189, w_022_5190, w_022_5191, w_022_5196, w_022_5197, w_022_5199, w_022_5200, w_022_5201, w_022_5202, w_022_5203, w_022_5208, w_022_5209, w_022_5215, w_022_5216, w_022_5217, w_022_5218, w_022_5221, w_022_5223, w_022_5226, w_022_5228, w_022_5230, w_022_5232, w_022_5233, w_022_5235, w_022_5237, w_022_5239, w_022_5241, w_022_5242, w_022_5246, w_022_5248, w_022_5249, w_022_5251, w_022_5252, w_022_5253, w_022_5254, w_022_5259, w_022_5260, w_022_5261, w_022_5268, w_022_5273, w_022_5274, w_022_5275, w_022_5276, w_022_5279, w_022_5280, w_022_5281, w_022_5284, w_022_5285, w_022_5287, w_022_5289, w_022_5294, w_022_5297, w_022_5299, w_022_5300, w_022_5301, w_022_5303, w_022_5305, w_022_5309, w_022_5311, w_022_5312, w_022_5313, w_022_5316, w_022_5317, w_022_5319, w_022_5322, w_022_5323, w_022_5326, w_022_5329, w_022_5330, w_022_5331, w_022_5332, w_022_5334, w_022_5335, w_022_5336, w_022_5337, w_022_5340, w_022_5342, w_022_5345, w_022_5347, w_022_5349, w_022_5350, w_022_5352, w_022_5354, w_022_5357, w_022_5360, w_022_5362, w_022_5364, w_022_5367, w_022_5369, w_022_5372, w_022_5373, w_022_5374, w_022_5375, w_022_5377, w_022_5378, w_022_5381, w_022_5382, w_022_5383, w_022_5385, w_022_5388, w_022_5392, w_022_5393, w_022_5396, w_022_5398, w_022_5399, w_022_5400, w_022_5401, w_022_5402, w_022_5403, w_022_5404, w_022_5405, w_022_5406, w_022_5408, w_022_5409, w_022_5410, w_022_5411, w_022_5412, w_022_5413, w_022_5416, w_022_5417, w_022_5418, w_022_5419, w_022_5420, w_022_5422, w_022_5423, w_022_5426, w_022_5429, w_022_5430, w_022_5432, w_022_5435, w_022_5436, w_022_5439, w_022_5442, w_022_5443, w_022_5444, w_022_5445, w_022_5447, w_022_5452, w_022_5453, w_022_5454, w_022_5455, w_022_5458, w_022_5460, w_022_5461, w_022_5462, w_022_5464, w_022_5465, w_022_5466, w_022_5467, w_022_5468, w_022_5469, w_022_5470, w_022_5471, w_022_5472, w_022_5473, w_022_5474, w_022_5478, w_022_5479, w_022_5480, w_022_5483, w_022_5484, w_022_5485, w_022_5486, w_022_5487, w_022_5488, w_022_5489, w_022_5490, w_022_5491, w_022_5492, w_022_5496, w_022_5497, w_022_5498, w_022_5499, w_022_5503, w_022_5504, w_022_5505, w_022_5506, w_022_5507, w_022_5509, w_022_5514, w_022_5515, w_022_5516, w_022_5517, w_022_5518, w_022_5520, w_022_5522, w_022_5523, w_022_5524, w_022_5526, w_022_5531, w_022_5532, w_022_5533, w_022_5536, w_022_5538, w_022_5539, w_022_5540, w_022_5542, w_022_5544, w_022_5545, w_022_5546, w_022_5547, w_022_5548, w_022_5550, w_022_5551, w_022_5553, w_022_5554, w_022_5555, w_022_5556, w_022_5557, w_022_5559, w_022_5560, w_022_5561, w_022_5562, w_022_5563, w_022_5564, w_022_5565, w_022_5566, w_022_5567, w_022_5569, w_022_5571, w_022_5572, w_022_5573, w_022_5575, w_022_5576, w_022_5577, w_022_5579, w_022_5582, w_022_5586, w_022_5589, w_022_5591, w_022_5593, w_022_5595, w_022_5596, w_022_5598, w_022_5599, w_022_5603, w_022_5604, w_022_5611, w_022_5612, w_022_5613, w_022_5614, w_022_5615, w_022_5616, w_022_5617, w_022_5618, w_022_5619, w_022_5620, w_022_5621, w_022_5624, w_022_5625, w_022_5627, w_022_5628, w_022_5629, w_022_5630, w_022_5631, w_022_5632, w_022_5633, w_022_5634, w_022_5635, w_022_5636, w_022_5640, w_022_5641, w_022_5646, w_022_5647, w_022_5648, w_022_5649, w_022_5655, w_022_5656, w_022_5657, w_022_5658, w_022_5660, w_022_5662, w_022_5663, w_022_5666, w_022_5667, w_022_5668, w_022_5669, w_022_5671, w_022_5674, w_022_5675, w_022_5676, w_022_5679, w_022_5681, w_022_5682, w_022_5683, w_022_5685, w_022_5686, w_022_5687, w_022_5688, w_022_5690, w_022_5691, w_022_5692, w_022_5693, w_022_5696, w_022_5699, w_022_5700, w_022_5701, w_022_5703, w_022_5705, w_022_5706, w_022_5709, w_022_5710, w_022_5713, w_022_5714, w_022_5715, w_022_5717, w_022_5720, w_022_5721, w_022_5723, w_022_5724, w_022_5725, w_022_5726, w_022_5729, w_022_5730, w_022_5732, w_022_5733, w_022_5734, w_022_5735, w_022_5736, w_022_5737, w_022_5738, w_022_5739, w_022_5740, w_022_5741, w_022_5743, w_022_5744, w_022_5748, w_022_5751, w_022_5752, w_022_5754, w_022_5756, w_022_5757, w_022_5761, w_022_5762, w_022_5764, w_022_5765, w_022_5766, w_022_5767, w_022_5769, w_022_5770, w_022_5774, w_022_5775, w_022_5777, w_022_5780, w_022_5781, w_022_5784, w_022_5788, w_022_5790, w_022_5793, w_022_5794, w_022_5795, w_022_5797, w_022_5798, w_022_5799, w_022_5801, w_022_5802, w_022_5803, w_022_5804, w_022_5805, w_022_5807, w_022_5810, w_022_5811, w_022_5812, w_022_5814, w_022_5816, w_022_5817, w_022_5818, w_022_5820, w_022_5821, w_022_5824, w_022_5826, w_022_5827, w_022_5828, w_022_5829, w_022_5830, w_022_5832, w_022_5833, w_022_5834, w_022_5835, w_022_5836, w_022_5837, w_022_5838, w_022_5840, w_022_5843, w_022_5846, w_022_5847, w_022_5848, w_022_5851, w_022_5854, w_022_5858, w_022_5859, w_022_5862, w_022_5865, w_022_5867, w_022_5868, w_022_5869, w_022_5870, w_022_5871, w_022_5872, w_022_5873, w_022_5874, w_022_5875, w_022_5878, w_022_5879, w_022_5880, w_022_5881, w_022_5882, w_022_5883, w_022_5885, w_022_5886, w_022_5888, w_022_5889, w_022_5890, w_022_5891, w_022_5892, w_022_5893, w_022_5897, w_022_5898, w_022_5899, w_022_5901, w_022_5902, w_022_5903, w_022_5904, w_022_5905, w_022_5907, w_022_5908, w_022_5909, w_022_5910, w_022_5914, w_022_5917, w_022_5921, w_022_5922, w_022_5923, w_022_5925, w_022_5926, w_022_5931, w_022_5932, w_022_5933, w_022_5937, w_022_5938, w_022_5940, w_022_5943, w_022_5944, w_022_5945, w_022_5946, w_022_5949, w_022_5954, w_022_5956, w_022_5958, w_022_5959, w_022_5960, w_022_5961, w_022_5962, w_022_5963, w_022_5965, w_022_5967, w_022_5969, w_022_5971, w_022_5972, w_022_5973, w_022_5974, w_022_5975, w_022_5977, w_022_5978, w_022_5979, w_022_5980, w_022_5981, w_022_5982, w_022_5984, w_022_5985, w_022_5988, w_022_5993, w_022_5996, w_022_5997, w_022_6000, w_022_6001, w_022_6003, w_022_6005, w_022_6008, w_022_6009, w_022_6010, w_022_6011, w_022_6012, w_022_6013, w_022_6014, w_022_6015, w_022_6016, w_022_6017, w_022_6022, w_022_6024, w_022_6027, w_022_6028, w_022_6029, w_022_6031, w_022_6034, w_022_6035, w_022_6036, w_022_6037, w_022_6038, w_022_6039, w_022_6040, w_022_6041, w_022_6043, w_022_6044, w_022_6046, w_022_6047, w_022_6048, w_022_6049, w_022_6051, w_022_6052, w_022_6054, w_022_6056, w_022_6057, w_022_6058, w_022_6059, w_022_6060, w_022_6064, w_022_6065, w_022_6066, w_022_6067, w_022_6069, w_022_6071, w_022_6075, w_022_6076, w_022_6077, w_022_6078, w_022_6079, w_022_6080, w_022_6082, w_022_6086, w_022_6087, w_022_6088, w_022_6089, w_022_6090, w_022_6091, w_022_6092, w_022_6093, w_022_6094, w_022_6097, w_022_6098, w_022_6099, w_022_6100, w_022_6101, w_022_6104, w_022_6107, w_022_6108, w_022_6109, w_022_6113, w_022_6114, w_022_6115, w_022_6116, w_022_6117, w_022_6119, w_022_6121, w_022_6122, w_022_6123, w_022_6124, w_022_6127, w_022_6128, w_022_6130, w_022_6133, w_022_6134, w_022_6135, w_022_6136, w_022_6137, w_022_6139, w_022_6141, w_022_6142, w_022_6143, w_022_6144, w_022_6145, w_022_6150, w_022_6152, w_022_6155, w_022_6159, w_022_6160, w_022_6161, w_022_6162, w_022_6163, w_022_6165, w_022_6167, w_022_6168, w_022_6169, w_022_6171, w_022_6172, w_022_6173, w_022_6175, w_022_6177, w_022_6178, w_022_6180, w_022_6181, w_022_6182, w_022_6185, w_022_6187, w_022_6188, w_022_6192, w_022_6194, w_022_6195, w_022_6197, w_022_6200, w_022_6202, w_022_6204, w_022_6205, w_022_6206, w_022_6207, w_022_6209, w_022_6210, w_022_6213, w_022_6214, w_022_6216, w_022_6217, w_022_6219, w_022_6220, w_022_6222, w_022_6223, w_022_6225, w_022_6226, w_022_6227, w_022_6230, w_022_6231, w_022_6232, w_022_6233, w_022_6235, w_022_6236, w_022_6238, w_022_6240, w_022_6242, w_022_6244, w_022_6245, w_022_6246, w_022_6248, w_022_6249, w_022_6250, w_022_6252, w_022_6253, w_022_6255, w_022_6256, w_022_6258, w_022_6263, w_022_6264, w_022_6265, w_022_6267, w_022_6270, w_022_6271, w_022_6272, w_022_6273, w_022_6274, w_022_6278, w_022_6279, w_022_6280, w_022_6282, w_022_6284, w_022_6290, w_022_6291, w_022_6292, w_022_6293, w_022_6295, w_022_6297, w_022_6299, w_022_6300, w_022_6301, w_022_6302, w_022_6303, w_022_6304, w_022_6306, w_022_6309, w_022_6311, w_022_6313, w_022_6315, w_022_6317, w_022_6319, w_022_6320, w_022_6321, w_022_6322, w_022_6323, w_022_6325, w_022_6326, w_022_6327, w_022_6330, w_022_6331, w_022_6333, w_022_6336, w_022_6337, w_022_6345, w_022_6348, w_022_6349, w_022_6352, w_022_6355, w_022_6356, w_022_6360, w_022_6363, w_022_6364, w_022_6365, w_022_6367, w_022_6369, w_022_6370, w_022_6371, w_022_6373, w_022_6374, w_022_6375, w_022_6376, w_022_6379, w_022_6380, w_022_6381, w_022_6382, w_022_6383, w_022_6385, w_022_6389, w_022_6390, w_022_6391, w_022_6395, w_022_6396, w_022_6397, w_022_6398, w_022_6403, w_022_6404, w_022_6406, w_022_6408, w_022_6409, w_022_6413, w_022_6417, w_022_6424, w_022_6425, w_022_6426, w_022_6427, w_022_6429, w_022_6430, w_022_6431, w_022_6432, w_022_6433, w_022_6434, w_022_6436, w_022_6437, w_022_6438, w_022_6439, w_022_6440, w_022_6446, w_022_6447, w_022_6448, w_022_6449, w_022_6451, w_022_6452, w_022_6453, w_022_6454, w_022_6455, w_022_6456, w_022_6459, w_022_6461, w_022_6462, w_022_6463, w_022_6464, w_022_6465, w_022_6466, w_022_6467, w_022_6468, w_022_6470, w_022_6471, w_022_6473, w_022_6475, w_022_6476, w_022_6477, w_022_6479, w_022_6482, w_022_6483, w_022_6484, w_022_6485, w_022_6486, w_022_6487, w_022_6488, w_022_6489, w_022_6494, w_022_6495, w_022_6497, w_022_6498, w_022_6499, w_022_6500, w_022_6501, w_022_6502, w_022_6503, w_022_6504, w_022_6508, w_022_6509, w_022_6510, w_022_6511, w_022_6514, w_022_6515, w_022_6516, w_022_6517, w_022_6518, w_022_6520, w_022_6521, w_022_6522, w_022_6523, w_022_6524, w_022_6525, w_022_6526, w_022_6528, w_022_6530, w_022_6531, w_022_6532, w_022_6533, w_022_6534, w_022_6538, w_022_6541, w_022_6542, w_022_6544, w_022_6546, w_022_6553, w_022_6554, w_022_6556, w_022_6557, w_022_6558, w_022_6559, w_022_6560, w_022_6562, w_022_6563, w_022_6566, w_022_6569, w_022_6572, w_022_6573, w_022_6574, w_022_6575, w_022_6578, w_022_6579, w_022_6580, w_022_6581, w_022_6582, w_022_6583, w_022_6586, w_022_6587, w_022_6588, w_022_6589, w_022_6590, w_022_6591, w_022_6594, w_022_6596, w_022_6597, w_022_6599, w_022_6601, w_022_6605, w_022_6606, w_022_6609, w_022_6611, w_022_6612, w_022_6613, w_022_6615, w_022_6616, w_022_6617, w_022_6618, w_022_6624, w_022_6625, w_022_6626, w_022_6630, w_022_6631, w_022_6632, w_022_6633, w_022_6635, w_022_6638, w_022_6642, w_022_6643, w_022_6644, w_022_6645, w_022_6646, w_022_6647, w_022_6650, w_022_6652, w_022_6654, w_022_6655, w_022_6656, w_022_6659, w_022_6660, w_022_6661, w_022_6662, w_022_6665, w_022_6668, w_022_6669, w_022_6671, w_022_6672, w_022_6674, w_022_6675, w_022_6677, w_022_6679, w_022_6680, w_022_6683, w_022_6684, w_022_6685, w_022_6687, w_022_6692, w_022_6693, w_022_6694, w_022_6695, w_022_6698, w_022_6699, w_022_6700, w_022_6703, w_022_6704, w_022_6705, w_022_6707, w_022_6711, w_022_6712, w_022_6713, w_022_6714, w_022_6715, w_022_6717, w_022_6718, w_022_6719, w_022_6721, w_022_6723, w_022_6727, w_022_6730, w_022_6731, w_022_6734, w_022_6735, w_022_6736, w_022_6737, w_022_6739, w_022_6740, w_022_6741, w_022_6742, w_022_6750, w_022_6752, w_022_6753, w_022_6755, w_022_6761, w_022_6762, w_022_6763, w_022_6765, w_022_6766, w_022_6767, w_022_6768, w_022_6770, w_022_6771, w_022_6773, w_022_6775, w_022_6776, w_022_6778, w_022_6779, w_022_6785, w_022_6786, w_022_6787, w_022_6789, w_022_6791, w_022_6793, w_022_6794, w_022_6797, w_022_6798, w_022_6799, w_022_6800, w_022_6803, w_022_6805, w_022_6806, w_022_6807, w_022_6809, w_022_6811, w_022_6813, w_022_6814, w_022_6816, w_022_6817, w_022_6818, w_022_6819, w_022_6820, w_022_6821, w_022_6822, w_022_6824, w_022_6827, w_022_6828, w_022_6829, w_022_6830, w_022_6831, w_022_6832, w_022_6833, w_022_6834, w_022_6835, w_022_6836, w_022_6843, w_022_6845, w_022_6846, w_022_6848, w_022_6849, w_022_6850, w_022_6851, w_022_6852, w_022_6854, w_022_6855, w_022_6856, w_022_6857, w_022_6858, w_022_6860, w_022_6861, w_022_6863, w_022_6864, w_022_6866, w_022_6868, w_022_6869, w_022_6871, w_022_6872, w_022_6874, w_022_6875, w_022_6876, w_022_6877, w_022_6878, w_022_6879, w_022_6880, w_022_6881, w_022_6884, w_022_6885, w_022_6887, w_022_6888, w_022_6892, w_022_6893, w_022_6894, w_022_6895, w_022_6898, w_022_6901, w_022_6903, w_022_6904, w_022_6905, w_022_6906, w_022_6907, w_022_6908, w_022_6909, w_022_6910, w_022_6911, w_022_6912, w_022_6913, w_022_6914, w_022_6916, w_022_6920, w_022_6923, w_022_6924, w_022_6925, w_022_6927, w_022_6928, w_022_6929, w_022_6931, w_022_6932, w_022_6933, w_022_6934, w_022_6935, w_022_6936, w_022_6937, w_022_6939, w_022_6942, w_022_6944, w_022_6947, w_022_6948, w_022_6950, w_022_6951, w_022_6952, w_022_6953, w_022_6954, w_022_6955, w_022_6957, w_022_6958, w_022_6959, w_022_6960, w_022_6961, w_022_6962, w_022_6963, w_022_6966, w_022_6968, w_022_6970, w_022_6971, w_022_6972, w_022_6973, w_022_6974, w_022_6976, w_022_6977, w_022_6978, w_022_6980, w_022_6981, w_022_6982, w_022_6984, w_022_6985, w_022_6987, w_022_6988, w_022_6990, w_022_6991, w_022_6993, w_022_6995, w_022_6996, w_022_6997, w_022_6998, w_022_7001, w_022_7002, w_022_7003, w_022_7005, w_022_7009, w_022_7010, w_022_7011, w_022_7012, w_022_7013, w_022_7014, w_022_7015, w_022_7018, w_022_7021, w_022_7022, w_022_7023, w_022_7024, w_022_7025, w_022_7026, w_022_7027, w_022_7028, w_022_7029, w_022_7030, w_022_7031, w_022_7032, w_022_7035, w_022_7036, w_022_7037, w_022_7038, w_022_7041, w_022_7042, w_022_7043, w_022_7045, w_022_7049, w_022_7050, w_022_7052, w_022_7053, w_022_7054, w_022_7056, w_022_7057, w_022_7060, w_022_7061, w_022_7062, w_022_7063, w_022_7064, w_022_7065, w_022_7067, w_022_7071, w_022_7072, w_022_7073, w_022_7074, w_022_7077, w_022_7078, w_022_7082, w_022_7086, w_022_7090, w_022_7091, w_022_7095, w_022_7096, w_022_7098, w_022_7099, w_022_7104, w_022_7105, w_022_7106, w_022_7107, w_022_7110, w_022_7111, w_022_7112, w_022_7114, w_022_7116, w_022_7117, w_022_7118, w_022_7120, w_022_7121, w_022_7122, w_022_7123, w_022_7124, w_022_7128, w_022_7129, w_022_7133, w_022_7134, w_022_7135, w_022_7138, w_022_7139, w_022_7140, w_022_7142, w_022_7143, w_022_7145, w_022_7146, w_022_7148, w_022_7154, w_022_7155, w_022_7156, w_022_7157, w_022_7158, w_022_7162, w_022_7165, w_022_7167, w_022_7168, w_022_7172, w_022_7173, w_022_7174, w_022_7175, w_022_7178, w_022_7182, w_022_7183, w_022_7187, w_022_7188, w_022_7190, w_022_7195, w_022_7196, w_022_7197, w_022_7198, w_022_7200, w_022_7201, w_022_7202, w_022_7204, w_022_7208, w_022_7209, w_022_7211, w_022_7212, w_022_7213, w_022_7216, w_022_7218, w_022_7219, w_022_7220, w_022_7221, w_022_7222, w_022_7223, w_022_7224, w_022_7225, w_022_7226, w_022_7228, w_022_7229, w_022_7232, w_022_7233, w_022_7237, w_022_7241, w_022_7243, w_022_7245, w_022_7247, w_022_7248, w_022_7249, w_022_7251, w_022_7253, w_022_7257, w_022_7259, w_022_7260, w_022_7261, w_022_7266, w_022_7267, w_022_7268, w_022_7269, w_022_7270, w_022_7271, w_022_7272, w_022_7273, w_022_7275, w_022_7277, w_022_7278, w_022_7279, w_022_7281, w_022_7282, w_022_7287, w_022_7288, w_022_7289, w_022_7291, w_022_7292, w_022_7293, w_022_7296, w_022_7297, w_022_7299, w_022_7301, w_022_7303, w_022_7306, w_022_7307, w_022_7309, w_022_7312, w_022_7314, w_022_7315, w_022_7316, w_022_7317, w_022_7320, w_022_7324, w_022_7325, w_022_7326, w_022_7328, w_022_7329, w_022_7333, w_022_7334, w_022_7335, w_022_7336, w_022_7337, w_022_7338, w_022_7340, w_022_7341, w_022_7342, w_022_7343, w_022_7344, w_022_7345, w_022_7346, w_022_7347, w_022_7348, w_022_7349, w_022_7351, w_022_7353, w_022_7354, w_022_7356, w_022_7357, w_022_7359, w_022_7360, w_022_7362, w_022_7364, w_022_7366, w_022_7370, w_022_7373, w_022_7374, w_022_7376, w_022_7378, w_022_7379, w_022_7382, w_022_7383, w_022_7387, w_022_7390, w_022_7392, w_022_7393, w_022_7395, w_022_7399, w_022_7400, w_022_7401, w_022_7402, w_022_7403, w_022_7405, w_022_7408, w_022_7409, w_022_7410, w_022_7411, w_022_7412, w_022_7413, w_022_7415, w_022_7418, w_022_7419, w_022_7420, w_022_7423, w_022_7425, w_022_7426, w_022_7427, w_022_7428, w_022_7429, w_022_7430, w_022_7432, w_022_7433, w_022_7434, w_022_7435, w_022_7436, w_022_7437, w_022_7438, w_022_7440, w_022_7441, w_022_7442, w_022_7444, w_022_7447, w_022_7448, w_022_7449, w_022_7452, w_022_7454, w_022_7458, w_022_7461, w_022_7463, w_022_7464, w_022_7465, w_022_7467, w_022_7468, w_022_7469, w_022_7470, w_022_7471, w_022_7473, w_022_7474, w_022_7475, w_022_7476, w_022_7479, w_022_7480, w_022_7482, w_022_7483, w_022_7485, w_022_7487, w_022_7488, w_022_7489, w_022_7490, w_022_7491, w_022_7492, w_022_7494, w_022_7495, w_022_7497, w_022_7498, w_022_7501, w_022_7502, w_022_7503, w_022_7504, w_022_7505, w_022_7508, w_022_7509, w_022_7510, w_022_7511, w_022_7512, w_022_7513, w_022_7514, w_022_7515, w_022_7516, w_022_7518, w_022_7519, w_022_7520, w_022_7521, w_022_7524, w_022_7527, w_022_7528, w_022_7530, w_022_7531, w_022_7536, w_022_7537, w_022_7538, w_022_7539, w_022_7540, w_022_7541, w_022_7543, w_022_7544, w_022_7545, w_022_7547, w_022_7550, w_022_7551, w_022_7553, w_022_7554, w_022_7556, w_022_7557, w_022_7558, w_022_7559, w_022_7560, w_022_7562, w_022_7565, w_022_7567, w_022_7568, w_022_7569, w_022_7570, w_022_7571, w_022_7575, w_022_7577, w_022_7578, w_022_7580, w_022_7581, w_022_7582, w_022_7584, w_022_7586, w_022_7587, w_022_7588, w_022_7589, w_022_7591, w_022_7592, w_022_7593, w_022_7595, w_022_7597, w_022_7599, w_022_7601, w_022_7602, w_022_7603, w_022_7604, w_022_7606, w_022_7607, w_022_7608, w_022_7609, w_022_7610, w_022_7612, w_022_7614, w_022_7617, w_022_7618, w_022_7619, w_022_7620, w_022_7622, w_022_7623, w_022_7624, w_022_7628, w_022_7632, w_022_7635, w_022_7636, w_022_7637, w_022_7639, w_022_7641, w_022_7644, w_022_7646, w_022_7648, w_022_7649, w_022_7650, w_022_7652, w_022_7654, w_022_7655, w_022_7656, w_022_7657, w_022_7658, w_022_7661, w_022_7662, w_022_7664, w_022_7666, w_022_7667, w_022_7669, w_022_7671, w_022_7672, w_022_7674, w_022_7675, w_022_7677, w_022_7678, w_022_7679, w_022_7681, w_022_7683, w_022_7684, w_022_7687, w_022_7690, w_022_7691, w_022_7694, w_022_7695, w_022_7696, w_022_7697, w_022_7699, w_022_7700, w_022_7701, w_022_7706, w_022_7707, w_022_7709, w_022_7710, w_022_7711, w_022_7713, w_022_7714, w_022_7715, w_022_7716, w_022_7717, w_022_7720, w_022_7721, w_022_7722, w_022_7723, w_022_7724, w_022_7726, w_022_7727, w_022_7729, w_022_7734, w_022_7735, w_022_7740, w_022_7742, w_022_7743, w_022_7745, w_022_7746, w_022_7747, w_022_7748, w_022_7749, w_022_7750, w_022_7751, w_022_7752, w_022_7753, w_022_7755, w_022_7756, w_022_7758, w_022_7759, w_022_7760, w_022_7761, w_022_7763, w_022_7765, w_022_7766, w_022_7768, w_022_7769, w_022_7770, w_022_7771, w_022_7773, w_022_7775, w_022_7777, w_022_7780, w_022_7781, w_022_7783, w_022_7785, w_022_7786, w_022_7787, w_022_7790, w_022_7791, w_022_7799, w_022_7801, w_022_7803, w_022_7805, w_022_7807, w_022_7808, w_022_7810, w_022_7811, w_022_7813, w_022_7815, w_022_7819, w_022_7821, w_022_7822, w_022_7824, w_022_7826, w_022_7827, w_022_7829, w_022_7831, w_022_7835, w_022_7837, w_022_7838, w_022_7839, w_022_7840, w_022_7842, w_022_7844, w_022_7846, w_022_7847, w_022_7848, w_022_7855, w_022_7858, w_022_7863, w_022_7865, w_022_7866, w_022_7867, w_022_7869, w_022_7871, w_022_7874, w_022_7876, w_022_7877, w_022_7879, w_022_7880, w_022_7881, w_022_7884, w_022_7885, w_022_7886, w_022_7887, w_022_7888, w_022_7890, w_022_7891, w_022_7892, w_022_7894, w_022_7898, w_022_7899, w_022_7900, w_022_7901, w_022_7908, w_022_7909, w_022_7910, w_022_7912, w_022_7915, w_022_7916, w_022_7917, w_022_7918, w_022_7919, w_022_7922, w_022_7923, w_022_7925, w_022_7926, w_022_7927, w_022_7928, w_022_7930, w_022_7932, w_022_7933, w_022_7934, w_022_7938, w_022_7939, w_022_7940, w_022_7944, w_022_7945, w_022_7946, w_022_7947, w_022_7948, w_022_7949, w_022_7950, w_022_7951, w_022_7952, w_022_7955, w_022_7956, w_022_7957, w_022_7960, w_022_7963, w_022_7964, w_022_7970, w_022_7971, w_022_7976, w_022_7977, w_022_7978, w_022_7979, w_022_7980, w_022_7983, w_022_7984, w_022_7988, w_022_7989, w_022_7990, w_022_7991, w_022_7992, w_022_7993, w_022_7995, w_022_7996, w_022_7997, w_022_7999, w_022_8000, w_022_8001, w_022_8002, w_022_8003, w_022_8004, w_022_8006, w_022_8007, w_022_8008, w_022_8011, w_022_8013, w_022_8015, w_022_8017, w_022_8018, w_022_8019, w_022_8020, w_022_8021, w_022_8023, w_022_8025, w_022_8027, w_022_8028, w_022_8029, w_022_8031, w_022_8033, w_022_8034, w_022_8036, w_022_8037, w_022_8038, w_022_8039, w_022_8040, w_022_8042, w_022_8043, w_022_8045, w_022_8048, w_022_8052, w_022_8053, w_022_8054, w_022_8055, w_022_8056, w_022_8057, w_022_8058, w_022_8059, w_022_8063, w_022_8064, w_022_8066, w_022_8068, w_022_8069, w_022_8071, w_022_8072, w_022_8073, w_022_8075, w_022_8077, w_022_8078, w_022_8079, w_022_8080, w_022_8081, w_022_8083, w_022_8086, w_022_8089, w_022_8092, w_022_8094, w_022_8095, w_022_8096, w_022_8098, w_022_8099, w_022_8103, w_022_8105, w_022_8107, w_022_8109, w_022_8110, w_022_8116, w_022_8117, w_022_8120, w_022_8122, w_022_8126, w_022_8127, w_022_8128, w_022_8131, w_022_8132, w_022_8136, w_022_8138, w_022_8139, w_022_8140, w_022_8147, w_022_8148, w_022_8149, w_022_8150, w_022_8152, w_022_8153, w_022_8154, w_022_8157, w_022_8158, w_022_8160, w_022_8161, w_022_8163, w_022_8164, w_022_8167, w_022_8168, w_022_8170, w_022_8171, w_022_8174, w_022_8175, w_022_8176, w_022_8177, w_022_8180, w_022_8181, w_022_8184, w_022_8185, w_022_8189, w_022_8190, w_022_8191, w_022_8193, w_022_8195, w_022_8196, w_022_8197, w_022_8199, w_022_8201, w_022_8202, w_022_8205, w_022_8208, w_022_8211, w_022_8212, w_022_8215, w_022_8216, w_022_8217, w_022_8218, w_022_8219, w_022_8220, w_022_8224, w_022_8226, w_022_8228, w_022_8229, w_022_8232, w_022_8233, w_022_8234, w_022_8237, w_022_8238, w_022_8239, w_022_8240, w_022_8241, w_022_8244, w_022_8245, w_022_8247, w_022_8248, w_022_8249, w_022_8250, w_022_8251, w_022_8252, w_022_8254, w_022_8255, w_022_8257, w_022_8258, w_022_8259, w_022_8261, w_022_8263, w_022_8264, w_022_8265, w_022_8266, w_022_8267, w_022_8269, w_022_8270, w_022_8272, w_022_8273, w_022_8274, w_022_8275, w_022_8276, w_022_8284, w_022_8286, w_022_8288, w_022_8290, w_022_8291, w_022_8292, w_022_8293, w_022_8294, w_022_8295, w_022_8297, w_022_8298, w_022_8300, w_022_8301, w_022_8305, w_022_8310, w_022_8311, w_022_8312, w_022_8314, w_022_8316, w_022_8317, w_022_8318, w_022_8319, w_022_8320, w_022_8321, w_022_8323, w_022_8324, w_022_8325, w_022_8326, w_022_8327, w_022_8329, w_022_8330, w_022_8332, w_022_8333, w_022_8335, w_022_8336, w_022_8337, w_022_8338, w_022_8340, w_022_8342, w_022_8345, w_022_8346, w_022_8347, w_022_8348, w_022_8349, w_022_8350, w_022_8351, w_022_8352, w_022_8353, w_022_8354, w_022_8355, w_022_8356, w_022_8360, w_022_8361, w_022_8362, w_022_8363, w_022_8364, w_022_8365, w_022_8366, w_022_8367, w_022_8369, w_022_8370, w_022_8371, w_022_8373, w_022_8374, w_022_8375, w_022_8377, w_022_8379, w_022_8381, w_022_8382, w_022_8384, w_022_8385, w_022_8387, w_022_8389, w_022_8391, w_022_8392, w_022_8394, w_022_8395, w_022_8398, w_022_8399, w_022_8400, w_022_8402, w_022_8404, w_022_8405, w_022_8407, w_022_8408, w_022_8410, w_022_8412, w_022_8413, w_022_8414, w_022_8415, w_022_8418, w_022_8420, w_022_8423, w_022_8424, w_022_8425, w_022_8427, w_022_8429, w_022_8430, w_022_8431, w_022_8435, w_022_8436, w_022_8437, w_022_8440, w_022_8442, w_022_8444, w_022_8445, w_022_8447, w_022_8448, w_022_8450, w_022_8454, w_022_8455, w_022_8457, w_022_8458, w_022_8461, w_022_8464, w_022_8468, w_022_8469, w_022_8471, w_022_8472, w_022_8473, w_022_8474, w_022_8475, w_022_8476, w_022_8477, w_022_8479, w_022_8480, w_022_8483, w_022_8484, w_022_8486, w_022_8487, w_022_8489, w_022_8491, w_022_8492, w_022_8493, w_022_8495, w_022_8496, w_022_8499, w_022_8500, w_022_8504, w_022_8506, w_022_8509, w_022_8513, w_022_8514, w_022_8517, w_022_8518, w_022_8519, w_022_8521, w_022_8524, w_022_8525, w_022_8526, w_022_8527, w_022_8528, w_022_8529, w_022_8530, w_022_8531, w_022_8533, w_022_8537, w_022_8539, w_022_8540, w_022_8542, w_022_8545, w_022_8546, w_022_8547, w_022_8548, w_022_8550, w_022_8551, w_022_8552, w_022_8553, w_022_8555, w_022_8556, w_022_8557, w_022_8559, w_022_8560, w_022_8561, w_022_8562, w_022_8564, w_022_8567, w_022_8568, w_022_8572, w_022_8575, w_022_8576, w_022_8577, w_022_8578, w_022_8579, w_022_8581, w_022_8582, w_022_8585, w_022_8589, w_022_8590, w_022_8591, w_022_8594, w_022_8595, w_022_8596, w_022_8597, w_022_8598, w_022_8599, w_022_8600, w_022_8602, w_022_8604, w_022_8605, w_022_8610, w_022_8613, w_022_8614, w_022_8615, w_022_8617, w_022_8619, w_022_8620, w_022_8621, w_022_8624, w_022_8627, w_022_8629, w_022_8630, w_022_8632, w_022_8633, w_022_8634, w_022_8635, w_022_8636, w_022_8637, w_022_8643, w_022_8644, w_022_8645, w_022_8650, w_022_8651, w_022_8652, w_022_8653, w_022_8654, w_022_8656, w_022_8658, w_022_8662, w_022_8663, w_022_8664, w_022_8665, w_022_8666, w_022_8667, w_022_8672, w_022_8674, w_022_8677, w_022_8678, w_022_8679, w_022_8681, w_022_8683, w_022_8685, w_022_8686, w_022_8687, w_022_8688, w_022_8689, w_022_8690, w_022_8691, w_022_8692, w_022_8693, w_022_8694, w_022_8695, w_022_8696, w_022_8699, w_022_8703, w_022_8705, w_022_8706, w_022_8707, w_022_8708, w_022_8709, w_022_8710, w_022_8712, w_022_8713, w_022_8715, w_022_8717, w_022_8718, w_022_8722, w_022_8727, w_022_8728, w_022_8729, w_022_8731, w_022_8734, w_022_8735, w_022_8736, w_022_8737, w_022_8740, w_022_8742, w_022_8743, w_022_8744, w_022_8745, w_022_8747, w_022_8748, w_022_8750, w_022_8751, w_022_8752, w_022_8754, w_022_8755, w_022_8756, w_022_8757, w_022_8758, w_022_8759, w_022_8761, w_022_8762, w_022_8765, w_022_8766, w_022_8767, w_022_8769, w_022_8770, w_022_8771, w_022_8773, w_022_8774, w_022_8775, w_022_8776, w_022_8777, w_022_8778, w_022_8779, w_022_8780, w_022_8781, w_022_8782, w_022_8783, w_022_8784, w_022_8787, w_022_8788, w_022_8789, w_022_8791, w_022_8792, w_022_8793, w_022_8794, w_022_8798, w_022_8799, w_022_8800, w_022_8801, w_022_8802, w_022_8803, w_022_8805, w_022_8806, w_022_8807, w_022_8808, w_022_8809, w_022_8810, w_022_8812, w_022_8813, w_022_8814, w_022_8815, w_022_8816, w_022_8820, w_022_8822, w_022_8824, w_022_8825, w_022_8826, w_022_8829, w_022_8830, w_022_8831, w_022_8834, w_022_8835, w_022_8840, w_022_8841, w_022_8842, w_022_8843, w_022_8844, w_022_8845, w_022_8847, w_022_8848, w_022_8857, w_022_8859, w_022_8861, w_022_8864, w_022_8865, w_022_8866, w_022_8868, w_022_8869, w_022_8870, w_022_8871, w_022_8876, w_022_8877, w_022_8878, w_022_8880, w_022_8881, w_022_8882, w_022_8883, w_022_8884, w_022_8886, w_022_8890, w_022_8891, w_022_8892, w_022_8893, w_022_8896, w_022_8897, w_022_8898, w_022_8899, w_022_8901, w_022_8902, w_022_8904, w_022_8905, w_022_8907, w_022_8910, w_022_8911, w_022_8913, w_022_8914, w_022_8915, w_022_8916, w_022_8920, w_022_8923, w_022_8924, w_022_8928, w_022_8929, w_022_8930, w_022_8933, w_022_8935, w_022_8937, w_022_8938, w_022_8942, w_022_8944, w_022_8945, w_022_8947, w_022_8949, w_022_8950, w_022_8951, w_022_8952, w_022_8953, w_022_8954, w_022_8955, w_022_8958, w_022_8960, w_022_8961, w_022_8962, w_022_8963, w_022_8965, w_022_8970, w_022_8971, w_022_8973, w_022_8975, w_022_8978, w_022_8980, w_022_8981, w_022_8982, w_022_8983, w_022_8985, w_022_8986, w_022_8989, w_022_8994, w_022_8996, w_022_8997, w_022_8998, w_022_9001, w_022_9004, w_022_9006, w_022_9007, w_022_9008, w_022_9009, w_022_9011, w_022_9012, w_022_9014, w_022_9015, w_022_9018, w_022_9020, w_022_9021, w_022_9026, w_022_9028, w_022_9029, w_022_9030, w_022_9031, w_022_9032, w_022_9035, w_022_9036, w_022_9037, w_022_9041, w_022_9042, w_022_9044, w_022_9045, w_022_9047, w_022_9050, w_022_9051, w_022_9052, w_022_9053, w_022_9054, w_022_9055, w_022_9056, w_022_9057, w_022_9058, w_022_9059, w_022_9060, w_022_9061, w_022_9062, w_022_9065, w_022_9066, w_022_9067, w_022_9069, w_022_9070, w_022_9072, w_022_9076, w_022_9077, w_022_9078, w_022_9079, w_022_9082, w_022_9085, w_022_9086, w_022_9089, w_022_9092, w_022_9093, w_022_9094, w_022_9095, w_022_9101, w_022_9102, w_022_9103, w_022_9105, w_022_9106, w_022_9109, w_022_9110, w_022_9112, w_022_9113, w_022_9114, w_022_9115, w_022_9117, w_022_9118, w_022_9121, w_022_9122, w_022_9123, w_022_9124, w_022_9126, w_022_9127, w_022_9129, w_022_9130, w_022_9131, w_022_9132, w_022_9133, w_022_9135, w_022_9138, w_022_9139, w_022_9141, w_022_9143, w_022_9144, w_022_9146, w_022_9147, w_022_9149, w_022_9150, w_022_9152, w_022_9153, w_022_9154, w_022_9156, w_022_9157, w_022_9158, w_022_9160, w_022_9163, w_022_9164, w_022_9165, w_022_9166, w_022_9167, w_022_9168, w_022_9169, w_022_9171, w_022_9172, w_022_9174, w_022_9176, w_022_9177, w_022_9178, w_022_9180, w_022_9183, w_022_9184, w_022_9185, w_022_9186, w_022_9187, w_022_9191, w_022_9192, w_022_9193, w_022_9194, w_022_9197, w_022_9198, w_022_9200, w_022_9201, w_022_9202, w_022_9203, w_022_9204, w_022_9206, w_022_9208, w_022_9211, w_022_9214, w_022_9215, w_022_9217, w_022_9218, w_022_9223, w_022_9224, w_022_9226, w_022_9227, w_022_9228, w_022_9230, w_022_9231, w_022_9233, w_022_9234, w_022_9238, w_022_9241, w_022_9242, w_022_9246, w_022_9247, w_022_9248, w_022_9249, w_022_9250, w_022_9251, w_022_9252, w_022_9254, w_022_9255, w_022_9256, w_022_9257, w_022_9258, w_022_9259, w_022_9261, w_022_9264, w_022_9265, w_022_9268, w_022_9269, w_022_9270, w_022_9271, w_022_9272, w_022_9274, w_022_9277, w_022_9280, w_022_9283, w_022_9285, w_022_9289, w_022_9290, w_022_9292, w_022_9298, w_022_9299, w_022_9301, w_022_9302, w_022_9304, w_022_9306, w_022_9309, w_022_9310, w_022_9312, w_022_9315, w_022_9316, w_022_9317, w_022_9318, w_022_9319, w_022_9321, w_022_9322, w_022_9324, w_022_9326, w_022_9327, w_022_9328, w_022_9329, w_022_9330, w_022_9331, w_022_9333, w_022_9334, w_022_9339, w_022_9340, w_022_9344, w_022_9345, w_022_9346, w_022_9348, w_022_9349, w_022_9354, w_022_9355, w_022_9356, w_022_9364, w_022_9366, w_022_9367, w_022_9369, w_022_9370, w_022_9371, w_022_9372, w_022_9373, w_022_9376, w_022_9377, w_022_9380, w_022_9382, w_022_9384, w_022_9385, w_022_9386, w_022_9390, w_022_9391, w_022_9392, w_022_9393, w_022_9394, w_022_9395, w_022_9396, w_022_9397, w_022_9398, w_022_9399, w_022_9400, w_022_9403, w_022_9409, w_022_9410, w_022_9411, w_022_9412, w_022_9416, w_022_9418, w_022_9419, w_022_9420, w_022_9421, w_022_9427, w_022_9428, w_022_9429, w_022_9430, w_022_9432, w_022_9433, w_022_9434, w_022_9436, w_022_9437, w_022_9438, w_022_9439, w_022_9440, w_022_9441, w_022_9442, w_022_9443, w_022_9444, w_022_9448, w_022_9449, w_022_9450, w_022_9452, w_022_9453, w_022_9455, w_022_9457, w_022_9462, w_022_9463, w_022_9470, w_022_9471, w_022_9473, w_022_9476, w_022_9478, w_022_9479, w_022_9481, w_022_9482, w_022_9483, w_022_9484, w_022_9486, w_022_9488, w_022_9489, w_022_9490, w_022_9493, w_022_9494, w_022_9495, w_022_9496, w_022_9497, w_022_9499, w_022_9500, w_022_9501, w_022_9503, w_022_9504, w_022_9506, w_022_9509, w_022_9511, w_022_9512, w_022_9513, w_022_9516, w_022_9517, w_022_9520, w_022_9522, w_022_9523, w_022_9524, w_022_9525, w_022_9526, w_022_9527, w_022_9530, w_022_9531, w_022_9534, w_022_9536, w_022_9537, w_022_9538, w_022_9540, w_022_9541, w_022_9542, w_022_9543, w_022_9544, w_022_9545, w_022_9547, w_022_9550, w_022_9553, w_022_9554, w_022_9555, w_022_9556, w_022_9559, w_022_9560, w_022_9562, w_022_9564, w_022_9565, w_022_9567, w_022_9572, w_022_9573, w_022_9575, w_022_9577, w_022_9578, w_022_9579, w_022_9580, w_022_9581, w_022_9582, w_022_9583, w_022_9584, w_022_9585, w_022_9586, w_022_9587, w_022_9589, w_022_9591, w_022_9592, w_022_9594, w_022_9595, w_022_9596, w_022_9597, w_022_9603, w_022_9604, w_022_9606, w_022_9608, w_022_9609, w_022_9611, w_022_9612, w_022_9613, w_022_9615, w_022_9616, w_022_9617, w_022_9618, w_022_9619, w_022_9620, w_022_9621, w_022_9623, w_022_9624, w_022_9627, w_022_9628, w_022_9629, w_022_9630, w_022_9631, w_022_9632, w_022_9633, w_022_9635, w_022_9637, w_022_9638, w_022_9639, w_022_9640, w_022_9642, w_022_9645, w_022_9647, w_022_9648, w_022_9650, w_022_9654, w_022_9655, w_022_9657, w_022_9658, w_022_9659, w_022_9661, w_022_9662, w_022_9663, w_022_9664, w_022_9665, w_022_9666, w_022_9668, w_022_9670, w_022_9671, w_022_9677, w_022_9679, w_022_9680, w_022_9681, w_022_9682, w_022_9683, w_022_9684, w_022_9685, w_022_9687, w_022_9688, w_022_9690, w_022_9691, w_022_9694, w_022_9695, w_022_9696, w_022_9697, w_022_9702, w_022_9704, w_022_9705, w_022_9707, w_022_9709, w_022_9712, w_022_9714, w_022_9715, w_022_9717, w_022_9718, w_022_9719, w_022_9723, w_022_9724, w_022_9725, w_022_9726, w_022_9727, w_022_9728, w_022_9729, w_022_9731, w_022_9732, w_022_9733, w_022_9736, w_022_9737, w_022_9739, w_022_9740, w_022_9741, w_022_9742, w_022_9744, w_022_9745, w_022_9746, w_022_9750, w_022_9751, w_022_9753, w_022_9754, w_022_9756, w_022_9758, w_022_9764, w_022_9766, w_022_9771, w_022_9773, w_022_9774, w_022_9776, w_022_9779, w_022_9780, w_022_9782, w_022_9783, w_022_9784, w_022_9785, w_022_9787, w_022_9791, w_022_9793, w_022_9795, w_022_9797, w_022_9798, w_022_9799, w_022_9800, w_022_9801, w_022_9802, w_022_9803, w_022_9804, w_022_9805, w_022_9806, w_022_9807, w_022_9808, w_022_9810, w_022_9811, w_022_9815, w_022_9817, w_022_9819, w_022_9823, w_022_9824, w_022_9825, w_022_9828, w_022_9829, w_022_9830, w_022_9833, w_022_9834, w_022_9835, w_022_9836, w_022_9837, w_022_9838, w_022_9839, w_022_9840, w_022_9841, w_022_9842, w_022_9843, w_022_9844, w_022_9846, w_022_9847, w_022_9848, w_022_9849, w_022_9850, w_022_9851, w_022_9852, w_022_9853, w_022_9854, w_022_9855, w_022_9856, w_022_9858, w_022_9861, w_022_9863, w_022_9864, w_022_9865, w_022_9867, w_022_9868, w_022_9869, w_022_9870, w_022_9871, w_022_9872, w_022_9874, w_022_9875, w_022_9876, w_022_9877, w_022_9879, w_022_9881, w_022_9882, w_022_9883, w_022_9884, w_022_9886, w_022_9887, w_022_9888, w_022_9890, w_022_9895, w_022_9896, w_022_9897, w_022_9900, w_022_9901, w_022_9903, w_022_9911, w_022_9914, w_022_9915, w_022_9917, w_022_9918, w_022_9919, w_022_9921, w_022_9922, w_022_9925, w_022_9926, w_022_9927, w_022_9930, w_022_9932, w_022_9933, w_022_9934, w_022_9935, w_022_9936, w_022_9937, w_022_9939, w_022_9940, w_022_9941, w_022_9943, w_022_9946, w_022_9948, w_022_9949, w_022_9950, w_022_9952, w_022_9953;
  wire w_023_000, w_023_001, w_023_002, w_023_003, w_023_004, w_023_005, w_023_007, w_023_008, w_023_009, w_023_010, w_023_011, w_023_012, w_023_014, w_023_017, w_023_018, w_023_019, w_023_020, w_023_022, w_023_023, w_023_024, w_023_025, w_023_026, w_023_027, w_023_029, w_023_030, w_023_031, w_023_032, w_023_035, w_023_036, w_023_037, w_023_038, w_023_040, w_023_041, w_023_042, w_023_045, w_023_046, w_023_047, w_023_048, w_023_050, w_023_051, w_023_052, w_023_053, w_023_054, w_023_055, w_023_056, w_023_057, w_023_058, w_023_059, w_023_060, w_023_061, w_023_062, w_023_063, w_023_065, w_023_066, w_023_069, w_023_070, w_023_073, w_023_074, w_023_075, w_023_076, w_023_077, w_023_078, w_023_079, w_023_081, w_023_082, w_023_083, w_023_085, w_023_086, w_023_089, w_023_091, w_023_092, w_023_093, w_023_094, w_023_095, w_023_097, w_023_098, w_023_099, w_023_100, w_023_101, w_023_103, w_023_104, w_023_105, w_023_106, w_023_107, w_023_109, w_023_110, w_023_112, w_023_114, w_023_115, w_023_116, w_023_117, w_023_118, w_023_119, w_023_120, w_023_121, w_023_122, w_023_123, w_023_125, w_023_128, w_023_129, w_023_130, w_023_131, w_023_133, w_023_134, w_023_135, w_023_137, w_023_138, w_023_139, w_023_140, w_023_141, w_023_143, w_023_144, w_023_145, w_023_147, w_023_148, w_023_149, w_023_150, w_023_151, w_023_152, w_023_153, w_023_154, w_023_155, w_023_156, w_023_157, w_023_160, w_023_161, w_023_162, w_023_163, w_023_164, w_023_165, w_023_166, w_023_167, w_023_168, w_023_169, w_023_170, w_023_171, w_023_172, w_023_174, w_023_176, w_023_177, w_023_178, w_023_180, w_023_181, w_023_183, w_023_184, w_023_185, w_023_186, w_023_187, w_023_188, w_023_189, w_023_190, w_023_191, w_023_192, w_023_193, w_023_195, w_023_196, w_023_197, w_023_198, w_023_199, w_023_200, w_023_201, w_023_202, w_023_203, w_023_204, w_023_205, w_023_206, w_023_207, w_023_208, w_023_209, w_023_210, w_023_211, w_023_212, w_023_214, w_023_215, w_023_216, w_023_217, w_023_218, w_023_219, w_023_220, w_023_221, w_023_222, w_023_223, w_023_224, w_023_225, w_023_226, w_023_227, w_023_228, w_023_229, w_023_230, w_023_231, w_023_232, w_023_233, w_023_234, w_023_235, w_023_236, w_023_238, w_023_239, w_023_240, w_023_241, w_023_242, w_023_243, w_023_244, w_023_245, w_023_246, w_023_247, w_023_248, w_023_249, w_023_252, w_023_253, w_023_254, w_023_255, w_023_256, w_023_257, w_023_258, w_023_259, w_023_260, w_023_261, w_023_264, w_023_266, w_023_267, w_023_268, w_023_269, w_023_270, w_023_272, w_023_273, w_023_274, w_023_275, w_023_278, w_023_279, w_023_280, w_023_281, w_023_282, w_023_283, w_023_284, w_023_285, w_023_286, w_023_289, w_023_291, w_023_292, w_023_293, w_023_294, w_023_295, w_023_296, w_023_297, w_023_298, w_023_299, w_023_300, w_023_301, w_023_304, w_023_305, w_023_306, w_023_307, w_023_308, w_023_310, w_023_311, w_023_313, w_023_314, w_023_315, w_023_316, w_023_319, w_023_320, w_023_321, w_023_322, w_023_323, w_023_324, w_023_325, w_023_327, w_023_328, w_023_329, w_023_330, w_023_331, w_023_332, w_023_333, w_023_334, w_023_335, w_023_336, w_023_338, w_023_339, w_023_340, w_023_341, w_023_342, w_023_343, w_023_344, w_023_347, w_023_348, w_023_351, w_023_352, w_023_353, w_023_354, w_023_355, w_023_357, w_023_358, w_023_360, w_023_361, w_023_362, w_023_363, w_023_365, w_023_366, w_023_367, w_023_368, w_023_369, w_023_370, w_023_372, w_023_373, w_023_374, w_023_375, w_023_376, w_023_377, w_023_378, w_023_379, w_023_381, w_023_382, w_023_383, w_023_384, w_023_385, w_023_386, w_023_387, w_023_388, w_023_389, w_023_390, w_023_391, w_023_392, w_023_393, w_023_394, w_023_395, w_023_396, w_023_398, w_023_400, w_023_401, w_023_402, w_023_403, w_023_404, w_023_405, w_023_406, w_023_407, w_023_408, w_023_409, w_023_410, w_023_411, w_023_412, w_023_413, w_023_414, w_023_415, w_023_417, w_023_419, w_023_420, w_023_422, w_023_423, w_023_424, w_023_425, w_023_426, w_023_428, w_023_429, w_023_430, w_023_431, w_023_432, w_023_433, w_023_434, w_023_435, w_023_436, w_023_437, w_023_438, w_023_439, w_023_440, w_023_441, w_023_442, w_023_443, w_023_444, w_023_445, w_023_446, w_023_448, w_023_449, w_023_450, w_023_451, w_023_452, w_023_453, w_023_455, w_023_456, w_023_457, w_023_458, w_023_459, w_023_460, w_023_461, w_023_462, w_023_464, w_023_466, w_023_467, w_023_468, w_023_470, w_023_471, w_023_472, w_023_473, w_023_474, w_023_475, w_023_476, w_023_477, w_023_478, w_023_479, w_023_480, w_023_481, w_023_482, w_023_483, w_023_486, w_023_488, w_023_490, w_023_494, w_023_495, w_023_497, w_023_498, w_023_500, w_023_501, w_023_502, w_023_503, w_023_505, w_023_506, w_023_507, w_023_509, w_023_510, w_023_511, w_023_513, w_023_514, w_023_515, w_023_517, w_023_518, w_023_524, w_023_527, w_023_531, w_023_533, w_023_536, w_023_538, w_023_539, w_023_541, w_023_542, w_023_543, w_023_545, w_023_546, w_023_547, w_023_549, w_023_550, w_023_551, w_023_552, w_023_554, w_023_555, w_023_556, w_023_557, w_023_558, w_023_559, w_023_562, w_023_564, w_023_565, w_023_566, w_023_567, w_023_568, w_023_572, w_023_576, w_023_578, w_023_579, w_023_581, w_023_584, w_023_585, w_023_587, w_023_588, w_023_589, w_023_591, w_023_598, w_023_599, w_023_600, w_023_601, w_023_602, w_023_604, w_023_605, w_023_606, w_023_607, w_023_609, w_023_610, w_023_611, w_023_613, w_023_614, w_023_616, w_023_620, w_023_622, w_023_623, w_023_624, w_023_625, w_023_626, w_023_627, w_023_628, w_023_629, w_023_632, w_023_634, w_023_636, w_023_638, w_023_640, w_023_641, w_023_643, w_023_644, w_023_646, w_023_647, w_023_653, w_023_655, w_023_658, w_023_659, w_023_660, w_023_661, w_023_664, w_023_668, w_023_669, w_023_670, w_023_671, w_023_672, w_023_673, w_023_675, w_023_676, w_023_677, w_023_678, w_023_681, w_023_684, w_023_685, w_023_686, w_023_687, w_023_688, w_023_689, w_023_692, w_023_693, w_023_695, w_023_698, w_023_700, w_023_702, w_023_703, w_023_704, w_023_705, w_023_706, w_023_707, w_023_711, w_023_712, w_023_713, w_023_716, w_023_717, w_023_718, w_023_719, w_023_720, w_023_721, w_023_723, w_023_725, w_023_729, w_023_731, w_023_732, w_023_734, w_023_736, w_023_738, w_023_739, w_023_742, w_023_743, w_023_745, w_023_746, w_023_748, w_023_749, w_023_753, w_023_755, w_023_758, w_023_759, w_023_760, w_023_761, w_023_762, w_023_763, w_023_765, w_023_766, w_023_767, w_023_769, w_023_773, w_023_774, w_023_776, w_023_777, w_023_780, w_023_783, w_023_784, w_023_785, w_023_787, w_023_789, w_023_793, w_023_795, w_023_796, w_023_797, w_023_798, w_023_799, w_023_800, w_023_801, w_023_803, w_023_804, w_023_805, w_023_809, w_023_811, w_023_812, w_023_816, w_023_817, w_023_818, w_023_820, w_023_821, w_023_823, w_023_824, w_023_830, w_023_832, w_023_833, w_023_834, w_023_835, w_023_836, w_023_837, w_023_838, w_023_840, w_023_841, w_023_843, w_023_847, w_023_849, w_023_851, w_023_853, w_023_854, w_023_858, w_023_859, w_023_860, w_023_862, w_023_863, w_023_864, w_023_866, w_023_867, w_023_868, w_023_871, w_023_872, w_023_873, w_023_874, w_023_875, w_023_878, w_023_879, w_023_880, w_023_881, w_023_882, w_023_884, w_023_886, w_023_891, w_023_892, w_023_893, w_023_896, w_023_898, w_023_899, w_023_900, w_023_901, w_023_902, w_023_906, w_023_907, w_023_912, w_023_913, w_023_914, w_023_917, w_023_918, w_023_919, w_023_921, w_023_922, w_023_924, w_023_928, w_023_930, w_023_931, w_023_932, w_023_935, w_023_936, w_023_937, w_023_938, w_023_939, w_023_941, w_023_943, w_023_944, w_023_945, w_023_948, w_023_949, w_023_950, w_023_951, w_023_952, w_023_953, w_023_954, w_023_955, w_023_957, w_023_961, w_023_962, w_023_964, w_023_966, w_023_967, w_023_968, w_023_972, w_023_973, w_023_974, w_023_976, w_023_979, w_023_980, w_023_981, w_023_982, w_023_983, w_023_985, w_023_986, w_023_987, w_023_988, w_023_991, w_023_994, w_023_997, w_023_998, w_023_999, w_023_1000, w_023_1001, w_023_1002, w_023_1005, w_023_1006, w_023_1008, w_023_1010, w_023_1011, w_023_1012, w_023_1013, w_023_1015, w_023_1016, w_023_1017, w_023_1018, w_023_1020, w_023_1021, w_023_1024, w_023_1025, w_023_1026, w_023_1029, w_023_1030, w_023_1031, w_023_1032, w_023_1033, w_023_1042, w_023_1043, w_023_1044, w_023_1045, w_023_1046, w_023_1048, w_023_1053, w_023_1054, w_023_1056, w_023_1057, w_023_1058, w_023_1060, w_023_1062, w_023_1065, w_023_1066, w_023_1067, w_023_1070, w_023_1071, w_023_1072, w_023_1074, w_023_1075, w_023_1076, w_023_1077, w_023_1078, w_023_1084, w_023_1085, w_023_1086, w_023_1087, w_023_1088, w_023_1089, w_023_1090, w_023_1092, w_023_1094, w_023_1095, w_023_1096, w_023_1097, w_023_1098, w_023_1099, w_023_1102, w_023_1104, w_023_1105, w_023_1106, w_023_1107, w_023_1108, w_023_1109, w_023_1110, w_023_1112, w_023_1113, w_023_1115, w_023_1116, w_023_1121, w_023_1124, w_023_1125, w_023_1126, w_023_1128, w_023_1130, w_023_1131, w_023_1132, w_023_1133, w_023_1136, w_023_1137, w_023_1139, w_023_1140, w_023_1141, w_023_1143, w_023_1145, w_023_1146, w_023_1148, w_023_1150, w_023_1153, w_023_1156, w_023_1157, w_023_1158, w_023_1159, w_023_1160, w_023_1161, w_023_1162, w_023_1167, w_023_1168, w_023_1169, w_023_1170, w_023_1171, w_023_1178, w_023_1179, w_023_1181, w_023_1184, w_023_1185, w_023_1188, w_023_1189, w_023_1190, w_023_1192, w_023_1196, w_023_1197, w_023_1200, w_023_1201, w_023_1202, w_023_1206, w_023_1207, w_023_1210, w_023_1211, w_023_1212, w_023_1214, w_023_1218, w_023_1220, w_023_1221, w_023_1223, w_023_1224, w_023_1225, w_023_1227, w_023_1228, w_023_1232, w_023_1233, w_023_1234, w_023_1235, w_023_1237, w_023_1241, w_023_1243, w_023_1246, w_023_1248, w_023_1254, w_023_1255, w_023_1258, w_023_1260, w_023_1262, w_023_1263, w_023_1267, w_023_1268, w_023_1269, w_023_1272, w_023_1273, w_023_1274, w_023_1275, w_023_1276, w_023_1277, w_023_1283, w_023_1285, w_023_1289, w_023_1292, w_023_1295, w_023_1299, w_023_1301, w_023_1302, w_023_1303, w_023_1304, w_023_1305, w_023_1306, w_023_1308, w_023_1309, w_023_1310, w_023_1311, w_023_1312, w_023_1314, w_023_1315, w_023_1316, w_023_1317, w_023_1319, w_023_1322, w_023_1323, w_023_1324, w_023_1325, w_023_1330, w_023_1331, w_023_1332, w_023_1333, w_023_1334, w_023_1336, w_023_1339, w_023_1342, w_023_1346, w_023_1347, w_023_1348, w_023_1349, w_023_1350, w_023_1351, w_023_1352, w_023_1354, w_023_1356, w_023_1358, w_023_1359, w_023_1360, w_023_1363, w_023_1364, w_023_1365, w_023_1366, w_023_1368, w_023_1369, w_023_1370, w_023_1378, w_023_1379, w_023_1380, w_023_1381, w_023_1382, w_023_1385, w_023_1387, w_023_1388, w_023_1391, w_023_1392, w_023_1393, w_023_1394, w_023_1395, w_023_1396, w_023_1397, w_023_1398, w_023_1400, w_023_1402, w_023_1403, w_023_1404, w_023_1406, w_023_1408, w_023_1409, w_023_1413, w_023_1415, w_023_1416, w_023_1418, w_023_1419, w_023_1420, w_023_1423, w_023_1424, w_023_1426, w_023_1428, w_023_1429, w_023_1431, w_023_1432, w_023_1435, w_023_1436, w_023_1438, w_023_1439, w_023_1440, w_023_1441, w_023_1442, w_023_1445, w_023_1446, w_023_1447, w_023_1448, w_023_1449, w_023_1451, w_023_1453, w_023_1454, w_023_1456, w_023_1457, w_023_1458, w_023_1459, w_023_1460, w_023_1462, w_023_1464, w_023_1465, w_023_1466, w_023_1468, w_023_1469, w_023_1470, w_023_1471, w_023_1472, w_023_1473, w_023_1475, w_023_1476, w_023_1481, w_023_1482, w_023_1485, w_023_1487, w_023_1489, w_023_1490, w_023_1491, w_023_1492, w_023_1496, w_023_1499, w_023_1502, w_023_1503, w_023_1504, w_023_1505, w_023_1507, w_023_1508, w_023_1510, w_023_1512, w_023_1513, w_023_1515, w_023_1519, w_023_1521, w_023_1523, w_023_1524, w_023_1525, w_023_1529, w_023_1530, w_023_1531, w_023_1532, w_023_1533, w_023_1534, w_023_1537, w_023_1538, w_023_1539, w_023_1540, w_023_1541, w_023_1543, w_023_1544, w_023_1547, w_023_1550, w_023_1551, w_023_1553, w_023_1554, w_023_1555, w_023_1558, w_023_1559, w_023_1560, w_023_1563, w_023_1565, w_023_1567, w_023_1568, w_023_1571, w_023_1572, w_023_1574, w_023_1575, w_023_1576, w_023_1580, w_023_1581, w_023_1582, w_023_1585, w_023_1586, w_023_1588, w_023_1589, w_023_1590, w_023_1592, w_023_1593, w_023_1595, w_023_1596, w_023_1597, w_023_1598, w_023_1599, w_023_1605, w_023_1606, w_023_1607, w_023_1608, w_023_1609, w_023_1612, w_023_1613, w_023_1615, w_023_1616, w_023_1618, w_023_1619, w_023_1621, w_023_1623, w_023_1624, w_023_1627, w_023_1628, w_023_1629, w_023_1630, w_023_1631, w_023_1632, w_023_1637, w_023_1638, w_023_1641, w_023_1642, w_023_1644, w_023_1646, w_023_1647, w_023_1649, w_023_1650, w_023_1651, w_023_1652, w_023_1653, w_023_1656, w_023_1657, w_023_1658, w_023_1659, w_023_1660, w_023_1661, w_023_1662, w_023_1663, w_023_1665, w_023_1666, w_023_1668, w_023_1669, w_023_1672, w_023_1674, w_023_1675, w_023_1677, w_023_1678, w_023_1679, w_023_1682, w_023_1683, w_023_1684, w_023_1685, w_023_1686, w_023_1687, w_023_1688, w_023_1689, w_023_1691, w_023_1693, w_023_1694, w_023_1695, w_023_1698, w_023_1699, w_023_1701, w_023_1702, w_023_1704, w_023_1705, w_023_1706, w_023_1707, w_023_1708, w_023_1711, w_023_1713, w_023_1714, w_023_1717, w_023_1718, w_023_1719, w_023_1720, w_023_1723, w_023_1724, w_023_1727, w_023_1729, w_023_1731, w_023_1732, w_023_1733, w_023_1734, w_023_1737, w_023_1738, w_023_1740, w_023_1741, w_023_1742, w_023_1743, w_023_1744, w_023_1745, w_023_1746, w_023_1748, w_023_1750, w_023_1751, w_023_1753, w_023_1754, w_023_1755, w_023_1756, w_023_1761, w_023_1762, w_023_1764, w_023_1765, w_023_1767, w_023_1768, w_023_1769, w_023_1771, w_023_1774, w_023_1775, w_023_1776, w_023_1777, w_023_1779, w_023_1781, w_023_1784, w_023_1785, w_023_1786, w_023_1787, w_023_1788, w_023_1789, w_023_1790, w_023_1791, w_023_1793, w_023_1794, w_023_1796, w_023_1797, w_023_1798, w_023_1800, w_023_1801, w_023_1802, w_023_1803, w_023_1806, w_023_1811, w_023_1812, w_023_1814, w_023_1815, w_023_1816, w_023_1817, w_023_1818, w_023_1821, w_023_1822, w_023_1823, w_023_1824, w_023_1827, w_023_1828, w_023_1830, w_023_1831, w_023_1832, w_023_1833, w_023_1834, w_023_1835, w_023_1836, w_023_1837, w_023_1838, w_023_1839, w_023_1840, w_023_1841, w_023_1842, w_023_1847, w_023_1848, w_023_1850, w_023_1851, w_023_1852, w_023_1855, w_023_1856, w_023_1857, w_023_1860, w_023_1861, w_023_1863, w_023_1866, w_023_1867, w_023_1868, w_023_1869, w_023_1870, w_023_1871, w_023_1872, w_023_1873, w_023_1875, w_023_1877, w_023_1878, w_023_1880, w_023_1881, w_023_1883, w_023_1884, w_023_1886, w_023_1891, w_023_1893, w_023_1895, w_023_1897, w_023_1898, w_023_1899, w_023_1900, w_023_1901, w_023_1903, w_023_1907, w_023_1908, w_023_1909, w_023_1911, w_023_1913, w_023_1915, w_023_1916, w_023_1921, w_023_1922, w_023_1923, w_023_1924, w_023_1928, w_023_1931, w_023_1932, w_023_1933, w_023_1934, w_023_1936, w_023_1941, w_023_1943, w_023_1944, w_023_1946, w_023_1947, w_023_1949, w_023_1951, w_023_1952, w_023_1953, w_023_1957, w_023_1960, w_023_1961, w_023_1962, w_023_1964, w_023_1966, w_023_1967, w_023_1969, w_023_1970, w_023_1973, w_023_1977, w_023_1978, w_023_1979, w_023_1980, w_023_1981, w_023_1983, w_023_1984, w_023_1985, w_023_1986, w_023_1987, w_023_1988, w_023_1989, w_023_1990, w_023_1992, w_023_1994, w_023_1995, w_023_1996, w_023_1998, w_023_2000, w_023_2002, w_023_2003, w_023_2007, w_023_2009, w_023_2015, w_023_2016, w_023_2021, w_023_2023, w_023_2024, w_023_2026, w_023_2029, w_023_2030, w_023_2031, w_023_2033, w_023_2039, w_023_2041, w_023_2042, w_023_2044, w_023_2045, w_023_2046, w_023_2047, w_023_2048, w_023_2049, w_023_2051, w_023_2052, w_023_2057, w_023_2061, w_023_2062, w_023_2063, w_023_2065, w_023_2066, w_023_2067, w_023_2068, w_023_2069, w_023_2073, w_023_2074, w_023_2076, w_023_2077, w_023_2078, w_023_2079, w_023_2080, w_023_2082, w_023_2086, w_023_2087, w_023_2088, w_023_2089, w_023_2090, w_023_2091, w_023_2093, w_023_2095, w_023_2096, w_023_2097, w_023_2099, w_023_2100, w_023_2101, w_023_2102, w_023_2103, w_023_2104, w_023_2106, w_023_2107, w_023_2108, w_023_2114, w_023_2117, w_023_2118, w_023_2119, w_023_2122, w_023_2124, w_023_2127, w_023_2128, w_023_2129, w_023_2132, w_023_2133, w_023_2134, w_023_2135, w_023_2138, w_023_2139, w_023_2142, w_023_2143, w_023_2144, w_023_2145, w_023_2147, w_023_2150, w_023_2151, w_023_2154, w_023_2155, w_023_2157, w_023_2158, w_023_2159, w_023_2161, w_023_2163, w_023_2165, w_023_2166, w_023_2167, w_023_2169, w_023_2171, w_023_2172, w_023_2175, w_023_2176, w_023_2177, w_023_2178, w_023_2179, w_023_2181, w_023_2183, w_023_2184, w_023_2189, w_023_2190, w_023_2191, w_023_2193, w_023_2196, w_023_2197, w_023_2198, w_023_2200, w_023_2201, w_023_2205, w_023_2206, w_023_2208, w_023_2209, w_023_2210, w_023_2211, w_023_2212, w_023_2217, w_023_2220, w_023_2223, w_023_2225, w_023_2227, w_023_2228, w_023_2230, w_023_2232, w_023_2233, w_023_2235, w_023_2236, w_023_2237, w_023_2238, w_023_2240, w_023_2243, w_023_2246, w_023_2247, w_023_2248, w_023_2250, w_023_2251, w_023_2252, w_023_2254, w_023_2255, w_023_2256, w_023_2258, w_023_2263, w_023_2265, w_023_2267, w_023_2270, w_023_2273, w_023_2274, w_023_2275, w_023_2276, w_023_2278, w_023_2281, w_023_2284, w_023_2285, w_023_2287, w_023_2288, w_023_2289, w_023_2290, w_023_2291, w_023_2294, w_023_2295, w_023_2297, w_023_2298, w_023_2299, w_023_2301, w_023_2303, w_023_2304, w_023_2305, w_023_2306, w_023_2309, w_023_2311, w_023_2312, w_023_2314, w_023_2315, w_023_2316, w_023_2318, w_023_2319, w_023_2322, w_023_2324, w_023_2327, w_023_2328, w_023_2331, w_023_2332, w_023_2334, w_023_2335, w_023_2336, w_023_2337, w_023_2338, w_023_2339, w_023_2340, w_023_2341, w_023_2342, w_023_2344, w_023_2348, w_023_2349, w_023_2350, w_023_2351, w_023_2352, w_023_2355, w_023_2360, w_023_2361, w_023_2364, w_023_2365, w_023_2366, w_023_2367, w_023_2368, w_023_2370, w_023_2371, w_023_2373, w_023_2378, w_023_2381, w_023_2382, w_023_2383, w_023_2384, w_023_2385, w_023_2386, w_023_2388, w_023_2389, w_023_2391, w_023_2392, w_023_2397, w_023_2400, w_023_2401, w_023_2404, w_023_2408, w_023_2409, w_023_2410, w_023_2412, w_023_2413, w_023_2414, w_023_2416, w_023_2417, w_023_2419, w_023_2421, w_023_2422, w_023_2424, w_023_2425, w_023_2427, w_023_2428, w_023_2429, w_023_2430, w_023_2431, w_023_2432, w_023_2433, w_023_2436, w_023_2438, w_023_2439, w_023_2440, w_023_2441, w_023_2442, w_023_2443, w_023_2444, w_023_2445, w_023_2446, w_023_2448, w_023_2449, w_023_2450, w_023_2451, w_023_2453, w_023_2455, w_023_2458, w_023_2459, w_023_2460, w_023_2463, w_023_2465, w_023_2467, w_023_2469, w_023_2472, w_023_2473, w_023_2474, w_023_2476, w_023_2477, w_023_2479, w_023_2480, w_023_2483, w_023_2488, w_023_2489, w_023_2490, w_023_2491, w_023_2493, w_023_2494, w_023_2497, w_023_2498, w_023_2499, w_023_2500, w_023_2501, w_023_2503, w_023_2504, w_023_2507, w_023_2508, w_023_2509, w_023_2511, w_023_2512, w_023_2514, w_023_2515, w_023_2518, w_023_2519, w_023_2523, w_023_2524, w_023_2525, w_023_2528, w_023_2529, w_023_2530, w_023_2531, w_023_2532, w_023_2534, w_023_2536, w_023_2538, w_023_2539, w_023_2541, w_023_2542, w_023_2545, w_023_2547, w_023_2550, w_023_2553, w_023_2558, w_023_2559, w_023_2561, w_023_2562, w_023_2563, w_023_2565, w_023_2566, w_023_2567, w_023_2568, w_023_2569, w_023_2572, w_023_2573, w_023_2579, w_023_2580, w_023_2581, w_023_2584, w_023_2587, w_023_2589, w_023_2590, w_023_2595, w_023_2597, w_023_2598, w_023_2599, w_023_2600, w_023_2602, w_023_2604, w_023_2605, w_023_2608, w_023_2609, w_023_2610, w_023_2611, w_023_2612, w_023_2613, w_023_2614, w_023_2617, w_023_2621, w_023_2623, w_023_2624, w_023_2626, w_023_2627, w_023_2631, w_023_2632, w_023_2634, w_023_2636, w_023_2638, w_023_2639, w_023_2640, w_023_2641, w_023_2643, w_023_2644, w_023_2646, w_023_2647, w_023_2648, w_023_2649, w_023_2650, w_023_2651, w_023_2653, w_023_2657, w_023_2660, w_023_2662, w_023_2663, w_023_2666, w_023_2667, w_023_2669, w_023_2672, w_023_2673, w_023_2674, w_023_2676, w_023_2677, w_023_2678, w_023_2679, w_023_2680, w_023_2681, w_023_2682, w_023_2684, w_023_2685, w_023_2686, w_023_2687, w_023_2690, w_023_2695, w_023_2696, w_023_2699, w_023_2700, w_023_2702, w_023_2705, w_023_2706, w_023_2707, w_023_2708, w_023_2710, w_023_2713, w_023_2714, w_023_2717, w_023_2718, w_023_2721, w_023_2723, w_023_2725, w_023_2726, w_023_2727, w_023_2729, w_023_2731, w_023_2734, w_023_2735, w_023_2736, w_023_2737, w_023_2739, w_023_2740, w_023_2743, w_023_2744, w_023_2746, w_023_2747, w_023_2748, w_023_2750, w_023_2752, w_023_2753, w_023_2754, w_023_2758, w_023_2759, w_023_2761, w_023_2762, w_023_2764, w_023_2765, w_023_2767, w_023_2768, w_023_2769, w_023_2772, w_023_2773, w_023_2774, w_023_2776, w_023_2780, w_023_2781, w_023_2783, w_023_2784, w_023_2785, w_023_2786, w_023_2787, w_023_2789, w_023_2790, w_023_2791, w_023_2792, w_023_2794, w_023_2796, w_023_2797, w_023_2800, w_023_2801, w_023_2805, w_023_2806, w_023_2807, w_023_2808, w_023_2810, w_023_2812, w_023_2813, w_023_2817, w_023_2818, w_023_2820, w_023_2821, w_023_2822, w_023_2823, w_023_2824, w_023_2825, w_023_2827, w_023_2829, w_023_2830, w_023_2831, w_023_2832, w_023_2833, w_023_2834, w_023_2838, w_023_2839, w_023_2841, w_023_2842, w_023_2844, w_023_2847, w_023_2848, w_023_2850, w_023_2852, w_023_2855, w_023_2856, w_023_2857, w_023_2858, w_023_2859, w_023_2860, w_023_2861, w_023_2863, w_023_2866, w_023_2870, w_023_2872, w_023_2874, w_023_2875, w_023_2876, w_023_2877, w_023_2879, w_023_2882, w_023_2883, w_023_2884, w_023_2886, w_023_2887, w_023_2889, w_023_2891, w_023_2893, w_023_2894, w_023_2895, w_023_2896, w_023_2897, w_023_2898, w_023_2899, w_023_2900, w_023_2901, w_023_2902, w_023_2903, w_023_2905, w_023_2906, w_023_2907, w_023_2911, w_023_2912, w_023_2913, w_023_2914, w_023_2917, w_023_2918, w_023_2919, w_023_2920, w_023_2922, w_023_2924, w_023_2925, w_023_2927, w_023_2929, w_023_2932, w_023_2941, w_023_2946, w_023_2949, w_023_2950, w_023_2951, w_023_2952, w_023_2954, w_023_2955, w_023_2957, w_023_2958, w_023_2959, w_023_2965, w_023_2966, w_023_2969, w_023_2971, w_023_2973, w_023_2974, w_023_2975, w_023_2978, w_023_2980, w_023_2981, w_023_2983, w_023_2984, w_023_2985, w_023_2990, w_023_2992, w_023_2994, w_023_2995, w_023_2996, w_023_2997, w_023_2998, w_023_2999, w_023_3000, w_023_3002, w_023_3003, w_023_3005, w_023_3006, w_023_3008, w_023_3009, w_023_3010, w_023_3012, w_023_3013, w_023_3014, w_023_3016, w_023_3017, w_023_3020, w_023_3022, w_023_3023, w_023_3024, w_023_3025, w_023_3026, w_023_3027, w_023_3028, w_023_3029, w_023_3032, w_023_3033, w_023_3034, w_023_3036, w_023_3038, w_023_3041, w_023_3042, w_023_3043, w_023_3045, w_023_3047, w_023_3049, w_023_3050, w_023_3052, w_023_3053, w_023_3054, w_023_3055, w_023_3058, w_023_3059, w_023_3060, w_023_3062, w_023_3066, w_023_3071, w_023_3072, w_023_3074, w_023_3075, w_023_3076, w_023_3077, w_023_3082, w_023_3083, w_023_3084, w_023_3085, w_023_3087, w_023_3089, w_023_3090, w_023_3094, w_023_3095, w_023_3101, w_023_3103, w_023_3106, w_023_3108, w_023_3109, w_023_3110, w_023_3114, w_023_3116, w_023_3118, w_023_3119, w_023_3121, w_023_3124, w_023_3127, w_023_3130, w_023_3133, w_023_3134, w_023_3135, w_023_3137, w_023_3139, w_023_3140, w_023_3142, w_023_3143, w_023_3144, w_023_3145, w_023_3147, w_023_3151, w_023_3152, w_023_3155, w_023_3158, w_023_3159, w_023_3163, w_023_3164, w_023_3166, w_023_3169, w_023_3171, w_023_3173, w_023_3174, w_023_3177, w_023_3181, w_023_3182, w_023_3184, w_023_3185, w_023_3186, w_023_3187, w_023_3188, w_023_3191, w_023_3192, w_023_3193, w_023_3194, w_023_3199, w_023_3200, w_023_3202, w_023_3205, w_023_3206, w_023_3207, w_023_3208, w_023_3210, w_023_3211, w_023_3212, w_023_3214, w_023_3216, w_023_3219, w_023_3221, w_023_3222, w_023_3223, w_023_3224, w_023_3225, w_023_3226, w_023_3227, w_023_3229, w_023_3231, w_023_3233, w_023_3236, w_023_3240, w_023_3241, w_023_3242, w_023_3243, w_023_3246, w_023_3248, w_023_3252, w_023_3253, w_023_3256, w_023_3258, w_023_3259, w_023_3262, w_023_3263, w_023_3265, w_023_3266, w_023_3267, w_023_3269, w_023_3271, w_023_3272, w_023_3273, w_023_3275, w_023_3276, w_023_3277, w_023_3280, w_023_3285, w_023_3287, w_023_3289, w_023_3291, w_023_3293, w_023_3295, w_023_3296, w_023_3297, w_023_3300, w_023_3304, w_023_3305, w_023_3307, w_023_3309, w_023_3310, w_023_3312, w_023_3313, w_023_3314, w_023_3315, w_023_3316, w_023_3319, w_023_3321, w_023_3323, w_023_3324, w_023_3325, w_023_3327, w_023_3328, w_023_3331, w_023_3332, w_023_3333, w_023_3334, w_023_3335, w_023_3336, w_023_3337, w_023_3339, w_023_3341, w_023_3342, w_023_3344, w_023_3345, w_023_3346, w_023_3347, w_023_3349, w_023_3354, w_023_3357, w_023_3358, w_023_3360, w_023_3361, w_023_3364, w_023_3367, w_023_3368, w_023_3371, w_023_3372, w_023_3373, w_023_3374, w_023_3375, w_023_3384, w_023_3385, w_023_3386, w_023_3388, w_023_3392, w_023_3393, w_023_3396, w_023_3399, w_023_3402, w_023_3403, w_023_3404, w_023_3405, w_023_3406, w_023_3407, w_023_3408, w_023_3409, w_023_3411, w_023_3413, w_023_3414, w_023_3416, w_023_3417, w_023_3418, w_023_3420, w_023_3422, w_023_3424, w_023_3426, w_023_3427, w_023_3429, w_023_3430, w_023_3431, w_023_3432, w_023_3433, w_023_3434, w_023_3435, w_023_3436, w_023_3437, w_023_3438, w_023_3441, w_023_3444, w_023_3445, w_023_3448, w_023_3450, w_023_3451, w_023_3452, w_023_3453, w_023_3454, w_023_3456, w_023_3457, w_023_3461, w_023_3462, w_023_3465, w_023_3467, w_023_3469, w_023_3471, w_023_3473, w_023_3475, w_023_3476, w_023_3478, w_023_3479, w_023_3480, w_023_3484, w_023_3486, w_023_3489, w_023_3491, w_023_3493, w_023_3494, w_023_3495, w_023_3496, w_023_3497, w_023_3498, w_023_3500, w_023_3501, w_023_3502, w_023_3503, w_023_3504, w_023_3505, w_023_3507, w_023_3508, w_023_3510, w_023_3511, w_023_3512, w_023_3513, w_023_3514, w_023_3516, w_023_3517, w_023_3518, w_023_3520, w_023_3521, w_023_3523, w_023_3527, w_023_3528, w_023_3530, w_023_3533, w_023_3535, w_023_3538, w_023_3540, w_023_3541, w_023_3542, w_023_3544, w_023_3545, w_023_3546, w_023_3548, w_023_3549, w_023_3553, w_023_3554, w_023_3555, w_023_3556, w_023_3557, w_023_3558, w_023_3559, w_023_3560, w_023_3561, w_023_3562, w_023_3563, w_023_3564, w_023_3565, w_023_3566, w_023_3567, w_023_3568, w_023_3572, w_023_3573, w_023_3575, w_023_3577, w_023_3580, w_023_3581, w_023_3582, w_023_3583, w_023_3584, w_023_3585, w_023_3588, w_023_3589, w_023_3590, w_023_3591, w_023_3592, w_023_3594, w_023_3595, w_023_3597, w_023_3598, w_023_3601, w_023_3603, w_023_3604, w_023_3605, w_023_3606, w_023_3607, w_023_3611, w_023_3612, w_023_3613, w_023_3614, w_023_3615, w_023_3616, w_023_3617, w_023_3620, w_023_3622, w_023_3623, w_023_3626, w_023_3628, w_023_3636, w_023_3642, w_023_3644, w_023_3645, w_023_3646, w_023_3647, w_023_3652, w_023_3653, w_023_3654, w_023_3655, w_023_3656, w_023_3657, w_023_3658, w_023_3659, w_023_3660, w_023_3665, w_023_3666, w_023_3668, w_023_3669, w_023_3670, w_023_3671, w_023_3672, w_023_3673, w_023_3674, w_023_3676, w_023_3677, w_023_3678, w_023_3681, w_023_3685, w_023_3686, w_023_3688, w_023_3689, w_023_3690, w_023_3693, w_023_3694, w_023_3696, w_023_3698, w_023_3699, w_023_3700, w_023_3703, w_023_3704, w_023_3705, w_023_3706, w_023_3707, w_023_3708, w_023_3709, w_023_3710, w_023_3711, w_023_3714, w_023_3715, w_023_3716, w_023_3717, w_023_3719, w_023_3720, w_023_3721, w_023_3725, w_023_3726, w_023_3727, w_023_3728, w_023_3729, w_023_3733, w_023_3734, w_023_3738, w_023_3739, w_023_3740, w_023_3742, w_023_3745, w_023_3746, w_023_3747, w_023_3748, w_023_3752, w_023_3754, w_023_3755, w_023_3756, w_023_3757, w_023_3758, w_023_3761, w_023_3762, w_023_3763, w_023_3765, w_023_3766, w_023_3767, w_023_3768, w_023_3770, w_023_3771, w_023_3772, w_023_3777, w_023_3778, w_023_3780, w_023_3781, w_023_3782, w_023_3783, w_023_3785, w_023_3786, w_023_3787, w_023_3788, w_023_3789, w_023_3790, w_023_3791, w_023_3794, w_023_3795, w_023_3798, w_023_3799, w_023_3800, w_023_3801, w_023_3802, w_023_3803, w_023_3804, w_023_3805, w_023_3806, w_023_3807, w_023_3808, w_023_3809, w_023_3814, w_023_3818, w_023_3820, w_023_3821, w_023_3825, w_023_3828, w_023_3829, w_023_3830, w_023_3831, w_023_3832, w_023_3842, w_023_3843, w_023_3844, w_023_3845, w_023_3846, w_023_3847, w_023_3848, w_023_3849, w_023_3851, w_023_3852, w_023_3854, w_023_3857, w_023_3858, w_023_3860, w_023_3861, w_023_3862, w_023_3865, w_023_3866, w_023_3868, w_023_3870, w_023_3873, w_023_3875, w_023_3876, w_023_3877, w_023_3878, w_023_3879, w_023_3882, w_023_3883, w_023_3884, w_023_3886, w_023_3887, w_023_3888, w_023_3890, w_023_3891, w_023_3894, w_023_3895, w_023_3896, w_023_3903, w_023_3904, w_023_3905, w_023_3906, w_023_3908, w_023_3909, w_023_3910, w_023_3911, w_023_3912, w_023_3914, w_023_3915, w_023_3916, w_023_3917, w_023_3918, w_023_3919, w_023_3920, w_023_3921, w_023_3922, w_023_3924, w_023_3926, w_023_3931, w_023_3932, w_023_3935, w_023_3936, w_023_3940, w_023_3943, w_023_3945, w_023_3946, w_023_3947, w_023_3949, w_023_3950, w_023_3951, w_023_3952, w_023_3953, w_023_3955, w_023_3956, w_023_3957, w_023_3961, w_023_3963, w_023_3965, w_023_3966, w_023_3967, w_023_3968, w_023_3969, w_023_3970, w_023_3973, w_023_3974, w_023_3975, w_023_3976, w_023_3978, w_023_3979, w_023_3982, w_023_3983, w_023_3985, w_023_3986, w_023_3987, w_023_3990, w_023_3991, w_023_3992, w_023_3994, w_023_3995, w_023_3998, w_023_4000, w_023_4003, w_023_4004, w_023_4005, w_023_4006, w_023_4009, w_023_4011, w_023_4014, w_023_4015, w_023_4017, w_023_4018, w_023_4020, w_023_4022, w_023_4023, w_023_4024, w_023_4027, w_023_4028, w_023_4029, w_023_4030, w_023_4031, w_023_4032, w_023_4033, w_023_4037, w_023_4038, w_023_4041, w_023_4042, w_023_4045, w_023_4047, w_023_4048, w_023_4049, w_023_4051, w_023_4052, w_023_4054, w_023_4055, w_023_4057, w_023_4061, w_023_4062, w_023_4064, w_023_4066, w_023_4068, w_023_4069, w_023_4070, w_023_4071, w_023_4072, w_023_4073, w_023_4074, w_023_4075, w_023_4076, w_023_4078, w_023_4081, w_023_4083, w_023_4084, w_023_4085, w_023_4086, w_023_4087, w_023_4088, w_023_4089, w_023_4090, w_023_4092, w_023_4093, w_023_4094, w_023_4095, w_023_4096, w_023_4099, w_023_4100, w_023_4101, w_023_4102, w_023_4103, w_023_4105, w_023_4107, w_023_4108, w_023_4109, w_023_4111, w_023_4112, w_023_4113, w_023_4116, w_023_4117, w_023_4118, w_023_4120, w_023_4121, w_023_4122, w_023_4125, w_023_4127, w_023_4128, w_023_4130, w_023_4132, w_023_4134, w_023_4135, w_023_4136, w_023_4137, w_023_4141, w_023_4142, w_023_4146, w_023_4147, w_023_4149, w_023_4152, w_023_4154, w_023_4155, w_023_4157, w_023_4159, w_023_4160, w_023_4162, w_023_4163, w_023_4165, w_023_4167, w_023_4172, w_023_4176, w_023_4177, w_023_4178, w_023_4179, w_023_4180, w_023_4181, w_023_4182, w_023_4184, w_023_4185, w_023_4186, w_023_4187, w_023_4190, w_023_4191, w_023_4193, w_023_4196, w_023_4197, w_023_4200, w_023_4202, w_023_4203, w_023_4204, w_023_4205, w_023_4206, w_023_4207, w_023_4208, w_023_4209, w_023_4214, w_023_4215, w_023_4216, w_023_4217, w_023_4220, w_023_4221, w_023_4222, w_023_4226, w_023_4228, w_023_4229, w_023_4231, w_023_4232, w_023_4234, w_023_4236, w_023_4237, w_023_4238, w_023_4239, w_023_4240, w_023_4242, w_023_4243, w_023_4245, w_023_4246, w_023_4247, w_023_4248, w_023_4251, w_023_4252, w_023_4253, w_023_4254, w_023_4255, w_023_4257, w_023_4258, w_023_4259, w_023_4261, w_023_4262, w_023_4266, w_023_4268, w_023_4270, w_023_4271, w_023_4272, w_023_4276, w_023_4277, w_023_4278, w_023_4279, w_023_4280, w_023_4281, w_023_4283, w_023_4284, w_023_4286, w_023_4289, w_023_4290, w_023_4291, w_023_4292, w_023_4293, w_023_4296, w_023_4297, w_023_4301, w_023_4302, w_023_4303, w_023_4305, w_023_4306, w_023_4307, w_023_4308, w_023_4309, w_023_4312, w_023_4315, w_023_4316, w_023_4317, w_023_4319, w_023_4321, w_023_4323, w_023_4324, w_023_4325, w_023_4327, w_023_4329, w_023_4330, w_023_4333, w_023_4336, w_023_4337, w_023_4338, w_023_4340, w_023_4341, w_023_4342, w_023_4343, w_023_4345, w_023_4346, w_023_4348, w_023_4349, w_023_4350, w_023_4352, w_023_4353, w_023_4354, w_023_4356, w_023_4358, w_023_4360, w_023_4361, w_023_4362, w_023_4363, w_023_4364, w_023_4365, w_023_4366, w_023_4367, w_023_4369, w_023_4370, w_023_4371, w_023_4372, w_023_4373, w_023_4374, w_023_4378, w_023_4379, w_023_4380, w_023_4381, w_023_4382, w_023_4383, w_023_4386, w_023_4388, w_023_4392, w_023_4393, w_023_4394, w_023_4395, w_023_4396, w_023_4400, w_023_4401, w_023_4404, w_023_4405, w_023_4407, w_023_4409, w_023_4412, w_023_4416, w_023_4418, w_023_4419, w_023_4420, w_023_4422, w_023_4423, w_023_4424, w_023_4425, w_023_4427, w_023_4428, w_023_4429, w_023_4430, w_023_4431, w_023_4432, w_023_4434, w_023_4435, w_023_4436, w_023_4437, w_023_4438, w_023_4439, w_023_4443, w_023_4445, w_023_4446, w_023_4449, w_023_4450, w_023_4451, w_023_4452, w_023_4453, w_023_4454, w_023_4456, w_023_4457, w_023_4458, w_023_4459, w_023_4461, w_023_4464, w_023_4466, w_023_4467, w_023_4468, w_023_4471, w_023_4472, w_023_4475, w_023_4477, w_023_4478, w_023_4481, w_023_4483, w_023_4484, w_023_4485, w_023_4486, w_023_4487, w_023_4488, w_023_4489, w_023_4490, w_023_4492, w_023_4494, w_023_4495, w_023_4496, w_023_4498, w_023_4500, w_023_4501, w_023_4503, w_023_4504, w_023_4505, w_023_4507, w_023_4509, w_023_4512, w_023_4515, w_023_4516, w_023_4517, w_023_4519, w_023_4520, w_023_4524, w_023_4526, w_023_4527, w_023_4528, w_023_4531, w_023_4532, w_023_4533, w_023_4534, w_023_4536, w_023_4538, w_023_4540, w_023_4545, w_023_4547, w_023_4548, w_023_4551, w_023_4553, w_023_4557, w_023_4558, w_023_4559, w_023_4560, w_023_4563, w_023_4564, w_023_4567, w_023_4568, w_023_4571, w_023_4573, w_023_4574, w_023_4575, w_023_4577, w_023_4578, w_023_4579, w_023_4580, w_023_4581, w_023_4582, w_023_4584, w_023_4586, w_023_4587, w_023_4588, w_023_4590, w_023_4591, w_023_4592, w_023_4593, w_023_4594, w_023_4595, w_023_4596, w_023_4598, w_023_4599, w_023_4600, w_023_4601, w_023_4602, w_023_4605, w_023_4610, w_023_4611, w_023_4613, w_023_4616, w_023_4619, w_023_4620, w_023_4622, w_023_4623, w_023_4624, w_023_4626, w_023_4627, w_023_4629, w_023_4630, w_023_4631, w_023_4633, w_023_4634, w_023_4635, w_023_4638, w_023_4639, w_023_4642, w_023_4643, w_023_4644, w_023_4645, w_023_4646, w_023_4647, w_023_4652, w_023_4655, w_023_4657, w_023_4659, w_023_4660, w_023_4661, w_023_4664, w_023_4665, w_023_4668, w_023_4669, w_023_4671, w_023_4674, w_023_4675, w_023_4678, w_023_4679, w_023_4680, w_023_4681, w_023_4682, w_023_4688, w_023_4689, w_023_4690, w_023_4695, w_023_4698, w_023_4699, w_023_4700, w_023_4701, w_023_4702, w_023_4703, w_023_4704, w_023_4706, w_023_4707, w_023_4709, w_023_4711, w_023_4715, w_023_4718, w_023_4719, w_023_4720, w_023_4722, w_023_4724, w_023_4725, w_023_4726, w_023_4727, w_023_4728, w_023_4729, w_023_4731, w_023_4733, w_023_4734, w_023_4735, w_023_4737, w_023_4738, w_023_4740, w_023_4741, w_023_4744, w_023_4745, w_023_4747, w_023_4749, w_023_4750, w_023_4751, w_023_4752, w_023_4753, w_023_4755, w_023_4756, w_023_4759, w_023_4760, w_023_4761, w_023_4762, w_023_4764, w_023_4765, w_023_4766, w_023_4767, w_023_4768, w_023_4769, w_023_4771, w_023_4772, w_023_4773, w_023_4774, w_023_4775, w_023_4777, w_023_4778, w_023_4780, w_023_4781, w_023_4782, w_023_4785, w_023_4786, w_023_4787, w_023_4790, w_023_4791, w_023_4794, w_023_4795, w_023_4797, w_023_4798, w_023_4799, w_023_4801, w_023_4804, w_023_4805, w_023_4806, w_023_4807, w_023_4808, w_023_4809, w_023_4810, w_023_4811, w_023_4815, w_023_4816, w_023_4817, w_023_4821, w_023_4822, w_023_4823, w_023_4824, w_023_4825, w_023_4826, w_023_4829, w_023_4830, w_023_4831, w_023_4832, w_023_4833, w_023_4834, w_023_4835, w_023_4836, w_023_4840, w_023_4841, w_023_4843, w_023_4844, w_023_4848, w_023_4849, w_023_4850, w_023_4852, w_023_4853, w_023_4857, w_023_4858, w_023_4859, w_023_4860, w_023_4861, w_023_4863, w_023_4865, w_023_4867, w_023_4868, w_023_4869, w_023_4870, w_023_4872, w_023_4873, w_023_4874, w_023_4876, w_023_4877, w_023_4879, w_023_4882, w_023_4884, w_023_4885, w_023_4887, w_023_4888, w_023_4889, w_023_4891, w_023_4892, w_023_4893, w_023_4894, w_023_4895, w_023_4896, w_023_4898, w_023_4901, w_023_4902, w_023_4903, w_023_4904, w_023_4905, w_023_4906, w_023_4907, w_023_4908, w_023_4910, w_023_4911, w_023_4912, w_023_4913, w_023_4914, w_023_4915, w_023_4916, w_023_4917, w_023_4919, w_023_4920, w_023_4921, w_023_4923, w_023_4925, w_023_4927, w_023_4928, w_023_4929, w_023_4931, w_023_4932, w_023_4934, w_023_4936, w_023_4937, w_023_4938, w_023_4939, w_023_4940, w_023_4944, w_023_4945, w_023_4947, w_023_4948, w_023_4949, w_023_4950, w_023_4951, w_023_4953, w_023_4954, w_023_4955, w_023_4956, w_023_4957, w_023_4958, w_023_4959, w_023_4960, w_023_4963, w_023_4967, w_023_4968, w_023_4969, w_023_4971, w_023_4972, w_023_4977, w_023_4979, w_023_4980, w_023_4982, w_023_4983, w_023_4986, w_023_4987, w_023_4988, w_023_4989, w_023_4990, w_023_4991, w_023_4992, w_023_4994, w_023_4995, w_023_4997, w_023_4998, w_023_4999, w_023_5001, w_023_5003, w_023_5004, w_023_5006, w_023_5009, w_023_5010, w_023_5014, w_023_5016, w_023_5017, w_023_5019, w_023_5020, w_023_5023, w_023_5025, w_023_5026, w_023_5027, w_023_5028, w_023_5031, w_023_5036, w_023_5037, w_023_5038, w_023_5039, w_023_5040, w_023_5044, w_023_5046, w_023_5047, w_023_5049, w_023_5050, w_023_5053, w_023_5054, w_023_5055, w_023_5056, w_023_5058, w_023_5059, w_023_5061, w_023_5062, w_023_5063, w_023_5066, w_023_5067, w_023_5069, w_023_5070, w_023_5072, w_023_5073, w_023_5075, w_023_5076, w_023_5077, w_023_5078, w_023_5081, w_023_5082, w_023_5083, w_023_5087, w_023_5088, w_023_5090, w_023_5091, w_023_5094, w_023_5095, w_023_5096, w_023_5097, w_023_5098, w_023_5099, w_023_5102, w_023_5103, w_023_5105, w_023_5106, w_023_5108, w_023_5111, w_023_5113, w_023_5114, w_023_5116, w_023_5117, w_023_5122, w_023_5123, w_023_5125, w_023_5126, w_023_5132, w_023_5133, w_023_5135, w_023_5136, w_023_5138, w_023_5142, w_023_5145, w_023_5146, w_023_5147, w_023_5148, w_023_5149, w_023_5153, w_023_5154, w_023_5155, w_023_5157, w_023_5158, w_023_5159, w_023_5160, w_023_5165, w_023_5169, w_023_5170, w_023_5172, w_023_5177, w_023_5179, w_023_5180, w_023_5182, w_023_5187, w_023_5188, w_023_5192, w_023_5193, w_023_5194, w_023_5195, w_023_5196, w_023_5197, w_023_5198, w_023_5200, w_023_5204, w_023_5209, w_023_5210, w_023_5211, w_023_5212, w_023_5215, w_023_5216, w_023_5217, w_023_5219, w_023_5223, w_023_5224, w_023_5225, w_023_5229, w_023_5231, w_023_5232, w_023_5233, w_023_5235, w_023_5236, w_023_5237, w_023_5238, w_023_5239, w_023_5241, w_023_5243, w_023_5244, w_023_5245, w_023_5246, w_023_5249, w_023_5250, w_023_5253, w_023_5254, w_023_5257, w_023_5258, w_023_5261, w_023_5263, w_023_5265, w_023_5266, w_023_5267, w_023_5270, w_023_5271, w_023_5272, w_023_5274, w_023_5275, w_023_5276, w_023_5279, w_023_5281, w_023_5284, w_023_5285, w_023_5286, w_023_5287, w_023_5288, w_023_5289, w_023_5290, w_023_5291, w_023_5294, w_023_5297, w_023_5298, w_023_5300, w_023_5301, w_023_5303, w_023_5305, w_023_5306, w_023_5308, w_023_5309, w_023_5310, w_023_5311, w_023_5312, w_023_5313, w_023_5314, w_023_5316, w_023_5317, w_023_5318, w_023_5319, w_023_5320, w_023_5321, w_023_5322, w_023_5323, w_023_5325, w_023_5327, w_023_5328, w_023_5329, w_023_5333, w_023_5334, w_023_5338, w_023_5339, w_023_5340, w_023_5342, w_023_5343, w_023_5345, w_023_5346, w_023_5348, w_023_5350, w_023_5353, w_023_5355, w_023_5357, w_023_5359, w_023_5360, w_023_5362, w_023_5363, w_023_5364, w_023_5365, w_023_5366, w_023_5367, w_023_5370, w_023_5371, w_023_5374, w_023_5376, w_023_5379, w_023_5382, w_023_5384, w_023_5386, w_023_5387, w_023_5390, w_023_5392, w_023_5394, w_023_5395, w_023_5397, w_023_5400, w_023_5403, w_023_5407, w_023_5410, w_023_5414, w_023_5415, w_023_5417, w_023_5418, w_023_5419, w_023_5421, w_023_5423, w_023_5424, w_023_5427, w_023_5429, w_023_5432, w_023_5433, w_023_5435, w_023_5437, w_023_5438, w_023_5439, w_023_5440, w_023_5442, w_023_5443, w_023_5444, w_023_5445, w_023_5448, w_023_5455, w_023_5456, w_023_5457, w_023_5459, w_023_5460, w_023_5461, w_023_5463, w_023_5467, w_023_5468, w_023_5469, w_023_5470, w_023_5471, w_023_5473, w_023_5474, w_023_5475, w_023_5476, w_023_5478, w_023_5479, w_023_5480, w_023_5484, w_023_5485, w_023_5487, w_023_5492, w_023_5493, w_023_5494, w_023_5498, w_023_5499, w_023_5500, w_023_5501, w_023_5502, w_023_5503, w_023_5505, w_023_5507, w_023_5510, w_023_5511, w_023_5513, w_023_5514, w_023_5515, w_023_5520, w_023_5521, w_023_5523, w_023_5527, w_023_5529, w_023_5530, w_023_5531, w_023_5532, w_023_5533, w_023_5534, w_023_5536, w_023_5537, w_023_5539, w_023_5541, w_023_5543, w_023_5546, w_023_5549, w_023_5550, w_023_5552, w_023_5553, w_023_5555, w_023_5556, w_023_5559, w_023_5560, w_023_5564, w_023_5567, w_023_5568, w_023_5569, w_023_5570, w_023_5571, w_023_5572, w_023_5575, w_023_5578, w_023_5580, w_023_5584, w_023_5587, w_023_5588, w_023_5589, w_023_5590, w_023_5592, w_023_5593, w_023_5595, w_023_5598, w_023_5599, w_023_5600, w_023_5601, w_023_5602, w_023_5604, w_023_5608, w_023_5610, w_023_5611, w_023_5612, w_023_5614, w_023_5615, w_023_5616, w_023_5619, w_023_5621, w_023_5622, w_023_5623, w_023_5624, w_023_5625, w_023_5626, w_023_5627, w_023_5630, w_023_5631, w_023_5632, w_023_5633, w_023_5634, w_023_5635, w_023_5636, w_023_5639, w_023_5640, w_023_5643, w_023_5644, w_023_5645, w_023_5646, w_023_5648, w_023_5649, w_023_5650, w_023_5651, w_023_5652, w_023_5654, w_023_5656, w_023_5657, w_023_5659, w_023_5660, w_023_5661, w_023_5662, w_023_5663, w_023_5664, w_023_5665, w_023_5667, w_023_5668, w_023_5671, w_023_5672, w_023_5673, w_023_5676, w_023_5679, w_023_5683, w_023_5684, w_023_5685, w_023_5686, w_023_5691, w_023_5692, w_023_5693, w_023_5694, w_023_5695, w_023_5696, w_023_5697, w_023_5699, w_023_5700, w_023_5703, w_023_5704, w_023_5707, w_023_5708, w_023_5709, w_023_5710, w_023_5711, w_023_5712, w_023_5713, w_023_5714, w_023_5715, w_023_5717, w_023_5718, w_023_5719, w_023_5721, w_023_5722, w_023_5723, w_023_5725, w_023_5726, w_023_5727, w_023_5728, w_023_5729, w_023_5730, w_023_5731, w_023_5733, w_023_5734, w_023_5735, w_023_5738, w_023_5739, w_023_5741, w_023_5743, w_023_5745, w_023_5746, w_023_5747, w_023_5749, w_023_5750, w_023_5752, w_023_5753, w_023_5758, w_023_5764, w_023_5765, w_023_5766, w_023_5767, w_023_5768, w_023_5770, w_023_5771, w_023_5773, w_023_5774, w_023_5776, w_023_5778, w_023_5780, w_023_5783, w_023_5787, w_023_5788, w_023_5789, w_023_5790, w_023_5791, w_023_5792, w_023_5793, w_023_5796, w_023_5802, w_023_5803, w_023_5804, w_023_5805, w_023_5806, w_023_5810, w_023_5811, w_023_5812, w_023_5813, w_023_5814, w_023_5816, w_023_5818, w_023_5819, w_023_5820, w_023_5822, w_023_5825, w_023_5827, w_023_5831, w_023_5832, w_023_5835, w_023_5840, w_023_5842, w_023_5844, w_023_5845, w_023_5846, w_023_5848, w_023_5852, w_023_5853, w_023_5854, w_023_5855, w_023_5857, w_023_5858, w_023_5861, w_023_5862, w_023_5863, w_023_5864, w_023_5867, w_023_5868, w_023_5869, w_023_5872, w_023_5873, w_023_5874, w_023_5876, w_023_5877, w_023_5879, w_023_5884, w_023_5886, w_023_5887, w_023_5888, w_023_5889, w_023_5891, w_023_5893, w_023_5894, w_023_5896, w_023_5897, w_023_5898, w_023_5899, w_023_5905, w_023_5906, w_023_5907, w_023_5909, w_023_5911, w_023_5913, w_023_5914, w_023_5915, w_023_5918, w_023_5920, w_023_5921, w_023_5923, w_023_5924, w_023_5925, w_023_5926, w_023_5929, w_023_5931, w_023_5932, w_023_5934, w_023_5935, w_023_5936, w_023_5937, w_023_5938, w_023_5939, w_023_5941, w_023_5942, w_023_5943, w_023_5944, w_023_5945, w_023_5948, w_023_5953, w_023_5954, w_023_5955, w_023_5956, w_023_5959, w_023_5960, w_023_5961, w_023_5962, w_023_5964, w_023_5965, w_023_5966, w_023_5968, w_023_5969, w_023_5972, w_023_5974, w_023_5978, w_023_5981, w_023_5983, w_023_5984, w_023_5986, w_023_5987, w_023_5988, w_023_5989, w_023_5990, w_023_5991, w_023_5992, w_023_5993, w_023_5997, w_023_5998, w_023_5999, w_023_6001, w_023_6002, w_023_6003, w_023_6004, w_023_6007, w_023_6009, w_023_6010, w_023_6012, w_023_6013, w_023_6014, w_023_6017, w_023_6020, w_023_6021, w_023_6023, w_023_6024, w_023_6025, w_023_6026, w_023_6027, w_023_6029, w_023_6031, w_023_6032, w_023_6033, w_023_6034, w_023_6035, w_023_6038, w_023_6039, w_023_6040, w_023_6041, w_023_6045, w_023_6046, w_023_6047, w_023_6050, w_023_6054, w_023_6057, w_023_6061, w_023_6062, w_023_6064, w_023_6065, w_023_6067, w_023_6068, w_023_6069, w_023_6071, w_023_6073, w_023_6074, w_023_6079, w_023_6081, w_023_6082, w_023_6085, w_023_6086, w_023_6087, w_023_6089, w_023_6092, w_023_6094, w_023_6096, w_023_6097, w_023_6098, w_023_6100, w_023_6101, w_023_6102, w_023_6103, w_023_6105, w_023_6107, w_023_6108, w_023_6109, w_023_6111, w_023_6112, w_023_6114, w_023_6115, w_023_6118, w_023_6119, w_023_6120, w_023_6121, w_023_6122, w_023_6123, w_023_6124, w_023_6125, w_023_6126, w_023_6127, w_023_6128, w_023_6129, w_023_6131, w_023_6132, w_023_6137, w_023_6139, w_023_6141, w_023_6144, w_023_6145, w_023_6148, w_023_6149, w_023_6150, w_023_6152, w_023_6154, w_023_6155, w_023_6157, w_023_6158, w_023_6163, w_023_6164, w_023_6165, w_023_6166, w_023_6167, w_023_6169, w_023_6170, w_023_6171, w_023_6172, w_023_6174, w_023_6179, w_023_6180, w_023_6181, w_023_6182, w_023_6185, w_023_6186, w_023_6187, w_023_6188, w_023_6189, w_023_6190, w_023_6191, w_023_6193, w_023_6194, w_023_6196, w_023_6197, w_023_6198, w_023_6199, w_023_6201, w_023_6202, w_023_6204, w_023_6207, w_023_6208, w_023_6209, w_023_6212, w_023_6213, w_023_6214, w_023_6215, w_023_6216, w_023_6218, w_023_6220, w_023_6221, w_023_6223, w_023_6224, w_023_6228, w_023_6229, w_023_6230, w_023_6233, w_023_6234, w_023_6235, w_023_6236, w_023_6237, w_023_6238, w_023_6240, w_023_6244, w_023_6246, w_023_6249, w_023_6250, w_023_6251, w_023_6252, w_023_6253, w_023_6254, w_023_6255, w_023_6256, w_023_6257, w_023_6259, w_023_6261, w_023_6263, w_023_6267, w_023_6268, w_023_6269, w_023_6272, w_023_6273, w_023_6274, w_023_6275, w_023_6276, w_023_6278, w_023_6281, w_023_6283, w_023_6284, w_023_6286, w_023_6287, w_023_6289, w_023_6295, w_023_6296, w_023_6298, w_023_6299, w_023_6301, w_023_6303, w_023_6305, w_023_6307, w_023_6310, w_023_6311, w_023_6313, w_023_6314, w_023_6315, w_023_6321, w_023_6324, w_023_6326, w_023_6328, w_023_6329, w_023_6330, w_023_6333, w_023_6334, w_023_6335, w_023_6336, w_023_6338, w_023_6340, w_023_6341, w_023_6343, w_023_6345, w_023_6349, w_023_6351, w_023_6352, w_023_6358, w_023_6359, w_023_6360, w_023_6362, w_023_6363, w_023_6365, w_023_6366, w_023_6367, w_023_6369, w_023_6372, w_023_6374, w_023_6376, w_023_6378, w_023_6379, w_023_6381, w_023_6383, w_023_6385, w_023_6386, w_023_6387, w_023_6388, w_023_6389, w_023_6390, w_023_6391, w_023_6392, w_023_6396, w_023_6397, w_023_6399, w_023_6400, w_023_6404, w_023_6407, w_023_6408, w_023_6409, w_023_6411, w_023_6412, w_023_6416, w_023_6417, w_023_6423, w_023_6424, w_023_6426, w_023_6427, w_023_6428, w_023_6430, w_023_6432, w_023_6433, w_023_6434, w_023_6435, w_023_6436, w_023_6437, w_023_6438, w_023_6439, w_023_6441, w_023_6442, w_023_6443, w_023_6444, w_023_6447, w_023_6453, w_023_6454, w_023_6457, w_023_6458, w_023_6459, w_023_6461, w_023_6462, w_023_6463, w_023_6466, w_023_6468, w_023_6470, w_023_6471, w_023_6473, w_023_6474, w_023_6475, w_023_6477, w_023_6479, w_023_6481, w_023_6483, w_023_6484, w_023_6485, w_023_6491, w_023_6493, w_023_6495, w_023_6498, w_023_6499, w_023_6500, w_023_6502, w_023_6503, w_023_6504, w_023_6505, w_023_6507, w_023_6508, w_023_6509, w_023_6510, w_023_6512, w_023_6513, w_023_6514, w_023_6517, w_023_6518, w_023_6519, w_023_6520, w_023_6522, w_023_6523, w_023_6524, w_023_6526, w_023_6527, w_023_6530, w_023_6531, w_023_6533, w_023_6534, w_023_6536, w_023_6538, w_023_6539, w_023_6542, w_023_6546, w_023_6548, w_023_6549, w_023_6551, w_023_6552, w_023_6554, w_023_6555, w_023_6557, w_023_6558, w_023_6560, w_023_6561, w_023_6562, w_023_6566, w_023_6567, w_023_6568, w_023_6569, w_023_6570, w_023_6573, w_023_6575, w_023_6576, w_023_6577, w_023_6578, w_023_6579, w_023_6580, w_023_6581, w_023_6589, w_023_6590, w_023_6592, w_023_6594, w_023_6595, w_023_6596, w_023_6597, w_023_6598, w_023_6600, w_023_6601, w_023_6602, w_023_6603, w_023_6604, w_023_6605, w_023_6610, w_023_6614, w_023_6615, w_023_6617, w_023_6618, w_023_6619, w_023_6620, w_023_6623, w_023_6624, w_023_6625, w_023_6626, w_023_6627, w_023_6629, w_023_6632, w_023_6636, w_023_6638, w_023_6641, w_023_6642, w_023_6643, w_023_6644, w_023_6645, w_023_6646, w_023_6647, w_023_6651, w_023_6652, w_023_6653, w_023_6655, w_023_6656, w_023_6658, w_023_6661, w_023_6664, w_023_6666, w_023_6667, w_023_6668, w_023_6669, w_023_6675, w_023_6680, w_023_6682, w_023_6683, w_023_6684, w_023_6685, w_023_6686, w_023_6687, w_023_6688, w_023_6689, w_023_6690, w_023_6692, w_023_6693, w_023_6694, w_023_6695, w_023_6696, w_023_6697, w_023_6699, w_023_6703, w_023_6706, w_023_6708, w_023_6709, w_023_6712, w_023_6713, w_023_6714, w_023_6715, w_023_6716, w_023_6717, w_023_6719, w_023_6721, w_023_6722, w_023_6723, w_023_6725, w_023_6728, w_023_6729, w_023_6730, w_023_6731, w_023_6735, w_023_6739, w_023_6740, w_023_6741, w_023_6742, w_023_6743, w_023_6746, w_023_6747, w_023_6749, w_023_6750, w_023_6751, w_023_6752, w_023_6753, w_023_6754, w_023_6759, w_023_6762, w_023_6763, w_023_6764, w_023_6767, w_023_6768, w_023_6770, w_023_6772, w_023_6773, w_023_6775, w_023_6776, w_023_6777, w_023_6780, w_023_6781, w_023_6782, w_023_6783, w_023_6784, w_023_6788, w_023_6790, w_023_6791, w_023_6793, w_023_6798, w_023_6800, w_023_6802, w_023_6803, w_023_6804, w_023_6805, w_023_6806, w_023_6807, w_023_6808, w_023_6810, w_023_6813, w_023_6814, w_023_6815, w_023_6816, w_023_6817, w_023_6819, w_023_6821, w_023_6823, w_023_6824, w_023_6826, w_023_6827, w_023_6829, w_023_6833, w_023_6834, w_023_6836, w_023_6837, w_023_6838, w_023_6839, w_023_6840, w_023_6841, w_023_6843, w_023_6844, w_023_6845, w_023_6846, w_023_6847, w_023_6848, w_023_6849, w_023_6851, w_023_6855, w_023_6856, w_023_6858, w_023_6859, w_023_6862, w_023_6863, w_023_6864, w_023_6865, w_023_6870, w_023_6871, w_023_6873, w_023_6874, w_023_6875, w_023_6877, w_023_6879, w_023_6880, w_023_6882, w_023_6883, w_023_6884, w_023_6885, w_023_6888, w_023_6892, w_023_6893, w_023_6894, w_023_6895, w_023_6897, w_023_6899, w_023_6900, w_023_6901, w_023_6903, w_023_6905, w_023_6909, w_023_6910, w_023_6914, w_023_6915, w_023_6917, w_023_6918, w_023_6919, w_023_6922, w_023_6923, w_023_6924, w_023_6925, w_023_6926, w_023_6927, w_023_6928, w_023_6929, w_023_6933, w_023_6934, w_023_6935, w_023_6936, w_023_6937, w_023_6939, w_023_6941, w_023_6945, w_023_6947, w_023_6950, w_023_6951, w_023_6955, w_023_6956, w_023_6957, w_023_6958, w_023_6959, w_023_6963, w_023_6967, w_023_6970, w_023_6971, w_023_6972, w_023_6973, w_023_6974, w_023_6977, w_023_6978, w_023_6979, w_023_6981, w_023_6983, w_023_6985, w_023_6987, w_023_6989, w_023_6991, w_023_6994, w_023_6997, w_023_6998, w_023_6999, w_023_7001, w_023_7002, w_023_7004, w_023_7005, w_023_7010, w_023_7013, w_023_7014, w_023_7018, w_023_7020, w_023_7022, w_023_7023, w_023_7024, w_023_7025, w_023_7026, w_023_7027, w_023_7028, w_023_7029, w_023_7030, w_023_7032, w_023_7033, w_023_7037, w_023_7038, w_023_7041, w_023_7043, w_023_7044, w_023_7046, w_023_7048, w_023_7049, w_023_7051, w_023_7053, w_023_7054, w_023_7055, w_023_7056, w_023_7057, w_023_7058, w_023_7059, w_023_7060, w_023_7061, w_023_7062, w_023_7063, w_023_7064, w_023_7065, w_023_7068, w_023_7069, w_023_7071, w_023_7075, w_023_7078, w_023_7080, w_023_7081, w_023_7082, w_023_7083, w_023_7085, w_023_7086, w_023_7087, w_023_7088, w_023_7092, w_023_7093, w_023_7094, w_023_7097, w_023_7099, w_023_7100, w_023_7101, w_023_7102, w_023_7105, w_023_7106, w_023_7109, w_023_7110, w_023_7112, w_023_7113, w_023_7114, w_023_7116, w_023_7119, w_023_7120, w_023_7121, w_023_7122, w_023_7125, w_023_7126, w_023_7128, w_023_7130, w_023_7131, w_023_7134, w_023_7136, w_023_7137, w_023_7138, w_023_7139, w_023_7140, w_023_7141, w_023_7146, w_023_7147, w_023_7150, w_023_7153, w_023_7154, w_023_7155, w_023_7156, w_023_7157, w_023_7158, w_023_7161, w_023_7163, w_023_7165, w_023_7167, w_023_7168, w_023_7171, w_023_7172, w_023_7173, w_023_7179, w_023_7181, w_023_7182, w_023_7184, w_023_7186, w_023_7187, w_023_7190, w_023_7191, w_023_7193, w_023_7201, w_023_7202, w_023_7206, w_023_7208, w_023_7210, w_023_7211, w_023_7212, w_023_7217, w_023_7218, w_023_7219, w_023_7220, w_023_7221, w_023_7222, w_023_7223, w_023_7224, w_023_7227, w_023_7230, w_023_7232, w_023_7233, w_023_7237, w_023_7240, w_023_7241, w_023_7242, w_023_7244, w_023_7245, w_023_7246, w_023_7248, w_023_7249, w_023_7250, w_023_7251, w_023_7254, w_023_7257, w_023_7258, w_023_7259, w_023_7261, w_023_7262, w_023_7264, w_023_7265, w_023_7267, w_023_7268, w_023_7269, w_023_7271, w_023_7272, w_023_7273, w_023_7274, w_023_7275, w_023_7276, w_023_7277, w_023_7278, w_023_7279, w_023_7280, w_023_7281, w_023_7282, w_023_7283, w_023_7284, w_023_7285, w_023_7287, w_023_7288, w_023_7289, w_023_7291, w_023_7293, w_023_7294, w_023_7295, w_023_7296, w_023_7297, w_023_7298, w_023_7299, w_023_7300, w_023_7303, w_023_7304, w_023_7305, w_023_7306, w_023_7307, w_023_7309, w_023_7310, w_023_7311, w_023_7313, w_023_7314, w_023_7318, w_023_7319, w_023_7321, w_023_7322, w_023_7323, w_023_7325, w_023_7328, w_023_7329, w_023_7331, w_023_7332, w_023_7333, w_023_7334, w_023_7335, w_023_7337, w_023_7341, w_023_7342, w_023_7344, w_023_7345, w_023_7346, w_023_7350, w_023_7352, w_023_7353, w_023_7356, w_023_7359, w_023_7360, w_023_7366, w_023_7367, w_023_7368, w_023_7369, w_023_7370, w_023_7371, w_023_7373, w_023_7374, w_023_7375, w_023_7376, w_023_7377, w_023_7378, w_023_7381, w_023_7382, w_023_7384, w_023_7386, w_023_7388, w_023_7390, w_023_7391, w_023_7392, w_023_7393, w_023_7394, w_023_7395, w_023_7396, w_023_7397, w_023_7398, w_023_7400, w_023_7403, w_023_7404, w_023_7405, w_023_7407, w_023_7408, w_023_7410, w_023_7415, w_023_7416, w_023_7417, w_023_7418, w_023_7419, w_023_7420, w_023_7424, w_023_7425, w_023_7426, w_023_7427, w_023_7428, w_023_7430, w_023_7431, w_023_7433, w_023_7435, w_023_7436, w_023_7438, w_023_7439, w_023_7442, w_023_7443, w_023_7444, w_023_7445, w_023_7446, w_023_7447, w_023_7455, w_023_7457, w_023_7459, w_023_7460, w_023_7461, w_023_7463, w_023_7465, w_023_7466, w_023_7467, w_023_7469, w_023_7473, w_023_7475, w_023_7476, w_023_7478, w_023_7481, w_023_7482, w_023_7484, w_023_7485, w_023_7486, w_023_7487, w_023_7488, w_023_7490, w_023_7491, w_023_7492, w_023_7493, w_023_7495, w_023_7498, w_023_7501, w_023_7502, w_023_7503, w_023_7505, w_023_7506, w_023_7507, w_023_7509, w_023_7510, w_023_7512, w_023_7514, w_023_7516, w_023_7519, w_023_7523, w_023_7524, w_023_7526, w_023_7527, w_023_7528, w_023_7530, w_023_7531, w_023_7532, w_023_7533, w_023_7534, w_023_7536, w_023_7537, w_023_7538, w_023_7539, w_023_7542, w_023_7543, w_023_7546, w_023_7548, w_023_7549, w_023_7550, w_023_7551, w_023_7555, w_023_7556, w_023_7558, w_023_7559, w_023_7560, w_023_7563, w_023_7564, w_023_7568, w_023_7569, w_023_7570, w_023_7571, w_023_7573, w_023_7574, w_023_7577, w_023_7578, w_023_7579, w_023_7580, w_023_7582, w_023_7583, w_023_7584, w_023_7585, w_023_7586, w_023_7587, w_023_7588, w_023_7590, w_023_7592, w_023_7594, w_023_7595, w_023_7596, w_023_7602, w_023_7604, w_023_7607, w_023_7609, w_023_7611, w_023_7612, w_023_7613, w_023_7616, w_023_7618, w_023_7620, w_023_7621, w_023_7622, w_023_7626, w_023_7627, w_023_7628, w_023_7629, w_023_7630, w_023_7631, w_023_7632, w_023_7633, w_023_7634, w_023_7635, w_023_7636, w_023_7642, w_023_7643, w_023_7644, w_023_7645, w_023_7646, w_023_7647, w_023_7649, w_023_7653, w_023_7654, w_023_7656, w_023_7657, w_023_7659, w_023_7660, w_023_7661, w_023_7662, w_023_7663, w_023_7664, w_023_7666, w_023_7669, w_023_7670, w_023_7675, w_023_7679, w_023_7681, w_023_7682, w_023_7684, w_023_7686, w_023_7687, w_023_7688, w_023_7690, w_023_7692, w_023_7695, w_023_7696, w_023_7697, w_023_7698, w_023_7699, w_023_7700, w_023_7702, w_023_7705, w_023_7706, w_023_7707, w_023_7708, w_023_7714, w_023_7717, w_023_7719, w_023_7723, w_023_7724, w_023_7725, w_023_7726, w_023_7728, w_023_7729, w_023_7733, w_023_7734, w_023_7735, w_023_7736, w_023_7737, w_023_7738, w_023_7739, w_023_7744, w_023_7745, w_023_7747, w_023_7748, w_023_7749, w_023_7750, w_023_7755, w_023_7756, w_023_7757, w_023_7758, w_023_7759, w_023_7760, w_023_7761, w_023_7763, w_023_7766, w_023_7767, w_023_7768, w_023_7769, w_023_7773, w_023_7774, w_023_7775, w_023_7776, w_023_7778, w_023_7779, w_023_7780, w_023_7783, w_023_7785, w_023_7787, w_023_7789, w_023_7790, w_023_7794, w_023_7795, w_023_7796, w_023_7798, w_023_7799, w_023_7800, w_023_7801, w_023_7803, w_023_7804, w_023_7805, w_023_7806, w_023_7811, w_023_7813, w_023_7814, w_023_7815, w_023_7816, w_023_7817, w_023_7818, w_023_7819, w_023_7820, w_023_7823, w_023_7824, w_023_7825, w_023_7827, w_023_7828, w_023_7829, w_023_7830, w_023_7831, w_023_7832, w_023_7837, w_023_7838, w_023_7839, w_023_7841, w_023_7842, w_023_7846, w_023_7847, w_023_7849, w_023_7850, w_023_7851, w_023_7853, w_023_7854, w_023_7855, w_023_7856, w_023_7857, w_023_7858, w_023_7859, w_023_7863, w_023_7865, w_023_7866, w_023_7867, w_023_7870, w_023_7871, w_023_7872, w_023_7873, w_023_7874, w_023_7876, w_023_7877, w_023_7878, w_023_7879, w_023_7880, w_023_7882, w_023_7883, w_023_7884, w_023_7886, w_023_7889, w_023_7890, w_023_7891, w_023_7893, w_023_7895, w_023_7896, w_023_7897, w_023_7898, w_023_7899, w_023_7900, w_023_7901, w_023_7902, w_023_7903, w_023_7904, w_023_7908, w_023_7910, w_023_7912, w_023_7913, w_023_7914, w_023_7915, w_023_7916, w_023_7918, w_023_7919, w_023_7920, w_023_7921, w_023_7922, w_023_7924, w_023_7928, w_023_7929, w_023_7931, w_023_7932, w_023_7933, w_023_7934, w_023_7935, w_023_7937, w_023_7938, w_023_7939, w_023_7940, w_023_7941, w_023_7943, w_023_7948, w_023_7949, w_023_7950, w_023_7952, w_023_7955, w_023_7958, w_023_7960, w_023_7962, w_023_7963, w_023_7964, w_023_7965, w_023_7967, w_023_7969, w_023_7970, w_023_7971, w_023_7972, w_023_7976, w_023_7977, w_023_7979, w_023_7980, w_023_7983, w_023_7984, w_023_7985, w_023_7989, w_023_7990, w_023_7992, w_023_7993, w_023_7994, w_023_7995, w_023_7996, w_023_7997, w_023_7999, w_023_8000, w_023_8001, w_023_8002, w_023_8004, w_023_8005, w_023_8008, w_023_8011, w_023_8013, w_023_8014, w_023_8017, w_023_8018, w_023_8019, w_023_8020, w_023_8021, w_023_8022, w_023_8024, w_023_8025, w_023_8027, w_023_8028, w_023_8029, w_023_8030, w_023_8032, w_023_8036, w_023_8041, w_023_8042, w_023_8043, w_023_8047, w_023_8049, w_023_8050, w_023_8051, w_023_8052, w_023_8054, w_023_8055, w_023_8057, w_023_8058, w_023_8061, w_023_8064, w_023_8065, w_023_8066, w_023_8068, w_023_8069, w_023_8070, w_023_8072, w_023_8075, w_023_8079, w_023_8081, w_023_8083, w_023_8086, w_023_8088, w_023_8090, w_023_8092, w_023_8093, w_023_8094, w_023_8096, w_023_8097, w_023_8098, w_023_8100, w_023_8103, w_023_8106, w_023_8107, w_023_8110, w_023_8111, w_023_8114, w_023_8115, w_023_8118, w_023_8119, w_023_8120, w_023_8122, w_023_8124, w_023_8125, w_023_8127, w_023_8129, w_023_8131, w_023_8132, w_023_8133, w_023_8134, w_023_8139, w_023_8141, w_023_8147, w_023_8148, w_023_8149, w_023_8150, w_023_8153, w_023_8154, w_023_8155, w_023_8156, w_023_8160, w_023_8161, w_023_8162, w_023_8164, w_023_8166, w_023_8167, w_023_8169, w_023_8170, w_023_8174, w_023_8176, w_023_8178, w_023_8179, w_023_8180, w_023_8182, w_023_8184, w_023_8187, w_023_8188, w_023_8189, w_023_8190, w_023_8191, w_023_8192, w_023_8193, w_023_8194, w_023_8196, w_023_8197, w_023_8198, w_023_8199, w_023_8200, w_023_8203, w_023_8204, w_023_8205, w_023_8209, w_023_8211, w_023_8213, w_023_8214, w_023_8219, w_023_8220, w_023_8227, w_023_8230, w_023_8231, w_023_8232, w_023_8234, w_023_8235, w_023_8236, w_023_8237, w_023_8238, w_023_8240, w_023_8241, w_023_8242, w_023_8244, w_023_8248, w_023_8250, w_023_8251, w_023_8252, w_023_8253, w_023_8255, w_023_8256, w_023_8257, w_023_8258, w_023_8259, w_023_8260, w_023_8261, w_023_8262, w_023_8263, w_023_8265, w_023_8270, w_023_8271, w_023_8273, w_023_8274, w_023_8275, w_023_8280, w_023_8283, w_023_8284, w_023_8285, w_023_8291, w_023_8292, w_023_8295, w_023_8296, w_023_8297, w_023_8299, w_023_8301, w_023_8304, w_023_8307, w_023_8308, w_023_8309, w_023_8310, w_023_8311, w_023_8314, w_023_8317, w_023_8318, w_023_8319, w_023_8322, w_023_8323, w_023_8325, w_023_8326, w_023_8328, w_023_8330, w_023_8331, w_023_8332, w_023_8333, w_023_8338, w_023_8339, w_023_8341, w_023_8343, w_023_8344, w_023_8345, w_023_8348, w_023_8351, w_023_8352, w_023_8355, w_023_8356, w_023_8357, w_023_8359, w_023_8361, w_023_8362, w_023_8363, w_023_8364, w_023_8365, w_023_8366, w_023_8368, w_023_8371, w_023_8373, w_023_8374, w_023_8375, w_023_8376, w_023_8377, w_023_8379, w_023_8381, w_023_8382, w_023_8383, w_023_8384, w_023_8386, w_023_8388, w_023_8390, w_023_8391, w_023_8392, w_023_8393, w_023_8395, w_023_8397, w_023_8400, w_023_8402, w_023_8403, w_023_8408, w_023_8410, w_023_8412, w_023_8414, w_023_8416, w_023_8417, w_023_8418, w_023_8421, w_023_8423, w_023_8425, w_023_8427, w_023_8428, w_023_8429, w_023_8433, w_023_8434, w_023_8436, w_023_8437, w_023_8439, w_023_8440, w_023_8442, w_023_8443, w_023_8445, w_023_8446, w_023_8447, w_023_8449, w_023_8451, w_023_8452, w_023_8453, w_023_8454, w_023_8455, w_023_8456, w_023_8459, w_023_8460, w_023_8462, w_023_8467, w_023_8470, w_023_8472, w_023_8475, w_023_8478, w_023_8480, w_023_8483, w_023_8485, w_023_8486, w_023_8490, w_023_8491, w_023_8492, w_023_8495, w_023_8496, w_023_8498, w_023_8499, w_023_8500, w_023_8504, w_023_8506, w_023_8510, w_023_8512, w_023_8513, w_023_8514, w_023_8515, w_023_8516, w_023_8517, w_023_8518, w_023_8520, w_023_8522, w_023_8524, w_023_8526, w_023_8528, w_023_8530, w_023_8531, w_023_8535, w_023_8536, w_023_8538, w_023_8542, w_023_8544, w_023_8545, w_023_8548, w_023_8549, w_023_8550, w_023_8552, w_023_8553, w_023_8554, w_023_8556, w_023_8557, w_023_8558, w_023_8560, w_023_8561, w_023_8562, w_023_8563, w_023_8565, w_023_8566, w_023_8567, w_023_8568, w_023_8569, w_023_8570, w_023_8571, w_023_8572, w_023_8573, w_023_8575, w_023_8576, w_023_8578, w_023_8579, w_023_8580, w_023_8581, w_023_8585, w_023_8586, w_023_8587, w_023_8589, w_023_8590, w_023_8591, w_023_8592, w_023_8594, w_023_8595, w_023_8596, w_023_8600, w_023_8601, w_023_8602, w_023_8605, w_023_8606, w_023_8609, w_023_8612, w_023_8615, w_023_8616, w_023_8617, w_023_8619, w_023_8621, w_023_8622, w_023_8623, w_023_8624, w_023_8627, w_023_8628, w_023_8629, w_023_8631, w_023_8632, w_023_8635, w_023_8636, w_023_8637, w_023_8639, w_023_8640, w_023_8641, w_023_8642, w_023_8643, w_023_8646, w_023_8648, w_023_8649, w_023_8650, w_023_8651, w_023_8652, w_023_8655, w_023_8656, w_023_8658, w_023_8659, w_023_8661, w_023_8666, w_023_8672, w_023_8673, w_023_8675, w_023_8676, w_023_8677, w_023_8680, w_023_8681, w_023_8682, w_023_8684, w_023_8688, w_023_8689, w_023_8691, w_023_8693, w_023_8694, w_023_8696, w_023_8699, w_023_8700, w_023_8701, w_023_8706, w_023_8707, w_023_8708, w_023_8709, w_023_8713, w_023_8714, w_023_8716, w_023_8718, w_023_8721, w_023_8722, w_023_8723, w_023_8724, w_023_8725, w_023_8728, w_023_8731, w_023_8735, w_023_8737, w_023_8739, w_023_8740, w_023_8741, w_023_8743, w_023_8744, w_023_8748, w_023_8749, w_023_8750, w_023_8752, w_023_8754, w_023_8755, w_023_8757, w_023_8761, w_023_8762, w_023_8763, w_023_8764, w_023_8766, w_023_8767, w_023_8768, w_023_8771, w_023_8772, w_023_8773, w_023_8774, w_023_8775, w_023_8776, w_023_8777, w_023_8779, w_023_8780, w_023_8781, w_023_8782, w_023_8783, w_023_8784, w_023_8785, w_023_8786, w_023_8790, w_023_8791, w_023_8792, w_023_8793, w_023_8794, w_023_8795, w_023_8796, w_023_8797, w_023_8798, w_023_8799, w_023_8800, w_023_8801, w_023_8804, w_023_8805, w_023_8806, w_023_8808, w_023_8809, w_023_8810, w_023_8811, w_023_8812, w_023_8813, w_023_8816, w_023_8817, w_023_8819, w_023_8820, w_023_8822, w_023_8824, w_023_8827, w_023_8829, w_023_8832, w_023_8833, w_023_8834, w_023_8835, w_023_8837, w_023_8841, w_023_8842, w_023_8843, w_023_8844, w_023_8849, w_023_8852, w_023_8853, w_023_8854, w_023_8855, w_023_8856, w_023_8857, w_023_8862, w_023_8863, w_023_8865, w_023_8868, w_023_8869, w_023_8871, w_023_8872, w_023_8875, w_023_8877, w_023_8878, w_023_8879, w_023_8881, w_023_8882, w_023_8884, w_023_8885, w_023_8887, w_023_8888, w_023_8889, w_023_8892, w_023_8898, w_023_8900, w_023_8902, w_023_8905, w_023_8906, w_023_8907, w_023_8908, w_023_8909, w_023_8911, w_023_8912, w_023_8914, w_023_8915, w_023_8918, w_023_8919, w_023_8920, w_023_8922, w_023_8926, w_023_8928, w_023_8929, w_023_8931, w_023_8933, w_023_8934, w_023_8936, w_023_8937, w_023_8938, w_023_8942, w_023_8944, w_023_8946, w_023_8947, w_023_8948, w_023_8951, w_023_8953, w_023_8955, w_023_8957, w_023_8958, w_023_8959, w_023_8960, w_023_8962, w_023_8966, w_023_8968, w_023_8971, w_023_8974, w_023_8976, w_023_8977, w_023_8978, w_023_8979, w_023_8981, w_023_8982, w_023_8984, w_023_8985, w_023_8988, w_023_8989, w_023_8990, w_023_8991, w_023_8992, w_023_8993, w_023_8994, w_023_8995, w_023_8996, w_023_8997, w_023_8998, w_023_9001, w_023_9004, w_023_9006, w_023_9007, w_023_9012, w_023_9013, w_023_9014, w_023_9016, w_023_9017, w_023_9019, w_023_9020, w_023_9021, w_023_9022, w_023_9025, w_023_9026, w_023_9027, w_023_9030, w_023_9031, w_023_9033, w_023_9035, w_023_9039, w_023_9040, w_023_9043, w_023_9044, w_023_9045, w_023_9046, w_023_9047, w_023_9048, w_023_9049, w_023_9051, w_023_9053, w_023_9054, w_023_9057, w_023_9058, w_023_9060, w_023_9061, w_023_9063, w_023_9064, w_023_9065, w_023_9066, w_023_9067, w_023_9068, w_023_9071, w_023_9072, w_023_9073, w_023_9075, w_023_9076, w_023_9077, w_023_9078, w_023_9079, w_023_9080, w_023_9081, w_023_9082, w_023_9083, w_023_9086, w_023_9087, w_023_9088, w_023_9089, w_023_9095, w_023_9097, w_023_9098, w_023_9102, w_023_9103, w_023_9104, w_023_9107, w_023_9109, w_023_9111, w_023_9112, w_023_9113, w_023_9116, w_023_9117, w_023_9118, w_023_9119, w_023_9120, w_023_9121, w_023_9122, w_023_9123, w_023_9127, w_023_9128, w_023_9132, w_023_9133, w_023_9136, w_023_9138, w_023_9139, w_023_9146, w_023_9147, w_023_9148, w_023_9149, w_023_9150, w_023_9152, w_023_9153, w_023_9156, w_023_9158, w_023_9159, w_023_9161, w_023_9165, w_023_9167, w_023_9169, w_023_9170, w_023_9171, w_023_9172, w_023_9173, w_023_9175, w_023_9176, w_023_9178, w_023_9179, w_023_9180, w_023_9184, w_023_9186, w_023_9188, w_023_9189, w_023_9190, w_023_9191, w_023_9192, w_023_9193, w_023_9199, w_023_9200, w_023_9201, w_023_9203, w_023_9205, w_023_9207, w_023_9209, w_023_9211, w_023_9212, w_023_9214, w_023_9215, w_023_9216, w_023_9218, w_023_9220, w_023_9221, w_023_9222, w_023_9224, w_023_9225, w_023_9227, w_023_9228, w_023_9229, w_023_9230, w_023_9231, w_023_9233, w_023_9235, w_023_9236, w_023_9237, w_023_9238, w_023_9239, w_023_9240, w_023_9242, w_023_9245, w_023_9246, w_023_9247, w_023_9249, w_023_9251, w_023_9255, w_023_9256, w_023_9258, w_023_9259, w_023_9260, w_023_9262, w_023_9263, w_023_9264, w_023_9268, w_023_9270, w_023_9272, w_023_9274, w_023_9275, w_023_9277, w_023_9281, w_023_9283, w_023_9287, w_023_9288, w_023_9289, w_023_9291, w_023_9294, w_023_9296, w_023_9297, w_023_9298, w_023_9299, w_023_9300, w_023_9301, w_023_9307, w_023_9308, w_023_9309, w_023_9311, w_023_9312, w_023_9313, w_023_9315, w_023_9317, w_023_9318, w_023_9319, w_023_9320, w_023_9321, w_023_9323, w_023_9327, w_023_9328, w_023_9329, w_023_9330, w_023_9331, w_023_9332, w_023_9333, w_023_9334, w_023_9335, w_023_9341, w_023_9342, w_023_9343, w_023_9345, w_023_9346, w_023_9349, w_023_9351, w_023_9352, w_023_9355, w_023_9356, w_023_9357, w_023_9361, w_023_9364, w_023_9366, w_023_9367, w_023_9368, w_023_9372, w_023_9373, w_023_9374, w_023_9375, w_023_9376, w_023_9377, w_023_9378, w_023_9380, w_023_9381, w_023_9382, w_023_9383, w_023_9385, w_023_9392, w_023_9395, w_023_9398, w_023_9402, w_023_9403, w_023_9404, w_023_9405, w_023_9406, w_023_9407, w_023_9408, w_023_9409, w_023_9410, w_023_9413, w_023_9416, w_023_9417, w_023_9418, w_023_9419, w_023_9420, w_023_9423, w_023_9426, w_023_9428, w_023_9431, w_023_9435, w_023_9437, w_023_9439, w_023_9440, w_023_9441, w_023_9442, w_023_9443, w_023_9446, w_023_9451, w_023_9452, w_023_9453, w_023_9454, w_023_9455, w_023_9457, w_023_9458, w_023_9460, w_023_9461, w_023_9462, w_023_9466, w_023_9467, w_023_9468, w_023_9469, w_023_9470, w_023_9471, w_023_9472, w_023_9474, w_023_9475, w_023_9476, w_023_9477, w_023_9478, w_023_9479, w_023_9481, w_023_9483;
  wire w_024_000, w_024_002, w_024_003, w_024_004, w_024_005, w_024_006, w_024_008, w_024_009, w_024_010, w_024_012, w_024_013, w_024_014, w_024_015, w_024_016, w_024_017, w_024_018, w_024_019, w_024_020, w_024_021, w_024_022, w_024_023, w_024_024, w_024_025, w_024_026, w_024_027, w_024_028, w_024_030, w_024_031, w_024_032, w_024_033, w_024_034, w_024_035, w_024_037, w_024_038, w_024_039, w_024_040, w_024_041, w_024_042, w_024_043, w_024_044, w_024_045, w_024_046, w_024_047, w_024_048, w_024_049, w_024_050, w_024_051, w_024_053, w_024_054, w_024_055, w_024_056, w_024_057, w_024_058, w_024_059, w_024_060, w_024_061, w_024_062, w_024_063, w_024_064, w_024_065, w_024_066, w_024_067, w_024_068, w_024_069, w_024_070, w_024_071, w_024_072, w_024_074, w_024_075, w_024_076, w_024_077, w_024_078, w_024_079, w_024_080, w_024_081, w_024_082, w_024_083, w_024_084, w_024_085, w_024_086, w_024_088, w_024_089, w_024_090, w_024_091, w_024_092, w_024_093, w_024_094, w_024_095, w_024_096, w_024_097, w_024_098, w_024_099, w_024_100, w_024_101, w_024_103, w_024_104, w_024_105, w_024_106, w_024_107, w_024_108, w_024_109, w_024_110, w_024_111, w_024_112, w_024_113, w_024_114, w_024_115, w_024_116, w_024_117, w_024_118, w_024_119, w_024_120, w_024_121, w_024_122, w_024_124, w_024_127, w_024_128, w_024_129, w_024_130, w_024_131, w_024_132, w_024_133, w_024_134, w_024_135, w_024_136, w_024_137, w_024_138, w_024_139, w_024_140, w_024_141, w_024_142, w_024_143, w_024_144, w_024_145, w_024_146, w_024_147, w_024_148, w_024_149, w_024_150, w_024_151, w_024_152, w_024_153, w_024_154, w_024_155, w_024_156, w_024_157, w_024_158, w_024_159, w_024_160, w_024_161, w_024_162, w_024_163, w_024_164, w_024_165, w_024_166, w_024_168, w_024_169, w_024_170, w_024_171, w_024_172, w_024_174, w_024_175, w_024_176, w_024_178, w_024_179, w_024_180, w_024_181, w_024_182, w_024_183, w_024_184, w_024_185, w_024_186, w_024_187, w_024_188, w_024_190, w_024_191, w_024_192, w_024_193, w_024_194, w_024_195, w_024_196, w_024_197, w_024_198, w_024_199, w_024_200, w_024_201, w_024_202, w_024_203, w_024_204, w_024_205, w_024_206, w_024_207, w_024_208, w_024_209, w_024_210, w_024_211, w_024_213, w_024_214, w_024_215, w_024_217, w_024_218, w_024_219, w_024_221, w_024_222, w_024_223, w_024_224, w_024_225, w_024_226, w_024_227, w_024_228, w_024_229, w_024_230, w_024_231, w_024_232, w_024_233, w_024_235, w_024_237, w_024_238, w_024_239, w_024_240, w_024_241, w_024_242, w_024_243, w_024_244, w_024_245, w_024_246, w_024_247, w_024_248, w_024_249, w_024_250, w_024_251, w_024_252, w_024_253, w_024_254, w_024_255, w_024_256, w_024_257, w_024_258, w_024_259, w_024_260, w_024_261, w_024_262, w_024_263, w_024_264, w_024_265, w_024_266, w_024_267, w_024_268, w_024_269, w_024_270, w_024_271, w_024_272, w_024_273, w_024_274, w_024_275, w_024_276, w_024_278, w_024_279, w_024_280, w_024_281, w_024_282, w_024_283, w_024_284, w_024_285, w_024_286, w_024_287, w_024_288, w_024_289, w_024_290, w_024_291, w_024_292, w_024_293, w_024_294, w_024_296, w_024_297, w_024_298, w_024_299, w_024_300, w_024_301, w_024_302, w_024_303, w_024_304, w_024_305, w_024_306, w_024_307, w_024_308, w_024_309, w_024_310, w_024_311, w_024_312, w_024_313, w_024_314, w_024_315, w_024_316, w_024_318, w_024_319, w_024_320, w_024_321, w_024_322, w_024_323, w_024_324, w_024_325, w_024_326, w_024_327, w_024_328, w_024_329, w_024_330, w_024_332, w_024_333, w_024_334, w_024_335, w_024_337, w_024_338, w_024_339, w_024_340, w_024_341, w_024_342, w_024_343, w_024_345, w_024_346, w_024_347, w_024_348, w_024_349, w_024_350, w_024_351, w_024_352, w_024_353, w_024_355, w_024_356, w_024_357, w_024_358, w_024_359, w_024_360, w_024_361, w_024_362, w_024_363, w_024_364, w_024_365, w_024_366, w_024_367, w_024_368, w_024_369, w_024_370, w_024_371, w_024_372, w_024_373, w_024_374, w_024_375, w_024_376, w_024_377, w_024_378, w_024_379, w_024_380, w_024_381, w_024_382, w_024_383, w_024_384, w_024_385, w_024_386, w_024_387, w_024_388, w_024_389, w_024_391, w_024_393, w_024_394, w_024_395, w_024_396, w_024_397, w_024_398, w_024_399, w_024_400, w_024_401, w_024_402, w_024_403, w_024_404, w_024_406, w_024_407, w_024_408, w_024_409, w_024_410, w_024_411, w_024_412, w_024_413, w_024_414, w_024_415, w_024_416, w_024_417, w_024_418, w_024_421, w_024_422, w_024_423, w_024_424, w_024_425, w_024_426, w_024_427, w_024_428, w_024_429, w_024_430, w_024_431, w_024_433, w_024_434, w_024_435, w_024_436, w_024_437, w_024_438, w_024_439, w_024_440, w_024_441, w_024_442, w_024_443, w_024_444, w_024_445, w_024_446, w_024_447, w_024_448, w_024_449, w_024_450, w_024_451, w_024_452, w_024_453, w_024_454, w_024_455, w_024_456, w_024_457, w_024_458, w_024_459, w_024_461, w_024_462, w_024_463, w_024_464, w_024_465, w_024_466, w_024_467, w_024_468, w_024_470, w_024_471, w_024_472, w_024_474, w_024_475, w_024_476, w_024_477, w_024_478, w_024_479, w_024_480, w_024_481, w_024_482, w_024_483, w_024_485, w_024_486, w_024_487, w_024_488, w_024_489, w_024_491, w_024_492, w_024_493, w_024_494, w_024_495, w_024_496, w_024_497, w_024_499, w_024_500, w_024_502, w_024_504, w_024_505, w_024_506, w_024_507, w_024_508, w_024_509, w_024_510, w_024_512, w_024_513, w_024_514, w_024_515, w_024_516, w_024_517, w_024_518, w_024_519, w_024_520, w_024_521, w_024_522, w_024_523, w_024_524, w_024_525, w_024_526, w_024_527, w_024_528, w_024_529, w_024_530, w_024_531, w_024_532, w_024_533, w_024_534, w_024_535, w_024_536, w_024_537, w_024_538, w_024_539, w_024_540, w_024_541, w_024_543, w_024_544, w_024_545, w_024_546, w_024_547, w_024_548, w_024_549, w_024_550, w_024_551, w_024_553, w_024_554, w_024_555, w_024_556, w_024_557, w_024_558, w_024_559, w_024_560, w_024_561, w_024_562, w_024_563, w_024_564, w_024_565, w_024_566, w_024_567, w_024_568, w_024_569, w_024_570, w_024_571, w_024_572, w_024_573, w_024_574, w_024_575, w_024_576, w_024_577, w_024_579, w_024_580, w_024_581, w_024_582, w_024_583, w_024_584, w_024_585, w_024_586, w_024_587, w_024_588, w_024_589, w_024_590, w_024_592, w_024_593, w_024_594, w_024_595, w_024_596, w_024_597, w_024_598, w_024_599, w_024_600, w_024_601, w_024_602, w_024_604, w_024_605, w_024_606, w_024_607, w_024_610, w_024_611, w_024_612, w_024_614, w_024_615, w_024_616, w_024_618, w_024_619, w_024_620, w_024_622, w_024_624, w_024_625, w_024_626, w_024_627, w_024_629, w_024_630, w_024_631, w_024_632, w_024_633, w_024_635, w_024_636, w_024_637, w_024_638, w_024_640, w_024_641, w_024_643, w_024_645, w_024_646, w_024_647, w_024_648, w_024_649, w_024_651, w_024_652, w_024_653, w_024_654, w_024_655, w_024_656, w_024_657, w_024_658, w_024_659, w_024_660, w_024_661, w_024_662, w_024_663, w_024_664, w_024_665, w_024_666, w_024_667, w_024_668, w_024_669, w_024_670, w_024_671, w_024_672, w_024_673, w_024_674, w_024_675, w_024_676, w_024_677, w_024_678, w_024_679, w_024_680, w_024_682, w_024_683, w_024_684, w_024_685, w_024_686, w_024_687, w_024_688, w_024_689, w_024_690, w_024_691, w_024_692, w_024_693, w_024_694, w_024_695, w_024_696, w_024_697, w_024_698, w_024_699, w_024_700, w_024_701, w_024_703, w_024_704, w_024_705, w_024_706, w_024_707, w_024_708, w_024_709, w_024_710, w_024_711, w_024_713, w_024_714, w_024_715, w_024_716, w_024_717, w_024_718, w_024_719, w_024_720, w_024_721, w_024_722, w_024_723, w_024_724, w_024_725, w_024_726, w_024_727, w_024_728, w_024_729, w_024_730, w_024_731, w_024_732, w_024_733, w_024_734, w_024_735, w_024_736, w_024_737, w_024_738, w_024_739, w_024_740, w_024_741, w_024_742, w_024_743, w_024_744, w_024_745, w_024_746, w_024_747, w_024_748, w_024_749, w_024_750, w_024_751, w_024_752, w_024_753, w_024_754, w_024_755, w_024_756, w_024_757, w_024_758, w_024_759, w_024_760, w_024_761, w_024_762, w_024_763, w_024_764, w_024_765, w_024_766, w_024_767, w_024_768, w_024_769, w_024_770, w_024_771, w_024_772, w_024_774, w_024_775, w_024_776, w_024_777, w_024_778, w_024_779, w_024_780, w_024_781, w_024_782, w_024_783, w_024_784, w_024_785, w_024_786, w_024_787, w_024_788, w_024_789, w_024_790, w_024_791, w_024_792, w_024_793, w_024_794, w_024_795, w_024_796, w_024_797, w_024_798, w_024_799, w_024_800, w_024_801, w_024_802, w_024_803, w_024_804, w_024_805, w_024_806, w_024_807, w_024_808, w_024_809, w_024_810, w_024_811, w_024_812, w_024_813, w_024_814, w_024_815, w_024_817, w_024_818, w_024_819, w_024_821, w_024_822, w_024_823, w_024_824, w_024_825, w_024_826, w_024_827, w_024_828, w_024_829, w_024_830, w_024_831, w_024_832, w_024_833, w_024_834, w_024_835, w_024_836, w_024_837, w_024_838, w_024_839, w_024_840, w_024_841, w_024_842, w_024_844, w_024_845, w_024_846, w_024_847, w_024_848, w_024_849, w_024_850, w_024_851, w_024_852, w_024_853, w_024_854, w_024_855, w_024_856, w_024_857, w_024_858, w_024_859, w_024_860, w_024_861, w_024_862, w_024_863, w_024_864, w_024_865, w_024_866, w_024_867, w_024_868, w_024_869, w_024_870, w_024_871, w_024_873, w_024_874, w_024_875, w_024_876, w_024_877, w_024_878, w_024_879, w_024_880, w_024_882, w_024_883, w_024_884, w_024_885, w_024_886, w_024_887, w_024_888, w_024_889, w_024_890, w_024_891, w_024_892, w_024_893, w_024_894, w_024_895, w_024_897, w_024_898, w_024_899, w_024_900, w_024_901, w_024_902, w_024_903, w_024_904, w_024_905, w_024_907, w_024_908, w_024_909, w_024_911, w_024_912, w_024_913, w_024_914, w_024_915, w_024_917, w_024_918, w_024_919, w_024_920, w_024_921, w_024_922, w_024_923, w_024_924, w_024_925, w_024_926, w_024_927, w_024_928, w_024_930, w_024_931, w_024_932, w_024_933, w_024_934, w_024_935, w_024_936, w_024_937, w_024_938, w_024_939, w_024_941, w_024_942, w_024_943, w_024_944, w_024_945, w_024_946, w_024_947, w_024_948, w_024_949, w_024_950, w_024_951, w_024_952, w_024_953, w_024_954, w_024_955, w_024_956, w_024_957, w_024_958, w_024_959, w_024_960, w_024_961, w_024_962, w_024_963, w_024_964, w_024_965, w_024_966, w_024_967, w_024_968, w_024_969, w_024_970, w_024_971, w_024_972, w_024_973, w_024_974, w_024_975, w_024_977, w_024_978, w_024_979, w_024_980, w_024_981, w_024_982, w_024_984, w_024_985, w_024_986, w_024_987, w_024_988, w_024_989, w_024_990, w_024_992, w_024_994, w_024_995, w_024_996, w_024_997, w_024_998, w_024_999, w_024_1002, w_024_1003, w_024_1004, w_024_1005, w_024_1006, w_024_1007, w_024_1008, w_024_1009, w_024_1010, w_024_1011, w_024_1012, w_024_1013, w_024_1014, w_024_1015, w_024_1016, w_024_1017, w_024_1018, w_024_1019, w_024_1020, w_024_1021, w_024_1022, w_024_1024, w_024_1025, w_024_1026, w_024_1027, w_024_1028, w_024_1029, w_024_1030, w_024_1031, w_024_1032, w_024_1033, w_024_1034, w_024_1035, w_024_1036, w_024_1037, w_024_1038, w_024_1039, w_024_1040, w_024_1041, w_024_1042, w_024_1043, w_024_1044, w_024_1045, w_024_1046, w_024_1047, w_024_1048, w_024_1049, w_024_1050, w_024_1051, w_024_1052, w_024_1053, w_024_1054, w_024_1055, w_024_1056, w_024_1057, w_024_1058, w_024_1059, w_024_1060, w_024_1061, w_024_1062, w_024_1063, w_024_1064, w_024_1065, w_024_1066, w_024_1067, w_024_1068, w_024_1070, w_024_1071, w_024_1072, w_024_1073, w_024_1074, w_024_1075, w_024_1076, w_024_1077, w_024_1078, w_024_1079, w_024_1080, w_024_1081, w_024_1082, w_024_1083, w_024_1084, w_024_1085, w_024_1086, w_024_1087, w_024_1088, w_024_1089, w_024_1090, w_024_1091, w_024_1092, w_024_1093, w_024_1095, w_024_1096, w_024_1097, w_024_1098, w_024_1099, w_024_1100, w_024_1102, w_024_1103, w_024_1104, w_024_1106, w_024_1107, w_024_1108, w_024_1109, w_024_1110, w_024_1111, w_024_1112, w_024_1113, w_024_1114, w_024_1115, w_024_1116, w_024_1118, w_024_1119, w_024_1120, w_024_1121, w_024_1123, w_024_1124, w_024_1126, w_024_1127, w_024_1128, w_024_1129, w_024_1130, w_024_1131, w_024_1132, w_024_1133, w_024_1134, w_024_1135, w_024_1136, w_024_1137, w_024_1138, w_024_1139, w_024_1140, w_024_1141, w_024_1142, w_024_1143, w_024_1144, w_024_1145, w_024_1146, w_024_1147, w_024_1148, w_024_1149, w_024_1150, w_024_1151, w_024_1153, w_024_1154, w_024_1155, w_024_1156, w_024_1159, w_024_1160, w_024_1161, w_024_1162, w_024_1163, w_024_1164, w_024_1165, w_024_1166, w_024_1167, w_024_1168, w_024_1169, w_024_1170, w_024_1171, w_024_1172, w_024_1173, w_024_1174, w_024_1175, w_024_1176, w_024_1177, w_024_1178, w_024_1179, w_024_1180, w_024_1181, w_024_1182, w_024_1183, w_024_1184, w_024_1185, w_024_1186, w_024_1187, w_024_1189, w_024_1190, w_024_1191, w_024_1192, w_024_1193, w_024_1194, w_024_1195, w_024_1196, w_024_1197, w_024_1199, w_024_1200, w_024_1201, w_024_1202, w_024_1203, w_024_1204, w_024_1205, w_024_1207, w_024_1209, w_024_1210, w_024_1211, w_024_1213, w_024_1214, w_024_1215, w_024_1216, w_024_1217, w_024_1218, w_024_1219, w_024_1220, w_024_1221, w_024_1222, w_024_1223, w_024_1224, w_024_1225, w_024_1226, w_024_1227, w_024_1228, w_024_1230, w_024_1231, w_024_1232, w_024_1233, w_024_1234, w_024_1235, w_024_1236, w_024_1237, w_024_1238, w_024_1240, w_024_1242, w_024_1243, w_024_1244, w_024_1245, w_024_1247, w_024_1248, w_024_1249, w_024_1250, w_024_1251, w_024_1252, w_024_1253, w_024_1254, w_024_1255, w_024_1256, w_024_1257, w_024_1258, w_024_1262, w_024_1263, w_024_1264, w_024_1265, w_024_1266, w_024_1267, w_024_1268, w_024_1269, w_024_1270, w_024_1271, w_024_1272, w_024_1273, w_024_1274, w_024_1275, w_024_1276, w_024_1277, w_024_1278, w_024_1279, w_024_1280, w_024_1281, w_024_1282, w_024_1284, w_024_1285, w_024_1287, w_024_1288, w_024_1289, w_024_1290, w_024_1291, w_024_1293, w_024_1294, w_024_1295, w_024_1296, w_024_1297, w_024_1298, w_024_1299, w_024_1300, w_024_1301, w_024_1302, w_024_1303, w_024_1304, w_024_1305, w_024_1309, w_024_1310, w_024_1311, w_024_1312, w_024_1313, w_024_1314, w_024_1315, w_024_1316, w_024_1317, w_024_1318, w_024_1319, w_024_1320, w_024_1321, w_024_1323, w_024_1324, w_024_1325, w_024_1326, w_024_1327, w_024_1328, w_024_1329, w_024_1330, w_024_1331, w_024_1332, w_024_1333, w_024_1334, w_024_1335, w_024_1336, w_024_1337, w_024_1338, w_024_1339, w_024_1340, w_024_1342, w_024_1343, w_024_1344, w_024_1345, w_024_1346, w_024_1348, w_024_1349, w_024_1350, w_024_1351, w_024_1352, w_024_1354, w_024_1355, w_024_1356, w_024_1358, w_024_1359, w_024_1361, w_024_1362, w_024_1363, w_024_1364, w_024_1365, w_024_1366, w_024_1369, w_024_1370, w_024_1372, w_024_1373, w_024_1374, w_024_1375, w_024_1376, w_024_1378, w_024_1379, w_024_1380, w_024_1381, w_024_1382, w_024_1383, w_024_1384, w_024_1385, w_024_1386, w_024_1387, w_024_1388, w_024_1389, w_024_1390, w_024_1391, w_024_1392, w_024_1393, w_024_1395, w_024_1396, w_024_1397, w_024_1398, w_024_1399, w_024_1400, w_024_1402, w_024_1403, w_024_1404, w_024_1405, w_024_1406, w_024_1407, w_024_1409, w_024_1410, w_024_1411, w_024_1413, w_024_1414, w_024_1415, w_024_1416, w_024_1419, w_024_1422, w_024_1423, w_024_1425, w_024_1426, w_024_1427, w_024_1428, w_024_1431, w_024_1432, w_024_1433, w_024_1434, w_024_1435, w_024_1436, w_024_1437, w_024_1438, w_024_1439, w_024_1440, w_024_1441, w_024_1442, w_024_1443, w_024_1444, w_024_1445, w_024_1446, w_024_1447, w_024_1448, w_024_1449, w_024_1450, w_024_1451, w_024_1452, w_024_1453, w_024_1454, w_024_1456, w_024_1457, w_024_1459, w_024_1460, w_024_1461, w_024_1462, w_024_1463, w_024_1464, w_024_1465, w_024_1466, w_024_1467, w_024_1468, w_024_1470, w_024_1471, w_024_1472, w_024_1474, w_024_1475, w_024_1477, w_024_1478, w_024_1480, w_024_1482, w_024_1483, w_024_1485, w_024_1486, w_024_1487, w_024_1488, w_024_1489, w_024_1490, w_024_1491, w_024_1492, w_024_1493, w_024_1494, w_024_1495, w_024_1496, w_024_1497, w_024_1498, w_024_1499, w_024_1501, w_024_1502, w_024_1503, w_024_1506, w_024_1507, w_024_1508, w_024_1509, w_024_1510, w_024_1511, w_024_1512, w_024_1513, w_024_1514, w_024_1515, w_024_1516, w_024_1519, w_024_1520, w_024_1521, w_024_1524, w_024_1525, w_024_1526, w_024_1527, w_024_1528, w_024_1529, w_024_1530, w_024_1531, w_024_1532, w_024_1533, w_024_1534, w_024_1535, w_024_1536, w_024_1538, w_024_1539, w_024_1541, w_024_1542, w_024_1543, w_024_1544, w_024_1545, w_024_1546, w_024_1549, w_024_1550, w_024_1551, w_024_1552, w_024_1553, w_024_1554, w_024_1555, w_024_1556, w_024_1558, w_024_1559, w_024_1560, w_024_1561, w_024_1562, w_024_1563, w_024_1564, w_024_1565, w_024_1566, w_024_1567, w_024_1568, w_024_1569, w_024_1570, w_024_1571, w_024_1572, w_024_1573, w_024_1574, w_024_1576, w_024_1578, w_024_1579, w_024_1580, w_024_1581, w_024_1582, w_024_1583, w_024_1584, w_024_1585, w_024_1586, w_024_1588, w_024_1589, w_024_1590, w_024_1591, w_024_1592, w_024_1594, w_024_1596, w_024_1598, w_024_1599, w_024_1600, w_024_1601, w_024_1602, w_024_1603, w_024_1604, w_024_1606, w_024_1607, w_024_1608, w_024_1612, w_024_1613, w_024_1614, w_024_1616, w_024_1617, w_024_1618, w_024_1619, w_024_1620, w_024_1621, w_024_1623, w_024_1624, w_024_1626, w_024_1627, w_024_1629, w_024_1630, w_024_1634, w_024_1635, w_024_1636, w_024_1637, w_024_1638, w_024_1639, w_024_1640, w_024_1641, w_024_1642, w_024_1643, w_024_1644, w_024_1645, w_024_1646, w_024_1647, w_024_1648, w_024_1649, w_024_1650, w_024_1651, w_024_1652, w_024_1653, w_024_1654, w_024_1655, w_024_1656, w_024_1657, w_024_1658, w_024_1659, w_024_1660, w_024_1661, w_024_1662, w_024_1663, w_024_1664, w_024_1667, w_024_1669, w_024_1672, w_024_1674, w_024_1675, w_024_1676, w_024_1679, w_024_1680, w_024_1681, w_024_1682, w_024_1683, w_024_1684, w_024_1685, w_024_1686, w_024_1688, w_024_1689, w_024_1692, w_024_1693, w_024_1694, w_024_1695, w_024_1696, w_024_1697, w_024_1698, w_024_1699, w_024_1700, w_024_1701, w_024_1702, w_024_1703, w_024_1704, w_024_1705, w_024_1706, w_024_1707, w_024_1708, w_024_1711, w_024_1712, w_024_1713, w_024_1714, w_024_1716, w_024_1717, w_024_1718, w_024_1719, w_024_1720, w_024_1721, w_024_1722, w_024_1723, w_024_1724, w_024_1725, w_024_1726, w_024_1727, w_024_1728, w_024_1729, w_024_1731, w_024_1732, w_024_1735, w_024_1737, w_024_1738, w_024_1739, w_024_1740, w_024_1742, w_024_1743, w_024_1744, w_024_1745, w_024_1746, w_024_1748, w_024_1749, w_024_1750, w_024_1751, w_024_1752, w_024_1753, w_024_1754, w_024_1755, w_024_1756, w_024_1757, w_024_1758, w_024_1759, w_024_1760, w_024_1761, w_024_1762, w_024_1763, w_024_1764, w_024_1766, w_024_1767, w_024_1769, w_024_1770, w_024_1771, w_024_1772, w_024_1773, w_024_1775, w_024_1776, w_024_1777, w_024_1778, w_024_1779, w_024_1780, w_024_1781, w_024_1782, w_024_1783, w_024_1785, w_024_1787, w_024_1788, w_024_1790, w_024_1792, w_024_1794, w_024_1795, w_024_1797, w_024_1798, w_024_1800, w_024_1801, w_024_1802, w_024_1803, w_024_1804, w_024_1806, w_024_1807, w_024_1809, w_024_1810, w_024_1811, w_024_1812, w_024_1813, w_024_1814, w_024_1815, w_024_1816, w_024_1818, w_024_1820, w_024_1824, w_024_1826, w_024_1827, w_024_1829, w_024_1830, w_024_1831, w_024_1832, w_024_1833, w_024_1834, w_024_1836, w_024_1837, w_024_1838, w_024_1839, w_024_1840, w_024_1841, w_024_1843, w_024_1844, w_024_1845, w_024_1846, w_024_1847, w_024_1849, w_024_1850, w_024_1851, w_024_1853, w_024_1854, w_024_1855, w_024_1857, w_024_1859, w_024_1860, w_024_1861, w_024_1862, w_024_1863, w_024_1865, w_024_1867, w_024_1868, w_024_1869, w_024_1870, w_024_1871, w_024_1872, w_024_1873, w_024_1874, w_024_1875, w_024_1876, w_024_1879, w_024_1880, w_024_1882, w_024_1884, w_024_1885, w_024_1886, w_024_1888, w_024_1889, w_024_1890, w_024_1891, w_024_1892, w_024_1893, w_024_1894, w_024_1896, w_024_1897, w_024_1899, w_024_1900, w_024_1901, w_024_1902, w_024_1903, w_024_1905, w_024_1906, w_024_1908, w_024_1909, w_024_1910, w_024_1911, w_024_1912, w_024_1913, w_024_1916, w_024_1917, w_024_1918, w_024_1919, w_024_1920, w_024_1921, w_024_1922, w_024_1923, w_024_1924, w_024_1925, w_024_1926, w_024_1927, w_024_1928, w_024_1929, w_024_1930, w_024_1931, w_024_1933, w_024_1935, w_024_1937, w_024_1938, w_024_1940, w_024_1942, w_024_1943, w_024_1944, w_024_1947, w_024_1948, w_024_1950, w_024_1951, w_024_1952, w_024_1954, w_024_1955, w_024_1957, w_024_1958, w_024_1959, w_024_1960, w_024_1961, w_024_1962, w_024_1964, w_024_1965, w_024_1966, w_024_1967, w_024_1969, w_024_1970, w_024_1971, w_024_1972, w_024_1973, w_024_1974, w_024_1977, w_024_1978, w_024_1980, w_024_1981, w_024_1982, w_024_1983, w_024_1984, w_024_1985, w_024_1986, w_024_1987, w_024_1988, w_024_1989, w_024_1990, w_024_1991, w_024_1993, w_024_1994, w_024_1995, w_024_1997, w_024_1998, w_024_2000, w_024_2001, w_024_2002, w_024_2003, w_024_2006, w_024_2008, w_024_2009, w_024_2010, w_024_2011, w_024_2013, w_024_2014, w_024_2016, w_024_2019, w_024_2021, w_024_2023, w_024_2024, w_024_2025, w_024_2026, w_024_2027, w_024_2028, w_024_2029, w_024_2030, w_024_2031, w_024_2032, w_024_2033, w_024_2034, w_024_2035, w_024_2036, w_024_2037, w_024_2038, w_024_2039, w_024_2040, w_024_2042, w_024_2044, w_024_2045, w_024_2046, w_024_2047, w_024_2048, w_024_2049, w_024_2050, w_024_2051, w_024_2052, w_024_2053, w_024_2054, w_024_2055, w_024_2058, w_024_2059, w_024_2060, w_024_2062, w_024_2063, w_024_2064, w_024_2065, w_024_2068, w_024_2069, w_024_2070, w_024_2071, w_024_2072, w_024_2073, w_024_2075, w_024_2076, w_024_2077, w_024_2078, w_024_2079, w_024_2080, w_024_2081, w_024_2082, w_024_2083, w_024_2084, w_024_2086, w_024_2087, w_024_2088, w_024_2089, w_024_2090, w_024_2091, w_024_2092, w_024_2093, w_024_2094, w_024_2097, w_024_2098, w_024_2099, w_024_2101, w_024_2102, w_024_2103, w_024_2104, w_024_2105, w_024_2106, w_024_2107, w_024_2108, w_024_2109, w_024_2110, w_024_2111, w_024_2113, w_024_2114, w_024_2116, w_024_2117, w_024_2118, w_024_2119, w_024_2120, w_024_2122, w_024_2123, w_024_2124, w_024_2125, w_024_2126, w_024_2129, w_024_2130, w_024_2132, w_024_2133, w_024_2134, w_024_2135, w_024_2136, w_024_2137, w_024_2138, w_024_2139, w_024_2140, w_024_2142, w_024_2143, w_024_2144, w_024_2145, w_024_2146, w_024_2148, w_024_2151, w_024_2153, w_024_2154, w_024_2155, w_024_2156, w_024_2157, w_024_2158, w_024_2159, w_024_2161, w_024_2162, w_024_2163, w_024_2164, w_024_2165, w_024_2166, w_024_2167, w_024_2168, w_024_2169, w_024_2171, w_024_2173, w_024_2174, w_024_2176, w_024_2177, w_024_2180, w_024_2181, w_024_2182, w_024_2185, w_024_2186, w_024_2187, w_024_2188, w_024_2189, w_024_2190, w_024_2191, w_024_2192, w_024_2193, w_024_2194, w_024_2195, w_024_2197, w_024_2199, w_024_2201, w_024_2202, w_024_2205, w_024_2206, w_024_2207, w_024_2208, w_024_2209, w_024_2210, w_024_2213, w_024_2214, w_024_2215, w_024_2216, w_024_2217, w_024_2218, w_024_2219, w_024_2220, w_024_2221, w_024_2222, w_024_2223, w_024_2225, w_024_2226, w_024_2227, w_024_2228, w_024_2229, w_024_2230, w_024_2231, w_024_2232, w_024_2233, w_024_2234, w_024_2235, w_024_2237, w_024_2238, w_024_2239, w_024_2240, w_024_2241, w_024_2242, w_024_2243, w_024_2245, w_024_2246, w_024_2247, w_024_2248, w_024_2249, w_024_2250, w_024_2251, w_024_2252, w_024_2254, w_024_2255, w_024_2256, w_024_2257, w_024_2258, w_024_2259, w_024_2260, w_024_2261, w_024_2262, w_024_2264, w_024_2266, w_024_2267, w_024_2270, w_024_2271, w_024_2272, w_024_2273, w_024_2274, w_024_2275, w_024_2276, w_024_2278, w_024_2279, w_024_2281, w_024_2283, w_024_2285, w_024_2286, w_024_2287, w_024_2289, w_024_2290, w_024_2291, w_024_2294, w_024_2295, w_024_2299, w_024_2300, w_024_2301, w_024_2302, w_024_2303, w_024_2304, w_024_2305, w_024_2306, w_024_2307, w_024_2309, w_024_2310, w_024_2312, w_024_2313, w_024_2314, w_024_2315, w_024_2317, w_024_2319, w_024_2320, w_024_2322, w_024_2323, w_024_2324, w_024_2325, w_024_2326, w_024_2327, w_024_2329, w_024_2330, w_024_2331, w_024_2332, w_024_2333, w_024_2335, w_024_2337, w_024_2338, w_024_2339, w_024_2340, w_024_2341, w_024_2343, w_024_2344, w_024_2345, w_024_2346, w_024_2347, w_024_2348, w_024_2349, w_024_2350, w_024_2351, w_024_2353, w_024_2355, w_024_2356, w_024_2357, w_024_2358, w_024_2359, w_024_2360, w_024_2361, w_024_2362, w_024_2363, w_024_2364, w_024_2366, w_024_2368, w_024_2370, w_024_2371, w_024_2372, w_024_2374, w_024_2377, w_024_2379, w_024_2380, w_024_2381, w_024_2382, w_024_2384, w_024_2385, w_024_2386, w_024_2387, w_024_2389, w_024_2390, w_024_2391, w_024_2392, w_024_2393, w_024_2394, w_024_2395, w_024_2397, w_024_2398, w_024_2399, w_024_2401, w_024_2402, w_024_2403, w_024_2404, w_024_2405, w_024_2407, w_024_2408, w_024_2409, w_024_2410, w_024_2412, w_024_2413, w_024_2414, w_024_2415, w_024_2416, w_024_2418, w_024_2419, w_024_2421, w_024_2422, w_024_2423, w_024_2424, w_024_2426, w_024_2427, w_024_2428, w_024_2429, w_024_2430, w_024_2433, w_024_2434, w_024_2435, w_024_2436, w_024_2437, w_024_2438, w_024_2439, w_024_2441, w_024_2442, w_024_2443, w_024_2445, w_024_2446, w_024_2447, w_024_2448, w_024_2449, w_024_2450, w_024_2451, w_024_2453, w_024_2454, w_024_2455, w_024_2456, w_024_2457, w_024_2458, w_024_2459, w_024_2461, w_024_2462, w_024_2463, w_024_2464, w_024_2465, w_024_2466, w_024_2467, w_024_2469, w_024_2470, w_024_2471, w_024_2473, w_024_2474, w_024_2475, w_024_2476, w_024_2477, w_024_2478, w_024_2479, w_024_2480, w_024_2481, w_024_2482, w_024_2483, w_024_2484, w_024_2485, w_024_2486, w_024_2490, w_024_2491, w_024_2492, w_024_2494, w_024_2495, w_024_2496, w_024_2497, w_024_2498, w_024_2499, w_024_2500, w_024_2501, w_024_2502, w_024_2503, w_024_2504, w_024_2505, w_024_2506, w_024_2507, w_024_2508, w_024_2509, w_024_2510, w_024_2511, w_024_2512, w_024_2514, w_024_2515, w_024_2517, w_024_2518, w_024_2519, w_024_2520, w_024_2523, w_024_2524, w_024_2525, w_024_2526, w_024_2527, w_024_2528, w_024_2529, w_024_2531, w_024_2532, w_024_2533, w_024_2534, w_024_2536, w_024_2538, w_024_2539, w_024_2540, w_024_2541, w_024_2543, w_024_2544, w_024_2545, w_024_2546, w_024_2547, w_024_2548, w_024_2549, w_024_2550, w_024_2551, w_024_2552, w_024_2553, w_024_2554, w_024_2555, w_024_2556, w_024_2557, w_024_2558, w_024_2560, w_024_2561, w_024_2562, w_024_2563, w_024_2565, w_024_2566, w_024_2567, w_024_2568, w_024_2570, w_024_2572, w_024_2573, w_024_2574, w_024_2575, w_024_2577, w_024_2578, w_024_2579, w_024_2580, w_024_2581, w_024_2582, w_024_2583, w_024_2585, w_024_2586, w_024_2587, w_024_2588, w_024_2591, w_024_2592, w_024_2593, w_024_2595, w_024_2596, w_024_2597, w_024_2598, w_024_2599, w_024_2600, w_024_2601, w_024_2602, w_024_2603, w_024_2605, w_024_2606, w_024_2607, w_024_2610, w_024_2611, w_024_2612, w_024_2613, w_024_2614, w_024_2615, w_024_2618, w_024_2619, w_024_2621, w_024_2624, w_024_2625, w_024_2626, w_024_2627, w_024_2628, w_024_2629, w_024_2630, w_024_2631, w_024_2632, w_024_2633, w_024_2634, w_024_2635, w_024_2637, w_024_2638, w_024_2640, w_024_2641, w_024_2642, w_024_2643, w_024_2644, w_024_2645, w_024_2646, w_024_2648, w_024_2649, w_024_2650, w_024_2651, w_024_2652, w_024_2653, w_024_2654, w_024_2655, w_024_2656, w_024_2657, w_024_2658, w_024_2660, w_024_2661, w_024_2662, w_024_2663, w_024_2664, w_024_2665, w_024_2666, w_024_2667, w_024_2669, w_024_2670, w_024_2671, w_024_2672, w_024_2673, w_024_2675, w_024_2676, w_024_2678, w_024_2679, w_024_2680, w_024_2681, w_024_2682, w_024_2683, w_024_2684, w_024_2685, w_024_2686, w_024_2688, w_024_2689, w_024_2690, w_024_2691, w_024_2692, w_024_2693, w_024_2696, w_024_2697, w_024_2698, w_024_2700, w_024_2701, w_024_2703, w_024_2704, w_024_2705, w_024_2706, w_024_2707, w_024_2708, w_024_2710, w_024_2711, w_024_2712, w_024_2713, w_024_2714, w_024_2715, w_024_2716, w_024_2718, w_024_2719, w_024_2721, w_024_2722, w_024_2723, w_024_2724, w_024_2725, w_024_2726, w_024_2727, w_024_2728, w_024_2729, w_024_2730, w_024_2731, w_024_2732, w_024_2733, w_024_2734, w_024_2735, w_024_2736, w_024_2737, w_024_2738, w_024_2739, w_024_2740, w_024_2741, w_024_2742, w_024_2743, w_024_2744, w_024_2745, w_024_2746, w_024_2747, w_024_2748, w_024_2749, w_024_2750, w_024_2752, w_024_2753, w_024_2754, w_024_2755, w_024_2756, w_024_2757, w_024_2758, w_024_2759, w_024_2761, w_024_2762, w_024_2763, w_024_2764, w_024_2765, w_024_2766, w_024_2767, w_024_2768, w_024_2769, w_024_2771, w_024_2773, w_024_2775, w_024_2776, w_024_2777, w_024_2778, w_024_2779, w_024_2780, w_024_2781, w_024_2782, w_024_2783, w_024_2785, w_024_2786, w_024_2787, w_024_2788, w_024_2789, w_024_2790, w_024_2791, w_024_2792, w_024_2793, w_024_2794, w_024_2795, w_024_2796, w_024_2797, w_024_2798, w_024_2799, w_024_2800, w_024_2801, w_024_2803, w_024_2804, w_024_2805, w_024_2806, w_024_2807, w_024_2809, w_024_2810, w_024_2813, w_024_2814, w_024_2817, w_024_2818, w_024_2819, w_024_2820, w_024_2821, w_024_2822, w_024_2823, w_024_2824, w_024_2825, w_024_2827, w_024_2828, w_024_2829, w_024_2830, w_024_2831, w_024_2832, w_024_2833, w_024_2835, w_024_2836, w_024_2837, w_024_2839, w_024_2840, w_024_2841, w_024_2842, w_024_2843, w_024_2845, w_024_2846, w_024_2849, w_024_2850, w_024_2851, w_024_2852, w_024_2853, w_024_2854, w_024_2856, w_024_2857, w_024_2858, w_024_2859, w_024_2860, w_024_2861, w_024_2862, w_024_2863, w_024_2864, w_024_2865, w_024_2866, w_024_2867, w_024_2868, w_024_2869, w_024_2871, w_024_2872, w_024_2873, w_024_2876, w_024_2877, w_024_2878, w_024_2879, w_024_2880, w_024_2881, w_024_2883, w_024_2884, w_024_2885, w_024_2886, w_024_2887, w_024_2888, w_024_2889, w_024_2891, w_024_2892, w_024_2894, w_024_2895, w_024_2896, w_024_2897, w_024_2899, w_024_2900, w_024_2901, w_024_2903, w_024_2904, w_024_2905, w_024_2907, w_024_2908, w_024_2909, w_024_2910, w_024_2911, w_024_2912, w_024_2913, w_024_2914, w_024_2915, w_024_2916, w_024_2917, w_024_2918, w_024_2919, w_024_2920, w_024_2921, w_024_2922, w_024_2923, w_024_2924, w_024_2925, w_024_2926, w_024_2928, w_024_2929, w_024_2930, w_024_2931, w_024_2932, w_024_2934, w_024_2936, w_024_2939, w_024_2940, w_024_2941, w_024_2942, w_024_2943, w_024_2944, w_024_2945, w_024_2946, w_024_2947, w_024_2948, w_024_2949, w_024_2950, w_024_2951, w_024_2952, w_024_2953, w_024_2954, w_024_2955, w_024_2956, w_024_2957, w_024_2958, w_024_2959, w_024_2960, w_024_2961, w_024_2962, w_024_2963, w_024_2965, w_024_2966, w_024_2967, w_024_2969, w_024_2971, w_024_2972, w_024_2973, w_024_2974, w_024_2975, w_024_2976, w_024_2977, w_024_2978, w_024_2979, w_024_2980, w_024_2981, w_024_2982, w_024_2983, w_024_2985, w_024_2986, w_024_2987, w_024_2988, w_024_2989, w_024_2990, w_024_2993, w_024_2994, w_024_2995, w_024_2998, w_024_2999, w_024_3000, w_024_3001, w_024_3002, w_024_3003, w_024_3004, w_024_3005, w_024_3007, w_024_3009, w_024_3010, w_024_3012, w_024_3013, w_024_3014, w_024_3015, w_024_3016, w_024_3017, w_024_3018, w_024_3019, w_024_3020, w_024_3021, w_024_3023, w_024_3024, w_024_3025, w_024_3026, w_024_3027, w_024_3028, w_024_3029, w_024_3030, w_024_3031, w_024_3032, w_024_3033, w_024_3034, w_024_3035, w_024_3036, w_024_3039, w_024_3041, w_024_3042, w_024_3043, w_024_3044, w_024_3045, w_024_3046, w_024_3047, w_024_3048, w_024_3050, w_024_3051, w_024_3052, w_024_3053, w_024_3055, w_024_3056, w_024_3057, w_024_3058, w_024_3059, w_024_3060, w_024_3061, w_024_3062, w_024_3064, w_024_3065, w_024_3067, w_024_3068, w_024_3069, w_024_3070, w_024_3071, w_024_3073, w_024_3074, w_024_3076, w_024_3077, w_024_3079, w_024_3080, w_024_3081, w_024_3082, w_024_3083, w_024_3084, w_024_3085, w_024_3086, w_024_3087, w_024_3088, w_024_3090, w_024_3091, w_024_3092, w_024_3094, w_024_3095, w_024_3096, w_024_3097, w_024_3098, w_024_3099, w_024_3100, w_024_3101, w_024_3102, w_024_3103, w_024_3104, w_024_3106, w_024_3107, w_024_3108, w_024_3111, w_024_3112, w_024_3113, w_024_3114, w_024_3115, w_024_3117, w_024_3118, w_024_3120, w_024_3121, w_024_3122, w_024_3123, w_024_3124, w_024_3125, w_024_3127, w_024_3129, w_024_3130, w_024_3132, w_024_3133, w_024_3134, w_024_3135, w_024_3136, w_024_3137, w_024_3138, w_024_3140, w_024_3141, w_024_3142, w_024_3143, w_024_3145, w_024_3146, w_024_3147, w_024_3148, w_024_3149, w_024_3150, w_024_3151, w_024_3153, w_024_3154, w_024_3155, w_024_3156, w_024_3157, w_024_3160, w_024_3161, w_024_3162, w_024_3163, w_024_3164, w_024_3165, w_024_3168, w_024_3170, w_024_3171, w_024_3173, w_024_3174, w_024_3175, w_024_3178, w_024_3179, w_024_3180, w_024_3181, w_024_3183, w_024_3184, w_024_3185, w_024_3186, w_024_3189, w_024_3190, w_024_3193, w_024_3194, w_024_3195, w_024_3196, w_024_3197, w_024_3198, w_024_3199, w_024_3200, w_024_3201, w_024_3204, w_024_3205, w_024_3207, w_024_3208, w_024_3209, w_024_3210, w_024_3211, w_024_3212, w_024_3213, w_024_3214, w_024_3215, w_024_3217, w_024_3218, w_024_3219, w_024_3220, w_024_3221, w_024_3223, w_024_3225, w_024_3226, w_024_3227, w_024_3228, w_024_3229, w_024_3230, w_024_3231, w_024_3233, w_024_3234, w_024_3235, w_024_3236, w_024_3237, w_024_3238, w_024_3239, w_024_3240, w_024_3244, w_024_3245, w_024_3246, w_024_3247, w_024_3248, w_024_3249, w_024_3250, w_024_3251, w_024_3252, w_024_3255, w_024_3256, w_024_3257, w_024_3258, w_024_3259, w_024_3261, w_024_3262, w_024_3263, w_024_3264, w_024_3265, w_024_3266, w_024_3267, w_024_3268, w_024_3269, w_024_3270, w_024_3271, w_024_3272, w_024_3273, w_024_3274, w_024_3275, w_024_3276, w_024_3277, w_024_3280, w_024_3282, w_024_3283, w_024_3284, w_024_3285, w_024_3286, w_024_3288, w_024_3290, w_024_3291, w_024_3293, w_024_3295, w_024_3296, w_024_3297, w_024_3298, w_024_3299, w_024_3300, w_024_3301, w_024_3302, w_024_3303, w_024_3304, w_024_3305, w_024_3308, w_024_3310, w_024_3311, w_024_3312, w_024_3313, w_024_3314, w_024_3315, w_024_3316, w_024_3317, w_024_3318, w_024_3319, w_024_3320, w_024_3321, w_024_3322, w_024_3323, w_024_3324, w_024_3325, w_024_3326, w_024_3327, w_024_3329, w_024_3330, w_024_3332, w_024_3334, w_024_3336, w_024_3337, w_024_3338, w_024_3339, w_024_3340, w_024_3341, w_024_3342, w_024_3343, w_024_3344, w_024_3345, w_024_3346, w_024_3347, w_024_3349, w_024_3350, w_024_3352, w_024_3354, w_024_3355, w_024_3356, w_024_3357, w_024_3358, w_024_3359, w_024_3360, w_024_3361, w_024_3362, w_024_3363, w_024_3366, w_024_3367, w_024_3368, w_024_3369, w_024_3370, w_024_3371, w_024_3372, w_024_3373, w_024_3374, w_024_3376, w_024_3378, w_024_3379, w_024_3380, w_024_3382, w_024_3385, w_024_3386, w_024_3389, w_024_3390, w_024_3392, w_024_3393, w_024_3394, w_024_3395, w_024_3396, w_024_3398, w_024_3399, w_024_3400, w_024_3401, w_024_3403, w_024_3404, w_024_3405, w_024_3406, w_024_3407, w_024_3408, w_024_3409, w_024_3410, w_024_3411, w_024_3412, w_024_3413, w_024_3414, w_024_3415, w_024_3416, w_024_3417, w_024_3418, w_024_3419, w_024_3420, w_024_3421, w_024_3422, w_024_3423, w_024_3424, w_024_3425, w_024_3426, w_024_3428, w_024_3429, w_024_3430, w_024_3431, w_024_3433, w_024_3434, w_024_3435, w_024_3436, w_024_3437, w_024_3438, w_024_3440, w_024_3441, w_024_3442, w_024_3443, w_024_3444, w_024_3445, w_024_3447, w_024_3448, w_024_3449, w_024_3451, w_024_3452, w_024_3455, w_024_3456, w_024_3457, w_024_3458, w_024_3460, w_024_3461, w_024_3463, w_024_3464, w_024_3465, w_024_3466, w_024_3467, w_024_3468, w_024_3469, w_024_3470, w_024_3471, w_024_3472, w_024_3473, w_024_3474, w_024_3475, w_024_3476, w_024_3477, w_024_3478, w_024_3479, w_024_3480, w_024_3481, w_024_3482, w_024_3483, w_024_3484, w_024_3485, w_024_3486, w_024_3488, w_024_3490, w_024_3493, w_024_3494, w_024_3495, w_024_3497, w_024_3498, w_024_3499, w_024_3500, w_024_3501, w_024_3502, w_024_3503, w_024_3504, w_024_3505, w_024_3506, w_024_3507, w_024_3508, w_024_3510, w_024_3513, w_024_3514, w_024_3516, w_024_3517, w_024_3518, w_024_3519, w_024_3520, w_024_3521, w_024_3522, w_024_3523, w_024_3526, w_024_3528, w_024_3529, w_024_3530, w_024_3531, w_024_3532, w_024_3533, w_024_3534, w_024_3535, w_024_3536, w_024_3537, w_024_3538, w_024_3539, w_024_3540, w_024_3541, w_024_3542, w_024_3543, w_024_3544, w_024_3545, w_024_3546, w_024_3547, w_024_3548, w_024_3549, w_024_3550, w_024_3551, w_024_3552, w_024_3553, w_024_3555, w_024_3556, w_024_3557, w_024_3558, w_024_3559, w_024_3560, w_024_3562, w_024_3563, w_024_3565, w_024_3566, w_024_3567, w_024_3568, w_024_3570, w_024_3572, w_024_3573, w_024_3575, w_024_3576, w_024_3577, w_024_3578, w_024_3579, w_024_3580, w_024_3581, w_024_3582, w_024_3584, w_024_3586, w_024_3587, w_024_3588, w_024_3589, w_024_3591, w_024_3592, w_024_3593, w_024_3595, w_024_3597, w_024_3598, w_024_3599, w_024_3600, w_024_3601, w_024_3602, w_024_3603, w_024_3604, w_024_3606, w_024_3608, w_024_3609, w_024_3610, w_024_3611, w_024_3612, w_024_3614, w_024_3615, w_024_3617, w_024_3618, w_024_3619, w_024_3620, w_024_3621, w_024_3622, w_024_3623, w_024_3624, w_024_3625, w_024_3626, w_024_3627, w_024_3628, w_024_3629, w_024_3631, w_024_3633, w_024_3634, w_024_3635, w_024_3636, w_024_3637, w_024_3639, w_024_3640, w_024_3641, w_024_3643, w_024_3644, w_024_3646, w_024_3647, w_024_3650, w_024_3651, w_024_3652, w_024_3653, w_024_3655, w_024_3656, w_024_3657, w_024_3659, w_024_3660, w_024_3661, w_024_3662, w_024_3664, w_024_3665, w_024_3666, w_024_3668, w_024_3669, w_024_3670, w_024_3671, w_024_3672, w_024_3674, w_024_3675, w_024_3677, w_024_3678, w_024_3679, w_024_3680, w_024_3681, w_024_3682, w_024_3683, w_024_3684, w_024_3685, w_024_3686, w_024_3687, w_024_3688, w_024_3689, w_024_3690, w_024_3693, w_024_3695, w_024_3697, w_024_3698, w_024_3699, w_024_3700, w_024_3701, w_024_3702, w_024_3703, w_024_3704, w_024_3705, w_024_3706, w_024_3707, w_024_3708, w_024_3710, w_024_3711, w_024_3712, w_024_3713, w_024_3714, w_024_3715, w_024_3716, w_024_3717, w_024_3718, w_024_3720, w_024_3722, w_024_3723, w_024_3724, w_024_3725, w_024_3726, w_024_3727, w_024_3728, w_024_3729, w_024_3730, w_024_3732, w_024_3734, w_024_3735, w_024_3736, w_024_3737, w_024_3738, w_024_3739, w_024_3743, w_024_3744, w_024_3746, w_024_3747, w_024_3749, w_024_3750, w_024_3751, w_024_3752, w_024_3753, w_024_3754, w_024_3755, w_024_3757, w_024_3759, w_024_3760, w_024_3762, w_024_3763, w_024_3764, w_024_3765, w_024_3766, w_024_3767, w_024_3769, w_024_3770, w_024_3771, w_024_3772, w_024_3774, w_024_3777, w_024_3780, w_024_3782, w_024_3783, w_024_3784, w_024_3785, w_024_3786, w_024_3787, w_024_3788, w_024_3791, w_024_3792, w_024_3793, w_024_3794, w_024_3795, w_024_3796, w_024_3797, w_024_3799, w_024_3800, w_024_3801, w_024_3802, w_024_3803, w_024_3804, w_024_3805, w_024_3806, w_024_3807, w_024_3808, w_024_3809, w_024_3810, w_024_3811, w_024_3813, w_024_3815, w_024_3816, w_024_3817, w_024_3819, w_024_3820, w_024_3821, w_024_3822, w_024_3823, w_024_3825, w_024_3826, w_024_3827, w_024_3828, w_024_3829, w_024_3830, w_024_3831, w_024_3833, w_024_3834, w_024_3835, w_024_3836, w_024_3837, w_024_3838, w_024_3840, w_024_3842, w_024_3843, w_024_3844, w_024_3845, w_024_3846, w_024_3848, w_024_3849, w_024_3850, w_024_3851, w_024_3853, w_024_3854, w_024_3855, w_024_3856, w_024_3857, w_024_3858, w_024_3860, w_024_3861, w_024_3862, w_024_3863, w_024_3864, w_024_3865, w_024_3866, w_024_3868, w_024_3869, w_024_3870, w_024_3871, w_024_3872, w_024_3874, w_024_3876, w_024_3877, w_024_3878, w_024_3879, w_024_3880, w_024_3881, w_024_3883, w_024_3884, w_024_3886, w_024_3887, w_024_3888, w_024_3889, w_024_3890, w_024_3891, w_024_3892, w_024_3893, w_024_3894, w_024_3895, w_024_3896, w_024_3897, w_024_3898, w_024_3899, w_024_3900, w_024_3902, w_024_3903, w_024_3904, w_024_3905, w_024_3906, w_024_3907, w_024_3908, w_024_3909, w_024_3910, w_024_3912, w_024_3913, w_024_3914, w_024_3915, w_024_3919, w_024_3920, w_024_3921, w_024_3922, w_024_3923, w_024_3924, w_024_3926, w_024_3927, w_024_3928, w_024_3929, w_024_3930, w_024_3931, w_024_3933, w_024_3934, w_024_3935, w_024_3936, w_024_3937, w_024_3938, w_024_3939, w_024_3941, w_024_3942, w_024_3943, w_024_3944, w_024_3945, w_024_3946, w_024_3947, w_024_3949, w_024_3950, w_024_3951, w_024_3952, w_024_3953, w_024_3955, w_024_3957, w_024_3958, w_024_3959, w_024_3960, w_024_3961, w_024_3962, w_024_3963, w_024_3964, w_024_3965, w_024_3966, w_024_3968, w_024_3969, w_024_3970, w_024_3972, w_024_3973, w_024_3974, w_024_3975, w_024_3976, w_024_3977, w_024_3978, w_024_3980, w_024_3982, w_024_3983, w_024_3984, w_024_3985, w_024_3986, w_024_3987, w_024_3988, w_024_3989, w_024_3990, w_024_3992, w_024_3993, w_024_3994, w_024_3995, w_024_3996, w_024_3997, w_024_3999, w_024_4000, w_024_4001, w_024_4002, w_024_4003, w_024_4004, w_024_4005, w_024_4006, w_024_4008, w_024_4009, w_024_4010, w_024_4011, w_024_4012, w_024_4013, w_024_4014, w_024_4015, w_024_4016, w_024_4017, w_024_4018, w_024_4019, w_024_4020, w_024_4022, w_024_4024, w_024_4025, w_024_4026, w_024_4027, w_024_4028, w_024_4030, w_024_4032, w_024_4033, w_024_4034, w_024_4035, w_024_4039, w_024_4040, w_024_4041, w_024_4042, w_024_4043, w_024_4044, w_024_4045, w_024_4047, w_024_4049, w_024_4050, w_024_4051, w_024_4052, w_024_4053, w_024_4056, w_024_4058, w_024_4059, w_024_4060, w_024_4061, w_024_4062, w_024_4064, w_024_4065, w_024_4066, w_024_4067, w_024_4068, w_024_4069, w_024_4070, w_024_4071, w_024_4072, w_024_4073, w_024_4074, w_024_4076, w_024_4077, w_024_4081, w_024_4082, w_024_4083, w_024_4084, w_024_4085, w_024_4086, w_024_4088, w_024_4090, w_024_4091, w_024_4092, w_024_4095, w_024_4096, w_024_4097, w_024_4098, w_024_4099, w_024_4100, w_024_4101, w_024_4103, w_024_4104, w_024_4107, w_024_4108, w_024_4109, w_024_4110, w_024_4112, w_024_4114, w_024_4115, w_024_4116, w_024_4117, w_024_4118, w_024_4119, w_024_4120, w_024_4121, w_024_4122, w_024_4123, w_024_4124, w_024_4125, w_024_4128, w_024_4130, w_024_4131, w_024_4132, w_024_4133, w_024_4134, w_024_4135, w_024_4136, w_024_4137, w_024_4138, w_024_4139, w_024_4140, w_024_4141, w_024_4142, w_024_4143, w_024_4146, w_024_4147, w_024_4148, w_024_4149, w_024_4150, w_024_4151, w_024_4152, w_024_4153, w_024_4154, w_024_4155, w_024_4156, w_024_4157, w_024_4158, w_024_4159, w_024_4161, w_024_4162, w_024_4163, w_024_4164, w_024_4165, w_024_4167, w_024_4168, w_024_4169, w_024_4170, w_024_4171, w_024_4172, w_024_4174, w_024_4175, w_024_4177, w_024_4179, w_024_4180, w_024_4181, w_024_4182, w_024_4183, w_024_4184, w_024_4185, w_024_4186, w_024_4187, w_024_4188, w_024_4189, w_024_4190, w_024_4191, w_024_4192, w_024_4193, w_024_4194, w_024_4195, w_024_4196, w_024_4197, w_024_4198, w_024_4199, w_024_4200, w_024_4201, w_024_4202, w_024_4204, w_024_4205, w_024_4206, w_024_4207, w_024_4208, w_024_4209, w_024_4210, w_024_4211, w_024_4212, w_024_4214, w_024_4215, w_024_4216, w_024_4217, w_024_4220, w_024_4221, w_024_4222, w_024_4224, w_024_4226, w_024_4227, w_024_4228, w_024_4229, w_024_4230, w_024_4231, w_024_4233, w_024_4234, w_024_4235, w_024_4236, w_024_4237, w_024_4238, w_024_4239, w_024_4240, w_024_4241, w_024_4242, w_024_4243, w_024_4244, w_024_4245, w_024_4246, w_024_4247, w_024_4248, w_024_4249, w_024_4250, w_024_4251, w_024_4252, w_024_4253, w_024_4256, w_024_4257, w_024_4258, w_024_4260, w_024_4261, w_024_4263, w_024_4264, w_024_4265, w_024_4266, w_024_4267, w_024_4268, w_024_4269, w_024_4270, w_024_4271, w_024_4272, w_024_4273, w_024_4275, w_024_4277, w_024_4278, w_024_4280, w_024_4281, w_024_4282, w_024_4284, w_024_4285, w_024_4286, w_024_4287, w_024_4288, w_024_4289, w_024_4292, w_024_4293, w_024_4294, w_024_4295, w_024_4296, w_024_4301, w_024_4302, w_024_4303, w_024_4304, w_024_4309, w_024_4310, w_024_4311, w_024_4312, w_024_4313, w_024_4314, w_024_4315, w_024_4317, w_024_4318, w_024_4319, w_024_4321, w_024_4322, w_024_4323, w_024_4325, w_024_4326, w_024_4327, w_024_4328, w_024_4329, w_024_4331, w_024_4332, w_024_4333, w_024_4334, w_024_4337, w_024_4339, w_024_4341, w_024_4342, w_024_4343, w_024_4344, w_024_4345, w_024_4346, w_024_4347, w_024_4348, w_024_4350, w_024_4351, w_024_4353, w_024_4354, w_024_4355, w_024_4356, w_024_4357, w_024_4358, w_024_4359;
  wire w_025_000, w_025_001, w_025_002, w_025_003, w_025_004, w_025_005, w_025_006, w_025_007, w_025_008, w_025_009, w_025_010, w_025_011, w_025_012, w_025_013, w_025_014, w_025_015, w_025_016, w_025_017, w_025_018, w_025_019, w_025_020, w_025_021, w_025_022, w_025_023, w_025_024, w_025_025, w_025_026, w_025_027, w_025_028, w_025_029, w_025_030, w_025_031, w_025_032, w_025_033, w_025_034, w_025_035, w_025_036, w_025_037, w_025_038, w_025_039, w_025_040, w_025_041, w_025_042, w_025_043, w_025_044, w_025_045, w_025_046, w_025_047, w_025_048, w_025_049, w_025_050, w_025_051, w_025_052, w_025_053, w_025_054, w_025_055, w_025_056, w_025_057, w_025_058, w_025_059, w_025_060, w_025_061, w_025_062, w_025_063, w_025_064, w_025_065, w_025_066, w_025_067, w_025_068, w_025_069, w_025_070, w_025_071, w_025_072, w_025_073, w_025_074, w_025_075, w_025_076, w_025_077, w_025_078, w_025_079, w_025_080, w_025_081, w_025_082, w_025_083, w_025_084, w_025_085, w_025_086, w_025_087, w_025_088, w_025_089, w_025_090, w_025_091, w_025_092, w_025_093, w_025_094, w_025_095, w_025_096, w_025_097, w_025_098, w_025_099, w_025_100, w_025_101, w_025_102, w_025_103, w_025_104, w_025_105, w_025_106, w_025_107, w_025_108, w_025_109, w_025_110, w_025_111, w_025_112, w_025_113, w_025_114, w_025_115, w_025_116, w_025_117, w_025_118, w_025_119, w_025_120, w_025_121, w_025_122, w_025_123, w_025_124, w_025_125, w_025_126, w_025_127, w_025_128, w_025_129, w_025_130, w_025_131, w_025_132, w_025_133, w_025_134, w_025_135, w_025_136, w_025_137, w_025_138, w_025_139, w_025_140, w_025_141, w_025_142, w_025_143, w_025_144, w_025_145, w_025_146, w_025_147, w_025_148, w_025_149, w_025_150, w_025_151, w_025_152, w_025_153, w_025_154, w_025_155, w_025_156, w_025_157, w_025_158, w_025_159, w_025_160, w_025_161, w_025_162, w_025_163, w_025_164, w_025_165, w_025_166, w_025_167, w_025_168, w_025_169, w_025_170, w_025_171, w_025_172, w_025_173, w_025_174, w_025_175, w_025_176, w_025_177, w_025_178, w_025_179, w_025_180, w_025_181, w_025_182, w_025_183, w_025_184, w_025_185, w_025_186, w_025_187, w_025_188, w_025_189, w_025_190, w_025_191, w_025_192, w_025_193, w_025_194, w_025_195, w_025_196, w_025_197, w_025_198, w_025_199, w_025_200, w_025_201, w_025_202, w_025_203, w_025_204, w_025_205, w_025_206, w_025_207, w_025_208, w_025_209, w_025_210, w_025_211, w_025_212, w_025_213, w_025_214, w_025_215, w_025_216, w_025_217, w_025_218, w_025_219, w_025_220, w_025_221, w_025_222, w_025_223, w_025_224, w_025_225, w_025_226, w_025_227, w_025_228, w_025_229, w_025_230, w_025_231, w_025_232, w_025_233, w_025_234, w_025_235, w_025_236, w_025_237, w_025_238, w_025_239, w_025_240, w_025_241, w_025_242, w_025_243, w_025_244, w_025_245, w_025_246, w_025_247, w_025_248, w_025_249, w_025_250, w_025_251, w_025_252, w_025_253, w_025_254, w_025_255, w_025_256, w_025_257, w_025_258, w_025_259, w_025_260, w_025_261, w_025_262, w_025_263, w_025_264, w_025_265, w_025_266, w_025_267, w_025_268, w_025_269, w_025_270, w_025_271, w_025_272, w_025_273, w_025_274, w_025_275, w_025_276, w_025_277, w_025_278, w_025_279, w_025_280, w_025_281, w_025_282, w_025_283, w_025_284, w_025_285, w_025_286, w_025_287, w_025_288, w_025_289, w_025_290, w_025_291, w_025_292, w_025_293, w_025_294, w_025_295, w_025_296, w_025_297, w_025_298, w_025_299, w_025_300, w_025_301, w_025_302, w_025_303, w_025_304, w_025_305, w_025_306, w_025_307, w_025_308, w_025_309, w_025_310, w_025_311, w_025_312, w_025_313, w_025_314, w_025_315, w_025_316, w_025_317, w_025_318, w_025_319, w_025_320, w_025_321, w_025_322, w_025_323, w_025_324, w_025_325, w_025_326, w_025_327, w_025_328, w_025_329, w_025_330, w_025_331, w_025_332, w_025_333, w_025_334, w_025_335, w_025_336, w_025_337, w_025_338, w_025_339, w_025_340, w_025_341, w_025_342, w_025_343, w_025_344, w_025_345, w_025_346, w_025_347, w_025_348, w_025_349, w_025_350, w_025_351, w_025_352, w_025_353, w_025_354, w_025_355, w_025_356, w_025_357, w_025_358, w_025_359, w_025_360, w_025_361, w_025_362, w_025_363, w_025_364, w_025_365, w_025_366, w_025_367, w_025_368, w_025_369, w_025_370, w_025_371, w_025_372, w_025_373, w_025_374, w_025_375, w_025_376, w_025_377, w_025_378, w_025_379, w_025_380, w_025_381, w_025_382, w_025_383, w_025_384, w_025_385, w_025_386, w_025_387, w_025_388, w_025_389, w_025_390, w_025_391, w_025_392, w_025_393, w_025_394, w_025_395, w_025_396, w_025_397, w_025_398, w_025_399, w_025_400, w_025_401, w_025_402, w_025_403, w_025_404, w_025_405, w_025_406, w_025_407, w_025_408, w_025_409, w_025_410, w_025_411, w_025_412, w_025_413, w_025_414, w_025_415, w_025_416, w_025_417, w_025_418, w_025_419, w_025_420, w_025_421, w_025_422, w_025_423, w_025_424, w_025_425, w_025_426, w_025_427, w_025_428, w_025_429, w_025_430, w_025_431, w_025_432, w_025_433, w_025_434, w_025_435, w_025_436, w_025_437, w_025_438, w_025_440, w_025_441, w_025_442, w_025_443, w_025_444, w_025_445, w_025_446, w_025_447, w_025_448, w_025_449, w_025_450, w_025_451, w_025_452, w_025_453, w_025_454, w_025_455, w_025_456, w_025_457, w_025_458, w_025_459, w_025_460, w_025_462, w_025_463, w_025_464, w_025_465, w_025_466, w_025_467, w_025_468, w_025_469, w_025_470, w_025_471, w_025_472, w_025_473, w_025_474, w_025_475, w_025_476, w_025_477, w_025_478, w_025_479, w_025_480, w_025_481, w_025_482, w_025_483, w_025_484, w_025_485, w_025_486, w_025_487, w_025_488, w_025_489, w_025_490, w_025_491, w_025_492, w_025_493, w_025_494, w_025_495, w_025_496, w_025_497, w_025_498, w_025_499, w_025_500, w_025_501, w_025_502, w_025_503, w_025_504, w_025_505, w_025_506, w_025_507, w_025_508, w_025_509, w_025_510, w_025_511, w_025_512, w_025_513, w_025_514, w_025_515, w_025_516, w_025_517, w_025_518, w_025_519, w_025_520, w_025_521, w_025_522, w_025_523, w_025_524, w_025_525, w_025_526, w_025_527, w_025_528, w_025_529, w_025_530, w_025_531, w_025_532, w_025_533, w_025_534, w_025_535, w_025_536, w_025_537, w_025_538, w_025_539, w_025_540, w_025_541, w_025_542, w_025_543, w_025_544, w_025_545, w_025_546, w_025_547, w_025_548, w_025_549, w_025_550, w_025_551, w_025_552, w_025_553, w_025_554, w_025_555, w_025_556, w_025_557, w_025_558, w_025_559, w_025_560, w_025_561, w_025_562, w_025_563, w_025_564, w_025_565, w_025_566, w_025_567, w_025_568, w_025_569, w_025_570, w_025_571, w_025_572, w_025_573, w_025_574, w_025_575, w_025_576, w_025_577, w_025_578, w_025_579, w_025_580, w_025_581, w_025_582, w_025_583, w_025_584, w_025_585, w_025_586, w_025_587, w_025_588, w_025_589, w_025_590, w_025_591, w_025_592, w_025_593, w_025_594, w_025_595, w_025_596, w_025_597, w_025_598, w_025_599, w_025_600, w_025_601, w_025_602, w_025_603, w_025_604, w_025_605, w_025_606, w_025_607, w_025_608, w_025_609, w_025_610, w_025_611, w_025_612, w_025_613, w_025_614, w_025_615, w_025_616, w_025_617, w_025_618, w_025_619, w_025_620, w_025_621, w_025_622, w_025_623, w_025_624, w_025_625, w_025_626, w_025_627, w_025_628, w_025_629, w_025_630, w_025_631, w_025_632, w_025_633, w_025_634, w_025_635, w_025_636, w_025_637, w_025_638, w_025_639, w_025_640, w_025_641, w_025_642, w_025_643, w_025_644, w_025_645, w_025_646, w_025_647, w_025_648, w_025_649, w_025_650, w_025_651, w_025_652, w_025_653, w_025_654, w_025_655, w_025_656, w_025_657, w_025_658, w_025_659, w_025_660, w_025_661, w_025_662, w_025_663, w_025_664, w_025_665, w_025_666, w_025_667, w_025_668, w_025_669, w_025_670, w_025_671, w_025_672, w_025_673, w_025_674, w_025_675, w_025_676, w_025_677, w_025_678, w_025_679, w_025_680, w_025_681, w_025_682, w_025_683, w_025_684, w_025_685, w_025_686, w_025_687, w_025_688, w_025_689, w_025_690, w_025_691, w_025_692, w_025_693, w_025_694, w_025_695, w_025_696, w_025_697, w_025_698, w_025_699, w_025_700, w_025_701, w_025_702, w_025_703, w_025_704, w_025_705, w_025_706, w_025_707, w_025_708, w_025_709, w_025_710, w_025_711, w_025_712, w_025_713, w_025_714, w_025_715, w_025_716, w_025_717, w_025_718, w_025_719, w_025_720, w_025_721, w_025_722, w_025_723, w_025_724, w_025_725, w_025_726, w_025_727, w_025_728, w_025_729, w_025_730, w_025_731, w_025_732, w_025_733, w_025_734, w_025_735, w_025_736, w_025_737, w_025_738, w_025_739, w_025_740, w_025_741, w_025_742, w_025_743, w_025_744, w_025_745, w_025_746, w_025_747, w_025_748, w_025_749, w_025_750, w_025_751, w_025_752, w_025_753, w_025_754, w_025_755, w_025_756, w_025_757, w_025_758, w_025_759, w_025_760, w_025_761, w_025_762, w_025_763, w_025_764, w_025_765, w_025_766, w_025_767, w_025_768, w_025_769, w_025_770, w_025_771, w_025_772, w_025_773, w_025_774, w_025_775, w_025_776, w_025_777, w_025_778, w_025_779, w_025_780, w_025_781, w_025_782, w_025_783, w_025_784, w_025_785, w_025_786, w_025_787, w_025_788, w_025_789, w_025_790, w_025_791, w_025_792, w_025_793, w_025_794, w_025_795, w_025_796, w_025_797, w_025_798, w_025_799, w_025_800, w_025_801, w_025_802, w_025_803, w_025_804, w_025_805, w_025_806, w_025_807, w_025_808, w_025_809, w_025_810, w_025_811, w_025_812, w_025_813, w_025_814, w_025_815, w_025_816, w_025_817, w_025_818, w_025_819, w_025_820, w_025_821, w_025_822, w_025_823, w_025_824, w_025_825, w_025_826, w_025_827, w_025_828, w_025_829, w_025_830, w_025_831, w_025_832, w_025_833, w_025_834, w_025_835, w_025_836, w_025_837, w_025_838, w_025_839, w_025_840, w_025_841, w_025_842, w_025_843, w_025_844, w_025_845, w_025_846, w_025_847, w_025_848, w_025_849, w_025_850, w_025_851, w_025_852, w_025_853, w_025_854, w_025_855, w_025_856, w_025_857, w_025_858, w_025_859, w_025_860, w_025_861, w_025_862, w_025_863, w_025_864, w_025_865, w_025_866, w_025_867, w_025_868, w_025_869, w_025_870, w_025_871, w_025_872, w_025_873, w_025_874, w_025_875, w_025_876, w_025_877, w_025_878, w_025_879, w_025_880, w_025_881, w_025_883, w_025_884, w_025_885, w_025_886, w_025_887, w_025_888, w_025_889, w_025_890, w_025_891, w_025_892, w_025_893, w_025_894, w_025_895, w_025_896, w_025_897, w_025_898, w_025_899, w_025_900, w_025_901, w_025_902, w_025_903, w_025_904, w_025_905, w_025_906, w_025_907, w_025_908, w_025_909, w_025_910, w_025_911, w_025_912, w_025_913, w_025_914, w_025_915, w_025_916, w_025_917, w_025_918, w_025_919, w_025_920, w_025_921, w_025_922, w_025_923, w_025_924, w_025_925, w_025_926, w_025_927, w_025_928, w_025_929, w_025_930, w_025_931, w_025_932, w_025_933, w_025_934, w_025_935, w_025_936, w_025_937, w_025_938, w_025_939, w_025_940, w_025_941, w_025_942, w_025_943, w_025_944, w_025_945, w_025_946, w_025_947, w_025_948, w_025_949, w_025_950, w_025_951, w_025_952, w_025_953, w_025_954, w_025_955, w_025_956, w_025_957, w_025_958, w_025_959, w_025_960, w_025_961, w_025_962, w_025_963, w_025_964, w_025_965, w_025_966, w_025_967, w_025_968, w_025_969, w_025_970, w_025_971, w_025_972, w_025_973, w_025_974, w_025_975, w_025_976, w_025_977, w_025_978, w_025_979, w_025_980, w_025_981, w_025_982, w_025_983, w_025_984, w_025_985, w_025_986, w_025_987, w_025_988, w_025_989, w_025_990, w_025_991, w_025_992, w_025_993, w_025_994, w_025_995, w_025_996, w_025_997, w_025_998, w_025_999, w_025_1000, w_025_1001, w_025_1002, w_025_1003, w_025_1004, w_025_1005, w_025_1006, w_025_1007, w_025_1008, w_025_1009, w_025_1010, w_025_1011, w_025_1012, w_025_1013, w_025_1014, w_025_1015, w_025_1016, w_025_1017, w_025_1018, w_025_1019, w_025_1020, w_025_1021, w_025_1022, w_025_1023, w_025_1024, w_025_1025, w_025_1026, w_025_1027, w_025_1028, w_025_1029, w_025_1030, w_025_1031, w_025_1032, w_025_1033, w_025_1034, w_025_1035, w_025_1036, w_025_1037, w_025_1038, w_025_1039, w_025_1040, w_025_1041, w_025_1042, w_025_1043, w_025_1044, w_025_1045, w_025_1046, w_025_1047, w_025_1048, w_025_1049, w_025_1050, w_025_1051, w_025_1052, w_025_1053, w_025_1054, w_025_1055, w_025_1056, w_025_1057, w_025_1058, w_025_1059, w_025_1060, w_025_1061, w_025_1062, w_025_1063, w_025_1064, w_025_1065, w_025_1066, w_025_1067, w_025_1068, w_025_1069, w_025_1070, w_025_1071, w_025_1072, w_025_1073, w_025_1074, w_025_1075, w_025_1076, w_025_1077, w_025_1078, w_025_1079, w_025_1080, w_025_1081, w_025_1082, w_025_1083, w_025_1084, w_025_1085, w_025_1086, w_025_1087, w_025_1088, w_025_1089, w_025_1090, w_025_1091, w_025_1092, w_025_1093, w_025_1094, w_025_1095, w_025_1096, w_025_1097, w_025_1098, w_025_1099, w_025_1100, w_025_1101, w_025_1102, w_025_1103, w_025_1104, w_025_1105, w_025_1106, w_025_1107, w_025_1108, w_025_1109, w_025_1110, w_025_1111, w_025_1112, w_025_1113, w_025_1114, w_025_1115, w_025_1116, w_025_1117, w_025_1118, w_025_1119, w_025_1120, w_025_1121, w_025_1122, w_025_1123, w_025_1124, w_025_1125, w_025_1126, w_025_1127, w_025_1128, w_025_1129, w_025_1130, w_025_1131, w_025_1132, w_025_1133, w_025_1134, w_025_1135, w_025_1136, w_025_1137, w_025_1138, w_025_1139, w_025_1140, w_025_1141, w_025_1142, w_025_1143, w_025_1144, w_025_1145, w_025_1146, w_025_1147, w_025_1148, w_025_1149, w_025_1150, w_025_1151, w_025_1152, w_025_1153, w_025_1154, w_025_1155, w_025_1156, w_025_1157, w_025_1158, w_025_1159, w_025_1160, w_025_1161, w_025_1162, w_025_1163, w_025_1164, w_025_1165, w_025_1166, w_025_1167, w_025_1168, w_025_1169, w_025_1170, w_025_1171, w_025_1172, w_025_1173, w_025_1174, w_025_1175, w_025_1176, w_025_1177, w_025_1178, w_025_1179, w_025_1180, w_025_1181, w_025_1182, w_025_1183, w_025_1184, w_025_1185, w_025_1186, w_025_1187, w_025_1188, w_025_1189, w_025_1190, w_025_1191, w_025_1192, w_025_1193, w_025_1194, w_025_1195, w_025_1196, w_025_1197, w_025_1198, w_025_1199, w_025_1200, w_025_1201, w_025_1202, w_025_1203, w_025_1204, w_025_1205, w_025_1206, w_025_1207, w_025_1208, w_025_1209, w_025_1210, w_025_1211, w_025_1212, w_025_1213, w_025_1214, w_025_1215, w_025_1216, w_025_1217, w_025_1218, w_025_1219, w_025_1220, w_025_1221, w_025_1222, w_025_1223, w_025_1224, w_025_1225, w_025_1226, w_025_1227, w_025_1228, w_025_1229, w_025_1230, w_025_1231, w_025_1232, w_025_1233, w_025_1234, w_025_1235, w_025_1236, w_025_1237, w_025_1238, w_025_1239, w_025_1240, w_025_1241, w_025_1242, w_025_1243, w_025_1244, w_025_1245, w_025_1246, w_025_1247, w_025_1248, w_025_1249, w_025_1250, w_025_1251, w_025_1252, w_025_1253, w_025_1254, w_025_1255, w_025_1256, w_025_1257, w_025_1258, w_025_1259, w_025_1260, w_025_1261, w_025_1262, w_025_1263, w_025_1264, w_025_1265, w_025_1266, w_025_1267, w_025_1268, w_025_1269, w_025_1270, w_025_1271, w_025_1272, w_025_1273, w_025_1274, w_025_1275, w_025_1276, w_025_1277, w_025_1278, w_025_1279, w_025_1280, w_025_1281, w_025_1282, w_025_1283, w_025_1284, w_025_1285, w_025_1286, w_025_1287, w_025_1288, w_025_1289, w_025_1290, w_025_1291, w_025_1292, w_025_1293, w_025_1294, w_025_1295, w_025_1296, w_025_1297;
  wire w_026_000, w_026_001, w_026_002, w_026_003, w_026_004, w_026_005, w_026_006, w_026_007, w_026_008, w_026_009, w_026_010, w_026_011, w_026_012, w_026_013, w_026_014, w_026_015, w_026_016, w_026_017, w_026_018, w_026_020, w_026_022, w_026_024, w_026_025, w_026_026, w_026_027, w_026_028, w_026_029, w_026_031, w_026_032, w_026_033, w_026_034, w_026_035, w_026_036, w_026_037, w_026_038, w_026_039, w_026_040, w_026_041, w_026_042, w_026_043, w_026_044, w_026_045, w_026_046, w_026_047, w_026_048, w_026_049, w_026_050, w_026_051, w_026_052, w_026_053, w_026_054, w_026_055, w_026_057, w_026_058, w_026_059, w_026_061, w_026_062, w_026_064, w_026_065, w_026_066, w_026_067, w_026_068, w_026_069, w_026_070, w_026_071, w_026_072, w_026_073, w_026_074, w_026_075, w_026_076, w_026_077, w_026_078, w_026_079, w_026_080, w_026_081, w_026_082, w_026_083, w_026_084, w_026_085, w_026_086, w_026_087, w_026_088, w_026_089, w_026_090, w_026_091, w_026_092, w_026_093, w_026_094, w_026_095, w_026_096, w_026_097, w_026_098, w_026_099, w_026_100, w_026_101, w_026_102, w_026_104, w_026_105, w_026_106, w_026_107, w_026_108, w_026_109, w_026_110, w_026_111, w_026_112, w_026_113, w_026_114, w_026_115, w_026_116, w_026_117, w_026_118, w_026_119, w_026_120, w_026_121, w_026_122, w_026_123, w_026_124, w_026_125, w_026_126, w_026_127, w_026_128, w_026_129, w_026_130, w_026_131, w_026_132, w_026_133, w_026_134, w_026_135, w_026_136, w_026_137, w_026_138, w_026_139, w_026_140, w_026_142, w_026_143, w_026_144, w_026_145, w_026_146, w_026_147, w_026_148, w_026_149, w_026_150, w_026_151, w_026_152, w_026_153, w_026_154, w_026_155, w_026_156, w_026_157, w_026_158, w_026_159, w_026_160, w_026_161, w_026_162, w_026_163, w_026_164, w_026_165, w_026_166, w_026_167, w_026_168, w_026_169, w_026_170, w_026_171, w_026_172, w_026_173, w_026_174, w_026_175, w_026_176, w_026_178, w_026_179, w_026_180, w_026_181, w_026_182, w_026_183, w_026_184, w_026_185, w_026_186, w_026_187, w_026_188, w_026_189, w_026_190, w_026_191, w_026_192, w_026_193, w_026_194, w_026_195, w_026_196, w_026_197, w_026_198, w_026_199, w_026_200, w_026_201, w_026_202, w_026_203, w_026_205, w_026_206, w_026_207, w_026_208, w_026_209, w_026_210, w_026_211, w_026_212, w_026_213, w_026_214, w_026_215, w_026_216, w_026_217, w_026_218, w_026_219, w_026_220, w_026_222, w_026_223, w_026_224, w_026_225, w_026_226, w_026_227, w_026_228, w_026_229, w_026_230, w_026_231, w_026_232, w_026_233, w_026_234, w_026_235, w_026_236, w_026_237, w_026_238, w_026_239, w_026_240, w_026_241, w_026_242, w_026_243, w_026_244, w_026_245, w_026_246, w_026_247, w_026_248, w_026_249, w_026_250, w_026_251, w_026_252, w_026_253, w_026_254, w_026_255, w_026_256, w_026_257, w_026_258, w_026_259, w_026_260, w_026_261, w_026_262, w_026_263, w_026_264, w_026_265, w_026_267, w_026_268, w_026_269, w_026_270, w_026_271, w_026_272, w_026_273, w_026_274, w_026_275, w_026_276, w_026_277, w_026_278, w_026_279, w_026_280, w_026_281, w_026_282, w_026_283, w_026_284, w_026_285, w_026_286, w_026_287, w_026_288, w_026_289, w_026_290, w_026_292, w_026_293, w_026_294, w_026_295, w_026_296, w_026_297, w_026_298, w_026_299, w_026_300, w_026_301, w_026_302, w_026_303, w_026_304, w_026_305, w_026_306, w_026_308, w_026_309, w_026_310, w_026_311, w_026_312, w_026_313, w_026_314, w_026_315, w_026_316, w_026_317, w_026_318, w_026_319, w_026_320, w_026_321, w_026_322, w_026_323, w_026_324, w_026_325, w_026_326, w_026_327, w_026_328, w_026_329, w_026_330, w_026_331, w_026_332, w_026_333, w_026_334, w_026_335, w_026_336, w_026_337, w_026_338, w_026_339, w_026_340, w_026_341, w_026_342, w_026_343, w_026_344, w_026_345, w_026_346, w_026_347, w_026_348, w_026_349, w_026_350, w_026_352, w_026_353, w_026_354, w_026_355, w_026_356, w_026_357, w_026_358, w_026_359, w_026_360, w_026_361, w_026_362, w_026_363, w_026_364, w_026_365, w_026_366, w_026_367, w_026_368, w_026_369, w_026_370, w_026_371, w_026_372, w_026_373, w_026_374, w_026_375, w_026_376, w_026_377, w_026_379, w_026_380, w_026_381, w_026_382, w_026_383, w_026_384, w_026_385, w_026_386, w_026_388, w_026_389, w_026_390, w_026_391, w_026_392, w_026_393, w_026_394, w_026_395, w_026_396, w_026_397, w_026_398, w_026_399, w_026_400, w_026_401, w_026_402, w_026_403, w_026_404, w_026_405, w_026_406, w_026_407, w_026_408, w_026_409, w_026_410, w_026_411, w_026_412, w_026_413, w_026_414, w_026_415, w_026_416, w_026_417, w_026_418, w_026_419, w_026_420, w_026_421, w_026_422, w_026_423, w_026_424, w_026_425, w_026_426, w_026_427, w_026_428, w_026_429, w_026_430, w_026_431, w_026_432, w_026_433, w_026_434, w_026_435, w_026_436, w_026_437, w_026_438, w_026_439, w_026_440, w_026_441, w_026_442, w_026_443, w_026_444, w_026_445, w_026_446, w_026_447, w_026_448, w_026_449, w_026_450, w_026_451, w_026_452, w_026_453, w_026_454, w_026_455, w_026_456, w_026_457, w_026_458, w_026_459, w_026_460, w_026_461, w_026_462, w_026_463, w_026_464, w_026_465, w_026_466, w_026_467, w_026_468, w_026_469, w_026_470, w_026_471, w_026_472, w_026_473, w_026_474, w_026_475, w_026_476, w_026_477, w_026_478, w_026_479, w_026_480, w_026_482, w_026_483, w_026_484, w_026_485, w_026_486, w_026_487, w_026_489, w_026_490, w_026_491, w_026_492, w_026_493, w_026_494, w_026_495, w_026_496, w_026_497, w_026_498, w_026_499, w_026_500, w_026_501, w_026_502, w_026_503, w_026_504, w_026_505, w_026_506, w_026_507, w_026_508, w_026_509, w_026_510, w_026_511, w_026_512, w_026_513, w_026_514, w_026_515, w_026_516, w_026_517, w_026_518, w_026_519, w_026_520, w_026_522, w_026_523, w_026_524, w_026_525, w_026_526, w_026_527, w_026_528, w_026_529, w_026_530, w_026_531, w_026_532, w_026_533, w_026_534, w_026_535, w_026_536, w_026_537, w_026_538, w_026_539, w_026_540, w_026_541, w_026_542, w_026_543, w_026_544, w_026_545, w_026_546, w_026_547, w_026_548, w_026_549, w_026_550, w_026_551, w_026_552, w_026_553, w_026_554, w_026_555, w_026_556, w_026_557, w_026_558, w_026_559, w_026_562, w_026_563, w_026_564, w_026_565, w_026_566, w_026_567, w_026_568, w_026_569, w_026_570, w_026_571, w_026_573, w_026_574, w_026_575, w_026_577, w_026_578, w_026_579, w_026_580, w_026_581, w_026_582, w_026_583, w_026_584, w_026_585, w_026_586, w_026_587, w_026_588, w_026_589, w_026_590, w_026_591, w_026_592, w_026_593, w_026_594, w_026_595, w_026_596, w_026_597, w_026_598, w_026_599, w_026_600, w_026_602, w_026_603, w_026_604, w_026_605, w_026_606, w_026_607, w_026_608, w_026_609, w_026_610, w_026_611, w_026_612, w_026_613, w_026_614, w_026_615, w_026_616, w_026_617, w_026_618, w_026_619, w_026_620, w_026_621, w_026_622, w_026_623, w_026_624, w_026_625, w_026_626, w_026_627, w_026_628, w_026_629, w_026_630, w_026_631, w_026_632, w_026_633, w_026_634, w_026_635, w_026_637, w_026_638, w_026_639, w_026_640, w_026_641, w_026_642, w_026_643, w_026_644, w_026_645, w_026_646, w_026_647, w_026_648, w_026_649, w_026_650, w_026_651, w_026_652, w_026_653, w_026_654, w_026_655, w_026_656, w_026_657, w_026_658, w_026_659, w_026_660, w_026_661, w_026_662, w_026_664, w_026_665, w_026_666, w_026_667, w_026_668, w_026_669, w_026_670, w_026_671, w_026_672, w_026_673, w_026_674, w_026_675, w_026_676, w_026_677, w_026_678, w_026_679, w_026_680, w_026_681, w_026_682, w_026_683, w_026_684, w_026_685, w_026_686, w_026_687, w_026_688, w_026_689, w_026_690, w_026_691, w_026_692, w_026_693, w_026_694, w_026_695, w_026_696, w_026_697, w_026_698, w_026_699, w_026_700, w_026_701, w_026_702, w_026_703, w_026_704, w_026_705, w_026_706, w_026_707, w_026_708, w_026_709, w_026_710, w_026_711, w_026_712, w_026_713, w_026_714, w_026_715, w_026_716, w_026_717, w_026_718, w_026_719, w_026_720, w_026_721, w_026_722, w_026_723, w_026_724, w_026_725, w_026_727, w_026_728, w_026_729, w_026_730, w_026_731, w_026_732, w_026_733, w_026_734, w_026_735, w_026_736, w_026_737, w_026_738, w_026_739, w_026_740, w_026_741, w_026_742, w_026_743, w_026_744, w_026_745, w_026_746, w_026_747, w_026_748, w_026_749, w_026_750, w_026_751, w_026_752, w_026_753, w_026_754, w_026_755, w_026_756, w_026_757, w_026_758, w_026_759, w_026_760, w_026_761, w_026_762, w_026_763, w_026_764, w_026_765, w_026_766, w_026_767, w_026_768, w_026_769, w_026_770, w_026_771, w_026_772, w_026_773, w_026_774, w_026_775, w_026_776, w_026_777, w_026_778, w_026_779, w_026_780, w_026_781, w_026_782, w_026_783, w_026_784, w_026_786, w_026_787, w_026_788, w_026_790, w_026_791, w_026_793, w_026_794, w_026_795, w_026_796, w_026_797, w_026_798, w_026_799, w_026_800, w_026_801, w_026_802, w_026_803, w_026_804, w_026_805, w_026_806, w_026_807, w_026_808, w_026_809, w_026_810, w_026_811, w_026_812, w_026_813, w_026_814, w_026_815, w_026_816, w_026_817, w_026_818, w_026_819, w_026_820, w_026_821, w_026_822, w_026_823, w_026_824, w_026_825, w_026_826, w_026_827, w_026_828, w_026_829, w_026_830, w_026_831, w_026_832, w_026_833, w_026_834, w_026_835, w_026_836, w_026_838, w_026_839, w_026_841, w_026_842, w_026_843, w_026_844, w_026_845, w_026_846, w_026_847, w_026_848, w_026_849, w_026_850, w_026_851, w_026_852, w_026_853, w_026_854, w_026_856, w_026_857, w_026_858, w_026_859, w_026_860, w_026_861, w_026_862, w_026_863, w_026_864, w_026_865, w_026_866, w_026_867, w_026_868, w_026_869, w_026_870, w_026_871, w_026_872, w_026_874, w_026_875, w_026_876, w_026_877, w_026_878, w_026_879, w_026_880, w_026_881, w_026_883, w_026_884, w_026_885, w_026_886, w_026_887, w_026_888, w_026_889, w_026_890, w_026_891, w_026_892, w_026_893, w_026_894, w_026_896, w_026_897, w_026_899, w_026_900, w_026_901, w_026_902, w_026_903, w_026_904, w_026_905, w_026_906, w_026_907, w_026_908, w_026_909, w_026_910, w_026_911, w_026_912, w_026_913, w_026_914, w_026_915, w_026_916, w_026_917, w_026_918, w_026_919, w_026_920, w_026_921, w_026_922, w_026_923, w_026_924, w_026_925, w_026_927, w_026_928, w_026_929, w_026_930, w_026_931, w_026_932, w_026_933, w_026_934, w_026_935, w_026_936, w_026_937, w_026_938, w_026_939, w_026_940, w_026_941, w_026_942, w_026_943, w_026_944, w_026_945, w_026_946, w_026_947, w_026_948, w_026_949, w_026_950, w_026_951, w_026_952, w_026_953, w_026_954, w_026_955, w_026_956, w_026_957, w_026_958, w_026_959, w_026_960, w_026_961, w_026_962, w_026_963, w_026_964, w_026_965, w_026_966, w_026_967, w_026_968, w_026_969, w_026_970, w_026_971, w_026_972, w_026_973, w_026_974, w_026_975, w_026_976, w_026_977, w_026_978, w_026_979, w_026_980, w_026_981, w_026_982, w_026_983, w_026_984, w_026_985, w_026_986, w_026_987, w_026_988, w_026_989, w_026_990, w_026_991, w_026_993, w_026_994, w_026_995, w_026_996, w_026_997, w_026_998, w_026_999, w_026_1000, w_026_1001, w_026_1002, w_026_1003, w_026_1004, w_026_1005, w_026_1006, w_026_1007, w_026_1009, w_026_1010, w_026_1011, w_026_1012, w_026_1013, w_026_1014, w_026_1016, w_026_1017, w_026_1018, w_026_1019, w_026_1020, w_026_1021, w_026_1022, w_026_1023, w_026_1024, w_026_1025, w_026_1026, w_026_1027, w_026_1028, w_026_1029, w_026_1030, w_026_1031, w_026_1032, w_026_1034, w_026_1035, w_026_1036, w_026_1037, w_026_1038, w_026_1039, w_026_1040, w_026_1041, w_026_1043, w_026_1044, w_026_1045, w_026_1046, w_026_1047, w_026_1048, w_026_1049, w_026_1050, w_026_1051, w_026_1052, w_026_1053, w_026_1054, w_026_1055, w_026_1056, w_026_1057, w_026_1058, w_026_1059, w_026_1060, w_026_1061, w_026_1062, w_026_1063, w_026_1064, w_026_1065, w_026_1066, w_026_1067, w_026_1068, w_026_1069, w_026_1070, w_026_1071, w_026_1072, w_026_1073, w_026_1074, w_026_1075, w_026_1076, w_026_1077, w_026_1078, w_026_1079, w_026_1080, w_026_1081, w_026_1082, w_026_1084, w_026_1085, w_026_1086, w_026_1087, w_026_1088, w_026_1089, w_026_1090, w_026_1091, w_026_1092, w_026_1093, w_026_1094, w_026_1095, w_026_1096, w_026_1097, w_026_1098, w_026_1099, w_026_1100, w_026_1101, w_026_1102, w_026_1103, w_026_1105, w_026_1106, w_026_1107, w_026_1108, w_026_1109, w_026_1110, w_026_1111, w_026_1112, w_026_1113, w_026_1114, w_026_1115, w_026_1116, w_026_1117, w_026_1119, w_026_1120, w_026_1121, w_026_1122, w_026_1123, w_026_1124, w_026_1125, w_026_1126, w_026_1127, w_026_1128, w_026_1129, w_026_1131, w_026_1132, w_026_1133, w_026_1134, w_026_1135, w_026_1136, w_026_1137, w_026_1138, w_026_1139, w_026_1140, w_026_1141, w_026_1142, w_026_1144, w_026_1145, w_026_1146, w_026_1147, w_026_1148, w_026_1149, w_026_1150, w_026_1151, w_026_1152, w_026_1153, w_026_1154, w_026_1155, w_026_1156, w_026_1157, w_026_1158, w_026_1159, w_026_1160, w_026_1161, w_026_1162, w_026_1163, w_026_1164, w_026_1165, w_026_1167, w_026_1168, w_026_1169, w_026_1170, w_026_1171, w_026_1172, w_026_1173, w_026_1174, w_026_1175, w_026_1176, w_026_1177, w_026_1178, w_026_1179, w_026_1180, w_026_1181, w_026_1182, w_026_1183, w_026_1184, w_026_1185, w_026_1186, w_026_1187, w_026_1188, w_026_1189, w_026_1190, w_026_1191, w_026_1192, w_026_1193, w_026_1194, w_026_1195, w_026_1196, w_026_1197, w_026_1198, w_026_1199, w_026_1200, w_026_1201, w_026_1202, w_026_1203, w_026_1204, w_026_1205, w_026_1206, w_026_1207, w_026_1208, w_026_1209, w_026_1210, w_026_1211, w_026_1212, w_026_1213, w_026_1214, w_026_1215, w_026_1216, w_026_1217, w_026_1218, w_026_1219, w_026_1220, w_026_1221, w_026_1222, w_026_1223, w_026_1224, w_026_1225, w_026_1227, w_026_1228, w_026_1229, w_026_1231, w_026_1232, w_026_1233, w_026_1234, w_026_1235, w_026_1236, w_026_1237, w_026_1238, w_026_1241, w_026_1243, w_026_1244, w_026_1245, w_026_1246, w_026_1247, w_026_1248, w_026_1249, w_026_1250, w_026_1251, w_026_1252, w_026_1253, w_026_1254, w_026_1255, w_026_1256, w_026_1257, w_026_1258, w_026_1260, w_026_1261, w_026_1262, w_026_1263, w_026_1264, w_026_1265, w_026_1266, w_026_1267, w_026_1268, w_026_1269, w_026_1270, w_026_1271, w_026_1272, w_026_1273, w_026_1274, w_026_1275, w_026_1276, w_026_1277, w_026_1278, w_026_1279, w_026_1280, w_026_1282, w_026_1283, w_026_1284, w_026_1285, w_026_1286, w_026_1287, w_026_1289, w_026_1290, w_026_1291, w_026_1292, w_026_1293, w_026_1294, w_026_1295, w_026_1296, w_026_1297, w_026_1298, w_026_1299, w_026_1300, w_026_1301, w_026_1302, w_026_1303, w_026_1304, w_026_1305, w_026_1306, w_026_1307, w_026_1308, w_026_1309, w_026_1311, w_026_1312, w_026_1314, w_026_1315, w_026_1316, w_026_1317, w_026_1318, w_026_1319, w_026_1320, w_026_1321, w_026_1322, w_026_1323, w_026_1324, w_026_1325, w_026_1327, w_026_1328, w_026_1329, w_026_1330, w_026_1331, w_026_1332, w_026_1333, w_026_1334, w_026_1335, w_026_1336, w_026_1337, w_026_1339, w_026_1340, w_026_1341, w_026_1342, w_026_1343, w_026_1344, w_026_1345, w_026_1346, w_026_1347, w_026_1348, w_026_1349, w_026_1350, w_026_1351, w_026_1352, w_026_1353, w_026_1354, w_026_1355, w_026_1356, w_026_1357, w_026_1358, w_026_1359, w_026_1360, w_026_1361, w_026_1362, w_026_1363, w_026_1364, w_026_1365, w_026_1366, w_026_1367, w_026_1368, w_026_1369, w_026_1372, w_026_1373, w_026_1374, w_026_1375, w_026_1376, w_026_1377, w_026_1379, w_026_1380, w_026_1381, w_026_1382, w_026_1383, w_026_1385, w_026_1386, w_026_1387, w_026_1388, w_026_1389, w_026_1390, w_026_1391, w_026_1392, w_026_1393, w_026_1394, w_026_1395, w_026_1396, w_026_1397, w_026_1398, w_026_1399, w_026_1400, w_026_1401, w_026_1402, w_026_1403, w_026_1404, w_026_1405, w_026_1406, w_026_1407, w_026_1408, w_026_1409, w_026_1410, w_026_1411, w_026_1412, w_026_1413, w_026_1414, w_026_1415, w_026_1416, w_026_1417, w_026_1418, w_026_1419, w_026_1420, w_026_1422, w_026_1423, w_026_1424, w_026_1425, w_026_1426, w_026_1427, w_026_1428, w_026_1429, w_026_1430, w_026_1431, w_026_1432, w_026_1433, w_026_1435, w_026_1436, w_026_1437, w_026_1439, w_026_1442, w_026_1443, w_026_1445, w_026_1446, w_026_1447, w_026_1448, w_026_1449, w_026_1450, w_026_1451, w_026_1452, w_026_1453, w_026_1454, w_026_1455, w_026_1456, w_026_1458, w_026_1459, w_026_1460, w_026_1461, w_026_1462, w_026_1463, w_026_1464, w_026_1465, w_026_1466, w_026_1467, w_026_1469, w_026_1470, w_026_1471, w_026_1472, w_026_1473, w_026_1474, w_026_1475, w_026_1476, w_026_1477, w_026_1478, w_026_1479, w_026_1480, w_026_1481, w_026_1482, w_026_1483, w_026_1484, w_026_1485, w_026_1486, w_026_1487, w_026_1488, w_026_1489, w_026_1490, w_026_1491, w_026_1492, w_026_1493, w_026_1494, w_026_1495, w_026_1496, w_026_1497, w_026_1498, w_026_1500, w_026_1501, w_026_1502, w_026_1503, w_026_1504, w_026_1505, w_026_1506, w_026_1507, w_026_1508, w_026_1509, w_026_1510, w_026_1511, w_026_1512, w_026_1514, w_026_1515, w_026_1516, w_026_1517, w_026_1518, w_026_1519, w_026_1520, w_026_1521, w_026_1522, w_026_1523, w_026_1525, w_026_1526, w_026_1527, w_026_1528, w_026_1529, w_026_1531, w_026_1532, w_026_1534, w_026_1535, w_026_1536, w_026_1537, w_026_1538, w_026_1539, w_026_1540, w_026_1541, w_026_1543, w_026_1544, w_026_1545, w_026_1546, w_026_1547, w_026_1548, w_026_1549, w_026_1550, w_026_1551, w_026_1552, w_026_1553, w_026_1554, w_026_1555, w_026_1556, w_026_1557, w_026_1558, w_026_1559, w_026_1560, w_026_1561, w_026_1562, w_026_1563, w_026_1564, w_026_1565, w_026_1566, w_026_1567, w_026_1568, w_026_1569, w_026_1571, w_026_1572, w_026_1575, w_026_1576, w_026_1577, w_026_1578, w_026_1579, w_026_1580, w_026_1581, w_026_1582, w_026_1583, w_026_1584, w_026_1585, w_026_1586, w_026_1587, w_026_1588, w_026_1589, w_026_1590, w_026_1591, w_026_1592, w_026_1593, w_026_1594, w_026_1595, w_026_1596, w_026_1597, w_026_1598, w_026_1599, w_026_1600, w_026_1602, w_026_1603, w_026_1604, w_026_1605, w_026_1606, w_026_1607, w_026_1608, w_026_1609, w_026_1610, w_026_1611, w_026_1612, w_026_1613, w_026_1614, w_026_1615, w_026_1616, w_026_1617, w_026_1618, w_026_1619, w_026_1620, w_026_1621, w_026_1622, w_026_1623, w_026_1624, w_026_1625, w_026_1627, w_026_1628, w_026_1629, w_026_1631, w_026_1632, w_026_1633, w_026_1634, w_026_1635, w_026_1636, w_026_1637, w_026_1638, w_026_1640, w_026_1641, w_026_1642, w_026_1643, w_026_1644, w_026_1645, w_026_1646, w_026_1647, w_026_1648, w_026_1649, w_026_1650, w_026_1651, w_026_1652, w_026_1653, w_026_1654, w_026_1656, w_026_1657, w_026_1658, w_026_1659, w_026_1660, w_026_1661, w_026_1662, w_026_1663, w_026_1664, w_026_1665, w_026_1666, w_026_1667, w_026_1668, w_026_1669, w_026_1670, w_026_1671, w_026_1672, w_026_1673, w_026_1674, w_026_1675, w_026_1676, w_026_1678, w_026_1679, w_026_1680, w_026_1681, w_026_1682, w_026_1683, w_026_1684, w_026_1685, w_026_1686, w_026_1687, w_026_1688, w_026_1689, w_026_1691, w_026_1693, w_026_1694, w_026_1695, w_026_1696, w_026_1697, w_026_1698, w_026_1699, w_026_1702, w_026_1703, w_026_1704, w_026_1705, w_026_1706, w_026_1707, w_026_1708, w_026_1709, w_026_1711, w_026_1713, w_026_1714, w_026_1715, w_026_1716, w_026_1717, w_026_1718, w_026_1719, w_026_1720, w_026_1724, w_026_1725, w_026_1727, w_026_1728, w_026_1729, w_026_1730, w_026_1731, w_026_1732, w_026_1733, w_026_1734, w_026_1735, w_026_1736, w_026_1737, w_026_1738, w_026_1739, w_026_1740, w_026_1741, w_026_1742, w_026_1743, w_026_1744, w_026_1745, w_026_1746, w_026_1747, w_026_1748, w_026_1749, w_026_1750, w_026_1751, w_026_1752, w_026_1753, w_026_1754, w_026_1755, w_026_1757, w_026_1758, w_026_1759, w_026_1760, w_026_1761, w_026_1762, w_026_1763, w_026_1764, w_026_1765, w_026_1766, w_026_1767, w_026_1768, w_026_1769, w_026_1770, w_026_1772, w_026_1773, w_026_1774, w_026_1775, w_026_1777, w_026_1778, w_026_1779, w_026_1780, w_026_1781, w_026_1782, w_026_1783, w_026_1784, w_026_1785, w_026_1786, w_026_1788, w_026_1789, w_026_1790, w_026_1791, w_026_1792, w_026_1793, w_026_1794, w_026_1795, w_026_1796, w_026_1798, w_026_1799, w_026_1800, w_026_1801, w_026_1802, w_026_1803, w_026_1805, w_026_1806, w_026_1807, w_026_1808, w_026_1809, w_026_1811, w_026_1812, w_026_1813, w_026_1814, w_026_1815, w_026_1817, w_026_1818, w_026_1819, w_026_1820, w_026_1821, w_026_1822, w_026_1823, w_026_1824, w_026_1826, w_026_1827, w_026_1828, w_026_1829, w_026_1830, w_026_1831, w_026_1832, w_026_1833, w_026_1834, w_026_1835, w_026_1836, w_026_1838, w_026_1839, w_026_1840, w_026_1841, w_026_1842, w_026_1843, w_026_1844, w_026_1845, w_026_1846, w_026_1847, w_026_1848, w_026_1849, w_026_1850, w_026_1852, w_026_1853, w_026_1854, w_026_1855, w_026_1856, w_026_1857, w_026_1858, w_026_1859, w_026_1860, w_026_1861, w_026_1862, w_026_1863, w_026_1864, w_026_1865, w_026_1866, w_026_1867, w_026_1868, w_026_1869, w_026_1870, w_026_1871, w_026_1872, w_026_1873, w_026_1874, w_026_1875, w_026_1876, w_026_1877, w_026_1879, w_026_1880, w_026_1881, w_026_1882, w_026_1883, w_026_1884, w_026_1885, w_026_1886, w_026_1887, w_026_1888, w_026_1889, w_026_1890, w_026_1891, w_026_1892, w_026_1894, w_026_1895, w_026_1896, w_026_1897, w_026_1898, w_026_1899, w_026_1900, w_026_1901, w_026_1902, w_026_1903, w_026_1904, w_026_1905, w_026_1907, w_026_1909, w_026_1910, w_026_1912, w_026_1913, w_026_1914, w_026_1915, w_026_1916, w_026_1917, w_026_1918, w_026_1919, w_026_1920, w_026_1921, w_026_1922, w_026_1923, w_026_1925, w_026_1926, w_026_1928, w_026_1929, w_026_1930, w_026_1931, w_026_1932, w_026_1933, w_026_1934, w_026_1935, w_026_1936, w_026_1937, w_026_1938, w_026_1939, w_026_1940, w_026_1941, w_026_1942, w_026_1943, w_026_1944, w_026_1945, w_026_1946, w_026_1947, w_026_1948, w_026_1949, w_026_1950, w_026_1951, w_026_1952, w_026_1953, w_026_1954, w_026_1955, w_026_1956, w_026_1957, w_026_1958, w_026_1959, w_026_1960, w_026_1961, w_026_1962, w_026_1963, w_026_1964, w_026_1966, w_026_1967, w_026_1968, w_026_1970, w_026_1971, w_026_1972, w_026_1974, w_026_1975, w_026_1977, w_026_1978, w_026_1979, w_026_1981, w_026_1983, w_026_1984, w_026_1985, w_026_1986, w_026_1987, w_026_1988, w_026_1989, w_026_1990, w_026_1991, w_026_1992, w_026_1993, w_026_1994, w_026_1995, w_026_1996, w_026_1998, w_026_1999, w_026_2000, w_026_2001, w_026_2002, w_026_2003, w_026_2004, w_026_2005, w_026_2006, w_026_2007, w_026_2008, w_026_2009, w_026_2012, w_026_2014, w_026_2015, w_026_2016, w_026_2017, w_026_2018, w_026_2019, w_026_2020, w_026_2021, w_026_2022, w_026_2023, w_026_2024, w_026_2025, w_026_2026, w_026_2027, w_026_2028, w_026_2029, w_026_2030, w_026_2031, w_026_2033, w_026_2034, w_026_2035, w_026_2036, w_026_2037, w_026_2039, w_026_2040, w_026_2041, w_026_2042, w_026_2043, w_026_2044, w_026_2045, w_026_2048, w_026_2049, w_026_2050, w_026_2051, w_026_2052, w_026_2054, w_026_2055, w_026_2056, w_026_2057, w_026_2058, w_026_2059, w_026_2060, w_026_2061, w_026_2062, w_026_2063, w_026_2064, w_026_2065, w_026_2066, w_026_2067, w_026_2068, w_026_2069, w_026_2070, w_026_2072, w_026_2073, w_026_2074, w_026_2075, w_026_2076, w_026_2077, w_026_2078, w_026_2079, w_026_2080, w_026_2081, w_026_2082, w_026_2083, w_026_2084, w_026_2085, w_026_2086, w_026_2087, w_026_2088, w_026_2089, w_026_2090, w_026_2091, w_026_2092, w_026_2093, w_026_2094, w_026_2095, w_026_2096, w_026_2097, w_026_2099, w_026_2100, w_026_2101, w_026_2102, w_026_2103, w_026_2104, w_026_2105, w_026_2106, w_026_2107, w_026_2108, w_026_2109, w_026_2110, w_026_2111, w_026_2112, w_026_2113, w_026_2114, w_026_2115, w_026_2116, w_026_2117, w_026_2118, w_026_2119, w_026_2120, w_026_2121, w_026_2122, w_026_2123, w_026_2124, w_026_2125, w_026_2126, w_026_2127, w_026_2128, w_026_2129, w_026_2130, w_026_2131, w_026_2132, w_026_2133, w_026_2134, w_026_2135, w_026_2136, w_026_2137, w_026_2138, w_026_2139, w_026_2140, w_026_2141, w_026_2142, w_026_2143, w_026_2144, w_026_2146, w_026_2147, w_026_2148, w_026_2149, w_026_2150, w_026_2151, w_026_2152, w_026_2153, w_026_2154, w_026_2155, w_026_2156, w_026_2157, w_026_2158, w_026_2160, w_026_2161, w_026_2162, w_026_2163, w_026_2164, w_026_2165, w_026_2166, w_026_2167, w_026_2168, w_026_2169, w_026_2170, w_026_2171, w_026_2172, w_026_2173, w_026_2174, w_026_2175, w_026_2176, w_026_2177, w_026_2178, w_026_2179, w_026_2180, w_026_2181, w_026_2182, w_026_2183, w_026_2184, w_026_2185, w_026_2186, w_026_2187, w_026_2189, w_026_2190, w_026_2191, w_026_2192, w_026_2193, w_026_2194, w_026_2195, w_026_2197, w_026_2198, w_026_2199, w_026_2201, w_026_2202, w_026_2203, w_026_2204, w_026_2205, w_026_2206, w_026_2207, w_026_2208, w_026_2209, w_026_2210, w_026_2211, w_026_2212, w_026_2213, w_026_2214, w_026_2215, w_026_2216, w_026_2217, w_026_2218, w_026_2219, w_026_2221, w_026_2222, w_026_2223, w_026_2224, w_026_2225, w_026_2226, w_026_2227, w_026_2228, w_026_2229, w_026_2230, w_026_2231, w_026_2232, w_026_2233, w_026_2234, w_026_2235, w_026_2236, w_026_2237, w_026_2238, w_026_2239, w_026_2240, w_026_2241, w_026_2242, w_026_2243, w_026_2244, w_026_2245, w_026_2246, w_026_2247, w_026_2248, w_026_2249, w_026_2250, w_026_2251, w_026_2252, w_026_2253, w_026_2255, w_026_2256, w_026_2257, w_026_2258, w_026_2259, w_026_2260, w_026_2262, w_026_2263, w_026_2264, w_026_2265, w_026_2266, w_026_2267, w_026_2268, w_026_2269, w_026_2270, w_026_2271, w_026_2272, w_026_2273, w_026_2274, w_026_2275, w_026_2276, w_026_2277, w_026_2278, w_026_2279, w_026_2280, w_026_2281, w_026_2282, w_026_2283, w_026_2284, w_026_2285, w_026_2286, w_026_2287, w_026_2288, w_026_2289, w_026_2290, w_026_2292, w_026_2293, w_026_2294, w_026_2295, w_026_2296, w_026_2298, w_026_2299, w_026_2300, w_026_2301, w_026_2302, w_026_2303, w_026_2305, w_026_2306, w_026_2307, w_026_2308, w_026_2309, w_026_2310, w_026_2312, w_026_2313, w_026_2314, w_026_2315, w_026_2316, w_026_2317, w_026_2319, w_026_2320, w_026_2321, w_026_2322, w_026_2323, w_026_2324, w_026_2326, w_026_2327, w_026_2328, w_026_2329, w_026_2330, w_026_2331, w_026_2332, w_026_2336, w_026_2337, w_026_2338, w_026_2339, w_026_2340, w_026_2341, w_026_2342, w_026_2344, w_026_2345, w_026_2346, w_026_2347, w_026_2348, w_026_2349, w_026_2351, w_026_2352, w_026_2353, w_026_2355, w_026_2356, w_026_2357, w_026_2358, w_026_2359, w_026_2360, w_026_2362, w_026_2363, w_026_2365, w_026_2366, w_026_2367, w_026_2368, w_026_2369, w_026_2370, w_026_2371, w_026_2372, w_026_2373, w_026_2374, w_026_2375, w_026_2376, w_026_2377, w_026_2378, w_026_2379, w_026_2380, w_026_2381, w_026_2382, w_026_2383, w_026_2386, w_026_2388, w_026_2389, w_026_2390, w_026_2391, w_026_2392, w_026_2394, w_026_2395, w_026_2396, w_026_2397, w_026_2398, w_026_2399, w_026_2400, w_026_2401, w_026_2402, w_026_2403, w_026_2404, w_026_2405, w_026_2406, w_026_2407, w_026_2408, w_026_2409, w_026_2410, w_026_2411, w_026_2412, w_026_2413, w_026_2414, w_026_2415, w_026_2416, w_026_2417, w_026_2418, w_026_2419, w_026_2420, w_026_2421, w_026_2422, w_026_2423, w_026_2425, w_026_2426, w_026_2427, w_026_2428, w_026_2429, w_026_2431, w_026_2432, w_026_2433, w_026_2434, w_026_2435, w_026_2436, w_026_2437, w_026_2438, w_026_2439, w_026_2440, w_026_2441, w_026_2442, w_026_2443, w_026_2444, w_026_2445, w_026_2446, w_026_2447, w_026_2449, w_026_2450, w_026_2451, w_026_2452, w_026_2453, w_026_2454, w_026_2455, w_026_2456, w_026_2457, w_026_2458, w_026_2459, w_026_2460, w_026_2461, w_026_2462, w_026_2463, w_026_2464, w_026_2465, w_026_2466, w_026_2467, w_026_2468, w_026_2469, w_026_2470, w_026_2471, w_026_2472, w_026_2473, w_026_2474, w_026_2475, w_026_2476, w_026_2477, w_026_2478, w_026_2479, w_026_2480, w_026_2481, w_026_2482, w_026_2483, w_026_2484, w_026_2485, w_026_2486, w_026_2487, w_026_2489, w_026_2490, w_026_2491, w_026_2492, w_026_2493, w_026_2494, w_026_2495, w_026_2496, w_026_2497, w_026_2498, w_026_2499, w_026_2500, w_026_2502, w_026_2503, w_026_2504, w_026_2505, w_026_2506, w_026_2507, w_026_2508, w_026_2509, w_026_2510, w_026_2511, w_026_2512, w_026_2513, w_026_2516, w_026_2517, w_026_2519, w_026_2520, w_026_2521, w_026_2522, w_026_2523, w_026_2524, w_026_2526, w_026_2527, w_026_2528, w_026_2529, w_026_2530, w_026_2531, w_026_2532, w_026_2533, w_026_2534, w_026_2535, w_026_2537, w_026_2538, w_026_2539, w_026_2540, w_026_2542, w_026_2543, w_026_2544, w_026_2545, w_026_2546, w_026_2547, w_026_2548, w_026_2549, w_026_2550, w_026_2551, w_026_2552, w_026_2553, w_026_2554, w_026_2555, w_026_2556, w_026_2557, w_026_2558, w_026_2559, w_026_2560, w_026_2561, w_026_2562, w_026_2563, w_026_2564, w_026_2565, w_026_2566, w_026_2567, w_026_2568, w_026_2569, w_026_2570, w_026_2571, w_026_2573, w_026_2575, w_026_2576, w_026_2577, w_026_2578, w_026_2579, w_026_2581, w_026_2582, w_026_2583, w_026_2584, w_026_2585, w_026_2586, w_026_2587, w_026_2588, w_026_2589, w_026_2590, w_026_2591, w_026_2592, w_026_2593, w_026_2594, w_026_2596, w_026_2597, w_026_2598, w_026_2599, w_026_2600, w_026_2601, w_026_2603, w_026_2604, w_026_2605, w_026_2606, w_026_2608, w_026_2609, w_026_2610, w_026_2611, w_026_2612, w_026_2613, w_026_2614, w_026_2615, w_026_2616, w_026_2617, w_026_2618, w_026_2619, w_026_2620, w_026_2621, w_026_2622, w_026_2623, w_026_2624, w_026_2625, w_026_2626, w_026_2628, w_026_2629, w_026_2630, w_026_2631, w_026_2632, w_026_2633, w_026_2634, w_026_2635, w_026_2636, w_026_2637, w_026_2638, w_026_2640, w_026_2641, w_026_2642, w_026_2643, w_026_2644, w_026_2645, w_026_2646, w_026_2647, w_026_2648, w_026_2649, w_026_2650, w_026_2651, w_026_2652, w_026_2653, w_026_2654, w_026_2655, w_026_2656, w_026_2657, w_026_2658, w_026_2659, w_026_2660, w_026_2662, w_026_2663, w_026_2664, w_026_2666, w_026_2667, w_026_2668, w_026_2670, w_026_2671, w_026_2672, w_026_2673, w_026_2674, w_026_2675, w_026_2676, w_026_2677, w_026_2678, w_026_2679, w_026_2680, w_026_2681, w_026_2682, w_026_2684, w_026_2685, w_026_2686, w_026_2687, w_026_2688, w_026_2689, w_026_2690, w_026_2691, w_026_2692, w_026_2693, w_026_2694, w_026_2695, w_026_2696, w_026_2697, w_026_2698, w_026_2699, w_026_2700, w_026_2701, w_026_2702, w_026_2703, w_026_2704, w_026_2705, w_026_2706, w_026_2707, w_026_2708, w_026_2709, w_026_2710, w_026_2711, w_026_2712, w_026_2713, w_026_2714, w_026_2715, w_026_2716, w_026_2717, w_026_2718, w_026_2719, w_026_2720, w_026_2721, w_026_2722, w_026_2723, w_026_2724, w_026_2725, w_026_2726, w_026_2727, w_026_2728, w_026_2729, w_026_2730, w_026_2732, w_026_2733, w_026_2734, w_026_2735, w_026_2736, w_026_2737, w_026_2738, w_026_2740, w_026_2741, w_026_2742, w_026_2743, w_026_2744, w_026_2745, w_026_2746, w_026_2747, w_026_2748, w_026_2749, w_026_2750, w_026_2751, w_026_2752, w_026_2753, w_026_2754, w_026_2755, w_026_2756, w_026_2758, w_026_2759, w_026_2760, w_026_2761, w_026_2762, w_026_2763, w_026_2764, w_026_2765, w_026_2766, w_026_2767, w_026_2768, w_026_2769, w_026_2770, w_026_2771, w_026_2772, w_026_2773, w_026_2775, w_026_2776, w_026_2777, w_026_2778, w_026_2779, w_026_2780, w_026_2781, w_026_2782, w_026_2785, w_026_2786, w_026_2787, w_026_2788, w_026_2789, w_026_2790, w_026_2791, w_026_2793, w_026_2794, w_026_2795, w_026_2796, w_026_2797, w_026_2798, w_026_2799, w_026_2800, w_026_2801, w_026_2802, w_026_2804, w_026_2805, w_026_2806, w_026_2807, w_026_2808, w_026_2809, w_026_2810, w_026_2812, w_026_2813, w_026_2814, w_026_2815, w_026_2816, w_026_2817, w_026_2818, w_026_2819, w_026_2820, w_026_2821, w_026_2822, w_026_2823, w_026_2824, w_026_2825, w_026_2826, w_026_2827, w_026_2828, w_026_2829, w_026_2830, w_026_2831, w_026_2832, w_026_2833, w_026_2834, w_026_2835, w_026_2836, w_026_2838, w_026_2839, w_026_2840, w_026_2842, w_026_2843, w_026_2844, w_026_2845, w_026_2846, w_026_2847, w_026_2848, w_026_2849, w_026_2850, w_026_2851, w_026_2853, w_026_2854, w_026_2856, w_026_2857, w_026_2858, w_026_2859, w_026_2860, w_026_2861, w_026_2863, w_026_2865, w_026_2866, w_026_2867, w_026_2868, w_026_2869, w_026_2871, w_026_2872, w_026_2873, w_026_2874, w_026_2877, w_026_2878, w_026_2879, w_026_2880, w_026_2881, w_026_2882, w_026_2884, w_026_2885, w_026_2886, w_026_2887, w_026_2888, w_026_2889, w_026_2890, w_026_2891, w_026_2892, w_026_2893, w_026_2894, w_026_2895, w_026_2896, w_026_2897, w_026_2898, w_026_2899, w_026_2900, w_026_2901, w_026_2902, w_026_2903, w_026_2904, w_026_2905, w_026_2906, w_026_2907, w_026_2908, w_026_2909, w_026_2910, w_026_2911, w_026_2912, w_026_2913, w_026_2914, w_026_2916, w_026_2917, w_026_2918, w_026_2919, w_026_2920, w_026_2921, w_026_2922, w_026_2924, w_026_2925, w_026_2926, w_026_2927, w_026_2928, w_026_2929;
  wire w_027_000, w_027_001, w_027_002, w_027_003, w_027_004, w_027_005, w_027_006, w_027_007, w_027_008, w_027_009, w_027_010, w_027_011, w_027_012, w_027_013, w_027_014, w_027_015, w_027_016, w_027_017, w_027_018, w_027_019, w_027_020, w_027_021, w_027_022, w_027_023, w_027_024, w_027_025, w_027_026, w_027_027, w_027_028, w_027_029, w_027_030, w_027_031, w_027_032, w_027_033, w_027_034, w_027_035, w_027_036, w_027_037, w_027_038, w_027_039, w_027_040, w_027_041, w_027_042, w_027_043, w_027_044, w_027_045, w_027_046, w_027_047, w_027_048, w_027_049, w_027_050, w_027_051, w_027_052, w_027_053, w_027_054, w_027_055, w_027_056, w_027_057, w_027_058, w_027_059, w_027_060, w_027_061, w_027_062, w_027_063, w_027_064, w_027_065, w_027_066, w_027_067, w_027_068, w_027_069, w_027_070, w_027_071, w_027_072, w_027_073, w_027_074, w_027_075, w_027_076, w_027_077, w_027_078, w_027_079, w_027_080, w_027_081, w_027_082, w_027_083, w_027_084, w_027_085, w_027_086, w_027_087, w_027_088, w_027_089, w_027_090, w_027_091, w_027_092, w_027_093, w_027_094, w_027_095, w_027_096, w_027_097, w_027_098, w_027_099, w_027_100, w_027_101, w_027_102, w_027_103, w_027_104, w_027_105, w_027_106, w_027_107, w_027_108, w_027_109, w_027_110, w_027_111, w_027_112, w_027_113, w_027_114, w_027_115, w_027_116, w_027_117, w_027_118, w_027_119, w_027_120, w_027_121, w_027_122, w_027_123, w_027_124, w_027_125, w_027_126, w_027_127, w_027_128, w_027_129, w_027_130, w_027_131, w_027_132, w_027_133, w_027_134, w_027_135, w_027_136, w_027_137, w_027_138, w_027_139, w_027_140, w_027_141, w_027_142, w_027_143, w_027_144, w_027_145, w_027_146, w_027_147, w_027_148, w_027_149, w_027_150, w_027_151, w_027_152, w_027_153, w_027_154, w_027_155, w_027_156, w_027_157, w_027_158, w_027_159, w_027_160, w_027_161, w_027_162, w_027_163, w_027_164, w_027_165, w_027_166, w_027_167, w_027_168, w_027_169, w_027_170, w_027_171, w_027_172, w_027_173, w_027_174, w_027_175, w_027_176, w_027_177, w_027_178, w_027_179, w_027_180, w_027_181, w_027_182, w_027_183, w_027_184, w_027_185, w_027_186, w_027_187, w_027_188, w_027_189, w_027_190, w_027_191, w_027_192, w_027_193, w_027_194, w_027_195, w_027_196, w_027_197, w_027_198, w_027_199, w_027_200, w_027_201, w_027_202, w_027_203, w_027_204, w_027_205, w_027_206, w_027_207, w_027_208, w_027_209, w_027_210, w_027_211, w_027_212, w_027_213, w_027_214, w_027_215, w_027_216, w_027_217, w_027_218, w_027_219, w_027_220, w_027_221, w_027_222, w_027_223, w_027_224, w_027_225, w_027_226, w_027_227, w_027_228, w_027_229, w_027_230, w_027_231, w_027_232, w_027_233, w_027_234, w_027_235, w_027_236, w_027_237, w_027_238, w_027_239, w_027_240, w_027_241, w_027_242, w_027_243, w_027_244, w_027_245, w_027_246, w_027_247, w_027_248, w_027_249, w_027_250, w_027_251, w_027_252, w_027_253, w_027_254, w_027_255, w_027_256, w_027_257, w_027_258, w_027_259, w_027_260, w_027_261, w_027_262, w_027_263, w_027_264, w_027_265, w_027_266, w_027_267, w_027_268, w_027_269, w_027_270, w_027_271, w_027_272, w_027_273, w_027_274, w_027_275, w_027_276, w_027_277, w_027_278, w_027_279, w_027_280, w_027_281, w_027_282, w_027_283, w_027_284, w_027_285, w_027_286, w_027_287, w_027_288, w_027_289, w_027_290, w_027_291, w_027_292, w_027_293, w_027_294, w_027_295, w_027_296, w_027_297, w_027_298, w_027_299, w_027_300, w_027_301, w_027_302, w_027_303, w_027_304, w_027_305, w_027_306, w_027_307, w_027_308, w_027_309, w_027_310, w_027_311, w_027_312, w_027_313, w_027_314, w_027_315, w_027_316, w_027_317, w_027_318, w_027_319, w_027_320, w_027_321, w_027_322, w_027_323, w_027_324, w_027_325, w_027_326, w_027_327, w_027_328, w_027_329, w_027_330, w_027_331, w_027_332, w_027_333, w_027_334, w_027_335, w_027_336, w_027_337, w_027_338, w_027_339, w_027_340, w_027_341, w_027_342, w_027_343, w_027_344, w_027_345, w_027_346, w_027_347, w_027_348, w_027_349, w_027_350, w_027_351, w_027_352, w_027_353, w_027_354, w_027_355, w_027_356, w_027_357, w_027_358, w_027_359, w_027_360, w_027_361, w_027_362;
  wire w_028_000, w_028_001, w_028_002, w_028_003, w_028_004, w_028_005, w_028_006, w_028_007, w_028_008, w_028_009, w_028_010, w_028_011, w_028_012, w_028_013, w_028_014, w_028_015, w_028_016, w_028_017, w_028_018, w_028_019, w_028_020, w_028_021, w_028_022, w_028_023, w_028_024, w_028_025, w_028_026, w_028_027, w_028_028, w_028_029, w_028_030, w_028_031, w_028_032, w_028_033, w_028_034, w_028_035, w_028_036, w_028_037, w_028_038, w_028_039, w_028_040, w_028_041, w_028_042, w_028_043, w_028_044, w_028_045, w_028_046, w_028_047, w_028_048, w_028_049, w_028_050, w_028_051, w_028_052, w_028_053, w_028_054, w_028_055, w_028_056, w_028_057, w_028_058, w_028_059, w_028_060, w_028_061, w_028_062, w_028_063, w_028_064, w_028_065, w_028_066, w_028_067, w_028_068, w_028_069, w_028_070, w_028_071, w_028_072, w_028_073, w_028_074, w_028_075, w_028_076, w_028_077, w_028_078, w_028_079, w_028_080, w_028_081, w_028_082, w_028_083, w_028_084, w_028_085, w_028_086, w_028_087, w_028_088, w_028_089, w_028_090, w_028_091, w_028_092, w_028_093, w_028_094, w_028_095, w_028_096, w_028_097, w_028_098, w_028_099, w_028_100, w_028_101, w_028_102, w_028_103, w_028_104, w_028_105, w_028_106, w_028_107, w_028_108, w_028_109, w_028_110, w_028_111, w_028_112, w_028_113, w_028_114, w_028_115, w_028_116, w_028_117, w_028_118, w_028_119, w_028_120, w_028_121, w_028_122, w_028_123, w_028_124, w_028_125, w_028_126, w_028_127, w_028_128, w_028_129, w_028_130, w_028_131, w_028_132, w_028_133, w_028_134, w_028_135, w_028_136, w_028_137, w_028_138, w_028_139, w_028_140, w_028_141, w_028_142, w_028_143, w_028_144, w_028_145, w_028_146, w_028_147, w_028_148, w_028_149, w_028_150, w_028_151, w_028_152, w_028_153, w_028_154, w_028_155, w_028_156, w_028_157, w_028_158, w_028_159, w_028_160, w_028_161, w_028_162, w_028_163, w_028_164, w_028_165, w_028_166, w_028_167, w_028_168, w_028_169, w_028_170, w_028_171, w_028_172, w_028_173, w_028_174, w_028_175, w_028_176, w_028_177, w_028_178, w_028_179, w_028_180, w_028_181, w_028_182, w_028_183, w_028_184, w_028_185, w_028_186, w_028_187, w_028_188, w_028_189, w_028_190, w_028_191, w_028_192, w_028_193, w_028_194, w_028_195, w_028_196, w_028_197, w_028_198, w_028_199, w_028_200, w_028_201, w_028_202, w_028_203, w_028_204, w_028_205, w_028_206, w_028_207, w_028_208, w_028_209, w_028_210, w_028_211, w_028_212, w_028_213, w_028_214, w_028_215, w_028_216, w_028_217, w_028_218, w_028_219, w_028_220, w_028_221, w_028_222, w_028_223, w_028_224, w_028_225, w_028_226, w_028_227, w_028_228, w_028_229, w_028_230, w_028_231, w_028_232, w_028_233, w_028_234, w_028_235, w_028_236, w_028_237, w_028_238, w_028_239, w_028_240, w_028_241, w_028_242, w_028_243, w_028_244, w_028_245, w_028_246, w_028_247, w_028_248, w_028_249, w_028_250, w_028_251, w_028_252, w_028_253, w_028_254, w_028_255, w_028_256, w_028_257, w_028_258, w_028_259, w_028_260, w_028_261, w_028_262, w_028_263, w_028_264, w_028_265, w_028_266, w_028_267, w_028_268, w_028_269, w_028_270, w_028_271, w_028_272, w_028_273, w_028_274, w_028_275, w_028_276, w_028_277, w_028_278, w_028_279, w_028_280, w_028_281, w_028_282, w_028_283, w_028_284, w_028_285, w_028_286, w_028_287, w_028_288, w_028_289, w_028_290, w_028_291, w_028_292, w_028_293, w_028_294, w_028_295, w_028_296, w_028_297, w_028_298, w_028_299, w_028_300, w_028_301, w_028_302, w_028_303, w_028_304, w_028_305, w_028_306, w_028_307, w_028_308, w_028_309, w_028_310, w_028_311, w_028_312, w_028_313, w_028_314, w_028_315, w_028_316, w_028_317, w_028_318, w_028_319, w_028_320, w_028_321, w_028_322, w_028_323, w_028_324, w_028_325, w_028_326, w_028_327, w_028_328, w_028_329, w_028_330, w_028_331, w_028_332, w_028_333, w_028_334, w_028_335, w_028_336, w_028_337, w_028_338, w_028_339, w_028_340, w_028_341, w_028_342, w_028_343, w_028_344, w_028_345, w_028_346, w_028_347, w_028_348, w_028_349, w_028_350, w_028_351, w_028_352, w_028_353, w_028_354, w_028_355, w_028_356, w_028_357, w_028_358, w_028_359, w_028_360, w_028_361, w_028_362, w_028_363, w_028_364, w_028_365, w_028_366, w_028_367, w_028_368, w_028_369, w_028_370, w_028_371, w_028_372, w_028_373, w_028_374, w_028_375, w_028_376, w_028_377, w_028_378, w_028_379, w_028_380, w_028_381, w_028_382, w_028_383, w_028_384, w_028_385, w_028_386, w_028_387, w_028_388, w_028_389, w_028_390, w_028_391, w_028_392, w_028_393, w_028_394, w_028_395, w_028_396, w_028_397, w_028_398, w_028_399, w_028_400, w_028_401, w_028_402, w_028_403, w_028_404, w_028_405, w_028_406, w_028_407, w_028_408, w_028_409, w_028_410, w_028_411, w_028_412, w_028_413, w_028_414, w_028_415, w_028_416, w_028_417, w_028_418, w_028_419, w_028_420, w_028_421, w_028_422, w_028_423, w_028_424, w_028_425, w_028_426, w_028_427, w_028_428, w_028_429, w_028_430, w_028_431, w_028_432, w_028_433, w_028_434, w_028_435, w_028_436, w_028_437, w_028_438, w_028_439, w_028_440, w_028_441, w_028_442, w_028_443, w_028_444, w_028_445, w_028_446, w_028_447, w_028_448, w_028_449, w_028_450, w_028_451, w_028_452, w_028_453, w_028_454, w_028_455, w_028_456, w_028_457, w_028_458, w_028_459, w_028_460, w_028_461, w_028_462, w_028_463, w_028_464, w_028_465, w_028_466, w_028_467, w_028_468, w_028_469, w_028_470, w_028_471, w_028_472, w_028_473, w_028_474, w_028_475, w_028_476, w_028_477, w_028_478, w_028_479, w_028_480, w_028_481, w_028_482, w_028_483, w_028_484, w_028_485, w_028_486, w_028_487, w_028_488, w_028_489, w_028_490, w_028_491, w_028_492, w_028_493, w_028_494, w_028_495, w_028_496, w_028_497, w_028_498, w_028_499, w_028_500, w_028_501, w_028_502, w_028_503, w_028_504, w_028_505, w_028_506, w_028_507, w_028_508, w_028_509, w_028_510, w_028_511, w_028_512, w_028_513, w_028_514, w_028_515, w_028_516, w_028_517, w_028_518, w_028_519, w_028_520, w_028_521, w_028_522, w_028_523, w_028_524, w_028_525, w_028_526, w_028_527, w_028_528, w_028_529, w_028_530, w_028_531, w_028_532, w_028_533, w_028_534, w_028_535, w_028_536, w_028_537, w_028_538, w_028_539, w_028_540, w_028_541, w_028_542, w_028_543, w_028_544, w_028_545, w_028_546, w_028_547, w_028_548, w_028_549, w_028_550, w_028_551, w_028_552, w_028_553, w_028_554, w_028_555, w_028_556, w_028_557, w_028_558, w_028_559, w_028_560, w_028_561, w_028_562, w_028_563, w_028_564, w_028_565, w_028_566, w_028_567, w_028_568, w_028_569, w_028_570, w_028_571, w_028_572, w_028_573, w_028_574, w_028_575, w_028_576, w_028_577, w_028_578, w_028_579, w_028_580, w_028_581, w_028_582, w_028_583, w_028_584, w_028_585, w_028_586, w_028_587, w_028_588, w_028_589, w_028_590, w_028_591, w_028_592, w_028_593, w_028_594, w_028_595, w_028_596, w_028_597, w_028_598, w_028_599, w_028_600, w_028_601, w_028_602, w_028_603, w_028_604, w_028_605, w_028_606, w_028_607, w_028_608, w_028_609, w_028_610, w_028_611, w_028_612, w_028_613, w_028_614, w_028_615, w_028_616, w_028_617, w_028_618, w_028_619, w_028_620, w_028_621, w_028_622, w_028_623, w_028_624, w_028_625, w_028_626, w_028_627, w_028_628, w_028_629, w_028_630, w_028_631, w_028_632, w_028_633, w_028_634, w_028_635, w_028_636, w_028_637, w_028_638, w_028_639, w_028_640, w_028_641, w_028_642, w_028_643, w_028_644, w_028_645, w_028_646, w_028_647, w_028_648, w_028_649, w_028_650, w_028_651, w_028_652, w_028_653, w_028_654, w_028_655, w_028_656, w_028_657, w_028_658, w_028_659, w_028_660, w_028_661, w_028_662, w_028_663, w_028_664, w_028_665, w_028_666, w_028_667, w_028_668, w_028_669, w_028_670, w_028_671, w_028_672, w_028_673, w_028_674, w_028_675, w_028_676, w_028_677, w_028_678, w_028_679, w_028_680, w_028_681, w_028_682, w_028_683, w_028_684, w_028_685, w_028_686, w_028_687, w_028_688;
  wire w_029_000, w_029_001, w_029_002, w_029_003, w_029_004, w_029_005, w_029_006, w_029_007, w_029_008, w_029_009, w_029_010, w_029_011, w_029_012, w_029_013, w_029_014, w_029_015, w_029_016, w_029_017, w_029_018, w_029_019, w_029_020, w_029_021, w_029_022, w_029_023, w_029_024, w_029_025, w_029_026, w_029_027, w_029_028, w_029_029, w_029_030, w_029_031, w_029_032, w_029_033, w_029_034, w_029_035, w_029_036, w_029_037, w_029_038, w_029_039, w_029_040, w_029_041, w_029_042, w_029_043, w_029_044, w_029_045, w_029_046, w_029_047, w_029_048, w_029_049, w_029_050, w_029_051, w_029_052, w_029_053, w_029_054, w_029_055, w_029_056, w_029_057, w_029_058, w_029_059, w_029_060, w_029_061, w_029_062, w_029_063, w_029_064, w_029_065, w_029_066, w_029_067, w_029_068, w_029_069, w_029_070, w_029_071, w_029_072, w_029_073, w_029_074, w_029_075, w_029_076, w_029_077, w_029_078, w_029_079, w_029_080, w_029_081, w_029_082, w_029_083, w_029_084, w_029_085, w_029_086, w_029_087, w_029_088, w_029_089, w_029_090, w_029_091, w_029_092, w_029_093, w_029_094, w_029_095, w_029_096, w_029_097, w_029_098, w_029_099, w_029_100, w_029_101, w_029_102, w_029_103, w_029_104, w_029_105, w_029_106, w_029_107, w_029_108, w_029_109, w_029_110, w_029_111, w_029_112, w_029_113, w_029_114, w_029_115, w_029_116, w_029_117, w_029_118, w_029_119, w_029_120, w_029_121, w_029_122, w_029_123, w_029_124, w_029_125, w_029_126, w_029_127, w_029_128, w_029_129, w_029_130, w_029_131, w_029_132, w_029_133, w_029_134, w_029_135, w_029_136, w_029_137, w_029_138, w_029_139, w_029_140, w_029_141, w_029_142, w_029_143, w_029_144, w_029_145, w_029_146, w_029_147, w_029_148, w_029_149, w_029_150, w_029_151, w_029_152, w_029_153, w_029_154, w_029_155, w_029_156, w_029_157, w_029_158, w_029_159, w_029_160, w_029_161, w_029_162, w_029_163, w_029_164, w_029_165, w_029_166, w_029_167, w_029_168, w_029_169, w_029_170, w_029_171, w_029_172, w_029_173, w_029_174, w_029_175, w_029_176, w_029_177, w_029_178, w_029_179, w_029_180, w_029_181, w_029_182, w_029_183, w_029_184, w_029_185, w_029_186, w_029_187, w_029_188, w_029_189, w_029_190, w_029_191, w_029_192, w_029_193, w_029_194, w_029_195, w_029_196, w_029_197, w_029_198, w_029_199, w_029_200, w_029_201, w_029_202, w_029_203, w_029_204, w_029_205, w_029_206, w_029_207, w_029_208, w_029_209, w_029_210, w_029_211, w_029_212, w_029_213, w_029_214, w_029_215, w_029_216, w_029_217, w_029_218, w_029_219, w_029_220, w_029_221, w_029_222, w_029_223, w_029_224, w_029_225, w_029_226, w_029_227, w_029_228, w_029_229, w_029_230, w_029_231, w_029_232, w_029_233, w_029_234, w_029_235, w_029_236, w_029_237, w_029_238, w_029_239, w_029_240, w_029_241, w_029_242, w_029_243, w_029_244, w_029_245, w_029_246, w_029_247, w_029_248, w_029_249, w_029_250, w_029_251, w_029_252, w_029_253, w_029_254, w_029_255, w_029_256, w_029_257, w_029_258, w_029_259, w_029_260, w_029_261, w_029_262, w_029_263, w_029_264, w_029_265, w_029_266, w_029_267, w_029_268, w_029_269, w_029_270, w_029_271, w_029_272, w_029_273, w_029_274, w_029_275, w_029_276, w_029_277, w_029_278, w_029_279, w_029_280, w_029_281, w_029_282, w_029_283, w_029_284, w_029_285, w_029_286, w_029_287, w_029_288, w_029_289, w_029_290, w_029_291, w_029_292, w_029_293, w_029_294, w_029_295, w_029_296, w_029_297, w_029_298, w_029_299, w_029_300, w_029_301, w_029_302, w_029_303, w_029_304, w_029_305, w_029_306, w_029_307, w_029_308, w_029_309, w_029_310, w_029_311, w_029_312, w_029_313, w_029_314, w_029_315, w_029_316, w_029_317, w_029_318, w_029_319, w_029_320, w_029_321, w_029_322, w_029_323, w_029_324, w_029_325, w_029_326, w_029_327, w_029_328, w_029_329, w_029_330, w_029_331, w_029_332, w_029_333, w_029_334, w_029_335, w_029_336, w_029_337, w_029_338, w_029_339, w_029_340, w_029_341, w_029_342, w_029_343, w_029_344, w_029_345, w_029_346, w_029_347, w_029_348, w_029_349, w_029_350, w_029_351, w_029_352, w_029_353, w_029_354, w_029_355, w_029_356, w_029_357, w_029_358, w_029_359, w_029_360, w_029_361, w_029_362, w_029_363, w_029_364, w_029_365, w_029_366, w_029_367, w_029_368, w_029_369, w_029_370, w_029_371, w_029_372, w_029_373, w_029_374, w_029_375, w_029_376, w_029_377, w_029_378, w_029_379, w_029_380, w_029_381, w_029_382, w_029_383, w_029_384, w_029_385, w_029_386, w_029_387, w_029_388, w_029_389, w_029_390, w_029_391, w_029_392, w_029_393, w_029_394, w_029_395, w_029_396, w_029_397, w_029_398, w_029_399, w_029_400, w_029_401, w_029_402, w_029_403, w_029_404, w_029_405, w_029_406, w_029_407, w_029_408, w_029_409, w_029_410, w_029_411, w_029_412, w_029_413, w_029_414, w_029_415, w_029_416, w_029_417, w_029_418, w_029_419, w_029_420, w_029_421, w_029_422, w_029_423, w_029_424, w_029_425, w_029_426, w_029_427, w_029_428, w_029_429, w_029_430, w_029_431, w_029_432, w_029_433, w_029_434, w_029_435, w_029_436, w_029_437, w_029_438, w_029_439, w_029_440, w_029_441, w_029_442, w_029_443, w_029_444, w_029_445, w_029_446, w_029_447, w_029_448, w_029_449, w_029_450, w_029_451, w_029_452, w_029_453, w_029_454, w_029_455, w_029_456, w_029_457, w_029_458, w_029_459, w_029_460, w_029_461, w_029_462, w_029_463, w_029_464, w_029_465, w_029_466, w_029_467, w_029_468, w_029_469, w_029_470, w_029_471, w_029_472, w_029_473, w_029_474, w_029_475, w_029_476, w_029_477, w_029_478, w_029_479, w_029_480, w_029_481, w_029_482, w_029_483, w_029_484, w_029_485, w_029_486, w_029_487, w_029_488, w_029_489, w_029_490, w_029_491, w_029_492, w_029_493, w_029_494, w_029_495, w_029_496, w_029_497, w_029_498, w_029_499, w_029_500, w_029_501, w_029_502, w_029_503, w_029_504, w_029_505, w_029_506, w_029_507, w_029_508, w_029_509, w_029_510, w_029_511, w_029_512, w_029_513, w_029_514, w_029_515, w_029_516, w_029_517, w_029_518, w_029_519, w_029_520, w_029_521, w_029_522, w_029_523, w_029_524, w_029_525, w_029_526, w_029_527, w_029_528, w_029_529, w_029_530, w_029_531, w_029_532, w_029_533, w_029_534, w_029_535, w_029_536, w_029_537, w_029_538, w_029_539, w_029_540, w_029_541, w_029_542, w_029_543, w_029_544, w_029_545, w_029_546, w_029_547, w_029_548, w_029_549, w_029_550, w_029_551, w_029_552, w_029_553, w_029_554, w_029_555, w_029_556, w_029_557, w_029_558, w_029_559, w_029_560, w_029_561, w_029_562, w_029_563, w_029_564, w_029_565, w_029_566, w_029_567, w_029_568, w_029_569, w_029_570, w_029_571, w_029_572, w_029_573, w_029_574, w_029_575, w_029_576, w_029_577, w_029_578, w_029_579, w_029_580, w_029_581, w_029_582, w_029_583, w_029_584, w_029_585, w_029_586, w_029_587;
  wire w_030_000, w_030_001, w_030_002, w_030_003, w_030_004, w_030_005, w_030_006, w_030_007, w_030_008, w_030_009, w_030_010, w_030_011, w_030_012, w_030_013, w_030_014, w_030_015, w_030_016, w_030_017, w_030_018, w_030_019, w_030_020, w_030_021, w_030_022, w_030_023, w_030_024, w_030_025, w_030_026, w_030_027, w_030_028, w_030_029, w_030_030, w_030_031, w_030_032, w_030_033, w_030_034, w_030_035, w_030_036, w_030_037, w_030_038, w_030_039, w_030_040, w_030_041, w_030_042, w_030_043, w_030_044, w_030_045, w_030_046, w_030_047, w_030_048, w_030_049, w_030_050, w_030_051, w_030_052, w_030_053, w_030_054, w_030_055, w_030_056, w_030_057, w_030_058, w_030_059, w_030_060, w_030_061, w_030_062, w_030_063, w_030_064, w_030_065, w_030_066, w_030_067, w_030_068, w_030_069, w_030_070, w_030_071, w_030_072, w_030_073, w_030_074, w_030_075, w_030_076, w_030_077, w_030_078, w_030_079, w_030_080, w_030_081, w_030_082, w_030_083, w_030_084, w_030_085, w_030_086, w_030_087, w_030_088, w_030_089, w_030_090, w_030_091, w_030_092, w_030_093, w_030_094, w_030_095, w_030_096, w_030_097, w_030_098, w_030_099, w_030_100, w_030_101, w_030_102, w_030_103, w_030_104, w_030_105, w_030_106, w_030_107, w_030_108, w_030_109, w_030_110, w_030_111, w_030_112, w_030_113, w_030_114, w_030_115, w_030_116, w_030_117, w_030_118, w_030_119, w_030_120, w_030_121, w_030_122, w_030_123, w_030_124, w_030_125, w_030_126, w_030_127, w_030_128, w_030_129, w_030_130, w_030_131, w_030_132, w_030_133, w_030_134, w_030_135, w_030_136, w_030_137, w_030_138, w_030_139, w_030_140, w_030_141, w_030_142, w_030_143, w_030_144, w_030_145, w_030_146, w_030_147, w_030_148, w_030_149, w_030_150, w_030_151, w_030_152, w_030_153, w_030_154, w_030_155, w_030_156, w_030_157, w_030_158, w_030_159, w_030_160, w_030_161, w_030_162, w_030_163, w_030_164, w_030_165, w_030_166, w_030_167, w_030_168, w_030_169, w_030_170, w_030_171, w_030_172, w_030_173, w_030_174, w_030_175, w_030_176, w_030_177, w_030_178, w_030_179, w_030_180, w_030_181, w_030_182, w_030_183, w_030_184, w_030_185, w_030_186, w_030_187, w_030_188, w_030_189, w_030_190, w_030_191, w_030_192, w_030_193, w_030_194, w_030_195, w_030_196, w_030_197, w_030_198, w_030_199, w_030_200, w_030_201, w_030_202, w_030_203, w_030_204, w_030_205, w_030_206, w_030_207, w_030_208, w_030_209, w_030_210, w_030_211, w_030_212, w_030_213, w_030_214, w_030_215, w_030_216, w_030_217, w_030_218, w_030_219, w_030_220, w_030_221, w_030_222, w_030_223, w_030_224, w_030_225, w_030_226, w_030_227, w_030_228, w_030_229, w_030_230, w_030_231, w_030_232, w_030_233, w_030_234, w_030_235, w_030_236, w_030_237, w_030_238, w_030_239, w_030_240, w_030_241, w_030_242, w_030_243, w_030_244, w_030_245, w_030_246, w_030_247, w_030_248, w_030_249, w_030_250, w_030_251, w_030_252, w_030_253, w_030_254, w_030_255, w_030_256, w_030_257, w_030_258, w_030_259, w_030_260, w_030_261, w_030_262, w_030_263, w_030_264, w_030_265, w_030_266, w_030_267, w_030_268, w_030_269, w_030_270, w_030_271, w_030_272, w_030_273, w_030_274, w_030_275, w_030_276, w_030_277, w_030_278, w_030_279, w_030_280, w_030_281, w_030_282, w_030_283, w_030_284, w_030_285, w_030_286, w_030_287, w_030_288, w_030_289, w_030_290, w_030_291, w_030_292, w_030_293, w_030_294, w_030_295, w_030_296, w_030_297, w_030_298, w_030_299, w_030_300, w_030_301, w_030_302, w_030_303, w_030_304, w_030_305, w_030_306, w_030_307, w_030_308, w_030_309, w_030_310, w_030_311, w_030_312, w_030_313, w_030_314, w_030_315, w_030_316, w_030_317, w_030_318, w_030_319, w_030_320, w_030_321, w_030_322, w_030_323, w_030_324, w_030_325, w_030_326, w_030_327, w_030_328, w_030_329, w_030_330, w_030_331, w_030_332, w_030_333, w_030_334, w_030_335, w_030_336, w_030_337, w_030_338, w_030_339, w_030_340, w_030_341, w_030_342, w_030_343, w_030_344, w_030_345, w_030_346, w_030_347, w_030_348, w_030_349, w_030_350, w_030_351, w_030_352, w_030_353, w_030_354, w_030_355, w_030_356, w_030_357, w_030_358, w_030_359, w_030_360, w_030_361, w_030_362, w_030_363, w_030_364, w_030_365, w_030_366, w_030_367, w_030_368, w_030_369, w_030_370, w_030_371, w_030_372, w_030_373, w_030_374, w_030_375, w_030_376, w_030_377, w_030_378, w_030_379, w_030_380, w_030_381, w_030_382, w_030_383, w_030_384, w_030_385, w_030_386, w_030_387, w_030_388, w_030_389, w_030_390, w_030_391, w_030_392, w_030_393, w_030_394, w_030_395, w_030_396, w_030_397, w_030_398, w_030_399, w_030_400, w_030_401, w_030_402, w_030_403, w_030_404, w_030_405, w_030_406, w_030_407, w_030_408, w_030_409, w_030_410, w_030_411, w_030_412, w_030_413, w_030_414, w_030_415, w_030_416, w_030_417, w_030_418, w_030_419, w_030_420, w_030_421, w_030_422, w_030_423, w_030_424, w_030_425, w_030_426, w_030_427, w_030_428, w_030_429, w_030_430, w_030_431, w_030_432, w_030_433, w_030_434, w_030_435, w_030_436, w_030_437, w_030_438, w_030_439, w_030_440, w_030_441, w_030_442, w_030_443, w_030_444, w_030_445, w_030_446, w_030_447, w_030_448, w_030_449, w_030_450, w_030_451, w_030_452, w_030_453, w_030_454, w_030_455, w_030_456, w_030_457, w_030_458, w_030_459, w_030_460, w_030_461, w_030_462, w_030_463, w_030_464, w_030_465, w_030_466, w_030_467, w_030_468, w_030_469, w_030_470, w_030_471, w_030_472, w_030_473, w_030_474, w_030_475, w_030_476, w_030_477, w_030_478, w_030_479, w_030_480, w_030_481, w_030_482, w_030_483, w_030_484, w_030_485, w_030_486, w_030_487, w_030_488, w_030_489, w_030_490, w_030_491, w_030_492, w_030_493, w_030_494, w_030_495, w_030_496, w_030_497, w_030_498, w_030_499, w_030_500, w_030_501, w_030_502, w_030_503, w_030_504, w_030_505, w_030_506, w_030_507, w_030_508, w_030_509, w_030_510, w_030_511, w_030_512, w_030_513, w_030_514, w_030_515, w_030_516, w_030_517, w_030_518, w_030_519, w_030_520, w_030_521, w_030_522, w_030_523, w_030_524, w_030_525, w_030_526, w_030_527, w_030_528, w_030_529, w_030_530, w_030_531, w_030_532, w_030_533, w_030_534, w_030_535, w_030_536, w_030_537, w_030_538, w_030_539, w_030_540, w_030_541, w_030_542, w_030_543, w_030_544, w_030_545, w_030_546, w_030_547, w_030_548, w_030_549, w_030_550, w_030_551, w_030_552, w_030_553, w_030_554, w_030_555, w_030_556;
  wire w_031_000, w_031_001, w_031_002, w_031_004, w_031_005, w_031_006, w_031_007, w_031_009, w_031_010, w_031_011, w_031_012, w_031_013, w_031_014, w_031_015, w_031_016, w_031_017, w_031_018, w_031_020, w_031_021, w_031_022, w_031_023, w_031_024, w_031_026, w_031_027, w_031_028, w_031_029, w_031_030, w_031_032, w_031_033, w_031_037, w_031_038, w_031_039, w_031_041, w_031_042, w_031_043, w_031_044, w_031_045, w_031_046, w_031_048, w_031_050, w_031_051, w_031_052, w_031_053, w_031_054, w_031_056, w_031_057, w_031_058, w_031_059, w_031_060, w_031_062, w_031_063, w_031_065, w_031_069, w_031_070, w_031_071, w_031_072, w_031_073, w_031_074, w_031_076, w_031_077, w_031_078, w_031_079, w_031_081, w_031_082, w_031_083, w_031_084, w_031_085, w_031_089, w_031_090, w_031_091, w_031_092, w_031_093, w_031_094, w_031_095, w_031_096, w_031_098, w_031_099, w_031_100, w_031_102, w_031_104, w_031_106, w_031_107, w_031_108, w_031_109, w_031_110, w_031_111, w_031_112, w_031_114, w_031_115, w_031_116, w_031_118, w_031_119, w_031_120, w_031_121, w_031_122, w_031_123, w_031_124, w_031_125, w_031_126, w_031_129, w_031_130, w_031_131, w_031_132, w_031_133, w_031_134, w_031_135, w_031_137, w_031_138, w_031_141, w_031_142, w_031_143, w_031_144, w_031_145, w_031_146, w_031_147, w_031_148, w_031_150, w_031_151, w_031_152, w_031_153, w_031_154, w_031_156, w_031_157, w_031_158, w_031_159, w_031_160, w_031_162, w_031_163, w_031_164, w_031_167, w_031_168, w_031_169, w_031_170, w_031_171, w_031_172, w_031_173, w_031_174, w_031_175, w_031_176, w_031_177, w_031_178, w_031_179, w_031_180, w_031_181, w_031_182, w_031_183, w_031_184, w_031_185, w_031_186, w_031_187, w_031_188, w_031_189, w_031_190, w_031_191, w_031_192, w_031_193, w_031_194, w_031_195, w_031_196, w_031_197, w_031_198, w_031_199, w_031_200, w_031_201, w_031_203, w_031_204, w_031_205, w_031_206, w_031_207, w_031_209, w_031_210, w_031_212, w_031_213, w_031_214, w_031_215, w_031_216, w_031_217, w_031_218, w_031_219, w_031_220, w_031_221, w_031_222, w_031_223, w_031_224, w_031_229, w_031_230, w_031_232, w_031_234, w_031_235, w_031_236, w_031_238, w_031_239, w_031_240, w_031_241, w_031_242, w_031_244, w_031_245, w_031_246, w_031_249, w_031_250, w_031_251, w_031_252, w_031_253, w_031_256, w_031_258, w_031_260, w_031_261, w_031_262, w_031_263, w_031_264, w_031_265, w_031_268, w_031_269, w_031_271, w_031_272, w_031_274, w_031_275, w_031_276, w_031_277, w_031_278, w_031_279, w_031_280, w_031_281, w_031_283, w_031_284, w_031_286, w_031_287, w_031_288, w_031_289, w_031_291, w_031_292, w_031_293, w_031_294, w_031_295, w_031_296, w_031_297, w_031_299, w_031_300, w_031_302, w_031_304, w_031_306, w_031_307, w_031_308, w_031_309, w_031_310, w_031_311, w_031_312, w_031_313, w_031_314, w_031_315, w_031_316, w_031_317, w_031_318, w_031_320, w_031_321, w_031_322, w_031_323, w_031_325, w_031_327, w_031_329, w_031_330, w_031_333, w_031_334, w_031_335, w_031_336, w_031_338, w_031_339, w_031_340, w_031_342, w_031_344, w_031_345, w_031_347, w_031_348, w_031_349, w_031_351, w_031_352, w_031_353, w_031_354, w_031_355, w_031_356, w_031_357, w_031_359, w_031_360, w_031_361, w_031_362, w_031_363, w_031_364, w_031_366, w_031_367, w_031_368, w_031_369, w_031_370, w_031_371, w_031_372, w_031_373, w_031_374, w_031_375, w_031_377, w_031_378, w_031_379, w_031_380, w_031_381, w_031_382, w_031_383, w_031_384, w_031_385, w_031_386, w_031_387, w_031_389, w_031_391, w_031_392, w_031_393, w_031_394, w_031_395, w_031_397, w_031_398, w_031_400, w_031_401, w_031_402, w_031_403, w_031_404, w_031_406, w_031_407, w_031_408, w_031_410, w_031_411, w_031_414, w_031_415, w_031_416, w_031_417, w_031_418, w_031_419, w_031_421, w_031_422, w_031_424, w_031_426, w_031_427, w_031_428, w_031_429, w_031_430, w_031_432, w_031_433, w_031_434, w_031_435, w_031_436, w_031_437, w_031_438, w_031_439, w_031_440, w_031_442, w_031_443, w_031_444, w_031_445, w_031_446, w_031_447, w_031_448, w_031_449, w_031_450, w_031_451, w_031_452, w_031_453, w_031_454, w_031_455, w_031_456, w_031_457, w_031_458, w_031_461, w_031_462, w_031_463, w_031_464, w_031_465, w_031_466, w_031_468, w_031_469, w_031_470, w_031_471, w_031_472, w_031_473, w_031_476, w_031_477, w_031_478, w_031_479, w_031_481, w_031_482, w_031_483, w_031_484, w_031_485, w_031_486, w_031_488, w_031_491, w_031_493, w_031_495, w_031_496, w_031_497, w_031_498, w_031_499, w_031_500, w_031_501, w_031_502, w_031_504, w_031_505, w_031_506, w_031_507, w_031_508, w_031_509, w_031_510, w_031_511, w_031_515, w_031_516, w_031_517, w_031_518, w_031_519, w_031_520, w_031_521, w_031_522, w_031_523, w_031_525, w_031_526, w_031_527, w_031_528, w_031_529, w_031_530, w_031_531, w_031_532, w_031_533, w_031_534, w_031_535, w_031_536, w_031_538, w_031_539, w_031_540, w_031_541, w_031_542, w_031_543, w_031_545, w_031_546, w_031_547, w_031_548, w_031_549, w_031_550, w_031_551, w_031_552, w_031_553, w_031_554, w_031_555, w_031_556, w_031_558, w_031_559, w_031_560, w_031_561, w_031_562, w_031_563, w_031_564, w_031_565, w_031_566, w_031_567, w_031_568, w_031_569, w_031_570, w_031_571, w_031_572, w_031_573, w_031_574, w_031_575, w_031_577, w_031_578, w_031_579, w_031_580, w_031_584, w_031_585, w_031_586, w_031_587, w_031_588, w_031_589, w_031_590, w_031_591, w_031_592, w_031_593, w_031_595, w_031_596, w_031_597, w_031_598, w_031_599, w_031_600, w_031_601, w_031_605, w_031_606, w_031_609, w_031_610, w_031_613, w_031_615, w_031_617, w_031_618, w_031_619, w_031_620, w_031_621, w_031_622, w_031_624, w_031_625, w_031_626, w_031_627, w_031_629, w_031_630, w_031_632, w_031_635, w_031_636, w_031_637, w_031_638, w_031_639, w_031_640, w_031_642, w_031_643, w_031_645, w_031_647, w_031_649, w_031_650, w_031_653, w_031_654, w_031_655, w_031_656, w_031_657, w_031_658, w_031_659, w_031_660, w_031_661, w_031_662, w_031_664, w_031_665, w_031_666, w_031_667, w_031_669, w_031_670, w_031_671, w_031_672, w_031_673, w_031_674, w_031_675, w_031_676, w_031_677, w_031_679, w_031_680, w_031_681, w_031_683, w_031_686, w_031_687, w_031_688, w_031_689, w_031_690, w_031_691, w_031_692, w_031_693, w_031_694, w_031_695, w_031_697, w_031_698, w_031_699, w_031_700, w_031_701, w_031_702, w_031_704, w_031_705, w_031_708, w_031_709, w_031_710, w_031_711, w_031_712, w_031_714, w_031_715, w_031_717, w_031_718, w_031_719, w_031_720, w_031_721, w_031_722, w_031_723, w_031_724, w_031_725, w_031_726, w_031_727, w_031_728, w_031_729, w_031_730, w_031_731, w_031_732, w_031_734, w_031_736, w_031_737, w_031_738, w_031_739, w_031_740, w_031_741, w_031_742, w_031_743, w_031_744, w_031_745, w_031_746, w_031_747, w_031_748, w_031_749, w_031_750, w_031_751, w_031_752, w_031_753, w_031_754, w_031_755, w_031_757, w_031_759, w_031_761, w_031_763, w_031_764, w_031_766, w_031_768, w_031_769, w_031_770, w_031_771, w_031_773, w_031_774, w_031_775, w_031_776, w_031_777, w_031_778, w_031_780, w_031_781, w_031_782, w_031_783, w_031_784, w_031_785, w_031_786, w_031_788, w_031_789, w_031_791, w_031_792, w_031_793, w_031_794, w_031_795, w_031_796, w_031_797, w_031_799, w_031_800, w_031_801, w_031_802, w_031_803, w_031_804, w_031_805, w_031_806, w_031_807, w_031_808, w_031_809, w_031_810, w_031_811, w_031_812, w_031_815, w_031_816, w_031_817, w_031_818, w_031_819, w_031_821, w_031_822, w_031_823, w_031_824, w_031_825, w_031_826, w_031_829, w_031_830, w_031_831, w_031_832, w_031_833, w_031_834, w_031_836, w_031_837, w_031_838, w_031_839, w_031_840, w_031_842, w_031_843, w_031_845, w_031_846, w_031_847, w_031_849, w_031_850, w_031_851, w_031_852, w_031_853, w_031_854, w_031_855, w_031_856, w_031_857, w_031_858, w_031_859, w_031_860, w_031_862, w_031_863, w_031_864, w_031_866, w_031_867, w_031_869, w_031_870, w_031_871, w_031_872, w_031_873, w_031_875, w_031_877, w_031_878, w_031_879, w_031_880, w_031_882, w_031_883, w_031_884, w_031_885, w_031_886, w_031_887, w_031_888, w_031_889, w_031_890, w_031_891, w_031_893, w_031_894, w_031_896, w_031_897, w_031_898, w_031_900, w_031_902, w_031_903, w_031_905, w_031_906, w_031_907, w_031_909, w_031_911, w_031_913, w_031_914, w_031_915, w_031_917, w_031_919, w_031_920, w_031_921, w_031_922, w_031_923, w_031_924, w_031_926, w_031_928, w_031_929, w_031_931, w_031_932, w_031_934, w_031_935, w_031_936, w_031_937, w_031_938, w_031_939, w_031_940, w_031_942, w_031_943, w_031_944, w_031_946, w_031_947, w_031_949, w_031_950, w_031_951, w_031_953, w_031_954, w_031_955, w_031_956, w_031_957, w_031_958, w_031_959, w_031_960, w_031_962, w_031_963, w_031_964, w_031_965, w_031_966, w_031_967, w_031_968, w_031_969, w_031_970, w_031_971, w_031_972, w_031_973, w_031_974, w_031_975, w_031_976, w_031_977, w_031_979, w_031_980, w_031_981, w_031_982, w_031_984, w_031_985, w_031_986, w_031_987, w_031_988, w_031_989, w_031_990, w_031_991, w_031_992, w_031_993, w_031_996, w_031_998, w_031_1000, w_031_1001, w_031_1002, w_031_1003, w_031_1004, w_031_1005, w_031_1006, w_031_1007, w_031_1008, w_031_1009, w_031_1010, w_031_1012, w_031_1013, w_031_1014, w_031_1015, w_031_1016, w_031_1018, w_031_1019, w_031_1020, w_031_1021, w_031_1022, w_031_1023, w_031_1024, w_031_1025, w_031_1026, w_031_1027, w_031_1028, w_031_1030, w_031_1031, w_031_1032, w_031_1034, w_031_1035, w_031_1036, w_031_1037, w_031_1039, w_031_1040, w_031_1041, w_031_1042, w_031_1044, w_031_1045, w_031_1048, w_031_1049, w_031_1050, w_031_1051, w_031_1052, w_031_1053, w_031_1055, w_031_1056, w_031_1057, w_031_1058, w_031_1059, w_031_1060, w_031_1061, w_031_1063, w_031_1064, w_031_1065, w_031_1066, w_031_1068, w_031_1069, w_031_1072, w_031_1073, w_031_1075, w_031_1076, w_031_1077, w_031_1078, w_031_1080, w_031_1082, w_031_1083, w_031_1084, w_031_1085, w_031_1086, w_031_1088, w_031_1089, w_031_1090, w_031_1091, w_031_1092, w_031_1093, w_031_1096, w_031_1097, w_031_1098, w_031_1099, w_031_1101, w_031_1102, w_031_1103, w_031_1104, w_031_1105, w_031_1106, w_031_1107, w_031_1108, w_031_1109, w_031_1110, w_031_1111, w_031_1112, w_031_1114, w_031_1116, w_031_1117, w_031_1118, w_031_1119, w_031_1120, w_031_1121, w_031_1123, w_031_1124, w_031_1125, w_031_1126, w_031_1127, w_031_1128, w_031_1129, w_031_1130, w_031_1131, w_031_1132, w_031_1133, w_031_1135, w_031_1136, w_031_1137, w_031_1138, w_031_1142, w_031_1143, w_031_1146, w_031_1147, w_031_1148, w_031_1149, w_031_1150, w_031_1152, w_031_1153, w_031_1155, w_031_1158, w_031_1159, w_031_1160, w_031_1162, w_031_1164, w_031_1165, w_031_1166, w_031_1167, w_031_1168, w_031_1170, w_031_1171, w_031_1174, w_031_1175, w_031_1176, w_031_1177, w_031_1178, w_031_1179, w_031_1181, w_031_1182, w_031_1183, w_031_1184, w_031_1185, w_031_1187, w_031_1188, w_031_1189, w_031_1190, w_031_1192, w_031_1193, w_031_1194, w_031_1195, w_031_1196, w_031_1197, w_031_1198, w_031_1199, w_031_1200, w_031_1201, w_031_1202, w_031_1203, w_031_1205, w_031_1206, w_031_1208, w_031_1209, w_031_1210, w_031_1211, w_031_1212, w_031_1213, w_031_1214, w_031_1215, w_031_1216, w_031_1217, w_031_1218, w_031_1219, w_031_1220, w_031_1221, w_031_1222, w_031_1223, w_031_1224, w_031_1225, w_031_1226, w_031_1227, w_031_1228, w_031_1229, w_031_1232, w_031_1233, w_031_1234, w_031_1235, w_031_1236, w_031_1237, w_031_1238, w_031_1239, w_031_1240, w_031_1241, w_031_1242, w_031_1243, w_031_1244, w_031_1245, w_031_1246, w_031_1247, w_031_1248, w_031_1249, w_031_1250, w_031_1251, w_031_1252, w_031_1253, w_031_1254, w_031_1255, w_031_1256, w_031_1258, w_031_1259, w_031_1260, w_031_1261, w_031_1262, w_031_1263, w_031_1264, w_031_1265, w_031_1266, w_031_1267, w_031_1268, w_031_1269, w_031_1270, w_031_1271, w_031_1272, w_031_1274, w_031_1276, w_031_1277, w_031_1278, w_031_1280, w_031_1281, w_031_1283, w_031_1284, w_031_1285, w_031_1286, w_031_1288, w_031_1290, w_031_1291, w_031_1292, w_031_1294, w_031_1295, w_031_1296, w_031_1298, w_031_1299, w_031_1300, w_031_1301, w_031_1302, w_031_1303, w_031_1304, w_031_1305, w_031_1306, w_031_1308, w_031_1309, w_031_1310, w_031_1311, w_031_1312, w_031_1313, w_031_1314, w_031_1316, w_031_1318, w_031_1319, w_031_1320, w_031_1321, w_031_1322, w_031_1323, w_031_1324, w_031_1326, w_031_1327, w_031_1329, w_031_1330, w_031_1331, w_031_1332, w_031_1333, w_031_1334, w_031_1335, w_031_1336, w_031_1337, w_031_1338, w_031_1339, w_031_1340, w_031_1341, w_031_1343, w_031_1344, w_031_1345, w_031_1346, w_031_1347, w_031_1348, w_031_1349, w_031_1350, w_031_1351, w_031_1352, w_031_1355, w_031_1356, w_031_1357, w_031_1359, w_031_1360, w_031_1361, w_031_1363, w_031_1364, w_031_1365, w_031_1366, w_031_1367, w_031_1369, w_031_1370, w_031_1372, w_031_1373, w_031_1374, w_031_1375, w_031_1376, w_031_1378, w_031_1379, w_031_1381, w_031_1382, w_031_1383, w_031_1384, w_031_1386, w_031_1387, w_031_1388, w_031_1389, w_031_1391, w_031_1392, w_031_1393, w_031_1394, w_031_1395, w_031_1396, w_031_1397, w_031_1399, w_031_1401, w_031_1404, w_031_1405, w_031_1406, w_031_1407, w_031_1408, w_031_1409, w_031_1410, w_031_1411, w_031_1412, w_031_1413, w_031_1414, w_031_1416, w_031_1417, w_031_1418, w_031_1419, w_031_1420, w_031_1421, w_031_1422, w_031_1424, w_031_1425, w_031_1427, w_031_1428, w_031_1430, w_031_1431, w_031_1432, w_031_1433, w_031_1434, w_031_1435, w_031_1436, w_031_1437, w_031_1440, w_031_1442, w_031_1443, w_031_1445, w_031_1446, w_031_1447, w_031_1448, w_031_1449, w_031_1450, w_031_1451, w_031_1452, w_031_1453, w_031_1456, w_031_1457, w_031_1458, w_031_1461, w_031_1462, w_031_1463, w_031_1464, w_031_1465, w_031_1466, w_031_1467, w_031_1468, w_031_1470, w_031_1471, w_031_1472, w_031_1473, w_031_1474, w_031_1475, w_031_1476, w_031_1479, w_031_1480, w_031_1481, w_031_1482, w_031_1484, w_031_1486, w_031_1487, w_031_1488, w_031_1490, w_031_1491, w_031_1492, w_031_1494, w_031_1495, w_031_1496, w_031_1499, w_031_1500, w_031_1501, w_031_1502, w_031_1503, w_031_1504, w_031_1505, w_031_1509, w_031_1510, w_031_1511, w_031_1512, w_031_1513, w_031_1514, w_031_1515, w_031_1516, w_031_1517, w_031_1519, w_031_1520, w_031_1521, w_031_1522, w_031_1523, w_031_1524, w_031_1525, w_031_1527, w_031_1528, w_031_1529, w_031_1530, w_031_1531, w_031_1533, w_031_1534, w_031_1535, w_031_1536, w_031_1537, w_031_1538, w_031_1540, w_031_1541, w_031_1543, w_031_1544, w_031_1545, w_031_1546, w_031_1547, w_031_1548, w_031_1550, w_031_1551, w_031_1552, w_031_1553, w_031_1554, w_031_1556, w_031_1557, w_031_1558, w_031_1559, w_031_1560, w_031_1561, w_031_1563, w_031_1564, w_031_1565, w_031_1566, w_031_1567, w_031_1568, w_031_1570, w_031_1571, w_031_1572, w_031_1573, w_031_1575, w_031_1577, w_031_1578, w_031_1579, w_031_1580, w_031_1581, w_031_1582, w_031_1583, w_031_1584, w_031_1585, w_031_1586, w_031_1587, w_031_1589, w_031_1591, w_031_1592, w_031_1594, w_031_1595, w_031_1596, w_031_1597, w_031_1598, w_031_1599, w_031_1600, w_031_1601, w_031_1602, w_031_1603, w_031_1604, w_031_1606, w_031_1607, w_031_1608, w_031_1610, w_031_1611, w_031_1612, w_031_1613, w_031_1614, w_031_1616, w_031_1617, w_031_1618, w_031_1619, w_031_1621, w_031_1622, w_031_1624, w_031_1626, w_031_1627, w_031_1628, w_031_1629, w_031_1630, w_031_1632, w_031_1633, w_031_1634, w_031_1636, w_031_1637, w_031_1639, w_031_1640, w_031_1641, w_031_1642, w_031_1643, w_031_1644, w_031_1645, w_031_1648, w_031_1649, w_031_1650, w_031_1651, w_031_1652, w_031_1653, w_031_1654, w_031_1656, w_031_1657, w_031_1658, w_031_1659, w_031_1660, w_031_1662, w_031_1664, w_031_1665, w_031_1666, w_031_1667, w_031_1670, w_031_1671, w_031_1672, w_031_1673, w_031_1674, w_031_1675, w_031_1677, w_031_1678, w_031_1679, w_031_1680, w_031_1683, w_031_1684, w_031_1685, w_031_1686, w_031_1687, w_031_1688, w_031_1689, w_031_1690, w_031_1691, w_031_1692, w_031_1694, w_031_1695, w_031_1696, w_031_1697, w_031_1698, w_031_1700, w_031_1701, w_031_1704, w_031_1705, w_031_1706, w_031_1708, w_031_1711, w_031_1712, w_031_1713, w_031_1714, w_031_1715, w_031_1717, w_031_1719, w_031_1720, w_031_1721, w_031_1722, w_031_1723, w_031_1725, w_031_1726, w_031_1727, w_031_1728, w_031_1729, w_031_1730, w_031_1731, w_031_1732, w_031_1734, w_031_1735, w_031_1736, w_031_1737, w_031_1738, w_031_1740, w_031_1741, w_031_1742, w_031_1744, w_031_1745, w_031_1747, w_031_1748, w_031_1750, w_031_1751, w_031_1753, w_031_1754, w_031_1755, w_031_1756, w_031_1758, w_031_1759, w_031_1760, w_031_1761, w_031_1762, w_031_1763, w_031_1764, w_031_1766, w_031_1767, w_031_1768, w_031_1769, w_031_1770, w_031_1772, w_031_1773, w_031_1774, w_031_1775, w_031_1776, w_031_1779, w_031_1780, w_031_1781, w_031_1783, w_031_1784, w_031_1785, w_031_1786, w_031_1787, w_031_1788, w_031_1790, w_031_1791, w_031_1794, w_031_1795, w_031_1797, w_031_1798, w_031_1799, w_031_1800, w_031_1801, w_031_1802, w_031_1803, w_031_1804, w_031_1805, w_031_1807, w_031_1809, w_031_1810, w_031_1811, w_031_1812, w_031_1813, w_031_1814, w_031_1815, w_031_1816, w_031_1817, w_031_1818, w_031_1819, w_031_1822, w_031_1824, w_031_1825, w_031_1826, w_031_1828, w_031_1829, w_031_1830, w_031_1831, w_031_1832, w_031_1833, w_031_1834, w_031_1835, w_031_1836, w_031_1839, w_031_1840, w_031_1841, w_031_1842, w_031_1843, w_031_1845, w_031_1847, w_031_1848, w_031_1850, w_031_1851, w_031_1853, w_031_1854, w_031_1855, w_031_1856, w_031_1857, w_031_1858, w_031_1859, w_031_1860, w_031_1861, w_031_1862, w_031_1863, w_031_1865, w_031_1867, w_031_1868, w_031_1869, w_031_1870, w_031_1871, w_031_1872, w_031_1873, w_031_1874, w_031_1876, w_031_1877, w_031_1878, w_031_1879, w_031_1880, w_031_1881, w_031_1882, w_031_1883, w_031_1884, w_031_1886, w_031_1887, w_031_1888, w_031_1889, w_031_1890, w_031_1891, w_031_1894, w_031_1895, w_031_1899, w_031_1900, w_031_1902, w_031_1904, w_031_1905, w_031_1906, w_031_1907, w_031_1909, w_031_1910, w_031_1911, w_031_1912, w_031_1913, w_031_1914, w_031_1916, w_031_1917, w_031_1918, w_031_1919, w_031_1920, w_031_1921, w_031_1922, w_031_1925, w_031_1926, w_031_1927, w_031_1928, w_031_1929, w_031_1931, w_031_1932, w_031_1933, w_031_1934, w_031_1935, w_031_1936, w_031_1937, w_031_1938, w_031_1939, w_031_1940, w_031_1941, w_031_1942, w_031_1943, w_031_1944, w_031_1946, w_031_1947, w_031_1948, w_031_1949, w_031_1950, w_031_1951, w_031_1952, w_031_1953, w_031_1954, w_031_1955, w_031_1957, w_031_1959, w_031_1961, w_031_1962, w_031_1963, w_031_1965, w_031_1966, w_031_1967, w_031_1968, w_031_1969, w_031_1970, w_031_1971, w_031_1972, w_031_1973, w_031_1976, w_031_1977, w_031_1978, w_031_1979, w_031_1980, w_031_1981, w_031_1982, w_031_1983, w_031_1984, w_031_1985, w_031_1986, w_031_1988, w_031_1989, w_031_1990, w_031_1993, w_031_1994, w_031_1995, w_031_1996, w_031_1997, w_031_1998, w_031_1999, w_031_2000, w_031_2001, w_031_2002, w_031_2003, w_031_2004, w_031_2005, w_031_2007, w_031_2008, w_031_2009, w_031_2010, w_031_2011, w_031_2012, w_031_2014, w_031_2015, w_031_2016, w_031_2017, w_031_2019, w_031_2020, w_031_2021, w_031_2024, w_031_2025, w_031_2026, w_031_2027, w_031_2028, w_031_2029, w_031_2030, w_031_2031, w_031_2032, w_031_2033, w_031_2034, w_031_2035, w_031_2036, w_031_2037, w_031_2040, w_031_2041, w_031_2043, w_031_2044, w_031_2045, w_031_2046, w_031_2047, w_031_2048, w_031_2049, w_031_2050, w_031_2051, w_031_2052, w_031_2053, w_031_2054, w_031_2055, w_031_2056, w_031_2057, w_031_2058, w_031_2060, w_031_2061, w_031_2063, w_031_2064, w_031_2065, w_031_2066, w_031_2067, w_031_2068, w_031_2069, w_031_2070, w_031_2074, w_031_2075, w_031_2076, w_031_2077, w_031_2079, w_031_2080, w_031_2082, w_031_2083, w_031_2085, w_031_2086, w_031_2089, w_031_2091, w_031_2094, w_031_2096, w_031_2100, w_031_2101, w_031_2106, w_031_2108, w_031_2109, w_031_2110, w_031_2111, w_031_2114, w_031_2115, w_031_2116, w_031_2119, w_031_2122, w_031_2125, w_031_2126, w_031_2127, w_031_2128, w_031_2129, w_031_2130, w_031_2133, w_031_2137, w_031_2138, w_031_2139, w_031_2140, w_031_2141, w_031_2144, w_031_2146, w_031_2147, w_031_2151, w_031_2153, w_031_2155, w_031_2159, w_031_2160, w_031_2161, w_031_2162, w_031_2163, w_031_2164, w_031_2165, w_031_2166, w_031_2167, w_031_2168, w_031_2172, w_031_2173, w_031_2176, w_031_2179, w_031_2180, w_031_2184, w_031_2185, w_031_2186, w_031_2188, w_031_2189, w_031_2190, w_031_2195, w_031_2197, w_031_2198, w_031_2202, w_031_2203, w_031_2204, w_031_2210, w_031_2212, w_031_2215, w_031_2217, w_031_2218, w_031_2219, w_031_2222, w_031_2225, w_031_2226, w_031_2229, w_031_2230, w_031_2232, w_031_2234, w_031_2238, w_031_2239, w_031_2248, w_031_2253, w_031_2256, w_031_2257, w_031_2258, w_031_2259, w_031_2260, w_031_2263, w_031_2264, w_031_2266, w_031_2267, w_031_2268, w_031_2269, w_031_2270, w_031_2271, w_031_2272, w_031_2273, w_031_2276, w_031_2277, w_031_2278, w_031_2280, w_031_2282, w_031_2285, w_031_2286, w_031_2287, w_031_2288, w_031_2291, w_031_2294, w_031_2295, w_031_2296, w_031_2298, w_031_2299, w_031_2301, w_031_2304, w_031_2305, w_031_2306, w_031_2307, w_031_2309, w_031_2310, w_031_2314, w_031_2315, w_031_2316, w_031_2317, w_031_2318, w_031_2320, w_031_2323, w_031_2325, w_031_2327, w_031_2328, w_031_2330, w_031_2333, w_031_2334, w_031_2339, w_031_2340, w_031_2341, w_031_2342, w_031_2346, w_031_2349, w_031_2350, w_031_2351, w_031_2352, w_031_2354, w_031_2355, w_031_2356, w_031_2357, w_031_2358, w_031_2361, w_031_2364, w_031_2366, w_031_2367, w_031_2368, w_031_2371, w_031_2372, w_031_2373, w_031_2374, w_031_2375, w_031_2376, w_031_2383, w_031_2384, w_031_2385, w_031_2386, w_031_2387, w_031_2388, w_031_2389, w_031_2390, w_031_2392, w_031_2394, w_031_2396, w_031_2397, w_031_2400, w_031_2401, w_031_2402, w_031_2404, w_031_2405, w_031_2406, w_031_2409, w_031_2410, w_031_2412, w_031_2413, w_031_2414, w_031_2416, w_031_2417, w_031_2420, w_031_2421, w_031_2422, w_031_2426, w_031_2427, w_031_2429, w_031_2430, w_031_2431, w_031_2433, w_031_2438, w_031_2441, w_031_2443, w_031_2444, w_031_2445, w_031_2449, w_031_2450, w_031_2451, w_031_2452, w_031_2456, w_031_2458, w_031_2459, w_031_2461, w_031_2462, w_031_2464, w_031_2465, w_031_2466, w_031_2468, w_031_2470, w_031_2472, w_031_2474, w_031_2477, w_031_2481, w_031_2486, w_031_2487, w_031_2488, w_031_2489, w_031_2491, w_031_2492, w_031_2495, w_031_2499, w_031_2504, w_031_2505, w_031_2507, w_031_2508, w_031_2511, w_031_2512, w_031_2513, w_031_2516, w_031_2518, w_031_2519, w_031_2520, w_031_2522, w_031_2523, w_031_2525, w_031_2526, w_031_2531, w_031_2533, w_031_2535, w_031_2538, w_031_2540, w_031_2543, w_031_2544, w_031_2546, w_031_2547, w_031_2548, w_031_2549, w_031_2551, w_031_2555, w_031_2557, w_031_2558, w_031_2561, w_031_2563, w_031_2565, w_031_2568, w_031_2569, w_031_2570, w_031_2571, w_031_2572, w_031_2573, w_031_2574, w_031_2576, w_031_2577, w_031_2578, w_031_2579, w_031_2580, w_031_2581, w_031_2583, w_031_2584, w_031_2589, w_031_2590, w_031_2592, w_031_2593, w_031_2595, w_031_2596, w_031_2597, w_031_2598, w_031_2599, w_031_2602, w_031_2604, w_031_2605, w_031_2606, w_031_2607, w_031_2610, w_031_2611, w_031_2612, w_031_2615, w_031_2617, w_031_2619, w_031_2621, w_031_2623, w_031_2626, w_031_2628, w_031_2630, w_031_2632, w_031_2636, w_031_2639, w_031_2641, w_031_2642, w_031_2644, w_031_2646, w_031_2648, w_031_2649, w_031_2650, w_031_2654, w_031_2655, w_031_2657, w_031_2660, w_031_2661, w_031_2662, w_031_2663, w_031_2664, w_031_2667, w_031_2670, w_031_2671, w_031_2672, w_031_2675, w_031_2676, w_031_2679, w_031_2680, w_031_2686, w_031_2687, w_031_2688, w_031_2690, w_031_2691, w_031_2692, w_031_2693, w_031_2695, w_031_2697, w_031_2699, w_031_2700, w_031_2702, w_031_2703, w_031_2706, w_031_2711, w_031_2712, w_031_2714, w_031_2718, w_031_2719, w_031_2720, w_031_2721, w_031_2722, w_031_2723, w_031_2724, w_031_2726, w_031_2727, w_031_2729, w_031_2730, w_031_2732, w_031_2733, w_031_2734, w_031_2735, w_031_2737, w_031_2739, w_031_2740, w_031_2741, w_031_2742, w_031_2743, w_031_2744, w_031_2745, w_031_2746, w_031_2747, w_031_2748, w_031_2750, w_031_2753, w_031_2755, w_031_2756, w_031_2757, w_031_2761, w_031_2762, w_031_2763, w_031_2765, w_031_2766, w_031_2767, w_031_2769, w_031_2770, w_031_2772, w_031_2773, w_031_2774, w_031_2776, w_031_2777, w_031_2778, w_031_2779, w_031_2780, w_031_2782, w_031_2783, w_031_2784, w_031_2785, w_031_2786, w_031_2789, w_031_2793, w_031_2794, w_031_2798, w_031_2799, w_031_2800, w_031_2802, w_031_2803, w_031_2804, w_031_2805, w_031_2806, w_031_2807, w_031_2808, w_031_2809, w_031_2811, w_031_2814, w_031_2819, w_031_2820, w_031_2822, w_031_2825, w_031_2826, w_031_2827, w_031_2828, w_031_2829, w_031_2831, w_031_2833, w_031_2835, w_031_2837, w_031_2840, w_031_2842, w_031_2845, w_031_2846, w_031_2847, w_031_2849, w_031_2851, w_031_2853, w_031_2856, w_031_2857, w_031_2859, w_031_2860, w_031_2861, w_031_2863, w_031_2864, w_031_2865, w_031_2866, w_031_2867, w_031_2868, w_031_2869, w_031_2871, w_031_2872, w_031_2882, w_031_2887, w_031_2888, w_031_2889, w_031_2896, w_031_2897, w_031_2899, w_031_2900, w_031_2901, w_031_2902, w_031_2903, w_031_2905, w_031_2909, w_031_2910, w_031_2911, w_031_2912, w_031_2913, w_031_2914, w_031_2917, w_031_2918, w_031_2921, w_031_2922, w_031_2923, w_031_2924, w_031_2925, w_031_2927, w_031_2929, w_031_2933, w_031_2934, w_031_2935, w_031_2936, w_031_2937, w_031_2939, w_031_2941, w_031_2946, w_031_2947, w_031_2949, w_031_2952, w_031_2961, w_031_2963, w_031_2964, w_031_2968, w_031_2969, w_031_2971, w_031_2972, w_031_2973, w_031_2979, w_031_2980, w_031_2981, w_031_2983, w_031_2986, w_031_2989, w_031_2990, w_031_2991, w_031_2992, w_031_2993, w_031_2999, w_031_3000, w_031_3001, w_031_3005, w_031_3006, w_031_3007, w_031_3009, w_031_3010, w_031_3011, w_031_3012, w_031_3015, w_031_3016, w_031_3018, w_031_3021, w_031_3023, w_031_3027, w_031_3028, w_031_3030, w_031_3033, w_031_3036, w_031_3037, w_031_3040, w_031_3041, w_031_3047, w_031_3048, w_031_3050, w_031_3051, w_031_3052, w_031_3053, w_031_3058, w_031_3060, w_031_3061, w_031_3062, w_031_3063, w_031_3065, w_031_3069, w_031_3070, w_031_3073, w_031_3074, w_031_3075, w_031_3077, w_031_3082, w_031_3083, w_031_3086, w_031_3087, w_031_3088, w_031_3092, w_031_3095, w_031_3097, w_031_3098, w_031_3102, w_031_3103, w_031_3106, w_031_3108, w_031_3110, w_031_3111, w_031_3114, w_031_3115, w_031_3116, w_031_3117, w_031_3118, w_031_3119, w_031_3120, w_031_3121, w_031_3124, w_031_3125, w_031_3127, w_031_3130, w_031_3132, w_031_3134, w_031_3135, w_031_3137, w_031_3140, w_031_3142, w_031_3146, w_031_3147, w_031_3148, w_031_3149, w_031_3151, w_031_3152, w_031_3157, w_031_3158, w_031_3159, w_031_3163, w_031_3166, w_031_3170, w_031_3171, w_031_3173, w_031_3175, w_031_3177, w_031_3178, w_031_3179, w_031_3180, w_031_3184, w_031_3185, w_031_3186, w_031_3190, w_031_3192, w_031_3193, w_031_3196, w_031_3198, w_031_3199, w_031_3200, w_031_3201, w_031_3204, w_031_3207, w_031_3211, w_031_3214, w_031_3215, w_031_3216, w_031_3217, w_031_3220, w_031_3222, w_031_3223, w_031_3225, w_031_3226, w_031_3229, w_031_3230, w_031_3233, w_031_3235, w_031_3236, w_031_3237, w_031_3238, w_031_3239, w_031_3241, w_031_3242, w_031_3243, w_031_3245, w_031_3246, w_031_3247, w_031_3249, w_031_3250, w_031_3251, w_031_3255, w_031_3260, w_031_3261, w_031_3263, w_031_3264, w_031_3265, w_031_3266, w_031_3267, w_031_3268, w_031_3269, w_031_3273, w_031_3275, w_031_3276, w_031_3278, w_031_3279, w_031_3285, w_031_3286, w_031_3287, w_031_3288, w_031_3289, w_031_3291, w_031_3292, w_031_3293, w_031_3294, w_031_3295, w_031_3297, w_031_3301, w_031_3307, w_031_3308, w_031_3310, w_031_3312, w_031_3313, w_031_3314, w_031_3317, w_031_3318, w_031_3320, w_031_3324, w_031_3325, w_031_3329, w_031_3330, w_031_3331, w_031_3332, w_031_3334, w_031_3336, w_031_3337, w_031_3341, w_031_3345, w_031_3346, w_031_3349, w_031_3350, w_031_3352, w_031_3353, w_031_3357, w_031_3358, w_031_3359, w_031_3362, w_031_3363, w_031_3364, w_031_3366, w_031_3368, w_031_3372, w_031_3373, w_031_3375, w_031_3376, w_031_3377, w_031_3379, w_031_3380, w_031_3381, w_031_3382, w_031_3383, w_031_3385, w_031_3386, w_031_3387, w_031_3388, w_031_3389, w_031_3390, w_031_3391, w_031_3394, w_031_3395, w_031_3397, w_031_3398, w_031_3399, w_031_3401, w_031_3402, w_031_3403, w_031_3404, w_031_3405, w_031_3407, w_031_3408, w_031_3409, w_031_3410, w_031_3411, w_031_3412, w_031_3413, w_031_3414, w_031_3415, w_031_3416, w_031_3417, w_031_3418, w_031_3420, w_031_3423, w_031_3424, w_031_3425, w_031_3426, w_031_3427, w_031_3428, w_031_3432, w_031_3434, w_031_3435, w_031_3436, w_031_3438, w_031_3439, w_031_3441, w_031_3442, w_031_3444, w_031_3447, w_031_3449, w_031_3450, w_031_3456, w_031_3457, w_031_3458, w_031_3459, w_031_3460, w_031_3461, w_031_3462, w_031_3463, w_031_3464, w_031_3465, w_031_3468, w_031_3469, w_031_3470, w_031_3472, w_031_3473, w_031_3476, w_031_3477, w_031_3480, w_031_3484, w_031_3488, w_031_3489, w_031_3490, w_031_3492, w_031_3493, w_031_3495, w_031_3496, w_031_3499, w_031_3500, w_031_3501, w_031_3503, w_031_3504, w_031_3506, w_031_3507, w_031_3508, w_031_3510, w_031_3512, w_031_3514, w_031_3515, w_031_3516, w_031_3518, w_031_3519, w_031_3522, w_031_3523, w_031_3524, w_031_3525, w_031_3526, w_031_3530, w_031_3531, w_031_3532, w_031_3533, w_031_3537, w_031_3538, w_031_3540, w_031_3543, w_031_3547, w_031_3549, w_031_3550, w_031_3551, w_031_3552, w_031_3553, w_031_3555, w_031_3557, w_031_3558, w_031_3559, w_031_3561, w_031_3563, w_031_3565, w_031_3566, w_031_3568, w_031_3571, w_031_3572, w_031_3574, w_031_3577, w_031_3579, w_031_3581, w_031_3583, w_031_3584, w_031_3585, w_031_3590, w_031_3593, w_031_3595, w_031_3596, w_031_3600, w_031_3601, w_031_3602, w_031_3603, w_031_3604, w_031_3605, w_031_3606, w_031_3607, w_031_3608, w_031_3609, w_031_3610, w_031_3613, w_031_3614, w_031_3615, w_031_3617, w_031_3619, w_031_3622, w_031_3624, w_031_3625, w_031_3626, w_031_3629, w_031_3632, w_031_3633, w_031_3635, w_031_3636, w_031_3638, w_031_3645, w_031_3650, w_031_3651, w_031_3653, w_031_3658, w_031_3662, w_031_3663, w_031_3665, w_031_3666, w_031_3667, w_031_3668, w_031_3669, w_031_3674, w_031_3676, w_031_3679, w_031_3680, w_031_3681, w_031_3682, w_031_3683, w_031_3684, w_031_3687, w_031_3688, w_031_3689, w_031_3690, w_031_3695, w_031_3697, w_031_3698, w_031_3700, w_031_3702, w_031_3703, w_031_3704, w_031_3705, w_031_3706, w_031_3708, w_031_3709, w_031_3710, w_031_3712, w_031_3713, w_031_3715, w_031_3720, w_031_3721, w_031_3722, w_031_3723, w_031_3725, w_031_3726, w_031_3727, w_031_3728, w_031_3730, w_031_3733, w_031_3734, w_031_3737, w_031_3738, w_031_3739, w_031_3741, w_031_3744, w_031_3747, w_031_3748, w_031_3750, w_031_3752, w_031_3753, w_031_3754, w_031_3757, w_031_3758, w_031_3759, w_031_3762, w_031_3763, w_031_3765, w_031_3766, w_031_3767, w_031_3768, w_031_3769, w_031_3773, w_031_3774, w_031_3775, w_031_3776, w_031_3777, w_031_3778, w_031_3781, w_031_3782, w_031_3783, w_031_3784, w_031_3785, w_031_3788, w_031_3794, w_031_3798, w_031_3801, w_031_3803, w_031_3804, w_031_3805, w_031_3806, w_031_3807, w_031_3808, w_031_3810, w_031_3811, w_031_3815, w_031_3818, w_031_3820, w_031_3821, w_031_3823, w_031_3826, w_031_3829, w_031_3830, w_031_3832, w_031_3835, w_031_3838, w_031_3839, w_031_3840, w_031_3841, w_031_3843, w_031_3846, w_031_3850, w_031_3851, w_031_3853, w_031_3854, w_031_3857, w_031_3858, w_031_3859, w_031_3861, w_031_3862, w_031_3863, w_031_3865, w_031_3866, w_031_3867, w_031_3869, w_031_3870, w_031_3873, w_031_3875, w_031_3878, w_031_3879, w_031_3883, w_031_3885, w_031_3886, w_031_3891, w_031_3892, w_031_3893, w_031_3895, w_031_3896, w_031_3897, w_031_3900, w_031_3901, w_031_3904, w_031_3907, w_031_3908, w_031_3909, w_031_3910, w_031_3911, w_031_3912, w_031_3914, w_031_3915, w_031_3917, w_031_3918, w_031_3919, w_031_3920, w_031_3927, w_031_3928, w_031_3932, w_031_3933, w_031_3934, w_031_3935, w_031_3936, w_031_3938, w_031_3941, w_031_3943, w_031_3944, w_031_3945, w_031_3947, w_031_3948, w_031_3949, w_031_3953, w_031_3954, w_031_3956, w_031_3957, w_031_3958, w_031_3959, w_031_3962, w_031_3965, w_031_3966, w_031_3967, w_031_3968, w_031_3970, w_031_3973, w_031_3974, w_031_3976, w_031_3979, w_031_3980, w_031_3981, w_031_3982, w_031_3983, w_031_3984, w_031_3985, w_031_3989, w_031_3990, w_031_3991, w_031_3995, w_031_3999, w_031_4002, w_031_4003, w_031_4005, w_031_4006, w_031_4007, w_031_4009, w_031_4010, w_031_4011, w_031_4013, w_031_4016, w_031_4019, w_031_4023, w_031_4026, w_031_4027, w_031_4035, w_031_4036, w_031_4038, w_031_4041, w_031_4044, w_031_4046, w_031_4049, w_031_4050, w_031_4051, w_031_4052, w_031_4054, w_031_4058, w_031_4059, w_031_4061, w_031_4062, w_031_4067, w_031_4070, w_031_4071, w_031_4072, w_031_4074, w_031_4076, w_031_4079, w_031_4081, w_031_4082, w_031_4084, w_031_4085, w_031_4087, w_031_4090, w_031_4092, w_031_4094, w_031_4098, w_031_4107, w_031_4109, w_031_4110, w_031_4111, w_031_4114, w_031_4115, w_031_4117, w_031_4120, w_031_4124, w_031_4126, w_031_4129, w_031_4131, w_031_4132, w_031_4134, w_031_4135, w_031_4137, w_031_4139, w_031_4140, w_031_4141, w_031_4143, w_031_4147, w_031_4152, w_031_4156, w_031_4157, w_031_4158, w_031_4160, w_031_4161, w_031_4162, w_031_4163, w_031_4164, w_031_4165, w_031_4166, w_031_4168, w_031_4171, w_031_4172, w_031_4173, w_031_4174, w_031_4175, w_031_4177, w_031_4178, w_031_4179, w_031_4183, w_031_4188, w_031_4189, w_031_4190, w_031_4191, w_031_4195, w_031_4196, w_031_4199, w_031_4200, w_031_4201, w_031_4203, w_031_4204, w_031_4205, w_031_4206, w_031_4207, w_031_4209, w_031_4213, w_031_4215, w_031_4216, w_031_4218, w_031_4219, w_031_4220, w_031_4221, w_031_4223, w_031_4224, w_031_4225, w_031_4226, w_031_4227, w_031_4229, w_031_4230, w_031_4234, w_031_4236, w_031_4239, w_031_4242, w_031_4243, w_031_4244, w_031_4247, w_031_4248, w_031_4249, w_031_4251, w_031_4255, w_031_4256, w_031_4257, w_031_4260, w_031_4261, w_031_4263, w_031_4265, w_031_4267, w_031_4269, w_031_4271, w_031_4272, w_031_4273, w_031_4275, w_031_4276, w_031_4280, w_031_4281, w_031_4284, w_031_4285, w_031_4286, w_031_4287, w_031_4288, w_031_4291, w_031_4292, w_031_4293, w_031_4294, w_031_4295, w_031_4296, w_031_4297, w_031_4298, w_031_4299, w_031_4301, w_031_4302, w_031_4305, w_031_4307, w_031_4308, w_031_4309, w_031_4315, w_031_4316, w_031_4317, w_031_4318, w_031_4319, w_031_4320, w_031_4321, w_031_4323, w_031_4326, w_031_4329, w_031_4332, w_031_4333, w_031_4334, w_031_4335, w_031_4336, w_031_4338, w_031_4346, w_031_4349, w_031_4350, w_031_4352, w_031_4353, w_031_4356, w_031_4360, w_031_4363, w_031_4365, w_031_4366, w_031_4367, w_031_4368, w_031_4369, w_031_4370, w_031_4372, w_031_4373, w_031_4374, w_031_4375, w_031_4376, w_031_4377, w_031_4379, w_031_4386, w_031_4387, w_031_4388, w_031_4389, w_031_4390, w_031_4391, w_031_4392, w_031_4393, w_031_4394, w_031_4395, w_031_4396, w_031_4397, w_031_4398, w_031_4399, w_031_4400, w_031_4404, w_031_4406, w_031_4410, w_031_4411, w_031_4415, w_031_4416, w_031_4417, w_031_4419, w_031_4421, w_031_4422, w_031_4424, w_031_4426, w_031_4427, w_031_4429, w_031_4430, w_031_4431, w_031_4432, w_031_4433, w_031_4434, w_031_4435, w_031_4437, w_031_4438, w_031_4439, w_031_4441, w_031_4444, w_031_4445, w_031_4447, w_031_4449, w_031_4454, w_031_4456, w_031_4457, w_031_4460, w_031_4462, w_031_4463, w_031_4464, w_031_4466, w_031_4468, w_031_4470, w_031_4475, w_031_4477, w_031_4480, w_031_4481, w_031_4482, w_031_4483, w_031_4484, w_031_4486, w_031_4488, w_031_4491, w_031_4495, w_031_4496, w_031_4497, w_031_4498, w_031_4499, w_031_4500, w_031_4502, w_031_4505, w_031_4507, w_031_4508, w_031_4511, w_031_4513, w_031_4516, w_031_4517, w_031_4519, w_031_4522, w_031_4524, w_031_4526, w_031_4527, w_031_4529, w_031_4530, w_031_4533, w_031_4535, w_031_4537, w_031_4538, w_031_4539, w_031_4540, w_031_4541, w_031_4542, w_031_4544, w_031_4545, w_031_4547, w_031_4549, w_031_4554, w_031_4555, w_031_4559, w_031_4561, w_031_4563, w_031_4564, w_031_4568, w_031_4573, w_031_4574, w_031_4575, w_031_4577, w_031_4578, w_031_4580, w_031_4582, w_031_4585, w_031_4586, w_031_4588, w_031_4589, w_031_4592, w_031_4593, w_031_4594, w_031_4596, w_031_4597, w_031_4601, w_031_4602, w_031_4604, w_031_4605, w_031_4610, w_031_4611, w_031_4612, w_031_4613, w_031_4615, w_031_4618, w_031_4622, w_031_4623, w_031_4625, w_031_4626, w_031_4627, w_031_4630, w_031_4631, w_031_4634, w_031_4635, w_031_4637, w_031_4638, w_031_4640, w_031_4641, w_031_4642, w_031_4643, w_031_4645, w_031_4646, w_031_4647, w_031_4648, w_031_4650, w_031_4652, w_031_4654, w_031_4662, w_031_4664, w_031_4665, w_031_4666, w_031_4667, w_031_4668, w_031_4671, w_031_4673, w_031_4675, w_031_4676, w_031_4679, w_031_4681, w_031_4684, w_031_4685, w_031_4686, w_031_4687, w_031_4688, w_031_4690, w_031_4691, w_031_4692, w_031_4693, w_031_4699, w_031_4701, w_031_4702, w_031_4703, w_031_4704, w_031_4705, w_031_4706, w_031_4707, w_031_4710, w_031_4711, w_031_4712, w_031_4713, w_031_4714, w_031_4715, w_031_4716, w_031_4717, w_031_4718, w_031_4719, w_031_4720, w_031_4721, w_031_4722, w_031_4723, w_031_4724, w_031_4725, w_031_4727, w_031_4729, w_031_4732, w_031_4734, w_031_4738, w_031_4739, w_031_4740, w_031_4743, w_031_4746, w_031_4747, w_031_4749, w_031_4751, w_031_4752, w_031_4754, w_031_4755, w_031_4756, w_031_4757, w_031_4760, w_031_4765, w_031_4766, w_031_4772, w_031_4773, w_031_4774, w_031_4775, w_031_4777, w_031_4778, w_031_4779, w_031_4780, w_031_4781, w_031_4783, w_031_4786, w_031_4790, w_031_4792, w_031_4793, w_031_4794, w_031_4797, w_031_4798, w_031_4802, w_031_4803, w_031_4805, w_031_4806, w_031_4807, w_031_4808, w_031_4809, w_031_4810, w_031_4811, w_031_4814, w_031_4816, w_031_4819, w_031_4820, w_031_4825, w_031_4827, w_031_4830, w_031_4832, w_031_4838, w_031_4842, w_031_4843, w_031_4844, w_031_4848, w_031_4849, w_031_4850, w_031_4854, w_031_4858, w_031_4860, w_031_4863, w_031_4864, w_031_4865, w_031_4866, w_031_4867, w_031_4868, w_031_4874, w_031_4875, w_031_4876, w_031_4877, w_031_4879, w_031_4884, w_031_4885, w_031_4886, w_031_4887, w_031_4889, w_031_4890, w_031_4892, w_031_4894, w_031_4896, w_031_4899, w_031_4901, w_031_4902, w_031_4903, w_031_4904, w_031_4905, w_031_4908, w_031_4913, w_031_4915, w_031_4916, w_031_4919, w_031_4920, w_031_4921, w_031_4923, w_031_4924, w_031_4933, w_031_4934, w_031_4936, w_031_4938, w_031_4939, w_031_4940, w_031_4942, w_031_4943, w_031_4944, w_031_4946, w_031_4947, w_031_4949, w_031_4953, w_031_4956, w_031_4957, w_031_4958, w_031_4959, w_031_4960, w_031_4961, w_031_4962, w_031_4963, w_031_4968, w_031_4969, w_031_4970, w_031_4971, w_031_4972, w_031_4974, w_031_4975, w_031_4977, w_031_4978, w_031_4980, w_031_4982, w_031_4983, w_031_4984, w_031_4987, w_031_4988, w_031_4990, w_031_4992, w_031_4994, w_031_4995, w_031_4996, w_031_4999, w_031_5002, w_031_5005, w_031_5006, w_031_5007, w_031_5008, w_031_5010, w_031_5011, w_031_5012, w_031_5013, w_031_5014, w_031_5015, w_031_5018, w_031_5019, w_031_5020, w_031_5024, w_031_5025, w_031_5026, w_031_5027, w_031_5029, w_031_5031, w_031_5032, w_031_5033, w_031_5034, w_031_5035, w_031_5037, w_031_5041, w_031_5042, w_031_5043, w_031_5044, w_031_5045, w_031_5048, w_031_5049, w_031_5050, w_031_5051, w_031_5053, w_031_5054, w_031_5055, w_031_5056, w_031_5057, w_031_5058, w_031_5061, w_031_5062, w_031_5065, w_031_5068, w_031_5069, w_031_5071, w_031_5072, w_031_5073, w_031_5074, w_031_5075, w_031_5078, w_031_5080, w_031_5081, w_031_5082, w_031_5083, w_031_5086, w_031_5089, w_031_5090, w_031_5093, w_031_5095, w_031_5096, w_031_5098, w_031_5101, w_031_5106, w_031_5107, w_031_5108, w_031_5110, w_031_5113, w_031_5114, w_031_5116, w_031_5117, w_031_5118, w_031_5119, w_031_5121, w_031_5122, w_031_5126, w_031_5130, w_031_5134, w_031_5136, w_031_5138, w_031_5140, w_031_5143, w_031_5144, w_031_5151, w_031_5152, w_031_5153, w_031_5156, w_031_5158, w_031_5160, w_031_5162, w_031_5163, w_031_5165, w_031_5167, w_031_5168, w_031_5169, w_031_5170, w_031_5172, w_031_5174, w_031_5177, w_031_5178, w_031_5179, w_031_5180, w_031_5182, w_031_5184, w_031_5186, w_031_5187, w_031_5190, w_031_5193, w_031_5194, w_031_5195, w_031_5196, w_031_5201, w_031_5202, w_031_5205, w_031_5208, w_031_5209, w_031_5210, w_031_5211, w_031_5212, w_031_5213, w_031_5214, w_031_5216, w_031_5217, w_031_5218, w_031_5220, w_031_5222, w_031_5224, w_031_5226, w_031_5227, w_031_5228, w_031_5232, w_031_5233, w_031_5234, w_031_5235, w_031_5236, w_031_5237, w_031_5239, w_031_5240, w_031_5241, w_031_5242, w_031_5243, w_031_5244, w_031_5246, w_031_5249, w_031_5250, w_031_5252, w_031_5254, w_031_5255, w_031_5256, w_031_5258, w_031_5259, w_031_5261, w_031_5262, w_031_5266, w_031_5268, w_031_5269, w_031_5270, w_031_5271, w_031_5272, w_031_5273, w_031_5274, w_031_5277, w_031_5280, w_031_5281, w_031_5283, w_031_5284, w_031_5285, w_031_5286, w_031_5287, w_031_5289, w_031_5290, w_031_5291, w_031_5292, w_031_5293, w_031_5294, w_031_5295, w_031_5296, w_031_5297, w_031_5303, w_031_5304, w_031_5306, w_031_5309, w_031_5311, w_031_5312, w_031_5316, w_031_5321, w_031_5325, w_031_5326, w_031_5331, w_031_5335, w_031_5336, w_031_5337, w_031_5338, w_031_5339, w_031_5340, w_031_5341, w_031_5342, w_031_5343, w_031_5345, w_031_5346, w_031_5349, w_031_5351, w_031_5353, w_031_5354, w_031_5355, w_031_5356, w_031_5361, w_031_5363, w_031_5364, w_031_5365, w_031_5369, w_031_5370, w_031_5375, w_031_5377, w_031_5378, w_031_5379, w_031_5380, w_031_5381, w_031_5382, w_031_5386, w_031_5388, w_031_5389, w_031_5391, w_031_5393, w_031_5396, w_031_5398, w_031_5399, w_031_5400, w_031_5401, w_031_5402, w_031_5404, w_031_5406, w_031_5408, w_031_5409, w_031_5413, w_031_5414, w_031_5417, w_031_5419, w_031_5424, w_031_5425, w_031_5426, w_031_5427, w_031_5428, w_031_5429, w_031_5430, w_031_5431, w_031_5437, w_031_5440, w_031_5441, w_031_5442, w_031_5445, w_031_5448, w_031_5455, w_031_5462, w_031_5463, w_031_5464, w_031_5465, w_031_5468, w_031_5470, w_031_5471, w_031_5472, w_031_5474, w_031_5475, w_031_5477, w_031_5478, w_031_5480, w_031_5481, w_031_5482, w_031_5484, w_031_5485, w_031_5486, w_031_5487, w_031_5488, w_031_5489, w_031_5491, w_031_5493, w_031_5495, w_031_5496, w_031_5499, w_031_5500, w_031_5501, w_031_5504, w_031_5505, w_031_5506, w_031_5507, w_031_5509, w_031_5510, w_031_5515, w_031_5520, w_031_5521, w_031_5522, w_031_5523, w_031_5524, w_031_5525, w_031_5526, w_031_5527, w_031_5528, w_031_5531, w_031_5533, w_031_5534, w_031_5536, w_031_5537, w_031_5541, w_031_5542, w_031_5545, w_031_5549, w_031_5550, w_031_5551, w_031_5552, w_031_5555, w_031_5557, w_031_5558, w_031_5561, w_031_5566, w_031_5567, w_031_5568, w_031_5570, w_031_5571, w_031_5572, w_031_5573, w_031_5574, w_031_5576, w_031_5577, w_031_5578, w_031_5580, w_031_5581, w_031_5584, w_031_5589, w_031_5591, w_031_5592, w_031_5596, w_031_5597, w_031_5598, w_031_5599, w_031_5600, w_031_5603, w_031_5605, w_031_5606, w_031_5610, w_031_5613, w_031_5617, w_031_5618, w_031_5619, w_031_5620, w_031_5623, w_031_5624, w_031_5625, w_031_5630, w_031_5631, w_031_5633, w_031_5634, w_031_5636, w_031_5637, w_031_5640, w_031_5642, w_031_5644, w_031_5646, w_031_5647, w_031_5648, w_031_5652, w_031_5655, w_031_5656, w_031_5662, w_031_5663, w_031_5664, w_031_5665, w_031_5666, w_031_5667, w_031_5668, w_031_5669, w_031_5671, w_031_5675, w_031_5676, w_031_5677, w_031_5678, w_031_5679, w_031_5680, w_031_5682, w_031_5683, w_031_5684, w_031_5685, w_031_5689, w_031_5690, w_031_5691, w_031_5692, w_031_5693, w_031_5694, w_031_5695, w_031_5698, w_031_5700, w_031_5701, w_031_5703, w_031_5705, w_031_5706, w_031_5707, w_031_5709, w_031_5716, w_031_5722, w_031_5723, w_031_5725, w_031_5726, w_031_5729, w_031_5732, w_031_5733, w_031_5734, w_031_5735, w_031_5736, w_031_5737, w_031_5738, w_031_5739, w_031_5742, w_031_5743, w_031_5744, w_031_5747, w_031_5748, w_031_5749, w_031_5750, w_031_5751, w_031_5752, w_031_5754, w_031_5755, w_031_5757, w_031_5759, w_031_5760, w_031_5761, w_031_5763, w_031_5764, w_031_5765, w_031_5767, w_031_5768, w_031_5773, w_031_5775, w_031_5776, w_031_5777, w_031_5779, w_031_5781, w_031_5782, w_031_5783, w_031_5786, w_031_5789, w_031_5790, w_031_5792, w_031_5793, w_031_5794, w_031_5795, w_031_5797, w_031_5798, w_031_5799, w_031_5802, w_031_5804, w_031_5805, w_031_5806, w_031_5807, w_031_5808, w_031_5810, w_031_5812, w_031_5813, w_031_5814, w_031_5815, w_031_5818, w_031_5820, w_031_5822, w_031_5824, w_031_5825, w_031_5831, w_031_5832, w_031_5833, w_031_5834, w_031_5836, w_031_5837, w_031_5838, w_031_5839, w_031_5840, w_031_5842, w_031_5848, w_031_5851, w_031_5854, w_031_5856, w_031_5859, w_031_5861, w_031_5862, w_031_5863, w_031_5866, w_031_5868, w_031_5872, w_031_5874, w_031_5876, w_031_5877, w_031_5879, w_031_5880, w_031_5881, w_031_5884, w_031_5886, w_031_5888, w_031_5890, w_031_5891, w_031_5892, w_031_5893, w_031_5894, w_031_5896, w_031_5897, w_031_5898, w_031_5899, w_031_5900, w_031_5902, w_031_5904, w_031_5905, w_031_5906, w_031_5907, w_031_5908, w_031_5911, w_031_5912, w_031_5913, w_031_5914, w_031_5915, w_031_5916, w_031_5917, w_031_5918, w_031_5920, w_031_5921, w_031_5924, w_031_5928, w_031_5929, w_031_5931, w_031_5932, w_031_5933, w_031_5935, w_031_5936, w_031_5938, w_031_5940, w_031_5941, w_031_5943, w_031_5947, w_031_5948, w_031_5951, w_031_5953, w_031_5954, w_031_5955, w_031_5957, w_031_5958, w_031_5959, w_031_5962, w_031_5963, w_031_5964, w_031_5965, w_031_5967, w_031_5968, w_031_5969, w_031_5970, w_031_5972, w_031_5974, w_031_5975, w_031_5976, w_031_5979, w_031_5980, w_031_5981, w_031_5982, w_031_5983, w_031_5987, w_031_5991, w_031_5993, w_031_5994, w_031_5995, w_031_5997, w_031_5998, w_031_6000, w_031_6001, w_031_6002, w_031_6005, w_031_6006, w_031_6007, w_031_6010, w_031_6012, w_031_6013, w_031_6014, w_031_6016, w_031_6019, w_031_6021, w_031_6022, w_031_6025, w_031_6026, w_031_6028, w_031_6032, w_031_6033, w_031_6036, w_031_6037, w_031_6039, w_031_6040, w_031_6041, w_031_6042, w_031_6047, w_031_6049, w_031_6051, w_031_6052, w_031_6054, w_031_6057, w_031_6058, w_031_6060, w_031_6061, w_031_6062, w_031_6063, w_031_6065, w_031_6068, w_031_6070, w_031_6072, w_031_6075, w_031_6076, w_031_6078, w_031_6079, w_031_6080, w_031_6081, w_031_6084, w_031_6085, w_031_6087, w_031_6088, w_031_6090, w_031_6092, w_031_6094, w_031_6095, w_031_6096, w_031_6098, w_031_6101, w_031_6102, w_031_6107, w_031_6109, w_031_6111, w_031_6112, w_031_6113, w_031_6114, w_031_6115, w_031_6117, w_031_6118, w_031_6119, w_031_6121, w_031_6122, w_031_6123, w_031_6125, w_031_6127, w_031_6128, w_031_6130, w_031_6132, w_031_6133, w_031_6136, w_031_6137, w_031_6138, w_031_6143, w_031_6144, w_031_6145, w_031_6146, w_031_6147, w_031_6150, w_031_6153, w_031_6154, w_031_6155, w_031_6156, w_031_6161, w_031_6162, w_031_6163, w_031_6165, w_031_6166, w_031_6169, w_031_6170, w_031_6172, w_031_6174, w_031_6175, w_031_6177, w_031_6180, w_031_6182, w_031_6183, w_031_6185, w_031_6186, w_031_6188, w_031_6190, w_031_6191, w_031_6192, w_031_6193, w_031_6195, w_031_6197, w_031_6199, w_031_6200, w_031_6202, w_031_6203, w_031_6205, w_031_6207, w_031_6208, w_031_6209, w_031_6212, w_031_6213, w_031_6214, w_031_6215, w_031_6217, w_031_6219, w_031_6223, w_031_6226, w_031_6230, w_031_6232, w_031_6233, w_031_6235, w_031_6237, w_031_6238, w_031_6242, w_031_6243, w_031_6244, w_031_6245, w_031_6248, w_031_6250, w_031_6251, w_031_6253, w_031_6257, w_031_6259, w_031_6261, w_031_6262, w_031_6263, w_031_6265, w_031_6267, w_031_6269, w_031_6273, w_031_6275, w_031_6276, w_031_6278, w_031_6279, w_031_6280, w_031_6281, w_031_6283, w_031_6284, w_031_6286, w_031_6287, w_031_6288, w_031_6289, w_031_6291, w_031_6293, w_031_6295, w_031_6301, w_031_6302, w_031_6303, w_031_6304, w_031_6306, w_031_6307, w_031_6309, w_031_6310, w_031_6311, w_031_6312, w_031_6313, w_031_6318, w_031_6319, w_031_6320, w_031_6321, w_031_6323, w_031_6325, w_031_6326, w_031_6330, w_031_6331, w_031_6333, w_031_6335, w_031_6336, w_031_6337, w_031_6339, w_031_6341, w_031_6342, w_031_6343, w_031_6346, w_031_6347, w_031_6348, w_031_6349, w_031_6354, w_031_6356, w_031_6357, w_031_6359, w_031_6360, w_031_6363, w_031_6366, w_031_6367, w_031_6368, w_031_6369, w_031_6371, w_031_6374, w_031_6375, w_031_6376, w_031_6377, w_031_6380, w_031_6381, w_031_6382, w_031_6384, w_031_6385, w_031_6386, w_031_6389, w_031_6390, w_031_6392, w_031_6393, w_031_6394, w_031_6395, w_031_6397, w_031_6398, w_031_6400, w_031_6401, w_031_6402, w_031_6404, w_031_6407, w_031_6408, w_031_6411, w_031_6413, w_031_6414, w_031_6415, w_031_6418, w_031_6419, w_031_6420, w_031_6421, w_031_6422, w_031_6423, w_031_6425, w_031_6426, w_031_6427, w_031_6429, w_031_6430, w_031_6434, w_031_6438, w_031_6440, w_031_6441, w_031_6442, w_031_6443, w_031_6444, w_031_6445, w_031_6446, w_031_6449, w_031_6450, w_031_6451, w_031_6452, w_031_6453, w_031_6456, w_031_6458, w_031_6461, w_031_6462, w_031_6463, w_031_6467, w_031_6469, w_031_6472, w_031_6473, w_031_6474, w_031_6475, w_031_6477, w_031_6482, w_031_6483, w_031_6484, w_031_6485, w_031_6486, w_031_6490, w_031_6491, w_031_6492, w_031_6494, w_031_6495, w_031_6496, w_031_6497, w_031_6498, w_031_6500, w_031_6503, w_031_6504, w_031_6507, w_031_6508, w_031_6511, w_031_6512, w_031_6516, w_031_6518, w_031_6519, w_031_6521, w_031_6523, w_031_6524, w_031_6529, w_031_6531, w_031_6534, w_031_6535, w_031_6536, w_031_6538, w_031_6539, w_031_6540, w_031_6541, w_031_6543, w_031_6544, w_031_6546, w_031_6547, w_031_6551, w_031_6554, w_031_6556, w_031_6558, w_031_6561, w_031_6563, w_031_6566, w_031_6569, w_031_6570, w_031_6572, w_031_6574, w_031_6575, w_031_6576, w_031_6578, w_031_6579, w_031_6580, w_031_6581, w_031_6583, w_031_6590, w_031_6592, w_031_6595, w_031_6596, w_031_6598, w_031_6601, w_031_6605, w_031_6609, w_031_6610, w_031_6611, w_031_6613, w_031_6615, w_031_6616, w_031_6617, w_031_6622, w_031_6623, w_031_6624, w_031_6625, w_031_6634, w_031_6635, w_031_6640, w_031_6642, w_031_6643, w_031_6645, w_031_6648, w_031_6650, w_031_6655, w_031_6656, w_031_6657, w_031_6659, w_031_6660, w_031_6662, w_031_6663, w_031_6664, w_031_6667, w_031_6668, w_031_6669, w_031_6670, w_031_6671, w_031_6672, w_031_6675, w_031_6677, w_031_6679, w_031_6681, w_031_6682, w_031_6683, w_031_6687, w_031_6689, w_031_6691, w_031_6693, w_031_6694, w_031_6696, w_031_6701, w_031_6702, w_031_6703, w_031_6708, w_031_6710, w_031_6711, w_031_6712, w_031_6716, w_031_6717, w_031_6718, w_031_6719, w_031_6720, w_031_6722, w_031_6723, w_031_6724, w_031_6726, w_031_6727, w_031_6728, w_031_6731, w_031_6735, w_031_6738, w_031_6743, w_031_6744, w_031_6745, w_031_6748, w_031_6749, w_031_6751, w_031_6753, w_031_6754, w_031_6757, w_031_6760, w_031_6762, w_031_6763, w_031_6765, w_031_6766, w_031_6767, w_031_6768, w_031_6769, w_031_6770, w_031_6772, w_031_6774, w_031_6777, w_031_6778, w_031_6779, w_031_6780, w_031_6781, w_031_6782, w_031_6785, w_031_6786, w_031_6787, w_031_6789, w_031_6791, w_031_6792, w_031_6793, w_031_6795, w_031_6796, w_031_6797, w_031_6798, w_031_6802, w_031_6806, w_031_6807, w_031_6809, w_031_6810, w_031_6811, w_031_6812, w_031_6814, w_031_6815, w_031_6817, w_031_6818, w_031_6819, w_031_6821, w_031_6822, w_031_6823, w_031_6824, w_031_6825, w_031_6826, w_031_6827, w_031_6829, w_031_6830, w_031_6833, w_031_6834, w_031_6835, w_031_6837, w_031_6839, w_031_6842, w_031_6843, w_031_6844, w_031_6845, w_031_6846, w_031_6847, w_031_6849, w_031_6851, w_031_6852, w_031_6853, w_031_6855, w_031_6856, w_031_6858, w_031_6860, w_031_6861, w_031_6862, w_031_6863, w_031_6865, w_031_6866, w_031_6868, w_031_6869, w_031_6872, w_031_6873, w_031_6874, w_031_6875, w_031_6876, w_031_6877, w_031_6878, w_031_6880, w_031_6883, w_031_6887, w_031_6888, w_031_6889, w_031_6892, w_031_6893, w_031_6896, w_031_6898, w_031_6899, w_031_6900, w_031_6901, w_031_6902, w_031_6903, w_031_6904, w_031_6906, w_031_6911, w_031_6912, w_031_6913, w_031_6915, w_031_6916, w_031_6919, w_031_6920, w_031_6921, w_031_6923, w_031_6924, w_031_6925, w_031_6927, w_031_6928, w_031_6929, w_031_6931, w_031_6932, w_031_6933, w_031_6934, w_031_6938, w_031_6939, w_031_6948, w_031_6951, w_031_6952, w_031_6953, w_031_6955, w_031_6956, w_031_6957, w_031_6959, w_031_6960, w_031_6961, w_031_6962, w_031_6964, w_031_6965, w_031_6966, w_031_6968, w_031_6969, w_031_6971, w_031_6973, w_031_6974, w_031_6976, w_031_6979, w_031_6981, w_031_6982, w_031_6985, w_031_6986, w_031_6987, w_031_6990, w_031_6992, w_031_6993, w_031_7001, w_031_7002, w_031_7003, w_031_7004, w_031_7005, w_031_7006, w_031_7007, w_031_7012, w_031_7013, w_031_7014, w_031_7015, w_031_7016, w_031_7018, w_031_7020, w_031_7021, w_031_7022, w_031_7025, w_031_7026, w_031_7028, w_031_7031, w_031_7032, w_031_7033, w_031_7034, w_031_7035, w_031_7038, w_031_7041, w_031_7043, w_031_7045, w_031_7048, w_031_7049, w_031_7050, w_031_7052, w_031_7055, w_031_7056, w_031_7058, w_031_7059, w_031_7060, w_031_7061, w_031_7062, w_031_7065, w_031_7068, w_031_7071, w_031_7072, w_031_7076, w_031_7078, w_031_7079, w_031_7081, w_031_7082, w_031_7083, w_031_7084, w_031_7085, w_031_7086, w_031_7087, w_031_7088, w_031_7089, w_031_7091, w_031_7096, w_031_7098, w_031_7099, w_031_7100, w_031_7101, w_031_7102, w_031_7105, w_031_7106, w_031_7108, w_031_7109, w_031_7110, w_031_7113, w_031_7114, w_031_7115, w_031_7116, w_031_7117, w_031_7119, w_031_7121, w_031_7123, w_031_7127, w_031_7128, w_031_7131, w_031_7132, w_031_7136, w_031_7138, w_031_7139, w_031_7140, w_031_7141, w_031_7142, w_031_7147, w_031_7148, w_031_7152, w_031_7153, w_031_7154, w_031_7155, w_031_7156, w_031_7158, w_031_7159, w_031_7167, w_031_7168, w_031_7169, w_031_7170, w_031_7171, w_031_7172, w_031_7174, w_031_7175, w_031_7176, w_031_7178, w_031_7180, w_031_7182, w_031_7184, w_031_7185, w_031_7186, w_031_7188, w_031_7189, w_031_7190, w_031_7191, w_031_7192, w_031_7193, w_031_7194, w_031_7196, w_031_7197, w_031_7198, w_031_7199, w_031_7201, w_031_7203, w_031_7204, w_031_7206, w_031_7209, w_031_7211, w_031_7215, w_031_7216, w_031_7217, w_031_7222, w_031_7223, w_031_7227, w_031_7228, w_031_7229, w_031_7230, w_031_7231, w_031_7232, w_031_7234, w_031_7237, w_031_7239, w_031_7240, w_031_7242, w_031_7243, w_031_7245, w_031_7247, w_031_7248, w_031_7251, w_031_7252, w_031_7255, w_031_7260, w_031_7261, w_031_7262, w_031_7263, w_031_7265, w_031_7266, w_031_7269, w_031_7274, w_031_7277, w_031_7278, w_031_7279, w_031_7282, w_031_7283, w_031_7284, w_031_7287, w_031_7292, w_031_7293, w_031_7294, w_031_7295, w_031_7301, w_031_7303, w_031_7304, w_031_7305, w_031_7307, w_031_7310, w_031_7316, w_031_7317, w_031_7319, w_031_7320, w_031_7321, w_031_7323, w_031_7324, w_031_7332, w_031_7334, w_031_7335, w_031_7337, w_031_7338, w_031_7339, w_031_7340, w_031_7341, w_031_7343, w_031_7344, w_031_7345, w_031_7348, w_031_7350, w_031_7353, w_031_7355, w_031_7357, w_031_7361, w_031_7363, w_031_7364, w_031_7365, w_031_7366, w_031_7368, w_031_7369, w_031_7370, w_031_7372, w_031_7374, w_031_7378, w_031_7380, w_031_7381, w_031_7382, w_031_7383, w_031_7386, w_031_7388, w_031_7389, w_031_7390, w_031_7391, w_031_7392, w_031_7394, w_031_7395, w_031_7396, w_031_7398, w_031_7399, w_031_7401, w_031_7402, w_031_7403, w_031_7406, w_031_7409, w_031_7411, w_031_7412, w_031_7414, w_031_7415, w_031_7416, w_031_7417, w_031_7418, w_031_7419, w_031_7421, w_031_7422, w_031_7423, w_031_7424, w_031_7427, w_031_7428, w_031_7429, w_031_7430, w_031_7431, w_031_7432, w_031_7434, w_031_7435, w_031_7436, w_031_7437, w_031_7438, w_031_7439, w_031_7440, w_031_7442, w_031_7445, w_031_7447, w_031_7448, w_031_7449, w_031_7452, w_031_7454, w_031_7456, w_031_7461, w_031_7463, w_031_7465, w_031_7466, w_031_7467, w_031_7468, w_031_7470, w_031_7472, w_031_7473, w_031_7474, w_031_7477, w_031_7478, w_031_7479, w_031_7488, w_031_7490, w_031_7491, w_031_7494, w_031_7498, w_031_7499, w_031_7501, w_031_7502, w_031_7503, w_031_7505, w_031_7506, w_031_7508, w_031_7510, w_031_7512, w_031_7513, w_031_7518, w_031_7520, w_031_7522, w_031_7523, w_031_7527, w_031_7528, w_031_7529, w_031_7530, w_031_7531, w_031_7532, w_031_7534, w_031_7536, w_031_7538, w_031_7539, w_031_7540, w_031_7542, w_031_7543, w_031_7544, w_031_7545, w_031_7546, w_031_7547, w_031_7549, w_031_7551, w_031_7553, w_031_7554, w_031_7558, w_031_7560, w_031_7561, w_031_7562, w_031_7564, w_031_7565, w_031_7567, w_031_7569, w_031_7570, w_031_7571, w_031_7573, w_031_7574, w_031_7575, w_031_7577, w_031_7578, w_031_7579, w_031_7580, w_031_7581, w_031_7584, w_031_7586, w_031_7587, w_031_7589, w_031_7590, w_031_7593, w_031_7594, w_031_7597, w_031_7598, w_031_7599, w_031_7602, w_031_7604, w_031_7605, w_031_7607, w_031_7608, w_031_7610, w_031_7611, w_031_7612, w_031_7613, w_031_7614, w_031_7615, w_031_7617, w_031_7620, w_031_7622, w_031_7624, w_031_7629, w_031_7630, w_031_7631, w_031_7632, w_031_7641, w_031_7642, w_031_7643, w_031_7644, w_031_7646, w_031_7651, w_031_7652, w_031_7653, w_031_7657, w_031_7658, w_031_7659, w_031_7661, w_031_7664, w_031_7666, w_031_7667, w_031_7668, w_031_7671, w_031_7672, w_031_7673, w_031_7676, w_031_7678, w_031_7679, w_031_7681, w_031_7682, w_031_7683, w_031_7684, w_031_7686, w_031_7688, w_031_7689, w_031_7690, w_031_7693, w_031_7694, w_031_7695, w_031_7697, w_031_7698, w_031_7699, w_031_7700, w_031_7702, w_031_7706, w_031_7707, w_031_7708, w_031_7709, w_031_7710, w_031_7711, w_031_7712, w_031_7713, w_031_7714, w_031_7715, w_031_7716, w_031_7718, w_031_7720, w_031_7723, w_031_7724, w_031_7726, w_031_7729, w_031_7730, w_031_7731, w_031_7732, w_031_7733, w_031_7735, w_031_7737, w_031_7738, w_031_7739, w_031_7740, w_031_7741, w_031_7745, w_031_7747, w_031_7748, w_031_7749, w_031_7752, w_031_7755, w_031_7757, w_031_7758, w_031_7759, w_031_7760, w_031_7761, w_031_7762, w_031_7763, w_031_7764, w_031_7767, w_031_7770, w_031_7771, w_031_7772, w_031_7773, w_031_7774, w_031_7776, w_031_7777, w_031_7780, w_031_7781, w_031_7782, w_031_7784, w_031_7785, w_031_7786, w_031_7788, w_031_7791, w_031_7792, w_031_7794, w_031_7795, w_031_7796, w_031_7798, w_031_7802, w_031_7803, w_031_7805, w_031_7806, w_031_7807, w_031_7811, w_031_7812, w_031_7813, w_031_7814, w_031_7816, w_031_7817, w_031_7818, w_031_7826, w_031_7827, w_031_7828, w_031_7829, w_031_7831, w_031_7832, w_031_7834, w_031_7836, w_031_7838, w_031_7840, w_031_7841, w_031_7842, w_031_7843, w_031_7844, w_031_7845, w_031_7846, w_031_7848, w_031_7849, w_031_7850, w_031_7852, w_031_7855, w_031_7857, w_031_7858, w_031_7860, w_031_7862, w_031_7865, w_031_7866, w_031_7867, w_031_7869, w_031_7872, w_031_7875, w_031_7876, w_031_7877, w_031_7880, w_031_7881, w_031_7882, w_031_7883, w_031_7884, w_031_7888, w_031_7891, w_031_7893, w_031_7894, w_031_7900, w_031_7901, w_031_7903, w_031_7904, w_031_7905, w_031_7912, w_031_7913;
  wire w_032_001, w_032_003, w_032_004, w_032_005, w_032_006, w_032_007, w_032_008, w_032_010, w_032_012, w_032_016, w_032_018, w_032_019, w_032_020, w_032_021, w_032_022, w_032_023, w_032_026, w_032_028, w_032_029, w_032_030, w_032_032, w_032_033, w_032_034, w_032_035, w_032_036, w_032_037, w_032_038, w_032_039, w_032_041, w_032_042, w_032_043, w_032_044, w_032_045, w_032_046, w_032_047, w_032_048, w_032_050, w_032_052, w_032_053, w_032_054, w_032_055, w_032_057, w_032_059, w_032_060, w_032_062, w_032_063, w_032_064, w_032_066, w_032_067, w_032_069, w_032_071, w_032_072, w_032_073, w_032_074, w_032_075, w_032_076, w_032_077, w_032_078, w_032_079, w_032_080, w_032_081, w_032_082, w_032_083, w_032_084, w_032_085, w_032_087, w_032_088, w_032_090, w_032_091, w_032_093, w_032_094, w_032_096, w_032_098, w_032_099, w_032_100, w_032_103, w_032_104, w_032_105, w_032_106, w_032_108, w_032_109, w_032_110, w_032_111, w_032_112, w_032_113, w_032_114, w_032_115, w_032_117, w_032_118, w_032_119, w_032_121, w_032_122, w_032_123, w_032_124, w_032_126, w_032_127, w_032_128, w_032_129, w_032_130, w_032_132, w_032_133, w_032_134, w_032_135, w_032_137, w_032_138, w_032_139, w_032_140, w_032_141, w_032_142, w_032_143, w_032_144, w_032_146, w_032_147, w_032_150, w_032_151, w_032_152, w_032_155, w_032_156, w_032_157, w_032_158, w_032_159, w_032_160, w_032_161, w_032_162, w_032_163, w_032_164, w_032_165, w_032_166, w_032_167, w_032_168, w_032_169, w_032_170, w_032_171, w_032_172, w_032_173, w_032_175, w_032_176, w_032_177, w_032_178, w_032_179, w_032_180, w_032_181, w_032_182, w_032_183, w_032_184, w_032_185, w_032_187, w_032_188, w_032_189, w_032_191, w_032_192, w_032_194, w_032_195, w_032_196, w_032_197, w_032_198, w_032_199, w_032_200, w_032_201, w_032_202, w_032_203, w_032_204, w_032_206, w_032_208, w_032_209, w_032_210, w_032_211, w_032_213, w_032_214, w_032_215, w_032_216, w_032_217, w_032_218, w_032_219, w_032_220, w_032_221, w_032_222, w_032_223, w_032_225, w_032_227, w_032_228, w_032_229, w_032_232, w_032_233, w_032_235, w_032_236, w_032_237, w_032_238, w_032_239, w_032_240, w_032_241, w_032_242, w_032_243, w_032_244, w_032_245, w_032_246, w_032_247, w_032_248, w_032_249, w_032_251, w_032_252, w_032_253, w_032_255, w_032_256, w_032_259, w_032_260, w_032_261, w_032_262, w_032_263, w_032_265, w_032_266, w_032_267, w_032_268, w_032_269, w_032_270, w_032_271, w_032_273, w_032_274, w_032_275, w_032_276, w_032_277, w_032_278, w_032_279, w_032_280, w_032_281, w_032_282, w_032_283, w_032_286, w_032_288, w_032_289, w_032_290, w_032_291, w_032_293, w_032_296, w_032_297, w_032_298, w_032_299, w_032_300, w_032_301, w_032_302, w_032_303, w_032_304, w_032_306, w_032_308, w_032_309, w_032_310, w_032_311, w_032_313, w_032_314, w_032_315, w_032_316, w_032_318, w_032_319, w_032_321, w_032_323, w_032_324, w_032_325, w_032_326, w_032_327, w_032_329, w_032_330, w_032_332, w_032_333, w_032_334, w_032_335, w_032_336, w_032_337, w_032_338, w_032_339, w_032_340, w_032_341, w_032_342, w_032_343, w_032_345, w_032_346, w_032_347, w_032_348, w_032_350, w_032_351, w_032_353, w_032_354, w_032_355, w_032_357, w_032_360, w_032_362, w_032_363, w_032_364, w_032_365, w_032_366, w_032_367, w_032_368, w_032_369, w_032_371, w_032_372, w_032_373, w_032_375, w_032_376, w_032_377, w_032_378, w_032_379, w_032_380, w_032_381, w_032_382, w_032_386, w_032_388, w_032_389, w_032_390, w_032_394, w_032_395, w_032_396, w_032_397, w_032_398, w_032_399, w_032_400, w_032_401, w_032_402, w_032_403, w_032_404, w_032_405, w_032_406, w_032_407, w_032_408, w_032_409, w_032_410, w_032_411, w_032_413, w_032_414, w_032_415, w_032_416, w_032_417, w_032_418, w_032_419, w_032_420, w_032_421, w_032_422, w_032_423, w_032_424, w_032_426, w_032_428, w_032_429, w_032_430, w_032_431, w_032_432, w_032_433, w_032_434, w_032_435, w_032_436, w_032_437, w_032_438, w_032_440, w_032_441, w_032_442, w_032_445, w_032_446, w_032_448, w_032_449, w_032_450, w_032_451, w_032_452, w_032_453, w_032_455, w_032_456, w_032_457, w_032_458, w_032_459, w_032_460, w_032_464, w_032_465, w_032_466, w_032_468, w_032_469, w_032_470, w_032_471, w_032_475, w_032_476, w_032_477, w_032_478, w_032_480, w_032_481, w_032_484, w_032_485, w_032_486, w_032_487, w_032_488, w_032_490, w_032_491, w_032_492, w_032_493, w_032_494, w_032_495, w_032_496, w_032_497, w_032_500, w_032_502, w_032_503, w_032_504, w_032_506, w_032_508, w_032_509, w_032_510, w_032_511, w_032_514, w_032_515, w_032_516, w_032_517, w_032_518, w_032_519, w_032_520, w_032_521, w_032_522, w_032_523, w_032_524, w_032_525, w_032_526, w_032_527, w_032_528, w_032_529, w_032_530, w_032_531, w_032_532, w_032_534, w_032_535, w_032_536, w_032_537, w_032_538, w_032_541, w_032_542, w_032_544, w_032_545, w_032_546, w_032_547, w_032_548, w_032_551, w_032_552, w_032_553, w_032_554, w_032_555, w_032_556, w_032_557, w_032_558, w_032_559, w_032_560, w_032_561, w_032_562, w_032_563, w_032_564, w_032_565, w_032_566, w_032_567, w_032_568, w_032_569, w_032_571, w_032_573, w_032_574, w_032_575, w_032_576, w_032_577, w_032_578, w_032_579, w_032_580, w_032_581, w_032_582, w_032_583, w_032_584, w_032_585, w_032_587, w_032_588, w_032_589, w_032_591, w_032_592, w_032_596, w_032_597, w_032_598, w_032_600, w_032_601, w_032_602, w_032_603, w_032_604, w_032_606, w_032_607, w_032_608, w_032_610, w_032_611, w_032_612, w_032_613, w_032_614, w_032_616, w_032_617, w_032_618, w_032_619, w_032_621, w_032_622, w_032_623, w_032_624, w_032_625, w_032_627, w_032_629, w_032_630, w_032_633, w_032_634, w_032_635, w_032_637, w_032_638, w_032_639, w_032_641, w_032_644, w_032_645, w_032_646, w_032_648, w_032_649, w_032_650, w_032_651, w_032_652, w_032_653, w_032_654, w_032_655, w_032_656, w_032_657, w_032_658, w_032_659, w_032_660, w_032_661, w_032_662, w_032_663, w_032_664, w_032_665, w_032_666, w_032_667, w_032_669, w_032_670, w_032_671, w_032_673, w_032_674, w_032_675, w_032_676, w_032_677, w_032_679, w_032_680, w_032_681, w_032_682, w_032_683, w_032_685, w_032_686, w_032_687, w_032_689, w_032_690, w_032_691, w_032_692, w_032_693, w_032_694, w_032_695, w_032_697, w_032_698, w_032_699, w_032_700, w_032_701, w_032_702, w_032_703, w_032_704, w_032_705, w_032_706, w_032_707, w_032_708, w_032_710, w_032_711, w_032_713, w_032_715, w_032_716, w_032_717, w_032_718, w_032_720, w_032_721, w_032_722, w_032_723, w_032_724, w_032_725, w_032_726, w_032_728, w_032_730, w_032_731, w_032_732, w_032_733, w_032_734, w_032_735, w_032_737, w_032_738, w_032_739, w_032_741, w_032_744, w_032_745, w_032_746, w_032_747, w_032_748, w_032_749, w_032_750, w_032_751, w_032_752, w_032_754, w_032_756, w_032_758, w_032_759, w_032_760, w_032_763, w_032_764, w_032_765, w_032_766, w_032_768, w_032_769, w_032_771, w_032_773, w_032_774, w_032_775, w_032_776, w_032_777, w_032_778, w_032_779, w_032_780, w_032_781, w_032_783, w_032_784, w_032_785, w_032_786, w_032_787, w_032_789, w_032_791, w_032_792, w_032_793, w_032_794, w_032_795, w_032_796, w_032_797, w_032_798, w_032_799, w_032_800, w_032_801, w_032_802, w_032_803, w_032_804, w_032_805, w_032_806, w_032_807, w_032_808, w_032_809, w_032_810, w_032_811, w_032_812, w_032_813, w_032_814, w_032_816, w_032_817, w_032_818, w_032_819, w_032_820, w_032_821, w_032_822, w_032_824, w_032_825, w_032_826, w_032_827, w_032_828, w_032_829, w_032_830, w_032_831, w_032_832, w_032_833, w_032_835, w_032_836, w_032_837, w_032_838, w_032_839, w_032_840, w_032_841, w_032_842, w_032_843, w_032_845, w_032_848, w_032_849, w_032_852, w_032_853, w_032_855, w_032_856, w_032_857, w_032_858, w_032_859, w_032_860, w_032_862, w_032_864, w_032_866, w_032_871, w_032_872, w_032_873, w_032_875, w_032_876, w_032_877, w_032_878, w_032_879, w_032_880, w_032_882, w_032_883, w_032_884, w_032_885, w_032_886, w_032_887, w_032_888, w_032_889, w_032_892, w_032_894, w_032_898, w_032_899, w_032_900, w_032_902, w_032_903, w_032_906, w_032_908, w_032_910, w_032_911, w_032_912, w_032_915, w_032_916, w_032_917, w_032_918, w_032_919, w_032_920, w_032_921, w_032_923, w_032_924, w_032_925, w_032_926, w_032_927, w_032_928, w_032_930, w_032_931, w_032_932, w_032_933, w_032_934, w_032_935, w_032_937, w_032_938, w_032_939, w_032_941, w_032_942, w_032_944, w_032_945, w_032_946, w_032_947, w_032_948, w_032_949, w_032_950, w_032_951, w_032_953, w_032_954, w_032_955, w_032_956, w_032_958, w_032_959, w_032_962, w_032_963, w_032_964, w_032_966, w_032_967, w_032_968, w_032_969, w_032_970, w_032_971, w_032_972, w_032_973, w_032_974, w_032_975, w_032_976, w_032_977, w_032_978, w_032_980, w_032_981, w_032_983, w_032_984, w_032_985, w_032_986, w_032_987, w_032_988, w_032_989, w_032_990, w_032_991, w_032_992, w_032_993, w_032_994, w_032_995, w_032_998, w_032_999, w_032_1000, w_032_1001, w_032_1002, w_032_1003, w_032_1004, w_032_1005, w_032_1006, w_032_1007, w_032_1008, w_032_1009, w_032_1010, w_032_1011, w_032_1012, w_032_1013, w_032_1014, w_032_1015, w_032_1016, w_032_1017, w_032_1019, w_032_1020, w_032_1021, w_032_1024, w_032_1025, w_032_1026, w_032_1028, w_032_1029, w_032_1030, w_032_1031, w_032_1032, w_032_1033, w_032_1035, w_032_1036, w_032_1039, w_032_1041, w_032_1043, w_032_1044, w_032_1045, w_032_1046, w_032_1047, w_032_1048, w_032_1049, w_032_1051, w_032_1054, w_032_1056, w_032_1057, w_032_1058, w_032_1060, w_032_1063, w_032_1064, w_032_1066, w_032_1067, w_032_1068, w_032_1069, w_032_1070, w_032_1071, w_032_1072, w_032_1073, w_032_1076, w_032_1077, w_032_1079, w_032_1080, w_032_1082, w_032_1083, w_032_1084, w_032_1085, w_032_1086, w_032_1088, w_032_1089, w_032_1090, w_032_1092, w_032_1093, w_032_1094, w_032_1095, w_032_1097, w_032_1098, w_032_1099, w_032_1100, w_032_1101, w_032_1102, w_032_1104, w_032_1105, w_032_1108, w_032_1109, w_032_1111, w_032_1113, w_032_1115, w_032_1116, w_032_1117, w_032_1120, w_032_1121, w_032_1122, w_032_1123, w_032_1124, w_032_1126, w_032_1127, w_032_1128, w_032_1129, w_032_1130, w_032_1131, w_032_1132, w_032_1133, w_032_1134, w_032_1135, w_032_1136, w_032_1137, w_032_1138, w_032_1139, w_032_1140, w_032_1141, w_032_1142, w_032_1143, w_032_1145, w_032_1146, w_032_1147, w_032_1148, w_032_1149, w_032_1150, w_032_1151, w_032_1152, w_032_1153, w_032_1154, w_032_1155, w_032_1157, w_032_1158, w_032_1159, w_032_1160, w_032_1161, w_032_1163, w_032_1164, w_032_1165, w_032_1166, w_032_1167, w_032_1168, w_032_1170, w_032_1173, w_032_1175, w_032_1176, w_032_1177, w_032_1178, w_032_1181, w_032_1182, w_032_1183, w_032_1184, w_032_1185, w_032_1186, w_032_1187, w_032_1189, w_032_1192, w_032_1194, w_032_1195, w_032_1196, w_032_1197, w_032_1198, w_032_1199, w_032_1200, w_032_1201, w_032_1202, w_032_1203, w_032_1204, w_032_1205, w_032_1207, w_032_1208, w_032_1209, w_032_1210, w_032_1211, w_032_1212, w_032_1213, w_032_1216, w_032_1217, w_032_1218, w_032_1220, w_032_1221, w_032_1224, w_032_1225, w_032_1226, w_032_1227, w_032_1228, w_032_1230, w_032_1231, w_032_1232, w_032_1233, w_032_1234, w_032_1235, w_032_1236, w_032_1238, w_032_1239, w_032_1240, w_032_1241, w_032_1243, w_032_1244, w_032_1245, w_032_1246, w_032_1248, w_032_1249, w_032_1250, w_032_1251, w_032_1252, w_032_1253, w_032_1256, w_032_1257, w_032_1258, w_032_1259, w_032_1261, w_032_1262, w_032_1264, w_032_1266, w_032_1269, w_032_1270, w_032_1271, w_032_1272, w_032_1273, w_032_1274, w_032_1275, w_032_1276, w_032_1277, w_032_1278, w_032_1279, w_032_1281, w_032_1282, w_032_1284, w_032_1285, w_032_1286, w_032_1288, w_032_1289, w_032_1291, w_032_1292, w_032_1293, w_032_1294, w_032_1296, w_032_1297, w_032_1298, w_032_1299, w_032_1300, w_032_1301, w_032_1305, w_032_1306, w_032_1307, w_032_1308, w_032_1309, w_032_1311, w_032_1312, w_032_1314, w_032_1315, w_032_1317, w_032_1318, w_032_1320, w_032_1321, w_032_1322, w_032_1324, w_032_1325, w_032_1327, w_032_1328, w_032_1329, w_032_1331, w_032_1332, w_032_1333, w_032_1334, w_032_1335, w_032_1336, w_032_1337, w_032_1338, w_032_1339, w_032_1340, w_032_1341, w_032_1342, w_032_1343, w_032_1344, w_032_1345, w_032_1346, w_032_1347, w_032_1348, w_032_1350, w_032_1351, w_032_1352, w_032_1354, w_032_1355, w_032_1356, w_032_1357, w_032_1359, w_032_1360, w_032_1362, w_032_1363, w_032_1364, w_032_1365, w_032_1366, w_032_1367, w_032_1368, w_032_1369, w_032_1370, w_032_1371, w_032_1372, w_032_1373, w_032_1374, w_032_1375, w_032_1376, w_032_1377, w_032_1378, w_032_1379, w_032_1380, w_032_1381, w_032_1383, w_032_1385, w_032_1386, w_032_1387, w_032_1388, w_032_1389, w_032_1390, w_032_1392, w_032_1393, w_032_1394, w_032_1396, w_032_1398, w_032_1399, w_032_1401, w_032_1402, w_032_1403, w_032_1405, w_032_1406, w_032_1408, w_032_1409, w_032_1410, w_032_1411, w_032_1412, w_032_1413, w_032_1414, w_032_1416, w_032_1417, w_032_1419, w_032_1420, w_032_1421, w_032_1422, w_032_1423, w_032_1424, w_032_1425, w_032_1426, w_032_1427, w_032_1428, w_032_1429, w_032_1430, w_032_1431, w_032_1432, w_032_1433, w_032_1434, w_032_1435, w_032_1436, w_032_1437, w_032_1438, w_032_1441, w_032_1442, w_032_1444, w_032_1445, w_032_1446, w_032_1447, w_032_1448, w_032_1449, w_032_1450, w_032_1451, w_032_1452, w_032_1453, w_032_1454, w_032_1456, w_032_1457, w_032_1458, w_032_1459, w_032_1460, w_032_1461, w_032_1462, w_032_1464, w_032_1465, w_032_1466, w_032_1467, w_032_1468, w_032_1469, w_032_1470, w_032_1471, w_032_1473, w_032_1474, w_032_1475, w_032_1476, w_032_1477, w_032_1479, w_032_1481, w_032_1482, w_032_1484, w_032_1485, w_032_1486, w_032_1487, w_032_1488, w_032_1490, w_032_1492, w_032_1493, w_032_1494, w_032_1495, w_032_1496, w_032_1497, w_032_1498, w_032_1499, w_032_1501, w_032_1502, w_032_1503, w_032_1504, w_032_1505, w_032_1506, w_032_1507, w_032_1508, w_032_1510, w_032_1511, w_032_1512, w_032_1513, w_032_1514, w_032_1516, w_032_1517, w_032_1518, w_032_1521, w_032_1522, w_032_1523, w_032_1527, w_032_1528, w_032_1529, w_032_1530, w_032_1531, w_032_1532, w_032_1533, w_032_1537, w_032_1538, w_032_1540, w_032_1541, w_032_1544, w_032_1546, w_032_1547, w_032_1548, w_032_1549, w_032_1550, w_032_1551, w_032_1552, w_032_1553, w_032_1555, w_032_1556, w_032_1557, w_032_1559, w_032_1560, w_032_1561, w_032_1562, w_032_1564, w_032_1565, w_032_1566, w_032_1567, w_032_1568, w_032_1569, w_032_1570, w_032_1571, w_032_1572, w_032_1575, w_032_1576, w_032_1577, w_032_1578, w_032_1579, w_032_1580, w_032_1581, w_032_1582, w_032_1583, w_032_1584, w_032_1587, w_032_1588, w_032_1589, w_032_1590, w_032_1592, w_032_1593, w_032_1596, w_032_1597, w_032_1598, w_032_1599, w_032_1600, w_032_1601, w_032_1602, w_032_1603, w_032_1604, w_032_1605, w_032_1606, w_032_1608, w_032_1609, w_032_1610, w_032_1611, w_032_1612, w_032_1613, w_032_1614, w_032_1615, w_032_1616, w_032_1617, w_032_1618, w_032_1619, w_032_1620, w_032_1621, w_032_1622, w_032_1623, w_032_1624, w_032_1626, w_032_1629, w_032_1630, w_032_1631, w_032_1632, w_032_1633, w_032_1634, w_032_1635, w_032_1637, w_032_1639, w_032_1642, w_032_1643, w_032_1644, w_032_1645, w_032_1647, w_032_1648, w_032_1649, w_032_1650, w_032_1651, w_032_1654, w_032_1655, w_032_1657, w_032_1658, w_032_1659, w_032_1660, w_032_1662, w_032_1663, w_032_1665, w_032_1666, w_032_1667, w_032_1668, w_032_1669, w_032_1670, w_032_1672, w_032_1673, w_032_1674, w_032_1675, w_032_1676, w_032_1678, w_032_1680, w_032_1681, w_032_1683, w_032_1685, w_032_1687, w_032_1689, w_032_1690, w_032_1691, w_032_1692, w_032_1693, w_032_1695, w_032_1697, w_032_1698, w_032_1700, w_032_1702, w_032_1703, w_032_1704, w_032_1705, w_032_1706, w_032_1707, w_032_1708, w_032_1710, w_032_1711, w_032_1712, w_032_1713, w_032_1714, w_032_1715, w_032_1716, w_032_1717, w_032_1718, w_032_1719, w_032_1720, w_032_1721, w_032_1724, w_032_1725, w_032_1726, w_032_1727, w_032_1728, w_032_1729, w_032_1731, w_032_1732, w_032_1733, w_032_1734, w_032_1736, w_032_1737, w_032_1738, w_032_1739, w_032_1740, w_032_1741, w_032_1742, w_032_1743, w_032_1744, w_032_1745, w_032_1748, w_032_1749, w_032_1750, w_032_1751, w_032_1752, w_032_1754, w_032_1755, w_032_1756, w_032_1757, w_032_1758, w_032_1759, w_032_1760, w_032_1762, w_032_1763, w_032_1764, w_032_1766, w_032_1767, w_032_1768, w_032_1769, w_032_1770, w_032_1771, w_032_1772, w_032_1773, w_032_1774, w_032_1775, w_032_1776, w_032_1777, w_032_1778, w_032_1781, w_032_1783, w_032_1784, w_032_1785, w_032_1786, w_032_1787, w_032_1788, w_032_1789, w_032_1790, w_032_1791, w_032_1792, w_032_1793, w_032_1794, w_032_1795, w_032_1796, w_032_1797, w_032_1798, w_032_1799, w_032_1800, w_032_1801, w_032_1802, w_032_1804, w_032_1805, w_032_1806, w_032_1807, w_032_1808, w_032_1810, w_032_1812, w_032_1813, w_032_1814, w_032_1817, w_032_1818, w_032_1819, w_032_1820, w_032_1822, w_032_1823, w_032_1824, w_032_1825, w_032_1826, w_032_1827, w_032_1828, w_032_1829, w_032_1830, w_032_1831, w_032_1833, w_032_1834, w_032_1835, w_032_1836, w_032_1837, w_032_1838, w_032_1839, w_032_1841, w_032_1842, w_032_1843, w_032_1844, w_032_1845, w_032_1846, w_032_1847, w_032_1848, w_032_1851, w_032_1852, w_032_1853, w_032_1855, w_032_1856, w_032_1857, w_032_1858, w_032_1859, w_032_1860, w_032_1861, w_032_1862, w_032_1865, w_032_1866, w_032_1868, w_032_1869, w_032_1870, w_032_1871, w_032_1872, w_032_1873, w_032_1874, w_032_1877, w_032_1879, w_032_1881, w_032_1882, w_032_1883, w_032_1884, w_032_1886, w_032_1888, w_032_1889, w_032_1890, w_032_1891, w_032_1892, w_032_1893, w_032_1894, w_032_1895, w_032_1896, w_032_1897, w_032_1898, w_032_1899, w_032_1901, w_032_1902, w_032_1903, w_032_1904, w_032_1905, w_032_1907, w_032_1908, w_032_1909, w_032_1911, w_032_1912, w_032_1913, w_032_1915, w_032_1916, w_032_1917, w_032_1918, w_032_1920, w_032_1922, w_032_1923, w_032_1924, w_032_1925, w_032_1926, w_032_1927, w_032_1928, w_032_1929, w_032_1930, w_032_1931, w_032_1932, w_032_1933, w_032_1934, w_032_1936, w_032_1937, w_032_1939, w_032_1942, w_032_1943, w_032_1945, w_032_1946, w_032_1948, w_032_1950, w_032_1951, w_032_1952, w_032_1953, w_032_1954, w_032_1955, w_032_1957, w_032_1958, w_032_1959, w_032_1960, w_032_1961, w_032_1962, w_032_1964, w_032_1965, w_032_1966, w_032_1967, w_032_1968, w_032_1969, w_032_1970, w_032_1971, w_032_1972, w_032_1973, w_032_1974, w_032_1976, w_032_1977, w_032_1978, w_032_1979, w_032_1980, w_032_1981, w_032_1982, w_032_1983, w_032_1984, w_032_1985, w_032_1986, w_032_1987, w_032_1988, w_032_1990, w_032_1991, w_032_1992, w_032_1993, w_032_1994, w_032_1995, w_032_1996, w_032_1997, w_032_1998, w_032_1999, w_032_2000, w_032_2001, w_032_2002, w_032_2003, w_032_2004, w_032_2006, w_032_2008, w_032_2009, w_032_2010, w_032_2012, w_032_2013, w_032_2014, w_032_2016, w_032_2017, w_032_2018, w_032_2019, w_032_2020, w_032_2021, w_032_2022, w_032_2023, w_032_2025, w_032_2026, w_032_2027, w_032_2028, w_032_2029, w_032_2030, w_032_2032, w_032_2033, w_032_2034, w_032_2036, w_032_2038, w_032_2039, w_032_2040, w_032_2041, w_032_2042, w_032_2043, w_032_2044, w_032_2046, w_032_2047, w_032_2048, w_032_2049, w_032_2050, w_032_2051, w_032_2053, w_032_2054, w_032_2056, w_032_2057, w_032_2058, w_032_2060, w_032_2061, w_032_2062, w_032_2063, w_032_2064, w_032_2066, w_032_2068, w_032_2072, w_032_2074, w_032_2075, w_032_2076, w_032_2077, w_032_2080, w_032_2081, w_032_2082, w_032_2085, w_032_2086, w_032_2087, w_032_2088, w_032_2090, w_032_2092, w_032_2093, w_032_2094, w_032_2095, w_032_2096, w_032_2097, w_032_2098, w_032_2099, w_032_2100, w_032_2102, w_032_2103, w_032_2104, w_032_2105, w_032_2106, w_032_2107, w_032_2108, w_032_2111, w_032_2112, w_032_2113, w_032_2114, w_032_2115, w_032_2116, w_032_2118, w_032_2120, w_032_2121, w_032_2122, w_032_2124, w_032_2125, w_032_2126, w_032_2127, w_032_2128, w_032_2132, w_032_2133, w_032_2134, w_032_2136, w_032_2137, w_032_2138, w_032_2139, w_032_2140, w_032_2141, w_032_2142, w_032_2144, w_032_2145, w_032_2146, w_032_2147, w_032_2148, w_032_2149, w_032_2150, w_032_2152, w_032_2153, w_032_2154, w_032_2155, w_032_2156, w_032_2157, w_032_2158, w_032_2159, w_032_2160, w_032_2161, w_032_2162, w_032_2163, w_032_2164, w_032_2165, w_032_2166, w_032_2167, w_032_2168, w_032_2170, w_032_2171, w_032_2172, w_032_2173, w_032_2175, w_032_2176, w_032_2177, w_032_2178, w_032_2179, w_032_2180, w_032_2181, w_032_2182, w_032_2183, w_032_2184, w_032_2186, w_032_2187, w_032_2188, w_032_2189, w_032_2190, w_032_2191, w_032_2192, w_032_2193, w_032_2194, w_032_2195, w_032_2198, w_032_2199, w_032_2200, w_032_2201, w_032_2202, w_032_2203, w_032_2204, w_032_2205, w_032_2206, w_032_2207, w_032_2208, w_032_2209, w_032_2210, w_032_2211, w_032_2212, w_032_2213, w_032_2214, w_032_2215, w_032_2217, w_032_2218, w_032_2219, w_032_2220, w_032_2221, w_032_2223, w_032_2224, w_032_2225, w_032_2226, w_032_2227, w_032_2228, w_032_2229, w_032_2230, w_032_2231, w_032_2232, w_032_2233, w_032_2234, w_032_2235, w_032_2237, w_032_2238, w_032_2239, w_032_2240, w_032_2241, w_032_2242, w_032_2245, w_032_2246, w_032_2247, w_032_2248, w_032_2251, w_032_2252, w_032_2253, w_032_2254, w_032_2256, w_032_2257, w_032_2258, w_032_2260, w_032_2261, w_032_2263, w_032_2264, w_032_2266, w_032_2267, w_032_2268, w_032_2269, w_032_2273, w_032_2274, w_032_2275, w_032_2276, w_032_2277, w_032_2278, w_032_2279, w_032_2281, w_032_2283, w_032_2284, w_032_2286, w_032_2289, w_032_2290, w_032_2291, w_032_2292, w_032_2293, w_032_2294, w_032_2295, w_032_2296, w_032_2297, w_032_2298, w_032_2299, w_032_2300, w_032_2301, w_032_2302, w_032_2303, w_032_2305, w_032_2306, w_032_2307, w_032_2308, w_032_2309, w_032_2311, w_032_2312, w_032_2314, w_032_2315, w_032_2316, w_032_2318, w_032_2320, w_032_2321, w_032_2322, w_032_2323, w_032_2324, w_032_2325, w_032_2326, w_032_2327, w_032_2329, w_032_2330, w_032_2332, w_032_2333, w_032_2334, w_032_2335, w_032_2336, w_032_2337, w_032_2338, w_032_2340, w_032_2342, w_032_2343, w_032_2345, w_032_2346, w_032_2347, w_032_2348, w_032_2349, w_032_2350, w_032_2351, w_032_2352, w_032_2353, w_032_2354, w_032_2355, w_032_2356, w_032_2357, w_032_2358, w_032_2359, w_032_2360, w_032_2361, w_032_2362, w_032_2363, w_032_2364, w_032_2365, w_032_2366, w_032_2367, w_032_2368, w_032_2369, w_032_2370, w_032_2371, w_032_2373, w_032_2375, w_032_2376, w_032_2377, w_032_2378, w_032_2379, w_032_2380, w_032_2381, w_032_2382, w_032_2384, w_032_2385, w_032_2386, w_032_2387, w_032_2388, w_032_2389, w_032_2391, w_032_2392, w_032_2394, w_032_2395, w_032_2396, w_032_2399, w_032_2400, w_032_2401, w_032_2403, w_032_2404, w_032_2405, w_032_2406, w_032_2407, w_032_2408, w_032_2409, w_032_2410, w_032_2411, w_032_2412, w_032_2413, w_032_2414, w_032_2415, w_032_2416, w_032_2417, w_032_2418, w_032_2419, w_032_2420, w_032_2423, w_032_2424, w_032_2426, w_032_2427, w_032_2428, w_032_2430, w_032_2431, w_032_2434, w_032_2435, w_032_2436, w_032_2438, w_032_2439, w_032_2440, w_032_2441, w_032_2446, w_032_2447, w_032_2449, w_032_2450, w_032_2451, w_032_2452, w_032_2453, w_032_2455, w_032_2456, w_032_2457, w_032_2458, w_032_2459, w_032_2460, w_032_2461, w_032_2462, w_032_2463, w_032_2464, w_032_2466, w_032_2467, w_032_2468, w_032_2469, w_032_2470, w_032_2471, w_032_2473, w_032_2474, w_032_2475, w_032_2478, w_032_2479, w_032_2480, w_032_2481, w_032_2482, w_032_2483, w_032_2484, w_032_2485, w_032_2486, w_032_2487, w_032_2488, w_032_2490, w_032_2492, w_032_2493, w_032_2494, w_032_2495, w_032_2496, w_032_2499, w_032_2500, w_032_2501, w_032_2502, w_032_2503, w_032_2504, w_032_2505, w_032_2506, w_032_2507, w_032_2508, w_032_2509, w_032_2510, w_032_2511, w_032_2514, w_032_2515, w_032_2516, w_032_2517, w_032_2518, w_032_2519, w_032_2520, w_032_2522, w_032_2523, w_032_2524, w_032_2525, w_032_2527, w_032_2531, w_032_2532, w_032_2533, w_032_2534, w_032_2537, w_032_2539, w_032_2540, w_032_2541, w_032_2542, w_032_2543, w_032_2545, w_032_2546, w_032_2547, w_032_2548, w_032_2549, w_032_2550, w_032_2551, w_032_2552, w_032_2553, w_032_2554, w_032_2555, w_032_2556, w_032_2560, w_032_2562, w_032_2563, w_032_2564, w_032_2566, w_032_2567, w_032_2569, w_032_2570, w_032_2571, w_032_2572, w_032_2573, w_032_2574, w_032_2575, w_032_2577, w_032_2578, w_032_2579, w_032_2580, w_032_2581, w_032_2582, w_032_2585, w_032_2586, w_032_2587, w_032_2589, w_032_2593, w_032_2594, w_032_2595, w_032_2596, w_032_2598, w_032_2599, w_032_2600, w_032_2601, w_032_2602, w_032_2603, w_032_2606, w_032_2607, w_032_2608, w_032_2609, w_032_2611, w_032_2613, w_032_2614, w_032_2615, w_032_2618, w_032_2619, w_032_2621, w_032_2622, w_032_2625, w_032_2626, w_032_2627, w_032_2628, w_032_2630, w_032_2631, w_032_2632, w_032_2633, w_032_2635, w_032_2636, w_032_2637, w_032_2638, w_032_2640, w_032_2641, w_032_2642, w_032_2643, w_032_2644, w_032_2646, w_032_2647, w_032_2648, w_032_2649, w_032_2650, w_032_2651, w_032_2652, w_032_2653, w_032_2655, w_032_2656, w_032_2657, w_032_2659, w_032_2660, w_032_2661, w_032_2662, w_032_2663, w_032_2665, w_032_2666, w_032_2669, w_032_2671, w_032_2672, w_032_2674, w_032_2675, w_032_2676, w_032_2678, w_032_2679, w_032_2681, w_032_2682, w_032_2683, w_032_2686, w_032_2687, w_032_2689, w_032_2690, w_032_2691, w_032_2692, w_032_2693, w_032_2694, w_032_2695, w_032_2696, w_032_2698, w_032_2699, w_032_2700, w_032_2701, w_032_2702, w_032_2703, w_032_2705, w_032_2706, w_032_2707, w_032_2708, w_032_2709, w_032_2710, w_032_2711, w_032_2713, w_032_2714, w_032_2715, w_032_2716, w_032_2718, w_032_2719, w_032_2721, w_032_2722, w_032_2723, w_032_2724, w_032_2727, w_032_2728, w_032_2729, w_032_2730, w_032_2732, w_032_2733, w_032_2734, w_032_2735, w_032_2736, w_032_2738, w_032_2739, w_032_2740, w_032_2742, w_032_2743, w_032_2745, w_032_2746, w_032_2747, w_032_2749, w_032_2751, w_032_2752, w_032_2753, w_032_2754, w_032_2755, w_032_2756, w_032_2757, w_032_2758, w_032_2759, w_032_2760, w_032_2761, w_032_2762, w_032_2763, w_032_2764, w_032_2765, w_032_2766, w_032_2767, w_032_2768, w_032_2769, w_032_2770, w_032_2771, w_032_2772, w_032_2773, w_032_2774, w_032_2775, w_032_2776, w_032_2778, w_032_2779, w_032_2780, w_032_2781, w_032_2783, w_032_2784, w_032_2786, w_032_2787, w_032_2788, w_032_2789, w_032_2790, w_032_2791, w_032_2792, w_032_2793, w_032_2795, w_032_2796, w_032_2798, w_032_2800, w_032_2802, w_032_2806, w_032_2807, w_032_2808, w_032_2810, w_032_2812, w_032_2813, w_032_2814, w_032_2815, w_032_2817, w_032_2818, w_032_2823, w_032_2824, w_032_2825, w_032_2826, w_032_2827, w_032_2830, w_032_2832, w_032_2833, w_032_2834, w_032_2835, w_032_2836, w_032_2838, w_032_2839, w_032_2840, w_032_2842, w_032_2843, w_032_2844, w_032_2845, w_032_2846, w_032_2847, w_032_2848, w_032_2849, w_032_2851, w_032_2852, w_032_2853, w_032_2854, w_032_2855, w_032_2856, w_032_2858, w_032_2859, w_032_2860, w_032_2861, w_032_2863, w_032_2864, w_032_2865, w_032_2866, w_032_2867, w_032_2868, w_032_2869, w_032_2870, w_032_2872, w_032_2873, w_032_2874, w_032_2875, w_032_2876, w_032_2877, w_032_2878, w_032_2879, w_032_2880, w_032_2881, w_032_2882, w_032_2884, w_032_2885, w_032_2886, w_032_2887, w_032_2888, w_032_2889, w_032_2890, w_032_2891, w_032_2892, w_032_2893, w_032_2894, w_032_2895, w_032_2896, w_032_2897, w_032_2899, w_032_2901, w_032_2902, w_032_2903, w_032_2904, w_032_2905, w_032_2906, w_032_2907, w_032_2908, w_032_2909, w_032_2911, w_032_2912, w_032_2913, w_032_2914, w_032_2915, w_032_2916, w_032_2917, w_032_2919, w_032_2920, w_032_2922, w_032_2923, w_032_2924, w_032_2926, w_032_2927, w_032_2928, w_032_2930, w_032_2931, w_032_2932, w_032_2934, w_032_2935, w_032_2937, w_032_2938, w_032_2939, w_032_2940, w_032_2942, w_032_2943, w_032_2944, w_032_2945, w_032_2946, w_032_2947, w_032_2948, w_032_2949, w_032_2950, w_032_2951, w_032_2952, w_032_2953, w_032_2954, w_032_2955, w_032_2956, w_032_2957, w_032_2958, w_032_2959, w_032_2960, w_032_2961, w_032_2963, w_032_2965, w_032_2966, w_032_2967, w_032_2968, w_032_2970, w_032_2971, w_032_2972, w_032_2974, w_032_2975, w_032_2976, w_032_2977, w_032_2978, w_032_2979, w_032_2980, w_032_2982, w_032_2985, w_032_2986, w_032_2988, w_032_2989, w_032_2990, w_032_2994, w_032_2996, w_032_2997, w_032_2998, w_032_3001, w_032_3002, w_032_3003, w_032_3004, w_032_3006, w_032_3007, w_032_3008, w_032_3010, w_032_3011, w_032_3013, w_032_3014, w_032_3015, w_032_3016, w_032_3017, w_032_3018, w_032_3019, w_032_3020, w_032_3022, w_032_3023, w_032_3024, w_032_3025, w_032_3026, w_032_3027, w_032_3030, w_032_3031, w_032_3032, w_032_3033, w_032_3035, w_032_3036, w_032_3039, w_032_3040, w_032_3041, w_032_3042, w_032_3043, w_032_3044, w_032_3045, w_032_3046, w_032_3047, w_032_3048, w_032_3050, w_032_3051, w_032_3052, w_032_3053, w_032_3054, w_032_3055, w_032_3056, w_032_3057, w_032_3059, w_032_3060, w_032_3061, w_032_3062, w_032_3063, w_032_3064, w_032_3065, w_032_3067, w_032_3068, w_032_3069, w_032_3070, w_032_3071, w_032_3072, w_032_3073, w_032_3074, w_032_3075, w_032_3076, w_032_3077, w_032_3078, w_032_3079, w_032_3081, w_032_3082, w_032_3083, w_032_3085, w_032_3086, w_032_3089, w_032_3090, w_032_3092, w_032_3094, w_032_3095, w_032_3096, w_032_3097, w_032_3098, w_032_3100, w_032_3103, w_032_3104, w_032_3105, w_032_3106, w_032_3107, w_032_3108, w_032_3109, w_032_3110, w_032_3111, w_032_3112, w_032_3113, w_032_3114, w_032_3115, w_032_3117, w_032_3118, w_032_3119, w_032_3120, w_032_3121, w_032_3122, w_032_3123, w_032_3124, w_032_3125, w_032_3126, w_032_3127, w_032_3128, w_032_3129, w_032_3130, w_032_3131, w_032_3132, w_032_3135, w_032_3138, w_032_3139, w_032_3140, w_032_3142, w_032_3143, w_032_3146, w_032_3147, w_032_3149, w_032_3151, w_032_3152, w_032_3153, w_032_3154, w_032_3157, w_032_3159, w_032_3160, w_032_3161, w_032_3162, w_032_3163, w_032_3164, w_032_3165, w_032_3166, w_032_3170, w_032_3172, w_032_3173, w_032_3174, w_032_3176, w_032_3177, w_032_3178, w_032_3181, w_032_3182, w_032_3186, w_032_3187, w_032_3190, w_032_3191, w_032_3192, w_032_3193, w_032_3194, w_032_3195, w_032_3197, w_032_3198, w_032_3199, w_032_3200, w_032_3201, w_032_3202, w_032_3203, w_032_3204, w_032_3205, w_032_3207, w_032_3208, w_032_3210, w_032_3211, w_032_3212, w_032_3213, w_032_3214, w_032_3215, w_032_3216, w_032_3217, w_032_3218, w_032_3219, w_032_3220, w_032_3221, w_032_3223, w_032_3224, w_032_3225, w_032_3227, w_032_3228, w_032_3229, w_032_3231, w_032_3232, w_032_3233, w_032_3235, w_032_3236, w_032_3237, w_032_3238, w_032_3241, w_032_3245, w_032_3248, w_032_3249, w_032_3251, w_032_3252, w_032_3253, w_032_3254, w_032_3255, w_032_3258, w_032_3259, w_032_3260, w_032_3261, w_032_3262, w_032_3263, w_032_3264, w_032_3265, w_032_3277, w_032_3278, w_032_3279, w_032_3280, w_032_3284, w_032_3285, w_032_3287, w_032_3289, w_032_3293, w_032_3297, w_032_3298, w_032_3299, w_032_3300, w_032_3301, w_032_3302, w_032_3303, w_032_3304, w_032_3308, w_032_3312, w_032_3313, w_032_3314, w_032_3315, w_032_3316, w_032_3317, w_032_3318, w_032_3321, w_032_3325, w_032_3327, w_032_3328, w_032_3330, w_032_3332, w_032_3335, w_032_3336, w_032_3339, w_032_3340, w_032_3341, w_032_3345, w_032_3347, w_032_3349, w_032_3350, w_032_3352, w_032_3353, w_032_3354, w_032_3356, w_032_3357, w_032_3358, w_032_3362, w_032_3364, w_032_3366, w_032_3369, w_032_3370, w_032_3371, w_032_3372, w_032_3374, w_032_3377, w_032_3381, w_032_3389, w_032_3390, w_032_3391, w_032_3392, w_032_3393, w_032_3394, w_032_3397, w_032_3398, w_032_3400, w_032_3402, w_032_3403, w_032_3404, w_032_3405, w_032_3406, w_032_3407, w_032_3408, w_032_3414, w_032_3416, w_032_3419, w_032_3420, w_032_3422, w_032_3425, w_032_3426, w_032_3427, w_032_3429, w_032_3430, w_032_3432, w_032_3436, w_032_3437, w_032_3438, w_032_3440, w_032_3443, w_032_3446, w_032_3447, w_032_3450, w_032_3453, w_032_3456, w_032_3458, w_032_3460, w_032_3461, w_032_3462, w_032_3463, w_032_3464, w_032_3465, w_032_3466, w_032_3467, w_032_3468, w_032_3470, w_032_3471, w_032_3473, w_032_3474, w_032_3475, w_032_3477, w_032_3478, w_032_3483, w_032_3487, w_032_3488, w_032_3489, w_032_3490, w_032_3492, w_032_3497, w_032_3500, w_032_3501, w_032_3503, w_032_3505, w_032_3507, w_032_3509, w_032_3514, w_032_3516, w_032_3518, w_032_3520, w_032_3521, w_032_3522, w_032_3524, w_032_3525, w_032_3527, w_032_3528, w_032_3529, w_032_3532, w_032_3533, w_032_3534, w_032_3535, w_032_3536, w_032_3537, w_032_3539, w_032_3540, w_032_3543, w_032_3544, w_032_3545, w_032_3549, w_032_3550, w_032_3554, w_032_3557, w_032_3558, w_032_3560, w_032_3564, w_032_3565, w_032_3567, w_032_3570, w_032_3571, w_032_3574, w_032_3575, w_032_3576, w_032_3577, w_032_3578, w_032_3579, w_032_3580, w_032_3582, w_032_3589, w_032_3590, w_032_3591, w_032_3592, w_032_3593, w_032_3594, w_032_3595, w_032_3596, w_032_3598, w_032_3603, w_032_3604, w_032_3606, w_032_3609, w_032_3610, w_032_3613, w_032_3615, w_032_3616, w_032_3620, w_032_3623, w_032_3624, w_032_3625, w_032_3626, w_032_3628, w_032_3632, w_032_3633, w_032_3634, w_032_3635, w_032_3636, w_032_3639, w_032_3644, w_032_3645, w_032_3652, w_032_3653, w_032_3654, w_032_3655, w_032_3656, w_032_3659, w_032_3660, w_032_3661, w_032_3662, w_032_3665, w_032_3666, w_032_3667, w_032_3672, w_032_3673, w_032_3674, w_032_3677, w_032_3678, w_032_3680, w_032_3681, w_032_3683, w_032_3684, w_032_3685, w_032_3687, w_032_3690, w_032_3692, w_032_3693, w_032_3695, w_032_3700, w_032_3705, w_032_3706, w_032_3709, w_032_3710, w_032_3711, w_032_3712, w_032_3714, w_032_3715, w_032_3717, w_032_3718, w_032_3721, w_032_3724, w_032_3726, w_032_3729, w_032_3731, w_032_3732, w_032_3733, w_032_3736, w_032_3737, w_032_3739, w_032_3742, w_032_3743, w_032_3746, w_032_3749, w_032_3751, w_032_3757, w_032_3758, w_032_3759, w_032_3760, w_032_3762, w_032_3766, w_032_3767, w_032_3768, w_032_3769, w_032_3773, w_032_3774, w_032_3776, w_032_3778, w_032_3779, w_032_3780, w_032_3781, w_032_3784, w_032_3785, w_032_3786, w_032_3787, w_032_3788, w_032_3790, w_032_3795, w_032_3800, w_032_3801, w_032_3802, w_032_3805, w_032_3806, w_032_3807, w_032_3808, w_032_3809, w_032_3813, w_032_3814, w_032_3818, w_032_3822, w_032_3824, w_032_3825, w_032_3829, w_032_3832, w_032_3833, w_032_3836, w_032_3837, w_032_3838, w_032_3841, w_032_3842, w_032_3843, w_032_3850, w_032_3852, w_032_3854, w_032_3855, w_032_3858, w_032_3865, w_032_3866, w_032_3867, w_032_3868, w_032_3870, w_032_3871, w_032_3872, w_032_3873, w_032_3875, w_032_3877, w_032_3878, w_032_3879, w_032_3881, w_032_3882, w_032_3883, w_032_3886, w_032_3889, w_032_3894, w_032_3897, w_032_3898, w_032_3899, w_032_3900, w_032_3901, w_032_3902, w_032_3903, w_032_3904, w_032_3905, w_032_3908, w_032_3909, w_032_3911, w_032_3912, w_032_3913, w_032_3917, w_032_3920, w_032_3924, w_032_3929, w_032_3930, w_032_3934, w_032_3935, w_032_3936, w_032_3938, w_032_3939, w_032_3943, w_032_3945, w_032_3948, w_032_3949, w_032_3950, w_032_3951, w_032_3953, w_032_3960, w_032_3961, w_032_3962, w_032_3963, w_032_3964, w_032_3966, w_032_3967, w_032_3969, w_032_3970, w_032_3971, w_032_3972, w_032_3975, w_032_3976, w_032_3977, w_032_3979, w_032_3981, w_032_3982, w_032_3984, w_032_3985, w_032_3986, w_032_3988, w_032_3989, w_032_3994, w_032_3995, w_032_3997, w_032_3998, w_032_4000, w_032_4001, w_032_4003, w_032_4004, w_032_4006, w_032_4008, w_032_4009, w_032_4010, w_032_4011, w_032_4012, w_032_4015, w_032_4017, w_032_4019, w_032_4020, w_032_4021, w_032_4022, w_032_4024, w_032_4025, w_032_4026, w_032_4030, w_032_4033, w_032_4035, w_032_4036, w_032_4038, w_032_4039, w_032_4040, w_032_4041, w_032_4042, w_032_4043, w_032_4044, w_032_4046, w_032_4047, w_032_4048, w_032_4049, w_032_4050, w_032_4056, w_032_4057, w_032_4058, w_032_4059, w_032_4060, w_032_4062, w_032_4063, w_032_4064, w_032_4070, w_032_4072, w_032_4073, w_032_4074, w_032_4076, w_032_4078, w_032_4080, w_032_4081, w_032_4087, w_032_4089, w_032_4090, w_032_4092, w_032_4093, w_032_4094, w_032_4097, w_032_4099, w_032_4102, w_032_4103, w_032_4106, w_032_4107, w_032_4108, w_032_4109, w_032_4111, w_032_4113, w_032_4114, w_032_4116, w_032_4117, w_032_4119, w_032_4121, w_032_4122, w_032_4123, w_032_4126, w_032_4133, w_032_4134, w_032_4136, w_032_4137, w_032_4139, w_032_4141, w_032_4143, w_032_4150, w_032_4151, w_032_4153, w_032_4156, w_032_4159, w_032_4160, w_032_4163, w_032_4164, w_032_4166, w_032_4168, w_032_4169, w_032_4171, w_032_4172, w_032_4173, w_032_4174, w_032_4175, w_032_4176, w_032_4177, w_032_4178, w_032_4179, w_032_4180, w_032_4183, w_032_4185, w_032_4186, w_032_4187, w_032_4188, w_032_4192, w_032_4196, w_032_4197, w_032_4199, w_032_4200, w_032_4201, w_032_4202, w_032_4203, w_032_4209, w_032_4210, w_032_4221, w_032_4223, w_032_4225, w_032_4227, w_032_4228, w_032_4229, w_032_4230, w_032_4232, w_032_4233, w_032_4238, w_032_4240, w_032_4241, w_032_4242, w_032_4243, w_032_4246, w_032_4250, w_032_4251, w_032_4252, w_032_4254, w_032_4257, w_032_4258, w_032_4259, w_032_4260, w_032_4261, w_032_4262, w_032_4263, w_032_4264, w_032_4265, w_032_4267, w_032_4270, w_032_4274, w_032_4276, w_032_4277, w_032_4278, w_032_4279, w_032_4280, w_032_4282, w_032_4285, w_032_4290, w_032_4293, w_032_4294, w_032_4297, w_032_4299, w_032_4300, w_032_4301, w_032_4304, w_032_4306, w_032_4307, w_032_4309, w_032_4314, w_032_4315, w_032_4317, w_032_4321, w_032_4323, w_032_4327, w_032_4328, w_032_4329, w_032_4330, w_032_4331, w_032_4335, w_032_4336, w_032_4338, w_032_4339, w_032_4345, w_032_4347, w_032_4348, w_032_4350, w_032_4352, w_032_4354, w_032_4358, w_032_4360, w_032_4361, w_032_4363, w_032_4370, w_032_4371, w_032_4374, w_032_4376, w_032_4378, w_032_4380, w_032_4382, w_032_4387, w_032_4389, w_032_4393, w_032_4394, w_032_4396, w_032_4398, w_032_4399, w_032_4400, w_032_4401, w_032_4402, w_032_4403, w_032_4406, w_032_4407, w_032_4409, w_032_4410, w_032_4412, w_032_4417, w_032_4420, w_032_4421, w_032_4422, w_032_4424, w_032_4425, w_032_4427, w_032_4429, w_032_4432, w_032_4433, w_032_4434, w_032_4435, w_032_4438, w_032_4439, w_032_4442, w_032_4443, w_032_4444, w_032_4445, w_032_4447, w_032_4450, w_032_4452, w_032_4453, w_032_4454, w_032_4455, w_032_4457, w_032_4459, w_032_4460, w_032_4461, w_032_4462, w_032_4463, w_032_4467, w_032_4470, w_032_4471, w_032_4472, w_032_4473, w_032_4474, w_032_4477, w_032_4478, w_032_4482, w_032_4483, w_032_4485, w_032_4486, w_032_4489, w_032_4490, w_032_4491, w_032_4494, w_032_4495, w_032_4497, w_032_4499, w_032_4500, w_032_4504, w_032_4506, w_032_4507, w_032_4512, w_032_4513, w_032_4514, w_032_4515, w_032_4516, w_032_4517, w_032_4518, w_032_4519, w_032_4522, w_032_4524, w_032_4525, w_032_4526, w_032_4528, w_032_4530, w_032_4532, w_032_4534, w_032_4536, w_032_4537, w_032_4538, w_032_4539, w_032_4540, w_032_4541, w_032_4545, w_032_4549, w_032_4551, w_032_4555, w_032_4556, w_032_4558, w_032_4559, w_032_4560, w_032_4563, w_032_4564, w_032_4568, w_032_4569, w_032_4571, w_032_4572, w_032_4573, w_032_4575, w_032_4578, w_032_4579, w_032_4581, w_032_4582, w_032_4584, w_032_4585, w_032_4586, w_032_4587, w_032_4588, w_032_4589, w_032_4590, w_032_4591, w_032_4594, w_032_4596, w_032_4597, w_032_4598, w_032_4601, w_032_4602, w_032_4604, w_032_4607, w_032_4608, w_032_4609, w_032_4610, w_032_4612, w_032_4613, w_032_4614, w_032_4615, w_032_4616, w_032_4617, w_032_4618, w_032_4619, w_032_4620, w_032_4621, w_032_4622, w_032_4625, w_032_4627, w_032_4629, w_032_4630, w_032_4631, w_032_4633, w_032_4634, w_032_4636, w_032_4640, w_032_4641, w_032_4642, w_032_4643, w_032_4645, w_032_4646, w_032_4647, w_032_4648, w_032_4649, w_032_4651, w_032_4654, w_032_4657, w_032_4663, w_032_4668, w_032_4670, w_032_4673, w_032_4677, w_032_4679, w_032_4680, w_032_4682, w_032_4684, w_032_4685, w_032_4687, w_032_4688, w_032_4689, w_032_4690, w_032_4691, w_032_4692, w_032_4696, w_032_4697, w_032_4699, w_032_4700, w_032_4702, w_032_4703, w_032_4704, w_032_4707, w_032_4709, w_032_4710, w_032_4712, w_032_4713, w_032_4715, w_032_4717, w_032_4718, w_032_4719, w_032_4720, w_032_4722, w_032_4726, w_032_4733, w_032_4734, w_032_4735, w_032_4739, w_032_4740, w_032_4741, w_032_4742, w_032_4745, w_032_4746, w_032_4749, w_032_4750, w_032_4751, w_032_4753, w_032_4756, w_032_4760, w_032_4762, w_032_4763, w_032_4765, w_032_4767, w_032_4768, w_032_4769, w_032_4770, w_032_4772, w_032_4773, w_032_4776, w_032_4779, w_032_4781, w_032_4784, w_032_4787, w_032_4792, w_032_4794, w_032_4795, w_032_4799, w_032_4803, w_032_4804, w_032_4806, w_032_4807, w_032_4809, w_032_4810, w_032_4811, w_032_4815, w_032_4817, w_032_4818, w_032_4819, w_032_4823, w_032_4824, w_032_4825, w_032_4828, w_032_4829, w_032_4837, w_032_4838, w_032_4840, w_032_4841, w_032_4842, w_032_4843, w_032_4845, w_032_4846, w_032_4847, w_032_4849, w_032_4850, w_032_4853, w_032_4854, w_032_4856, w_032_4857, w_032_4861, w_032_4863, w_032_4865, w_032_4866, w_032_4868, w_032_4869, w_032_4870, w_032_4874, w_032_4875, w_032_4876, w_032_4877, w_032_4879, w_032_4881, w_032_4882, w_032_4883, w_032_4884, w_032_4886, w_032_4887, w_032_4888, w_032_4891, w_032_4892, w_032_4894, w_032_4896, w_032_4898, w_032_4902, w_032_4904, w_032_4906, w_032_4907, w_032_4908, w_032_4909, w_032_4910, w_032_4912, w_032_4913, w_032_4914, w_032_4915, w_032_4916, w_032_4917, w_032_4918, w_032_4921, w_032_4922, w_032_4924, w_032_4926, w_032_4929, w_032_4930, w_032_4931, w_032_4932, w_032_4933, w_032_4935, w_032_4936, w_032_4937, w_032_4938, w_032_4941, w_032_4942, w_032_4944, w_032_4945, w_032_4947, w_032_4949, w_032_4950, w_032_4952, w_032_4954, w_032_4955, w_032_4957, w_032_4959, w_032_4960, w_032_4964, w_032_4965, w_032_4968, w_032_4969, w_032_4972, w_032_4974, w_032_4980, w_032_4984, w_032_4985, w_032_4986, w_032_4987, w_032_4990, w_032_4995, w_032_4996, w_032_5000, w_032_5001, w_032_5002, w_032_5004, w_032_5005, w_032_5006, w_032_5007, w_032_5010, w_032_5011, w_032_5012, w_032_5014, w_032_5015, w_032_5018, w_032_5021, w_032_5022, w_032_5023, w_032_5026, w_032_5027, w_032_5028, w_032_5029, w_032_5031, w_032_5032, w_032_5034, w_032_5036, w_032_5038, w_032_5042, w_032_5044, w_032_5045, w_032_5047, w_032_5051, w_032_5052, w_032_5056, w_032_5059, w_032_5060, w_032_5061, w_032_5062, w_032_5063, w_032_5064, w_032_5066, w_032_5067, w_032_5068, w_032_5070, w_032_5072, w_032_5077, w_032_5079, w_032_5080, w_032_5081, w_032_5082, w_032_5086, w_032_5087, w_032_5090, w_032_5091, w_032_5093, w_032_5094, w_032_5095, w_032_5096, w_032_5098, w_032_5101, w_032_5104, w_032_5108, w_032_5110, w_032_5111, w_032_5120, w_032_5123, w_032_5125, w_032_5127, w_032_5128, w_032_5130, w_032_5133, w_032_5134, w_032_5135, w_032_5136, w_032_5138, w_032_5142, w_032_5143, w_032_5145, w_032_5147, w_032_5148, w_032_5151, w_032_5152, w_032_5153, w_032_5154, w_032_5156, w_032_5157, w_032_5158, w_032_5161, w_032_5162, w_032_5164, w_032_5165, w_032_5170, w_032_5171, w_032_5173, w_032_5174, w_032_5178, w_032_5180, w_032_5183, w_032_5184, w_032_5188, w_032_5190, w_032_5191, w_032_5192, w_032_5196, w_032_5197, w_032_5198, w_032_5199, w_032_5202, w_032_5203, w_032_5204, w_032_5205, w_032_5207, w_032_5208, w_032_5210, w_032_5216, w_032_5217, w_032_5219, w_032_5220, w_032_5221, w_032_5222, w_032_5232, w_032_5233, w_032_5235, w_032_5236, w_032_5237, w_032_5246, w_032_5248, w_032_5251, w_032_5252, w_032_5253, w_032_5254, w_032_5257, w_032_5262, w_032_5264, w_032_5267, w_032_5268, w_032_5272, w_032_5276, w_032_5278, w_032_5279, w_032_5280, w_032_5281, w_032_5283, w_032_5284, w_032_5285, w_032_5286, w_032_5292, w_032_5293, w_032_5296, w_032_5297, w_032_5300, w_032_5301, w_032_5302, w_032_5303, w_032_5307, w_032_5309, w_032_5310, w_032_5311, w_032_5316, w_032_5317, w_032_5318, w_032_5319, w_032_5320, w_032_5322, w_032_5324, w_032_5325, w_032_5327, w_032_5328, w_032_5329, w_032_5335, w_032_5336, w_032_5338, w_032_5340, w_032_5341, w_032_5342, w_032_5343, w_032_5346, w_032_5348, w_032_5349, w_032_5351, w_032_5353, w_032_5354, w_032_5362, w_032_5363, w_032_5364, w_032_5366, w_032_5367, w_032_5368, w_032_5369, w_032_5370, w_032_5371, w_032_5373, w_032_5374, w_032_5376, w_032_5378, w_032_5379, w_032_5381, w_032_5382, w_032_5383, w_032_5385, w_032_5386, w_032_5387, w_032_5388, w_032_5389, w_032_5390, w_032_5392, w_032_5394, w_032_5396, w_032_5398, w_032_5400, w_032_5401, w_032_5402, w_032_5410, w_032_5411, w_032_5412, w_032_5414, w_032_5415, w_032_5417, w_032_5418, w_032_5419, w_032_5420, w_032_5422, w_032_5424, w_032_5425, w_032_5426, w_032_5429, w_032_5432, w_032_5433, w_032_5434, w_032_5437, w_032_5438, w_032_5439, w_032_5442, w_032_5443, w_032_5446, w_032_5447, w_032_5450, w_032_5452, w_032_5453, w_032_5454, w_032_5455, w_032_5456, w_032_5457, w_032_5458, w_032_5459, w_032_5460, w_032_5462, w_032_5463, w_032_5465, w_032_5467, w_032_5468, w_032_5469, w_032_5470, w_032_5472, w_032_5473, w_032_5477, w_032_5478, w_032_5480, w_032_5482, w_032_5484, w_032_5486, w_032_5488, w_032_5489, w_032_5492, w_032_5493, w_032_5494, w_032_5495, w_032_5496, w_032_5498, w_032_5499, w_032_5500, w_032_5502, w_032_5503, w_032_5506, w_032_5507, w_032_5510, w_032_5512, w_032_5513, w_032_5514, w_032_5515, w_032_5516, w_032_5524, w_032_5525, w_032_5526, w_032_5527, w_032_5528, w_032_5531, w_032_5532, w_032_5533, w_032_5535, w_032_5539, w_032_5540, w_032_5544, w_032_5545, w_032_5546, w_032_5549, w_032_5550, w_032_5551, w_032_5552, w_032_5553, w_032_5554, w_032_5556, w_032_5558, w_032_5560, w_032_5561, w_032_5566, w_032_5567, w_032_5571, w_032_5572, w_032_5576, w_032_5577, w_032_5578, w_032_5580, w_032_5583, w_032_5584, w_032_5585, w_032_5586, w_032_5588, w_032_5589, w_032_5592, w_032_5593, w_032_5596, w_032_5597, w_032_5598, w_032_5600, w_032_5601, w_032_5602, w_032_5603, w_032_5606, w_032_5609, w_032_5610, w_032_5612, w_032_5614, w_032_5616, w_032_5621, w_032_5623, w_032_5626, w_032_5632, w_032_5633, w_032_5635, w_032_5636, w_032_5638, w_032_5640, w_032_5641, w_032_5642, w_032_5644, w_032_5646, w_032_5647, w_032_5651, w_032_5653, w_032_5655, w_032_5656, w_032_5657, w_032_5660, w_032_5664, w_032_5667, w_032_5669, w_032_5670, w_032_5671, w_032_5672, w_032_5677, w_032_5679, w_032_5681, w_032_5683, w_032_5689, w_032_5690, w_032_5693, w_032_5694, w_032_5695, w_032_5697, w_032_5698, w_032_5699, w_032_5700, w_032_5702, w_032_5703, w_032_5704, w_032_5705, w_032_5706, w_032_5710, w_032_5712, w_032_5713, w_032_5714, w_032_5717, w_032_5719, w_032_5721, w_032_5724, w_032_5727, w_032_5728, w_032_5729, w_032_5731, w_032_5734, w_032_5737, w_032_5740, w_032_5741, w_032_5742, w_032_5743, w_032_5744, w_032_5747, w_032_5748, w_032_5752, w_032_5754, w_032_5755, w_032_5756, w_032_5757, w_032_5758, w_032_5759, w_032_5760, w_032_5761, w_032_5762, w_032_5764, w_032_5766, w_032_5767, w_032_5769, w_032_5771, w_032_5772, w_032_5773, w_032_5775, w_032_5776, w_032_5779, w_032_5781, w_032_5783, w_032_5786, w_032_5787, w_032_5788, w_032_5789, w_032_5791, w_032_5792, w_032_5793, w_032_5794, w_032_5795, w_032_5796, w_032_5797, w_032_5799, w_032_5800, w_032_5801, w_032_5802, w_032_5807, w_032_5808, w_032_5809, w_032_5810, w_032_5812, w_032_5815, w_032_5816, w_032_5819, w_032_5820, w_032_5822, w_032_5823, w_032_5824, w_032_5826, w_032_5828, w_032_5830, w_032_5831, w_032_5832, w_032_5833, w_032_5834, w_032_5837, w_032_5838, w_032_5840, w_032_5841, w_032_5843, w_032_5845, w_032_5847, w_032_5848, w_032_5851, w_032_5852, w_032_5855, w_032_5856, w_032_5857, w_032_5858, w_032_5860, w_032_5861, w_032_5863, w_032_5864, w_032_5865, w_032_5866, w_032_5867, w_032_5868, w_032_5869, w_032_5872, w_032_5876, w_032_5877, w_032_5879, w_032_5880, w_032_5882, w_032_5883, w_032_5884, w_032_5885, w_032_5890, w_032_5892, w_032_5893, w_032_5894, w_032_5895, w_032_5897, w_032_5901, w_032_5904, w_032_5905, w_032_5906, w_032_5912, w_032_5913, w_032_5914, w_032_5915, w_032_5916, w_032_5917, w_032_5919, w_032_5920, w_032_5921, w_032_5922, w_032_5923, w_032_5924, w_032_5926, w_032_5928, w_032_5929, w_032_5930, w_032_5931, w_032_5932, w_032_5935, w_032_5937, w_032_5939, w_032_5943, w_032_5944, w_032_5945, w_032_5946, w_032_5948, w_032_5949, w_032_5951, w_032_5952, w_032_5954, w_032_5955, w_032_5957, w_032_5958, w_032_5960, w_032_5961, w_032_5962, w_032_5966, w_032_5967, w_032_5968, w_032_5970, w_032_5971, w_032_5972, w_032_5974, w_032_5988, w_032_5990, w_032_5991, w_032_5992, w_032_5993, w_032_5996, w_032_5998, w_032_6000, w_032_6001, w_032_6002, w_032_6003, w_032_6005, w_032_6006, w_032_6007, w_032_6009, w_032_6010, w_032_6012, w_032_6013, w_032_6014, w_032_6017, w_032_6019, w_032_6020, w_032_6021, w_032_6022, w_032_6025, w_032_6026, w_032_6028, w_032_6029, w_032_6030, w_032_6031, w_032_6034, w_032_6035, w_032_6040, w_032_6042, w_032_6043, w_032_6045, w_032_6046, w_032_6047, w_032_6048, w_032_6050, w_032_6052, w_032_6053, w_032_6054, w_032_6056, w_032_6057, w_032_6058, w_032_6060, w_032_6063, w_032_6065, w_032_6067, w_032_6068, w_032_6070, w_032_6073, w_032_6075, w_032_6076, w_032_6078, w_032_6079, w_032_6081, w_032_6082, w_032_6083, w_032_6084, w_032_6085, w_032_6089, w_032_6093, w_032_6096, w_032_6097, w_032_6100, w_032_6101, w_032_6104, w_032_6107, w_032_6108, w_032_6115, w_032_6117, w_032_6121, w_032_6122, w_032_6123, w_032_6124, w_032_6131, w_032_6133, w_032_6134, w_032_6137, w_032_6139, w_032_6142, w_032_6144, w_032_6147, w_032_6150, w_032_6151, w_032_6152, w_032_6153, w_032_6155, w_032_6157, w_032_6158, w_032_6159, w_032_6160, w_032_6161, w_032_6162, w_032_6168, w_032_6171, w_032_6172, w_032_6173, w_032_6176, w_032_6179, w_032_6180, w_032_6181, w_032_6182, w_032_6186, w_032_6188, w_032_6189, w_032_6190, w_032_6191, w_032_6193, w_032_6194, w_032_6195, w_032_6197, w_032_6198, w_032_6199, w_032_6202, w_032_6203, w_032_6204, w_032_6205, w_032_6207, w_032_6210, w_032_6212, w_032_6213, w_032_6214, w_032_6218, w_032_6220, w_032_6222, w_032_6223, w_032_6224, w_032_6226, w_032_6227, w_032_6228, w_032_6229, w_032_6230, w_032_6232, w_032_6236, w_032_6238, w_032_6241, w_032_6244, w_032_6247, w_032_6248, w_032_6250, w_032_6251, w_032_6252, w_032_6254, w_032_6255, w_032_6258, w_032_6260, w_032_6263, w_032_6264, w_032_6268, w_032_6269, w_032_6274, w_032_6276, w_032_6277, w_032_6280, w_032_6281, w_032_6283, w_032_6285, w_032_6288, w_032_6289, w_032_6296, w_032_6298, w_032_6299, w_032_6303, w_032_6305, w_032_6306, w_032_6307, w_032_6309, w_032_6310, w_032_6311, w_032_6312, w_032_6313, w_032_6314, w_032_6316, w_032_6318, w_032_6319, w_032_6324, w_032_6326, w_032_6327, w_032_6328, w_032_6329, w_032_6330, w_032_6331, w_032_6332, w_032_6333, w_032_6334, w_032_6335, w_032_6336, w_032_6338, w_032_6339, w_032_6341, w_032_6344, w_032_6347, w_032_6352, w_032_6355, w_032_6356, w_032_6357, w_032_6359, w_032_6360, w_032_6361, w_032_6362, w_032_6363, w_032_6364, w_032_6367, w_032_6369, w_032_6370, w_032_6373, w_032_6376, w_032_6377, w_032_6378, w_032_6379, w_032_6380, w_032_6384, w_032_6386, w_032_6387, w_032_6389, w_032_6391, w_032_6392, w_032_6393, w_032_6395, w_032_6398, w_032_6402, w_032_6404, w_032_6405, w_032_6407, w_032_6409, w_032_6412, w_032_6415, w_032_6417, w_032_6418, w_032_6423, w_032_6424, w_032_6426, w_032_6427, w_032_6428, w_032_6431, w_032_6432, w_032_6433, w_032_6437, w_032_6439, w_032_6442, w_032_6446, w_032_6449, w_032_6450, w_032_6452, w_032_6455, w_032_6460, w_032_6462, w_032_6463, w_032_6464, w_032_6465, w_032_6466, w_032_6467, w_032_6469, w_032_6470, w_032_6472, w_032_6474, w_032_6475, w_032_6482, w_032_6484, w_032_6485, w_032_6486, w_032_6490, w_032_6492, w_032_6493, w_032_6495, w_032_6496, w_032_6497, w_032_6500, w_032_6501, w_032_6502, w_032_6503, w_032_6504, w_032_6506, w_032_6507, w_032_6509, w_032_6510, w_032_6513, w_032_6514, w_032_6515, w_032_6516, w_032_6517, w_032_6519, w_032_6520, w_032_6521, w_032_6522, w_032_6523, w_032_6524, w_032_6527, w_032_6529, w_032_6532, w_032_6536, w_032_6537, w_032_6538, w_032_6539, w_032_6540, w_032_6543, w_032_6544, w_032_6545, w_032_6546, w_032_6547, w_032_6549, w_032_6550, w_032_6552, w_032_6553, w_032_6554, w_032_6555, w_032_6557, w_032_6560, w_032_6566, w_032_6567, w_032_6569, w_032_6579, w_032_6580, w_032_6581, w_032_6582, w_032_6585, w_032_6586, w_032_6587, w_032_6588, w_032_6589, w_032_6590, w_032_6593, w_032_6594, w_032_6595, w_032_6596, w_032_6599, w_032_6600, w_032_6601, w_032_6603, w_032_6604, w_032_6605, w_032_6610, w_032_6612, w_032_6614, w_032_6615, w_032_6616, w_032_6617, w_032_6619, w_032_6621, w_032_6624, w_032_6625, w_032_6626, w_032_6627, w_032_6634, w_032_6635, w_032_6637, w_032_6643, w_032_6645, w_032_6646, w_032_6649, w_032_6651, w_032_6654, w_032_6656, w_032_6659, w_032_6661, w_032_6662, w_032_6663, w_032_6665, w_032_6667, w_032_6668, w_032_6674, w_032_6679, w_032_6680, w_032_6684, w_032_6686, w_032_6688, w_032_6689, w_032_6691, w_032_6692, w_032_6694, w_032_6695, w_032_6696, w_032_6698, w_032_6699, w_032_6701, w_032_6702, w_032_6703, w_032_6704, w_032_6705, w_032_6708, w_032_6710, w_032_6713, w_032_6714, w_032_6715, w_032_6718, w_032_6719, w_032_6720, w_032_6721, w_032_6723, w_032_6725, w_032_6726, w_032_6727;
  wire w_033_000, w_033_001, w_033_002, w_033_003, w_033_004, w_033_005, w_033_006, w_033_007, w_033_008, w_033_009, w_033_010, w_033_011, w_033_012, w_033_013, w_033_014, w_033_016, w_033_017, w_033_018, w_033_019, w_033_020, w_033_022, w_033_023, w_033_024, w_033_025, w_033_026, w_033_027, w_033_028, w_033_029, w_033_030, w_033_031, w_033_032, w_033_033, w_033_034, w_033_035, w_033_036, w_033_037, w_033_038, w_033_039, w_033_040, w_033_041, w_033_042, w_033_043, w_033_044, w_033_045, w_033_046, w_033_047, w_033_048, w_033_049, w_033_050, w_033_051, w_033_052, w_033_053, w_033_054, w_033_055, w_033_056, w_033_058, w_033_060, w_033_061, w_033_062, w_033_063, w_033_064, w_033_065, w_033_066, w_033_067, w_033_068, w_033_069, w_033_070, w_033_071, w_033_072, w_033_073, w_033_074, w_033_075, w_033_076, w_033_077, w_033_078, w_033_079, w_033_080, w_033_081, w_033_082, w_033_083, w_033_084, w_033_085, w_033_086, w_033_087, w_033_089, w_033_090, w_033_091, w_033_092, w_033_094, w_033_096, w_033_097, w_033_098, w_033_099, w_033_100, w_033_102, w_033_103, w_033_104, w_033_105, w_033_106, w_033_107, w_033_108, w_033_109, w_033_110, w_033_111, w_033_112, w_033_113, w_033_114, w_033_115, w_033_116, w_033_118, w_033_119, w_033_123, w_033_124, w_033_125, w_033_126, w_033_127, w_033_128, w_033_129, w_033_130, w_033_131, w_033_132, w_033_133, w_033_134, w_033_135, w_033_136, w_033_137, w_033_138, w_033_139, w_033_140, w_033_141, w_033_142, w_033_143, w_033_144, w_033_145, w_033_146, w_033_148, w_033_149, w_033_150, w_033_151, w_033_152, w_033_154, w_033_155, w_033_156, w_033_157, w_033_158, w_033_159, w_033_160, w_033_161, w_033_162, w_033_163, w_033_164, w_033_165, w_033_166, w_033_167, w_033_168, w_033_169, w_033_170, w_033_171, w_033_172, w_033_174, w_033_175, w_033_176, w_033_178, w_033_179, w_033_180, w_033_181, w_033_182, w_033_183, w_033_184, w_033_185, w_033_186, w_033_187, w_033_188, w_033_189, w_033_191, w_033_193, w_033_194, w_033_195, w_033_196, w_033_197, w_033_198, w_033_200, w_033_201, w_033_202, w_033_203, w_033_204, w_033_205, w_033_207, w_033_208, w_033_209, w_033_210, w_033_211, w_033_212, w_033_213, w_033_214, w_033_215, w_033_216, w_033_217, w_033_218, w_033_219, w_033_220, w_033_221, w_033_222, w_033_223, w_033_224, w_033_225, w_033_227, w_033_228, w_033_230, w_033_231, w_033_232, w_033_233, w_033_234, w_033_235, w_033_236, w_033_237, w_033_238, w_033_239, w_033_240, w_033_242, w_033_243, w_033_244, w_033_245, w_033_246, w_033_247, w_033_248, w_033_249, w_033_250, w_033_251, w_033_252, w_033_253, w_033_254, w_033_256, w_033_257, w_033_258, w_033_259, w_033_260, w_033_261, w_033_262, w_033_263, w_033_264, w_033_265, w_033_266, w_033_267, w_033_268, w_033_269, w_033_270, w_033_271, w_033_272, w_033_274, w_033_275, w_033_276, w_033_277, w_033_278, w_033_280, w_033_281, w_033_283, w_033_284, w_033_285, w_033_286, w_033_288, w_033_289, w_033_290, w_033_292, w_033_293, w_033_294, w_033_295, w_033_297, w_033_298, w_033_300, w_033_301, w_033_302, w_033_303, w_033_304, w_033_305, w_033_306, w_033_307, w_033_308, w_033_309, w_033_311, w_033_312, w_033_313, w_033_314, w_033_315, w_033_316, w_033_317, w_033_318, w_033_319, w_033_320, w_033_321, w_033_323, w_033_324, w_033_326, w_033_328, w_033_329, w_033_330, w_033_331, w_033_332, w_033_333, w_033_334, w_033_335, w_033_336, w_033_337, w_033_338, w_033_339, w_033_340, w_033_341, w_033_342, w_033_343, w_033_344, w_033_345, w_033_346, w_033_347, w_033_348, w_033_349, w_033_350, w_033_351, w_033_352, w_033_354, w_033_355, w_033_356, w_033_357, w_033_359, w_033_361, w_033_363, w_033_364, w_033_365, w_033_366, w_033_367, w_033_368, w_033_370, w_033_372, w_033_373, w_033_374, w_033_375, w_033_377, w_033_378, w_033_379, w_033_380, w_033_381, w_033_382, w_033_383, w_033_384, w_033_385, w_033_386, w_033_387, w_033_388, w_033_389, w_033_390, w_033_391, w_033_392, w_033_393, w_033_394, w_033_395, w_033_397, w_033_398, w_033_399, w_033_400, w_033_401, w_033_402, w_033_403, w_033_404, w_033_406, w_033_407, w_033_408, w_033_411, w_033_412, w_033_413, w_033_414, w_033_415, w_033_416, w_033_418, w_033_419, w_033_420, w_033_421, w_033_422, w_033_423, w_033_424, w_033_425, w_033_426, w_033_427, w_033_428, w_033_430, w_033_431, w_033_432, w_033_433, w_033_434, w_033_435, w_033_436, w_033_437, w_033_438, w_033_439, w_033_440, w_033_441, w_033_442, w_033_443, w_033_444, w_033_445, w_033_446, w_033_447, w_033_448, w_033_449, w_033_450, w_033_451, w_033_452, w_033_453, w_033_454, w_033_456, w_033_457, w_033_458, w_033_459, w_033_460, w_033_461, w_033_462, w_033_463, w_033_464, w_033_465, w_033_466, w_033_467, w_033_468, w_033_469, w_033_470, w_033_471, w_033_472, w_033_473, w_033_474, w_033_475, w_033_476, w_033_477, w_033_478, w_033_479, w_033_480, w_033_481, w_033_483, w_033_484, w_033_485, w_033_486, w_033_487, w_033_488, w_033_489, w_033_490, w_033_491, w_033_492, w_033_493, w_033_495, w_033_496, w_033_497, w_033_498, w_033_499, w_033_500, w_033_502, w_033_503, w_033_504, w_033_505, w_033_506, w_033_507, w_033_508, w_033_509, w_033_510, w_033_511, w_033_513, w_033_514, w_033_515, w_033_516, w_033_517, w_033_518, w_033_519, w_033_521, w_033_522, w_033_523, w_033_524, w_033_525, w_033_526, w_033_527, w_033_528, w_033_529, w_033_530, w_033_531, w_033_532, w_033_533, w_033_534, w_033_535, w_033_536, w_033_537, w_033_538, w_033_539, w_033_540, w_033_542, w_033_543, w_033_544, w_033_545, w_033_546, w_033_547, w_033_548, w_033_549, w_033_550, w_033_551, w_033_552, w_033_553, w_033_554, w_033_555, w_033_556, w_033_557, w_033_558, w_033_559, w_033_560, w_033_561, w_033_563, w_033_564, w_033_566, w_033_567, w_033_568, w_033_569, w_033_570, w_033_571, w_033_572, w_033_573, w_033_574, w_033_576, w_033_577, w_033_578, w_033_581, w_033_582, w_033_583, w_033_584, w_033_585, w_033_586, w_033_587, w_033_588, w_033_589, w_033_590, w_033_591, w_033_592, w_033_593, w_033_594, w_033_595, w_033_596, w_033_598, w_033_599, w_033_600, w_033_601, w_033_603, w_033_604, w_033_605, w_033_606, w_033_607, w_033_608, w_033_609, w_033_610, w_033_611, w_033_612, w_033_613, w_033_615, w_033_616, w_033_617, w_033_618, w_033_619, w_033_620, w_033_621, w_033_622, w_033_623, w_033_624, w_033_625, w_033_626, w_033_627, w_033_628, w_033_629, w_033_630, w_033_631, w_033_632, w_033_633, w_033_634, w_033_635, w_033_636, w_033_638, w_033_639, w_033_640, w_033_641, w_033_642, w_033_643, w_033_645, w_033_647, w_033_648, w_033_649, w_033_650, w_033_651, w_033_652, w_033_653, w_033_654, w_033_656, w_033_657, w_033_658, w_033_659, w_033_660, w_033_661, w_033_662, w_033_663, w_033_664, w_033_665, w_033_666, w_033_667, w_033_668, w_033_669, w_033_670, w_033_671, w_033_672, w_033_673, w_033_674, w_033_676, w_033_677, w_033_678, w_033_679, w_033_680, w_033_681, w_033_682, w_033_683, w_033_684, w_033_685, w_033_686, w_033_687, w_033_688, w_033_690, w_033_691, w_033_693, w_033_694, w_033_695, w_033_696, w_033_698, w_033_699, w_033_700, w_033_701, w_033_703, w_033_704, w_033_706, w_033_707, w_033_708, w_033_709, w_033_710, w_033_711, w_033_712, w_033_713, w_033_715, w_033_716, w_033_717, w_033_718, w_033_719, w_033_721, w_033_722, w_033_723, w_033_724, w_033_726, w_033_727, w_033_730, w_033_731, w_033_732, w_033_733, w_033_735, w_033_736, w_033_737, w_033_738, w_033_739, w_033_741, w_033_742, w_033_743, w_033_744, w_033_745, w_033_746, w_033_747, w_033_749, w_033_750, w_033_751, w_033_752, w_033_753, w_033_754, w_033_755, w_033_756, w_033_758, w_033_760, w_033_761, w_033_762, w_033_763, w_033_764, w_033_766, w_033_767, w_033_768, w_033_769, w_033_770, w_033_771, w_033_772, w_033_773, w_033_774, w_033_775, w_033_776, w_033_777, w_033_778, w_033_779, w_033_780, w_033_781, w_033_782, w_033_783, w_033_784, w_033_785, w_033_786, w_033_787, w_033_788, w_033_789, w_033_790, w_033_791, w_033_792, w_033_793, w_033_794, w_033_796, w_033_797, w_033_798, w_033_799, w_033_801, w_033_802, w_033_803, w_033_804, w_033_805, w_033_806, w_033_807, w_033_808, w_033_809, w_033_810, w_033_811, w_033_812, w_033_813, w_033_814, w_033_815, w_033_817, w_033_818, w_033_819, w_033_821, w_033_822, w_033_823, w_033_824, w_033_825, w_033_826, w_033_827, w_033_828, w_033_829, w_033_830, w_033_831, w_033_832, w_033_833, w_033_834, w_033_836, w_033_837, w_033_838, w_033_839, w_033_840, w_033_841, w_033_842, w_033_843, w_033_844, w_033_845, w_033_846, w_033_847, w_033_848, w_033_849, w_033_850, w_033_851, w_033_852, w_033_853, w_033_854, w_033_855, w_033_856, w_033_857, w_033_858, w_033_859, w_033_860, w_033_861, w_033_862, w_033_863, w_033_864, w_033_865, w_033_866, w_033_867, w_033_868, w_033_869, w_033_870, w_033_871, w_033_872, w_033_873, w_033_874, w_033_875, w_033_876, w_033_877, w_033_878, w_033_879, w_033_880, w_033_881, w_033_882, w_033_883, w_033_886, w_033_887, w_033_888, w_033_890, w_033_891, w_033_892, w_033_893, w_033_894, w_033_895, w_033_896, w_033_897, w_033_898, w_033_899, w_033_900, w_033_901, w_033_902, w_033_903, w_033_904, w_033_905, w_033_906, w_033_907, w_033_908, w_033_909, w_033_910, w_033_912, w_033_913, w_033_914, w_033_915, w_033_916, w_033_917, w_033_918, w_033_919, w_033_920, w_033_921, w_033_922, w_033_923, w_033_924, w_033_925, w_033_926, w_033_927, w_033_929, w_033_930, w_033_931, w_033_932, w_033_933, w_033_934, w_033_935, w_033_938, w_033_940, w_033_941, w_033_942, w_033_943, w_033_945, w_033_946, w_033_949, w_033_950, w_033_951, w_033_953, w_033_954, w_033_955, w_033_957, w_033_958, w_033_959, w_033_960, w_033_961, w_033_962, w_033_963, w_033_965, w_033_966, w_033_967, w_033_968, w_033_969, w_033_970, w_033_971, w_033_972, w_033_973, w_033_975, w_033_976, w_033_977, w_033_978, w_033_979, w_033_980, w_033_981, w_033_982, w_033_983, w_033_984, w_033_985, w_033_986, w_033_987, w_033_988, w_033_989, w_033_990, w_033_991, w_033_992, w_033_993, w_033_995, w_033_997, w_033_998, w_033_999, w_033_1000, w_033_1001, w_033_1002, w_033_1003, w_033_1004, w_033_1005, w_033_1006, w_033_1007, w_033_1009, w_033_1010, w_033_1012, w_033_1013, w_033_1015, w_033_1016, w_033_1018, w_033_1019, w_033_1020, w_033_1021, w_033_1023, w_033_1024, w_033_1025, w_033_1026, w_033_1027, w_033_1028, w_033_1029, w_033_1030, w_033_1031, w_033_1032, w_033_1033, w_033_1034, w_033_1036, w_033_1037, w_033_1038, w_033_1039, w_033_1040, w_033_1041, w_033_1042, w_033_1043, w_033_1044, w_033_1045, w_033_1046, w_033_1047, w_033_1048, w_033_1049, w_033_1050, w_033_1051, w_033_1052, w_033_1053, w_033_1054, w_033_1055, w_033_1056, w_033_1058, w_033_1059, w_033_1060, w_033_1061, w_033_1062, w_033_1063, w_033_1065, w_033_1066, w_033_1067, w_033_1069, w_033_1070, w_033_1071, w_033_1072, w_033_1073, w_033_1074, w_033_1075, w_033_1076, w_033_1078, w_033_1079, w_033_1080, w_033_1081, w_033_1082, w_033_1083, w_033_1084, w_033_1085, w_033_1086, w_033_1087, w_033_1088, w_033_1089, w_033_1090, w_033_1091, w_033_1092, w_033_1093, w_033_1094, w_033_1095, w_033_1096, w_033_1097, w_033_1099, w_033_1100, w_033_1102, w_033_1103, w_033_1104, w_033_1106, w_033_1107, w_033_1109, w_033_1110, w_033_1111, w_033_1112, w_033_1113, w_033_1114, w_033_1115, w_033_1116, w_033_1117, w_033_1118, w_033_1119, w_033_1120, w_033_1121, w_033_1122, w_033_1123, w_033_1124, w_033_1125, w_033_1126, w_033_1127, w_033_1128, w_033_1129, w_033_1130, w_033_1131, w_033_1132, w_033_1133, w_033_1134, w_033_1135, w_033_1136, w_033_1137, w_033_1138, w_033_1139, w_033_1140, w_033_1141, w_033_1142, w_033_1144, w_033_1145, w_033_1146, w_033_1147, w_033_1148, w_033_1149, w_033_1150, w_033_1152, w_033_1153, w_033_1154, w_033_1155, w_033_1156, w_033_1158, w_033_1159, w_033_1160, w_033_1161, w_033_1162, w_033_1163, w_033_1164, w_033_1165, w_033_1166, w_033_1167, w_033_1168, w_033_1171, w_033_1172, w_033_1173, w_033_1174, w_033_1175, w_033_1177, w_033_1178, w_033_1179, w_033_1180, w_033_1181, w_033_1182, w_033_1183, w_033_1184, w_033_1185, w_033_1186, w_033_1187, w_033_1190, w_033_1191, w_033_1192, w_033_1193, w_033_1194, w_033_1195, w_033_1196, w_033_1198, w_033_1199, w_033_1201, w_033_1202, w_033_1203, w_033_1204, w_033_1205, w_033_1207, w_033_1208, w_033_1209, w_033_1210, w_033_1211, w_033_1212, w_033_1213, w_033_1214, w_033_1216, w_033_1217, w_033_1218, w_033_1219, w_033_1220, w_033_1221, w_033_1222, w_033_1223, w_033_1224, w_033_1225, w_033_1226, w_033_1227, w_033_1228, w_033_1229, w_033_1230, w_033_1231, w_033_1232, w_033_1234, w_033_1235, w_033_1236, w_033_1237, w_033_1239, w_033_1240, w_033_1241, w_033_1242, w_033_1243, w_033_1244, w_033_1245, w_033_1246, w_033_1247, w_033_1248, w_033_1249, w_033_1250, w_033_1251, w_033_1252, w_033_1253, w_033_1255, w_033_1256, w_033_1257, w_033_1258, w_033_1259, w_033_1260, w_033_1261, w_033_1262, w_033_1263, w_033_1264, w_033_1265, w_033_1266, w_033_1268, w_033_1269, w_033_1270, w_033_1271, w_033_1272, w_033_1273, w_033_1275, w_033_1276, w_033_1277, w_033_1278, w_033_1279, w_033_1280, w_033_1281, w_033_1282, w_033_1284, w_033_1285, w_033_1286, w_033_1287, w_033_1288, w_033_1289, w_033_1290, w_033_1291, w_033_1292, w_033_1293, w_033_1294, w_033_1295, w_033_1296, w_033_1297, w_033_1299, w_033_1300, w_033_1301, w_033_1302, w_033_1303, w_033_1304, w_033_1305, w_033_1306, w_033_1307, w_033_1308, w_033_1309, w_033_1310, w_033_1311, w_033_1312, w_033_1313, w_033_1314, w_033_1317, w_033_1318, w_033_1319, w_033_1320, w_033_1321, w_033_1322, w_033_1323, w_033_1324, w_033_1325, w_033_1326, w_033_1327, w_033_1328, w_033_1329, w_033_1330, w_033_1331, w_033_1332, w_033_1333, w_033_1334, w_033_1335, w_033_1336, w_033_1338, w_033_1339, w_033_1340, w_033_1342, w_033_1343, w_033_1344, w_033_1346, w_033_1347, w_033_1348, w_033_1349, w_033_1350, w_033_1351, w_033_1352, w_033_1354, w_033_1355, w_033_1356, w_033_1357, w_033_1358, w_033_1359, w_033_1360, w_033_1361, w_033_1362, w_033_1363, w_033_1364, w_033_1366, w_033_1367, w_033_1368, w_033_1369, w_033_1370, w_033_1371, w_033_1372, w_033_1373, w_033_1374, w_033_1375, w_033_1376, w_033_1377, w_033_1379, w_033_1381, w_033_1382, w_033_1383, w_033_1384, w_033_1385, w_033_1386, w_033_1387, w_033_1388, w_033_1389, w_033_1390, w_033_1391, w_033_1392, w_033_1393, w_033_1394, w_033_1395, w_033_1397, w_033_1398, w_033_1399, w_033_1400, w_033_1401, w_033_1402, w_033_1403, w_033_1404, w_033_1405, w_033_1406, w_033_1407, w_033_1408, w_033_1409, w_033_1410, w_033_1411, w_033_1413, w_033_1414, w_033_1415, w_033_1416, w_033_1417, w_033_1418, w_033_1419, w_033_1420, w_033_1421, w_033_1422, w_033_1423, w_033_1424, w_033_1425, w_033_1426, w_033_1427, w_033_1428, w_033_1429, w_033_1430, w_033_1431, w_033_1433, w_033_1434, w_033_1435, w_033_1436, w_033_1437, w_033_1438, w_033_1440, w_033_1442, w_033_1443, w_033_1444, w_033_1446, w_033_1447, w_033_1448, w_033_1449, w_033_1450, w_033_1451, w_033_1452, w_033_1453, w_033_1454, w_033_1456, w_033_1457, w_033_1458, w_033_1459, w_033_1460, w_033_1461, w_033_1462, w_033_1464, w_033_1465, w_033_1466, w_033_1467, w_033_1469, w_033_1470, w_033_1471, w_033_1472, w_033_1473, w_033_1474, w_033_1475, w_033_1476, w_033_1477, w_033_1478, w_033_1480, w_033_1481, w_033_1482, w_033_1483, w_033_1484, w_033_1485, w_033_1486, w_033_1488, w_033_1489, w_033_1490, w_033_1491, w_033_1492, w_033_1493, w_033_1494, w_033_1495, w_033_1497, w_033_1498, w_033_1499, w_033_1500, w_033_1501, w_033_1502, w_033_1503, w_033_1504, w_033_1505, w_033_1506, w_033_1507, w_033_1508, w_033_1509, w_033_1510, w_033_1511, w_033_1512, w_033_1513, w_033_1514, w_033_1515, w_033_1517, w_033_1518, w_033_1519, w_033_1520, w_033_1521, w_033_1522, w_033_1523, w_033_1524, w_033_1525, w_033_1526, w_033_1527, w_033_1528, w_033_1529, w_033_1530, w_033_1531, w_033_1532, w_033_1533, w_033_1534, w_033_1536, w_033_1537, w_033_1538, w_033_1539, w_033_1540, w_033_1541, w_033_1542, w_033_1543, w_033_1544, w_033_1545, w_033_1546, w_033_1547, w_033_1548, w_033_1550, w_033_1551, w_033_1552, w_033_1553, w_033_1554, w_033_1555, w_033_1556, w_033_1557, w_033_1558, w_033_1559, w_033_1560, w_033_1561, w_033_1562, w_033_1563, w_033_1565, w_033_1566, w_033_1567, w_033_1568, w_033_1569, w_033_1570, w_033_1571, w_033_1572, w_033_1573, w_033_1574, w_033_1575, w_033_1576, w_033_1577, w_033_1578, w_033_1579, w_033_1580, w_033_1581, w_033_1582, w_033_1584, w_033_1586, w_033_1588, w_033_1590, w_033_1592, w_033_1594, w_033_1595, w_033_1596, w_033_1597, w_033_1598, w_033_1600, w_033_1601, w_033_1602, w_033_1603, w_033_1605, w_033_1606, w_033_1607, w_033_1608, w_033_1609, w_033_1610, w_033_1611, w_033_1612, w_033_1613, w_033_1614, w_033_1615, w_033_1616, w_033_1618, w_033_1619, w_033_1620, w_033_1621, w_033_1622, w_033_1623, w_033_1624, w_033_1625, w_033_1626, w_033_1628, w_033_1629, w_033_1630, w_033_1631, w_033_1632, w_033_1633, w_033_1634, w_033_1635, w_033_1636, w_033_1637, w_033_1638, w_033_1639, w_033_1640, w_033_1641, w_033_1642, w_033_1644, w_033_1645, w_033_1646, w_033_1647, w_033_1649, w_033_1650, w_033_1651, w_033_1652, w_033_1653, w_033_1654, w_033_1655, w_033_1656, w_033_1657, w_033_1658, w_033_1659, w_033_1660, w_033_1661, w_033_1662, w_033_1664, w_033_1665, w_033_1666, w_033_1667, w_033_1668, w_033_1669, w_033_1670, w_033_1671, w_033_1672, w_033_1673, w_033_1675, w_033_1676, w_033_1677, w_033_1678, w_033_1679, w_033_1680, w_033_1681, w_033_1682, w_033_1683, w_033_1684, w_033_1685, w_033_1686, w_033_1687, w_033_1688, w_033_1689, w_033_1690, w_033_1693, w_033_1694, w_033_1695, w_033_1696, w_033_1697, w_033_1698, w_033_1699, w_033_1700, w_033_1701, w_033_1702, w_033_1703, w_033_1704, w_033_1705, w_033_1706, w_033_1707, w_033_1708, w_033_1709, w_033_1710, w_033_1711, w_033_1712, w_033_1713, w_033_1714, w_033_1715, w_033_1716, w_033_1717, w_033_1719, w_033_1720, w_033_1721, w_033_1722, w_033_1723, w_033_1724, w_033_1725, w_033_1726, w_033_1727, w_033_1728, w_033_1729, w_033_1730, w_033_1731, w_033_1732, w_033_1733, w_033_1734, w_033_1735, w_033_1736, w_033_1737, w_033_1738, w_033_1739, w_033_1740, w_033_1741, w_033_1744, w_033_1745, w_033_1746, w_033_1747, w_033_1749, w_033_1750, w_033_1751, w_033_1752, w_033_1753, w_033_1755, w_033_1756, w_033_1757, w_033_1758, w_033_1759, w_033_1760, w_033_1761, w_033_1763, w_033_1764, w_033_1765, w_033_1766, w_033_1768, w_033_1769, w_033_1770, w_033_1772, w_033_1773, w_033_1774, w_033_1775, w_033_1776, w_033_1777, w_033_1778, w_033_1779, w_033_1780, w_033_1781, w_033_1782, w_033_1783, w_033_1785, w_033_1787, w_033_1788, w_033_1789, w_033_1790, w_033_1791, w_033_1792, w_033_1793, w_033_1794, w_033_1795, w_033_1796, w_033_1797, w_033_1798, w_033_1800, w_033_1801, w_033_1803, w_033_1804, w_033_1805, w_033_1806, w_033_1807, w_033_1808, w_033_1810, w_033_1811, w_033_1812, w_033_1813, w_033_1814, w_033_1816, w_033_1817, w_033_1818, w_033_1819, w_033_1820, w_033_1821, w_033_1822, w_033_1827, w_033_1828, w_033_1829, w_033_1830, w_033_1831, w_033_1832, w_033_1834, w_033_1835, w_033_1836, w_033_1837, w_033_1838, w_033_1839, w_033_1840, w_033_1841, w_033_1842, w_033_1843, w_033_1844, w_033_1845, w_033_1846, w_033_1847, w_033_1848, w_033_1849, w_033_1850, w_033_1851, w_033_1852, w_033_1853, w_033_1854, w_033_1855, w_033_1856, w_033_1857, w_033_1858, w_033_1860, w_033_1861, w_033_1862, w_033_1863, w_033_1864, w_033_1865, w_033_1866, w_033_1867, w_033_1868, w_033_1869, w_033_1870, w_033_1871, w_033_1872, w_033_1874, w_033_1875, w_033_1876, w_033_1877, w_033_1879, w_033_1880, w_033_1881, w_033_1882, w_033_1883, w_033_1884, w_033_1885, w_033_1886, w_033_1887, w_033_1889, w_033_1890, w_033_1892, w_033_1893, w_033_1894, w_033_1895, w_033_1896, w_033_1897, w_033_1898, w_033_1900, w_033_1901, w_033_1902, w_033_1903, w_033_1904, w_033_1905, w_033_1906, w_033_1907, w_033_1909, w_033_1910, w_033_1911, w_033_1912, w_033_1913, w_033_1914, w_033_1915, w_033_1916, w_033_1917, w_033_1918, w_033_1919, w_033_1920, w_033_1921, w_033_1923, w_033_1926, w_033_1927, w_033_1928, w_033_1929, w_033_1932, w_033_1933, w_033_1935, w_033_1936, w_033_1937, w_033_1938, w_033_1942, w_033_1943, w_033_1945, w_033_1946, w_033_1947, w_033_1948, w_033_1949, w_033_1950, w_033_1951, w_033_1952, w_033_1954, w_033_1955, w_033_1956, w_033_1957, w_033_1958, w_033_1960, w_033_1961, w_033_1962, w_033_1963, w_033_1965, w_033_1966, w_033_1967, w_033_1968, w_033_1969, w_033_1970, w_033_1971, w_033_1972, w_033_1973, w_033_1974, w_033_1975, w_033_1976, w_033_1977, w_033_1978, w_033_1979, w_033_1980, w_033_1981, w_033_1982, w_033_1983, w_033_1984, w_033_1985, w_033_1986, w_033_1987, w_033_1990, w_033_1991, w_033_1992, w_033_1993, w_033_1995, w_033_1996, w_033_1997, w_033_1998, w_033_1999, w_033_2000, w_033_2001, w_033_2002, w_033_2003, w_033_2004, w_033_2005, w_033_2006, w_033_2007, w_033_2008, w_033_2009, w_033_2010, w_033_2011, w_033_2012, w_033_2013, w_033_2014, w_033_2016, w_033_2017, w_033_2018, w_033_2019, w_033_2020, w_033_2021, w_033_2022, w_033_2023, w_033_2024, w_033_2025, w_033_2026, w_033_2027, w_033_2028, w_033_2029, w_033_2030, w_033_2031, w_033_2032, w_033_2033, w_033_2034, w_033_2036, w_033_2038, w_033_2039, w_033_2040, w_033_2041, w_033_2042, w_033_2044, w_033_2045, w_033_2046, w_033_2047, w_033_2048, w_033_2049, w_033_2050, w_033_2051, w_033_2052, w_033_2054, w_033_2055, w_033_2056, w_033_2058, w_033_2059, w_033_2060, w_033_2061, w_033_2062, w_033_2063, w_033_2064, w_033_2065, w_033_2066, w_033_2067, w_033_2068, w_033_2069, w_033_2070, w_033_2071, w_033_2072, w_033_2073, w_033_2074, w_033_2076, w_033_2077, w_033_2078, w_033_2080, w_033_2081, w_033_2084, w_033_2085, w_033_2086, w_033_2088, w_033_2089, w_033_2090, w_033_2091, w_033_2092, w_033_2093, w_033_2094, w_033_2095, w_033_2096, w_033_2097, w_033_2098, w_033_2099, w_033_2100, w_033_2102, w_033_2103, w_033_2104, w_033_2105, w_033_2106, w_033_2107, w_033_2108, w_033_2110, w_033_2111, w_033_2112, w_033_2113, w_033_2114, w_033_2115, w_033_2116, w_033_2117, w_033_2118, w_033_2120, w_033_2121, w_033_2122, w_033_2123, w_033_2124, w_033_2126, w_033_2127, w_033_2128, w_033_2129, w_033_2130, w_033_2131, w_033_2132, w_033_2133, w_033_2135, w_033_2136, w_033_2137, w_033_2138, w_033_2139, w_033_2140, w_033_2141, w_033_2142, w_033_2143, w_033_2144, w_033_2145, w_033_2146, w_033_2147, w_033_2148, w_033_2149, w_033_2150, w_033_2151, w_033_2152, w_033_2153, w_033_2154, w_033_2155, w_033_2156, w_033_2157, w_033_2158, w_033_2159, w_033_2160, w_033_2161, w_033_2162, w_033_2163, w_033_2164, w_033_2165, w_033_2166, w_033_2167, w_033_2169, w_033_2170, w_033_2171, w_033_2173, w_033_2174, w_033_2175, w_033_2176, w_033_2177, w_033_2179, w_033_2180, w_033_2181, w_033_2182, w_033_2183, w_033_2184, w_033_2185, w_033_2186, w_033_2187, w_033_2188, w_033_2189, w_033_2190, w_033_2191, w_033_2192, w_033_2193, w_033_2194, w_033_2195, w_033_2196, w_033_2197, w_033_2199, w_033_2200, w_033_2201, w_033_2202, w_033_2203, w_033_2204, w_033_2205, w_033_2206, w_033_2207, w_033_2210, w_033_2211, w_033_2212, w_033_2213, w_033_2215, w_033_2216, w_033_2218, w_033_2219, w_033_2220, w_033_2222, w_033_2223, w_033_2224, w_033_2225, w_033_2227, w_033_2228, w_033_2229, w_033_2230, w_033_2231, w_033_2232, w_033_2233, w_033_2234, w_033_2237, w_033_2238, w_033_2239, w_033_2240, w_033_2241, w_033_2242, w_033_2243, w_033_2244, w_033_2248, w_033_2249, w_033_2250, w_033_2252, w_033_2253, w_033_2254, w_033_2255, w_033_2257, w_033_2258, w_033_2259, w_033_2260, w_033_2261, w_033_2262, w_033_2263, w_033_2264, w_033_2265, w_033_2266, w_033_2267, w_033_2268, w_033_2269, w_033_2270, w_033_2271, w_033_2272, w_033_2274, w_033_2275, w_033_2276, w_033_2278, w_033_2279, w_033_2281, w_033_2282, w_033_2283, w_033_2284, w_033_2285, w_033_2286, w_033_2287, w_033_2288, w_033_2289, w_033_2290, w_033_2291, w_033_2292, w_033_2293, w_033_2294, w_033_2295, w_033_2296, w_033_2297, w_033_2298, w_033_2299, w_033_2300, w_033_2301, w_033_2302, w_033_2303, w_033_2304, w_033_2305, w_033_2306, w_033_2307, w_033_2308, w_033_2309, w_033_2310, w_033_2311, w_033_2312, w_033_2314, w_033_2316, w_033_2317, w_033_2319, w_033_2320, w_033_2321, w_033_2322, w_033_2323, w_033_2324, w_033_2325, w_033_2326, w_033_2327, w_033_2328, w_033_2329, w_033_2330, w_033_2331, w_033_2332, w_033_2333, w_033_2334, w_033_2336, w_033_2337, w_033_2338, w_033_2339, w_033_2340, w_033_2341, w_033_2342, w_033_2344, w_033_2345, w_033_2346, w_033_2347, w_033_2348, w_033_2349, w_033_2351, w_033_2352, w_033_2353, w_033_2354, w_033_2355, w_033_2356, w_033_2357, w_033_2358, w_033_2359, w_033_2360, w_033_2361, w_033_2362, w_033_2363, w_033_2364, w_033_2365, w_033_2366, w_033_2367, w_033_2368, w_033_2369, w_033_2370, w_033_2371, w_033_2372, w_033_2373, w_033_2374, w_033_2375, w_033_2376, w_033_2377, w_033_2378, w_033_2379, w_033_2380, w_033_2381, w_033_2382, w_033_2383, w_033_2384, w_033_2385, w_033_2387, w_033_2388, w_033_2389, w_033_2390, w_033_2391, w_033_2392, w_033_2393, w_033_2394, w_033_2395, w_033_2396, w_033_2397, w_033_2399, w_033_2400, w_033_2401, w_033_2402, w_033_2403, w_033_2404, w_033_2405, w_033_2408, w_033_2409, w_033_2410, w_033_2411, w_033_2412, w_033_2413, w_033_2414, w_033_2415, w_033_2417, w_033_2418, w_033_2419, w_033_2420, w_033_2421, w_033_2422, w_033_2423, w_033_2424, w_033_2425, w_033_2426, w_033_2427, w_033_2428, w_033_2429, w_033_2430, w_033_2431, w_033_2432, w_033_2433, w_033_2434, w_033_2435, w_033_2436, w_033_2437, w_033_2438, w_033_2439, w_033_2440, w_033_2441, w_033_2442, w_033_2443, w_033_2444, w_033_2445, w_033_2447, w_033_2448, w_033_2449, w_033_2450, w_033_2451, w_033_2452, w_033_2453, w_033_2454, w_033_2455, w_033_2456, w_033_2457, w_033_2458, w_033_2459, w_033_2460, w_033_2461, w_033_2462, w_033_2464, w_033_2465, w_033_2466, w_033_2467, w_033_2468, w_033_2469, w_033_2470, w_033_2471, w_033_2473, w_033_2474, w_033_2475, w_033_2476, w_033_2477, w_033_2478, w_033_2481, w_033_2482, w_033_2484, w_033_2485, w_033_2486, w_033_2487, w_033_2488, w_033_2490, w_033_2492, w_033_2493, w_033_2494, w_033_2495, w_033_2496, w_033_2497, w_033_2498, w_033_2499, w_033_2500, w_033_2502, w_033_2503, w_033_2504, w_033_2505, w_033_2506, w_033_2507, w_033_2508, w_033_2509, w_033_2510, w_033_2512, w_033_2513, w_033_2514, w_033_2515, w_033_2517, w_033_2518, w_033_2519, w_033_2520, w_033_2521, w_033_2523, w_033_2524, w_033_2525, w_033_2526, w_033_2527, w_033_2528, w_033_2529, w_033_2530, w_033_2531, w_033_2532, w_033_2533, w_033_2534, w_033_2535, w_033_2536, w_033_2538, w_033_2539, w_033_2540, w_033_2541, w_033_2542, w_033_2543, w_033_2544, w_033_2545, w_033_2546, w_033_2547, w_033_2548, w_033_2549, w_033_2551, w_033_2552, w_033_2553, w_033_2554, w_033_2555, w_033_2556, w_033_2557, w_033_2558, w_033_2559, w_033_2560, w_033_2561, w_033_2562, w_033_2563, w_033_2564, w_033_2565, w_033_2566, w_033_2567, w_033_2568, w_033_2569, w_033_2570, w_033_2571, w_033_2573, w_033_2575, w_033_2576, w_033_2577, w_033_2578, w_033_2579, w_033_2580, w_033_2581, w_033_2582, w_033_2583, w_033_2584, w_033_2585, w_033_2586, w_033_2587, w_033_2588, w_033_2589, w_033_2590, w_033_2591, w_033_2592, w_033_2593, w_033_2594, w_033_2595, w_033_2596, w_033_2597, w_033_2598, w_033_2599, w_033_2600, w_033_2601, w_033_2603, w_033_2604, w_033_2605, w_033_2607, w_033_2608, w_033_2610, w_033_2613, w_033_2614, w_033_2615, w_033_2616, w_033_2617, w_033_2618, w_033_2619, w_033_2621, w_033_2622, w_033_2623, w_033_2624, w_033_2625, w_033_2626, w_033_2627, w_033_2628, w_033_2629, w_033_2630, w_033_2631, w_033_2632, w_033_2633, w_033_2634, w_033_2635, w_033_2636, w_033_2637, w_033_2638, w_033_2639, w_033_2640, w_033_2641, w_033_2642, w_033_2643, w_033_2644, w_033_2645, w_033_2646, w_033_2647, w_033_2650, w_033_2651, w_033_2652, w_033_2653, w_033_2654, w_033_2655, w_033_2656, w_033_2657, w_033_2658, w_033_2659, w_033_2660, w_033_2661, w_033_2662, w_033_2663, w_033_2665, w_033_2666, w_033_2667, w_033_2668, w_033_2669, w_033_2671, w_033_2672, w_033_2673, w_033_2674, w_033_2675, w_033_2676, w_033_2677, w_033_2678, w_033_2679, w_033_2680, w_033_2681, w_033_2682, w_033_2684, w_033_2685, w_033_2686, w_033_2687, w_033_2688, w_033_2689, w_033_2690, w_033_2691, w_033_2692, w_033_2694, w_033_2695, w_033_2696, w_033_2697, w_033_2699, w_033_2700, w_033_2701, w_033_2702, w_033_2703, w_033_2704, w_033_2705, w_033_2706, w_033_2707, w_033_2709, w_033_2710, w_033_2711, w_033_2712, w_033_2714, w_033_2715, w_033_2716, w_033_2717, w_033_2718, w_033_2719, w_033_2722, w_033_2724, w_033_2726, w_033_2727, w_033_2728, w_033_2729, w_033_2730, w_033_2731, w_033_2732, w_033_2733, w_033_2734, w_033_2735, w_033_2737, w_033_2738, w_033_2739, w_033_2740, w_033_2741, w_033_2742, w_033_2743, w_033_2744, w_033_2745, w_033_2746, w_033_2747, w_033_2748, w_033_2749, w_033_2750, w_033_2751, w_033_2753, w_033_2754, w_033_2755, w_033_2757, w_033_2760, w_033_2761, w_033_2762, w_033_2765, w_033_2767, w_033_2768, w_033_2769, w_033_2770, w_033_2771, w_033_2773, w_033_2774, w_033_2775, w_033_2776, w_033_2777, w_033_2778, w_033_2779, w_033_2780, w_033_2781, w_033_2782, w_033_2784, w_033_2785, w_033_2787, w_033_2788, w_033_2789, w_033_2791, w_033_2793, w_033_2795, w_033_2797, w_033_2798, w_033_2799, w_033_2800, w_033_2801, w_033_2802, w_033_2803, w_033_2805, w_033_2806, w_033_2808, w_033_2809, w_033_2810, w_033_2811, w_033_2812, w_033_2813, w_033_2814, w_033_2817, w_033_2818, w_033_2820, w_033_2822, w_033_2823, w_033_2824, w_033_2825, w_033_2826, w_033_2827, w_033_2830, w_033_2831, w_033_2833, w_033_2834, w_033_2837, w_033_2838, w_033_2839, w_033_2840, w_033_2841, w_033_2842, w_033_2844, w_033_2846, w_033_2847, w_033_2848, w_033_2849, w_033_2851, w_033_2852, w_033_2854, w_033_2855, w_033_2857, w_033_2859, w_033_2860, w_033_2861, w_033_2862, w_033_2864, w_033_2865, w_033_2866, w_033_2867, w_033_2869, w_033_2871, w_033_2873, w_033_2874, w_033_2875, w_033_2876, w_033_2877, w_033_2880, w_033_2882, w_033_2883, w_033_2885, w_033_2886, w_033_2888, w_033_2889, w_033_2890, w_033_2891, w_033_2892, w_033_2894, w_033_2895, w_033_2896, w_033_2897, w_033_2898, w_033_2902, w_033_2903, w_033_2904, w_033_2905, w_033_2906, w_033_2908, w_033_2909, w_033_2910, w_033_2911, w_033_2912, w_033_2913, w_033_2914, w_033_2915, w_033_2916, w_033_2917, w_033_2918, w_033_2919, w_033_2921, w_033_2922, w_033_2923, w_033_2925, w_033_2926, w_033_2927, w_033_2928, w_033_2929, w_033_2931, w_033_2932, w_033_2933, w_033_2935, w_033_2936, w_033_2937, w_033_2938, w_033_2939, w_033_2940, w_033_2941, w_033_2942, w_033_2943, w_033_2944, w_033_2945, w_033_2946, w_033_2947, w_033_2948, w_033_2950, w_033_2953, w_033_2955, w_033_2956, w_033_2957, w_033_2958, w_033_2960, w_033_2961, w_033_2962, w_033_2964, w_033_2967, w_033_2968, w_033_2969, w_033_2970, w_033_2971, w_033_2972, w_033_2973, w_033_2974, w_033_2975, w_033_2976, w_033_2977, w_033_2980, w_033_2981, w_033_2983, w_033_2984, w_033_2985, w_033_2986, w_033_2989, w_033_2990, w_033_2991, w_033_2992, w_033_2995, w_033_2996, w_033_2997, w_033_2998, w_033_3000, w_033_3001, w_033_3002, w_033_3003, w_033_3004, w_033_3005, w_033_3006, w_033_3008, w_033_3009, w_033_3011, w_033_3012, w_033_3013, w_033_3014, w_033_3015, w_033_3021, w_033_3022, w_033_3023, w_033_3024, w_033_3025, w_033_3028, w_033_3029, w_033_3030, w_033_3031, w_033_3032, w_033_3033, w_033_3034, w_033_3035, w_033_3036, w_033_3037, w_033_3038, w_033_3039, w_033_3040, w_033_3041, w_033_3042, w_033_3043, w_033_3044, w_033_3045, w_033_3046, w_033_3047, w_033_3048, w_033_3049, w_033_3050, w_033_3051, w_033_3052, w_033_3053, w_033_3054, w_033_3058, w_033_3060, w_033_3061, w_033_3062, w_033_3063, w_033_3064, w_033_3065, w_033_3066, w_033_3067, w_033_3069, w_033_3070, w_033_3071, w_033_3072, w_033_3073, w_033_3074, w_033_3078, w_033_3080, w_033_3082, w_033_3085, w_033_3086, w_033_3088, w_033_3089, w_033_3090, w_033_3091, w_033_3092, w_033_3093, w_033_3094, w_033_3096, w_033_3097, w_033_3098, w_033_3100, w_033_3102, w_033_3104, w_033_3105, w_033_3106, w_033_3107, w_033_3109, w_033_3110, w_033_3111, w_033_3112, w_033_3113, w_033_3114, w_033_3115, w_033_3117, w_033_3118, w_033_3119, w_033_3120, w_033_3121, w_033_3122, w_033_3124, w_033_3125, w_033_3126, w_033_3128, w_033_3130, w_033_3131, w_033_3132, w_033_3133, w_033_3134, w_033_3135, w_033_3136, w_033_3137, w_033_3140, w_033_3141, w_033_3144, w_033_3146, w_033_3147, w_033_3148, w_033_3149, w_033_3150, w_033_3151, w_033_3152, w_033_3153, w_033_3154, w_033_3155, w_033_3157, w_033_3158, w_033_3159, w_033_3160, w_033_3162, w_033_3163, w_033_3164, w_033_3165, w_033_3166, w_033_3167, w_033_3168, w_033_3169, w_033_3170, w_033_3171, w_033_3172, w_033_3173, w_033_3175, w_033_3176, w_033_3177, w_033_3178, w_033_3180, w_033_3181, w_033_3182, w_033_3183, w_033_3184, w_033_3185, w_033_3186, w_033_3188, w_033_3189, w_033_3191, w_033_3192, w_033_3193, w_033_3194, w_033_3196, w_033_3197, w_033_3198, w_033_3199, w_033_3200, w_033_3201, w_033_3202, w_033_3204, w_033_3205, w_033_3206, w_033_3207, w_033_3208, w_033_3210, w_033_3212, w_033_3214, w_033_3216, w_033_3217, w_033_3218, w_033_3219, w_033_3220, w_033_3221, w_033_3222, w_033_3223, w_033_3225, w_033_3226, w_033_3227, w_033_3228, w_033_3229, w_033_3230, w_033_3231, w_033_3233, w_033_3234, w_033_3236, w_033_3237, w_033_3238, w_033_3239, w_033_3242, w_033_3243, w_033_3244, w_033_3246, w_033_3247, w_033_3249, w_033_3250, w_033_3251, w_033_3252, w_033_3253, w_033_3254, w_033_3255, w_033_3257, w_033_3258, w_033_3259, w_033_3262, w_033_3264, w_033_3266, w_033_3267, w_033_3268, w_033_3270, w_033_3272, w_033_3273, w_033_3275, w_033_3276, w_033_3277, w_033_3278, w_033_3279, w_033_3280, w_033_3281, w_033_3282, w_033_3283, w_033_3284, w_033_3285, w_033_3286, w_033_3289, w_033_3290, w_033_3292, w_033_3293, w_033_3295, w_033_3298, w_033_3299, w_033_3301, w_033_3302, w_033_3304, w_033_3305, w_033_3306, w_033_3307, w_033_3309, w_033_3310, w_033_3311, w_033_3312, w_033_3314, w_033_3315, w_033_3317, w_033_3319, w_033_3320, w_033_3322, w_033_3323, w_033_3324, w_033_3325, w_033_3327, w_033_3328, w_033_3331, w_033_3332, w_033_3333, w_033_3334, w_033_3335, w_033_3336, w_033_3338, w_033_3339, w_033_3340, w_033_3341, w_033_3342, w_033_3345, w_033_3348, w_033_3349, w_033_3351, w_033_3352, w_033_3353, w_033_3354, w_033_3355, w_033_3356, w_033_3357, w_033_3358, w_033_3359, w_033_3360, w_033_3361, w_033_3362, w_033_3363, w_033_3364, w_033_3365, w_033_3366, w_033_3368, w_033_3369, w_033_3370, w_033_3371, w_033_3372, w_033_3373, w_033_3374, w_033_3375, w_033_3376, w_033_3377, w_033_3378, w_033_3379, w_033_3380, w_033_3383, w_033_3384, w_033_3385, w_033_3387, w_033_3389, w_033_3390, w_033_3391, w_033_3392, w_033_3395, w_033_3396, w_033_3397, w_033_3398, w_033_3399, w_033_3400, w_033_3402, w_033_3403, w_033_3404, w_033_3405, w_033_3407, w_033_3408, w_033_3409, w_033_3410, w_033_3411, w_033_3412, w_033_3413, w_033_3414, w_033_3415, w_033_3417, w_033_3418, w_033_3420, w_033_3421, w_033_3423, w_033_3424, w_033_3425, w_033_3426, w_033_3428, w_033_3430, w_033_3431, w_033_3432, w_033_3433, w_033_3434, w_033_3435, w_033_3438, w_033_3439, w_033_3440, w_033_3441, w_033_3442, w_033_3443, w_033_3444, w_033_3445, w_033_3446, w_033_3448, w_033_3449, w_033_3450, w_033_3452, w_033_3454, w_033_3455, w_033_3457, w_033_3458, w_033_3459, w_033_3460, w_033_3461, w_033_3462, w_033_3463, w_033_3464, w_033_3465, w_033_3466, w_033_3467, w_033_3468, w_033_3470, w_033_3471, w_033_3472, w_033_3473, w_033_3474, w_033_3475, w_033_3476, w_033_3477, w_033_3478, w_033_3480, w_033_3481, w_033_3482, w_033_3483, w_033_3486, w_033_3487, w_033_3488, w_033_3489, w_033_3490, w_033_3492, w_033_3493, w_033_3495, w_033_3496, w_033_3497, w_033_3499, w_033_3500, w_033_3501, w_033_3502, w_033_3503, w_033_3505, w_033_3506, w_033_3507, w_033_3508, w_033_3509, w_033_3511, w_033_3513, w_033_3514, w_033_3515, w_033_3516, w_033_3517, w_033_3518, w_033_3519, w_033_3520, w_033_3521, w_033_3522, w_033_3523, w_033_3524, w_033_3526, w_033_3527, w_033_3528, w_033_3529, w_033_3530, w_033_3532, w_033_3533, w_033_3534, w_033_3535, w_033_3536, w_033_3537, w_033_3538, w_033_3539, w_033_3540, w_033_3541, w_033_3542, w_033_3543, w_033_3544, w_033_3549, w_033_3551, w_033_3552, w_033_3553, w_033_3554, w_033_3555, w_033_3556, w_033_3557, w_033_3559, w_033_3560, w_033_3561, w_033_3562, w_033_3565, w_033_3566, w_033_3567, w_033_3569, w_033_3571, w_033_3573, w_033_3574, w_033_3575, w_033_3576, w_033_3577, w_033_3578, w_033_3579, w_033_3580, w_033_3581, w_033_3583, w_033_3584, w_033_3586, w_033_3587, w_033_3588, w_033_3589, w_033_3593, w_033_3594, w_033_3596, w_033_3597, w_033_3598, w_033_3599, w_033_3600, w_033_3601, w_033_3602, w_033_3603, w_033_3605, w_033_3606, w_033_3607, w_033_3608, w_033_3609, w_033_3610, w_033_3611, w_033_3613, w_033_3614, w_033_3616, w_033_3618, w_033_3620, w_033_3621, w_033_3622, w_033_3623, w_033_3624, w_033_3625, w_033_3626, w_033_3629, w_033_3630, w_033_3631, w_033_3632, w_033_3633, w_033_3634, w_033_3635, w_033_3638, w_033_3639, w_033_3640;
  wire w_034_000, w_034_001, w_034_002, w_034_003, w_034_004, w_034_005, w_034_006, w_034_007, w_034_008, w_034_011, w_034_012, w_034_013, w_034_014, w_034_015, w_034_016, w_034_017, w_034_018, w_034_019, w_034_020, w_034_021, w_034_022, w_034_024, w_034_025, w_034_026, w_034_027, w_034_028, w_034_029, w_034_030, w_034_031, w_034_032, w_034_033, w_034_035, w_034_036, w_034_037, w_034_038, w_034_039, w_034_040, w_034_041, w_034_043, w_034_047, w_034_048, w_034_049, w_034_050, w_034_051, w_034_052, w_034_053, w_034_054, w_034_055, w_034_056, w_034_057, w_034_058, w_034_060, w_034_061, w_034_062, w_034_063, w_034_064, w_034_065, w_034_066, w_034_067, w_034_069, w_034_070, w_034_071, w_034_072, w_034_073, w_034_074, w_034_077, w_034_078, w_034_080, w_034_082, w_034_083, w_034_085, w_034_086, w_034_087, w_034_089, w_034_090, w_034_093, w_034_094, w_034_095, w_034_097, w_034_098, w_034_099, w_034_100, w_034_101, w_034_102, w_034_103, w_034_104, w_034_105, w_034_106, w_034_107, w_034_108, w_034_109, w_034_110, w_034_111, w_034_112, w_034_113, w_034_114, w_034_115, w_034_117, w_034_118, w_034_119, w_034_120, w_034_121, w_034_124, w_034_125, w_034_126, w_034_127, w_034_128, w_034_130, w_034_131, w_034_134, w_034_135, w_034_136, w_034_137, w_034_138, w_034_141, w_034_142, w_034_143, w_034_144, w_034_145, w_034_146, w_034_147, w_034_148, w_034_149, w_034_150, w_034_152, w_034_155, w_034_156, w_034_159, w_034_160, w_034_161, w_034_162, w_034_163, w_034_164, w_034_165, w_034_166, w_034_167, w_034_169, w_034_170, w_034_171, w_034_173, w_034_174, w_034_175, w_034_176, w_034_177, w_034_178, w_034_179, w_034_180, w_034_181, w_034_182, w_034_184, w_034_185, w_034_187, w_034_188, w_034_189, w_034_190, w_034_191, w_034_193, w_034_194, w_034_196, w_034_197, w_034_198, w_034_199, w_034_200, w_034_201, w_034_202, w_034_203, w_034_204, w_034_205, w_034_206, w_034_207, w_034_208, w_034_210, w_034_211, w_034_212, w_034_213, w_034_214, w_034_215, w_034_217, w_034_218, w_034_219, w_034_220, w_034_221, w_034_222, w_034_223, w_034_225, w_034_226, w_034_227, w_034_229, w_034_230, w_034_231, w_034_233, w_034_235, w_034_236, w_034_239, w_034_240, w_034_241, w_034_242, w_034_243, w_034_244, w_034_245, w_034_246, w_034_248, w_034_249, w_034_250, w_034_252, w_034_254, w_034_255, w_034_256, w_034_257, w_034_260, w_034_261, w_034_262, w_034_263, w_034_264, w_034_265, w_034_269, w_034_270, w_034_271, w_034_272, w_034_273, w_034_274, w_034_275, w_034_276, w_034_278, w_034_279, w_034_280, w_034_281, w_034_282, w_034_283, w_034_285, w_034_287, w_034_288, w_034_289, w_034_290, w_034_291, w_034_292, w_034_295, w_034_296, w_034_297, w_034_298, w_034_300, w_034_301, w_034_302, w_034_304, w_034_305, w_034_306, w_034_307, w_034_308, w_034_309, w_034_310, w_034_312, w_034_313, w_034_315, w_034_317, w_034_318, w_034_319, w_034_321, w_034_323, w_034_324, w_034_325, w_034_326, w_034_327, w_034_328, w_034_329, w_034_330, w_034_331, w_034_332, w_034_333, w_034_335, w_034_337, w_034_338, w_034_339, w_034_340, w_034_341, w_034_342, w_034_343, w_034_344, w_034_346, w_034_347, w_034_349, w_034_350, w_034_351, w_034_352, w_034_353, w_034_354, w_034_356, w_034_359, w_034_360, w_034_361, w_034_362, w_034_363, w_034_365, w_034_367, w_034_369, w_034_370, w_034_372, w_034_373, w_034_374, w_034_375, w_034_376, w_034_377, w_034_379, w_034_381, w_034_382, w_034_383, w_034_385, w_034_386, w_034_387, w_034_388, w_034_389, w_034_390, w_034_391, w_034_393, w_034_394, w_034_395, w_034_397, w_034_403, w_034_404, w_034_405, w_034_406, w_034_408, w_034_410, w_034_412, w_034_413, w_034_414, w_034_416, w_034_417, w_034_418, w_034_419, w_034_421, w_034_422, w_034_423, w_034_426, w_034_427, w_034_428, w_034_430, w_034_431, w_034_432, w_034_433, w_034_434, w_034_436, w_034_437, w_034_440, w_034_442, w_034_443, w_034_445, w_034_447, w_034_448, w_034_449, w_034_451, w_034_452, w_034_453, w_034_454, w_034_455, w_034_456, w_034_457, w_034_458, w_034_459, w_034_460, w_034_461, w_034_462, w_034_463, w_034_464, w_034_466, w_034_467, w_034_468, w_034_469, w_034_470, w_034_471, w_034_472, w_034_476, w_034_477, w_034_478, w_034_479, w_034_480, w_034_481, w_034_482, w_034_483, w_034_484, w_034_487, w_034_488, w_034_489, w_034_491, w_034_492, w_034_493, w_034_494, w_034_497, w_034_498, w_034_499, w_034_501, w_034_502, w_034_504, w_034_505, w_034_506, w_034_507, w_034_508, w_034_510, w_034_511, w_034_512, w_034_513, w_034_514, w_034_515, w_034_516, w_034_517, w_034_519, w_034_521, w_034_522, w_034_523, w_034_524, w_034_525, w_034_527, w_034_529, w_034_530, w_034_531, w_034_532, w_034_533, w_034_534, w_034_535, w_034_536, w_034_538, w_034_539, w_034_540, w_034_541, w_034_542, w_034_543, w_034_544, w_034_545, w_034_546, w_034_547, w_034_548, w_034_549, w_034_550, w_034_551, w_034_552, w_034_554, w_034_555, w_034_557, w_034_558, w_034_559, w_034_560, w_034_561, w_034_564, w_034_565, w_034_566, w_034_568, w_034_569, w_034_573, w_034_574, w_034_575, w_034_576, w_034_578, w_034_580, w_034_581, w_034_582, w_034_583, w_034_584, w_034_585, w_034_586, w_034_587, w_034_588, w_034_589, w_034_590, w_034_592, w_034_593, w_034_594, w_034_596, w_034_597, w_034_598, w_034_599, w_034_601, w_034_603, w_034_605, w_034_607, w_034_609, w_034_610, w_034_612, w_034_613, w_034_614, w_034_615, w_034_616, w_034_617, w_034_619, w_034_620, w_034_621, w_034_622, w_034_623, w_034_624, w_034_626, w_034_628, w_034_629, w_034_630, w_034_631, w_034_632, w_034_634, w_034_636, w_034_638, w_034_639, w_034_640, w_034_641, w_034_643, w_034_644, w_034_645, w_034_647, w_034_648, w_034_649, w_034_650, w_034_651, w_034_654, w_034_655, w_034_656, w_034_657, w_034_658, w_034_659, w_034_660, w_034_661, w_034_662, w_034_664, w_034_665, w_034_666, w_034_667, w_034_668, w_034_669, w_034_670, w_034_671, w_034_672, w_034_674, w_034_675, w_034_676, w_034_679, w_034_680, w_034_681, w_034_682, w_034_684, w_034_686, w_034_687, w_034_688, w_034_690, w_034_691, w_034_692, w_034_694, w_034_695, w_034_697, w_034_698, w_034_699, w_034_700, w_034_701, w_034_702, w_034_703, w_034_704, w_034_705, w_034_707, w_034_708, w_034_709, w_034_710, w_034_711, w_034_712, w_034_713, w_034_714, w_034_715, w_034_716, w_034_718, w_034_719, w_034_721, w_034_722, w_034_723, w_034_724, w_034_726, w_034_727, w_034_728, w_034_729, w_034_730, w_034_731, w_034_732, w_034_733, w_034_734, w_034_736, w_034_737, w_034_738, w_034_739, w_034_740, w_034_741, w_034_742, w_034_743, w_034_744, w_034_745, w_034_747, w_034_748, w_034_749, w_034_750, w_034_751, w_034_752, w_034_753, w_034_754, w_034_755, w_034_756, w_034_757, w_034_758, w_034_760, w_034_762, w_034_764, w_034_765, w_034_766, w_034_767, w_034_768, w_034_769, w_034_770, w_034_771, w_034_772, w_034_773, w_034_775, w_034_780, w_034_781, w_034_782, w_034_783, w_034_785, w_034_786, w_034_787, w_034_790, w_034_791, w_034_793, w_034_794, w_034_795, w_034_796, w_034_797, w_034_798, w_034_799, w_034_800, w_034_801, w_034_803, w_034_805, w_034_806, w_034_807, w_034_808, w_034_809, w_034_810, w_034_811, w_034_813, w_034_814, w_034_817, w_034_818, w_034_819, w_034_820, w_034_821, w_034_824, w_034_827, w_034_828, w_034_829, w_034_830, w_034_831, w_034_832, w_034_833, w_034_834, w_034_835, w_034_836, w_034_838, w_034_840, w_034_841, w_034_843, w_034_844, w_034_845, w_034_846, w_034_847, w_034_848, w_034_849, w_034_850, w_034_852, w_034_854, w_034_855, w_034_856, w_034_857, w_034_858, w_034_859, w_034_860, w_034_861, w_034_862, w_034_864, w_034_865, w_034_866, w_034_867, w_034_868, w_034_869, w_034_870, w_034_871, w_034_873, w_034_874, w_034_875, w_034_876, w_034_877, w_034_878, w_034_879, w_034_880, w_034_881, w_034_882, w_034_884, w_034_885, w_034_886, w_034_889, w_034_892, w_034_894, w_034_896, w_034_897, w_034_898, w_034_899, w_034_900, w_034_901, w_034_904, w_034_906, w_034_907, w_034_908, w_034_909, w_034_910, w_034_911, w_034_912, w_034_913, w_034_914, w_034_915, w_034_916, w_034_917, w_034_918, w_034_919, w_034_920, w_034_922, w_034_923, w_034_924, w_034_925, w_034_926, w_034_927, w_034_929, w_034_930, w_034_931, w_034_932, w_034_934, w_034_935, w_034_936, w_034_937, w_034_939, w_034_940, w_034_943, w_034_944, w_034_945, w_034_946, w_034_949, w_034_950, w_034_951, w_034_952, w_034_953, w_034_954, w_034_955, w_034_957, w_034_959, w_034_961, w_034_962, w_034_963, w_034_964, w_034_965, w_034_967, w_034_968, w_034_969, w_034_970, w_034_973, w_034_974, w_034_975, w_034_976, w_034_977, w_034_981, w_034_982, w_034_984, w_034_986, w_034_987, w_034_988, w_034_990, w_034_991, w_034_992, w_034_995, w_034_996, w_034_997, w_034_999, w_034_1000, w_034_1001, w_034_1002, w_034_1003, w_034_1004, w_034_1006, w_034_1007, w_034_1008, w_034_1009, w_034_1012, w_034_1013, w_034_1014, w_034_1015, w_034_1016, w_034_1017, w_034_1018, w_034_1019, w_034_1020, w_034_1021, w_034_1022, w_034_1023, w_034_1024, w_034_1025, w_034_1026, w_034_1027, w_034_1029, w_034_1030, w_034_1031, w_034_1033, w_034_1034, w_034_1035, w_034_1037, w_034_1038, w_034_1039, w_034_1040, w_034_1041, w_034_1042, w_034_1043, w_034_1044, w_034_1045, w_034_1046, w_034_1047, w_034_1048, w_034_1049, w_034_1051, w_034_1053, w_034_1056, w_034_1057, w_034_1058, w_034_1059, w_034_1060, w_034_1061, w_034_1063, w_034_1064, w_034_1065, w_034_1066, w_034_1067, w_034_1068, w_034_1069, w_034_1070, w_034_1071, w_034_1074, w_034_1075, w_034_1076, w_034_1077, w_034_1078, w_034_1079, w_034_1082, w_034_1083, w_034_1084, w_034_1085, w_034_1086, w_034_1089, w_034_1090, w_034_1091, w_034_1092, w_034_1093, w_034_1094, w_034_1096, w_034_1097, w_034_1098, w_034_1100, w_034_1104, w_034_1105, w_034_1107, w_034_1108, w_034_1109, w_034_1110, w_034_1111, w_034_1112, w_034_1114, w_034_1115, w_034_1116, w_034_1117, w_034_1118, w_034_1119, w_034_1120, w_034_1123, w_034_1125, w_034_1126, w_034_1127, w_034_1128, w_034_1129, w_034_1130, w_034_1131, w_034_1132, w_034_1133, w_034_1135, w_034_1137, w_034_1138, w_034_1139, w_034_1141, w_034_1143, w_034_1144, w_034_1145, w_034_1146, w_034_1148, w_034_1150, w_034_1152, w_034_1153, w_034_1154, w_034_1156, w_034_1159, w_034_1162, w_034_1166, w_034_1170, w_034_1172, w_034_1173, w_034_1174, w_034_1175, w_034_1176, w_034_1178, w_034_1180, w_034_1181, w_034_1182, w_034_1184, w_034_1185, w_034_1187, w_034_1188, w_034_1189, w_034_1190, w_034_1191, w_034_1192, w_034_1193, w_034_1194, w_034_1195, w_034_1196, w_034_1198, w_034_1199, w_034_1200, w_034_1201, w_034_1202, w_034_1205, w_034_1206, w_034_1207, w_034_1208, w_034_1209, w_034_1210, w_034_1211, w_034_1212, w_034_1213, w_034_1214, w_034_1216, w_034_1217, w_034_1218, w_034_1220, w_034_1221, w_034_1223, w_034_1224, w_034_1225, w_034_1226, w_034_1227, w_034_1229, w_034_1231, w_034_1234, w_034_1235, w_034_1238, w_034_1239, w_034_1240, w_034_1241, w_034_1242, w_034_1243, w_034_1244, w_034_1245, w_034_1247, w_034_1248, w_034_1249, w_034_1250, w_034_1252, w_034_1253, w_034_1254, w_034_1255, w_034_1256, w_034_1258, w_034_1259, w_034_1260, w_034_1261, w_034_1262, w_034_1265, w_034_1267, w_034_1268, w_034_1269, w_034_1271, w_034_1272, w_034_1274, w_034_1275, w_034_1276, w_034_1277, w_034_1278, w_034_1279, w_034_1281, w_034_1282, w_034_1283, w_034_1284, w_034_1285, w_034_1287, w_034_1288, w_034_1291, w_034_1292, w_034_1294, w_034_1295, w_034_1296, w_034_1297, w_034_1300, w_034_1303, w_034_1305, w_034_1306, w_034_1307, w_034_1308, w_034_1309, w_034_1310, w_034_1311, w_034_1312, w_034_1313, w_034_1314, w_034_1315, w_034_1316, w_034_1317, w_034_1318, w_034_1319, w_034_1320, w_034_1322, w_034_1323, w_034_1324, w_034_1325, w_034_1326, w_034_1327, w_034_1328, w_034_1329, w_034_1330, w_034_1331, w_034_1332, w_034_1333, w_034_1334, w_034_1335, w_034_1336, w_034_1337, w_034_1338, w_034_1339, w_034_1340, w_034_1341, w_034_1342, w_034_1343, w_034_1345, w_034_1346, w_034_1347, w_034_1348, w_034_1349, w_034_1351, w_034_1352, w_034_1353, w_034_1354, w_034_1355, w_034_1356, w_034_1357, w_034_1358, w_034_1359, w_034_1362, w_034_1363, w_034_1365, w_034_1366, w_034_1367, w_034_1368, w_034_1370, w_034_1371, w_034_1372, w_034_1373, w_034_1375, w_034_1376, w_034_1377, w_034_1378, w_034_1379, w_034_1380, w_034_1381, w_034_1382, w_034_1385, w_034_1386, w_034_1387, w_034_1388, w_034_1389, w_034_1390, w_034_1391, w_034_1392, w_034_1393, w_034_1394, w_034_1395, w_034_1396, w_034_1397, w_034_1398, w_034_1399, w_034_1400, w_034_1401, w_034_1404, w_034_1405, w_034_1408, w_034_1409, w_034_1411, w_034_1413, w_034_1414, w_034_1417, w_034_1418, w_034_1419, w_034_1420, w_034_1421, w_034_1422, w_034_1424, w_034_1426, w_034_1427, w_034_1428, w_034_1429, w_034_1430, w_034_1431, w_034_1432, w_034_1434, w_034_1435, w_034_1436, w_034_1437, w_034_1438, w_034_1439, w_034_1441, w_034_1442, w_034_1443, w_034_1444, w_034_1445, w_034_1446, w_034_1448, w_034_1449, w_034_1450, w_034_1451, w_034_1452, w_034_1453, w_034_1454, w_034_1455, w_034_1457, w_034_1458, w_034_1459, w_034_1460, w_034_1461, w_034_1462, w_034_1463, w_034_1466, w_034_1469, w_034_1470, w_034_1471, w_034_1472, w_034_1473, w_034_1474, w_034_1475, w_034_1477, w_034_1479, w_034_1480, w_034_1481, w_034_1482, w_034_1484, w_034_1485, w_034_1486, w_034_1487, w_034_1488, w_034_1489, w_034_1490, w_034_1492, w_034_1494, w_034_1495, w_034_1496, w_034_1497, w_034_1499, w_034_1500, w_034_1501, w_034_1502, w_034_1503, w_034_1504, w_034_1505, w_034_1506, w_034_1507, w_034_1508, w_034_1509, w_034_1510, w_034_1511, w_034_1512, w_034_1513, w_034_1514, w_034_1515, w_034_1516, w_034_1517, w_034_1518, w_034_1519, w_034_1522, w_034_1524, w_034_1525, w_034_1526, w_034_1529, w_034_1530, w_034_1531, w_034_1532, w_034_1533, w_034_1534, w_034_1536, w_034_1537, w_034_1538, w_034_1539, w_034_1541, w_034_1542, w_034_1543, w_034_1546, w_034_1547, w_034_1548, w_034_1549, w_034_1550, w_034_1553, w_034_1554, w_034_1555, w_034_1556, w_034_1557, w_034_1558, w_034_1559, w_034_1561, w_034_1562, w_034_1564, w_034_1565, w_034_1566, w_034_1567, w_034_1568, w_034_1569, w_034_1570, w_034_1571, w_034_1572, w_034_1573, w_034_1574, w_034_1576, w_034_1577, w_034_1578, w_034_1579, w_034_1580, w_034_1581, w_034_1582, w_034_1583, w_034_1584, w_034_1586, w_034_1587, w_034_1588, w_034_1589, w_034_1590, w_034_1592, w_034_1593, w_034_1594, w_034_1595, w_034_1596, w_034_1600, w_034_1602, w_034_1603, w_034_1605, w_034_1606, w_034_1607, w_034_1609, w_034_1612, w_034_1613, w_034_1615, w_034_1617, w_034_1619, w_034_1620, w_034_1621, w_034_1622, w_034_1624, w_034_1625, w_034_1626, w_034_1627, w_034_1628, w_034_1629, w_034_1630, w_034_1631, w_034_1632, w_034_1634, w_034_1635, w_034_1637, w_034_1638, w_034_1639, w_034_1640, w_034_1641, w_034_1643, w_034_1644, w_034_1645, w_034_1646, w_034_1647, w_034_1648, w_034_1649, w_034_1651, w_034_1652, w_034_1653, w_034_1654, w_034_1655, w_034_1656, w_034_1658, w_034_1659, w_034_1660, w_034_1661, w_034_1662, w_034_1667, w_034_1670, w_034_1671, w_034_1672, w_034_1673, w_034_1674, w_034_1675, w_034_1676, w_034_1677, w_034_1678, w_034_1680, w_034_1681, w_034_1682, w_034_1684, w_034_1685, w_034_1686, w_034_1687, w_034_1688, w_034_1689, w_034_1690, w_034_1691, w_034_1692, w_034_1693, w_034_1698, w_034_1699, w_034_1700, w_034_1701, w_034_1702, w_034_1703, w_034_1704, w_034_1705, w_034_1706, w_034_1707, w_034_1708, w_034_1710, w_034_1711, w_034_1712, w_034_1713, w_034_1714, w_034_1715, w_034_1716, w_034_1717, w_034_1718, w_034_1719, w_034_1721, w_034_1722, w_034_1723, w_034_1724, w_034_1725, w_034_1727, w_034_1728, w_034_1729, w_034_1731, w_034_1732, w_034_1734, w_034_1735, w_034_1737, w_034_1739, w_034_1740, w_034_1741, w_034_1742, w_034_1743, w_034_1744, w_034_1745, w_034_1746, w_034_1747, w_034_1749, w_034_1750, w_034_1751, w_034_1752, w_034_1753, w_034_1754, w_034_1757, w_034_1758, w_034_1760, w_034_1761, w_034_1762, w_034_1763, w_034_1764, w_034_1766, w_034_1768, w_034_1770, w_034_1772, w_034_1773, w_034_1774, w_034_1775, w_034_1776, w_034_1777, w_034_1778, w_034_1779, w_034_1780, w_034_1784, w_034_1786, w_034_1787, w_034_1789, w_034_1791, w_034_1793, w_034_1794, w_034_1796, w_034_1797, w_034_1799, w_034_1800, w_034_1801, w_034_1802, w_034_1803, w_034_1804, w_034_1806, w_034_1807, w_034_1808, w_034_1810, w_034_1813, w_034_1814, w_034_1815, w_034_1816, w_034_1817, w_034_1818, w_034_1819, w_034_1820, w_034_1821, w_034_1823, w_034_1824, w_034_1825, w_034_1827, w_034_1828, w_034_1830, w_034_1831, w_034_1835, w_034_1836, w_034_1837, w_034_1840, w_034_1841, w_034_1844, w_034_1845, w_034_1848, w_034_1849, w_034_1850, w_034_1851, w_034_1852, w_034_1855, w_034_1856, w_034_1857, w_034_1858, w_034_1859, w_034_1860, w_034_1861, w_034_1862, w_034_1863, w_034_1864, w_034_1865, w_034_1867, w_034_1868, w_034_1870, w_034_1871, w_034_1872, w_034_1874, w_034_1875, w_034_1876, w_034_1878, w_034_1880, w_034_1881, w_034_1883, w_034_1886, w_034_1887, w_034_1888, w_034_1890, w_034_1891, w_034_1892, w_034_1893, w_034_1895, w_034_1896, w_034_1897, w_034_1898, w_034_1899, w_034_1900, w_034_1901, w_034_1902, w_034_1903, w_034_1904, w_034_1905, w_034_1908, w_034_1910, w_034_1911, w_034_1913, w_034_1914, w_034_1915, w_034_1916, w_034_1918, w_034_1919, w_034_1921, w_034_1922, w_034_1923, w_034_1924, w_034_1930, w_034_1931, w_034_1932, w_034_1933, w_034_1934, w_034_1935, w_034_1937, w_034_1938, w_034_1940, w_034_1941, w_034_1946, w_034_1947, w_034_1949, w_034_1950, w_034_1951, w_034_1953, w_034_1954, w_034_1955, w_034_1956, w_034_1957, w_034_1960, w_034_1962, w_034_1963, w_034_1964, w_034_1965, w_034_1966, w_034_1967, w_034_1968, w_034_1969, w_034_1971, w_034_1972, w_034_1973, w_034_1974, w_034_1975, w_034_1976, w_034_1977, w_034_1978, w_034_1980, w_034_1981, w_034_1982, w_034_1984, w_034_1985, w_034_1986, w_034_1987, w_034_1990, w_034_1992, w_034_1993, w_034_1995, w_034_1997, w_034_1998, w_034_1999, w_034_2002, w_034_2004, w_034_2005, w_034_2006, w_034_2007, w_034_2008, w_034_2009, w_034_2012, w_034_2013, w_034_2015, w_034_2017, w_034_2018, w_034_2019, w_034_2023, w_034_2025, w_034_2026, w_034_2027, w_034_2029, w_034_2030, w_034_2031, w_034_2032, w_034_2033, w_034_2034, w_034_2035, w_034_2036, w_034_2038, w_034_2039, w_034_2040, w_034_2041, w_034_2042, w_034_2043, w_034_2044, w_034_2045, w_034_2046, w_034_2047, w_034_2048, w_034_2051, w_034_2052, w_034_2053, w_034_2054, w_034_2056, w_034_2057, w_034_2061, w_034_2062, w_034_2063, w_034_2065, w_034_2068, w_034_2069, w_034_2070, w_034_2071, w_034_2072, w_034_2075, w_034_2076, w_034_2077, w_034_2078, w_034_2079, w_034_2080, w_034_2081, w_034_2082, w_034_2083, w_034_2084, w_034_2085, w_034_2086, w_034_2087, w_034_2088, w_034_2089, w_034_2090, w_034_2091, w_034_2092, w_034_2093, w_034_2094, w_034_2095, w_034_2097, w_034_2098, w_034_2099, w_034_2101, w_034_2102, w_034_2103, w_034_2104, w_034_2105, w_034_2106, w_034_2107, w_034_2108, w_034_2109, w_034_2110, w_034_2111, w_034_2112, w_034_2113, w_034_2114, w_034_2115, w_034_2116, w_034_2117, w_034_2118, w_034_2120, w_034_2121, w_034_2122, w_034_2124, w_034_2125, w_034_2126, w_034_2128, w_034_2129, w_034_2130, w_034_2131, w_034_2132, w_034_2134, w_034_2135, w_034_2136, w_034_2139, w_034_2140, w_034_2141, w_034_2142, w_034_2143, w_034_2144, w_034_2145, w_034_2146, w_034_2148, w_034_2150, w_034_2151, w_034_2152, w_034_2154, w_034_2155, w_034_2156, w_034_2158, w_034_2159, w_034_2160, w_034_2161, w_034_2162, w_034_2163, w_034_2164, w_034_2165, w_034_2167, w_034_2168, w_034_2169, w_034_2170, w_034_2171, w_034_2172, w_034_2173, w_034_2176, w_034_2177, w_034_2178, w_034_2179, w_034_2180, w_034_2181, w_034_2182, w_034_2183, w_034_2184, w_034_2186, w_034_2187, w_034_2188, w_034_2189, w_034_2190, w_034_2191, w_034_2192, w_034_2194, w_034_2195, w_034_2196, w_034_2199, w_034_2201, w_034_2202, w_034_2203, w_034_2204, w_034_2206, w_034_2208, w_034_2210, w_034_2211, w_034_2212, w_034_2213, w_034_2215, w_034_2216, w_034_2217, w_034_2218, w_034_2219, w_034_2221, w_034_2223, w_034_2224, w_034_2227, w_034_2228, w_034_2229, w_034_2230, w_034_2234, w_034_2235, w_034_2236, w_034_2237, w_034_2238, w_034_2240, w_034_2241, w_034_2242, w_034_2243, w_034_2245, w_034_2246, w_034_2247, w_034_2248, w_034_2253, w_034_2254, w_034_2255, w_034_2256, w_034_2257, w_034_2258, w_034_2259, w_034_2261, w_034_2262, w_034_2263, w_034_2265, w_034_2266, w_034_2267, w_034_2268, w_034_2269, w_034_2270, w_034_2271, w_034_2272, w_034_2273, w_034_2274, w_034_2275, w_034_2276, w_034_2277, w_034_2278, w_034_2279, w_034_2282, w_034_2283, w_034_2284, w_034_2285, w_034_2286, w_034_2287, w_034_2288, w_034_2289, w_034_2290, w_034_2291, w_034_2292, w_034_2293, w_034_2294, w_034_2296, w_034_2297, w_034_2298, w_034_2299, w_034_2300, w_034_2301, w_034_2302, w_034_2303, w_034_2304, w_034_2305, w_034_2306, w_034_2307, w_034_2308, w_034_2309, w_034_2311, w_034_2312, w_034_2313, w_034_2314, w_034_2316, w_034_2317, w_034_2318, w_034_2320, w_034_2321, w_034_2322, w_034_2324, w_034_2325, w_034_2326, w_034_2327, w_034_2328, w_034_2329, w_034_2332, w_034_2334, w_034_2335, w_034_2336, w_034_2337, w_034_2339, w_034_2340, w_034_2341, w_034_2342, w_034_2343, w_034_2344, w_034_2345, w_034_2346, w_034_2348, w_034_2351, w_034_2352, w_034_2353, w_034_2354, w_034_2356, w_034_2357, w_034_2359, w_034_2360, w_034_2361, w_034_2362, w_034_2363, w_034_2364, w_034_2365, w_034_2366, w_034_2368, w_034_2369, w_034_2370, w_034_2373, w_034_2374, w_034_2375, w_034_2377, w_034_2378, w_034_2379, w_034_2380, w_034_2381, w_034_2382, w_034_2383, w_034_2384, w_034_2385, w_034_2386, w_034_2387, w_034_2389, w_034_2390, w_034_2391, w_034_2392, w_034_2394, w_034_2395, w_034_2396, w_034_2397, w_034_2398, w_034_2399, w_034_2400, w_034_2401, w_034_2402, w_034_2403, w_034_2405, w_034_2406, w_034_2407, w_034_2408, w_034_2410, w_034_2412, w_034_2413, w_034_2414, w_034_2415, w_034_2416, w_034_2417, w_034_2419, w_034_2420, w_034_2421, w_034_2424, w_034_2426, w_034_2428, w_034_2429, w_034_2430, w_034_2434, w_034_2435, w_034_2436, w_034_2437, w_034_2438, w_034_2439, w_034_2440, w_034_2441, w_034_2443, w_034_2444, w_034_2446, w_034_2447, w_034_2449, w_034_2450, w_034_2451, w_034_2452, w_034_2453, w_034_2454, w_034_2455, w_034_2456, w_034_2457, w_034_2459, w_034_2460, w_034_2462, w_034_2463, w_034_2464, w_034_2465, w_034_2466, w_034_2467, w_034_2468, w_034_2471, w_034_2472, w_034_2473, w_034_2475, w_034_2477, w_034_2478, w_034_2482, w_034_2483, w_034_2484, w_034_2486, w_034_2488, w_034_2489, w_034_2492, w_034_2493, w_034_2494, w_034_2495, w_034_2496, w_034_2497, w_034_2498, w_034_2501, w_034_2505, w_034_2506, w_034_2507, w_034_2508, w_034_2509, w_034_2510, w_034_2511, w_034_2512, w_034_2514, w_034_2515, w_034_2516, w_034_2517, w_034_2518, w_034_2519, w_034_2520, w_034_2521, w_034_2522, w_034_2523, w_034_2525, w_034_2527, w_034_2528, w_034_2529, w_034_2530, w_034_2531, w_034_2532, w_034_2533, w_034_2534, w_034_2535, w_034_2537, w_034_2538, w_034_2539, w_034_2540, w_034_2541, w_034_2544, w_034_2545, w_034_2546, w_034_2547, w_034_2548, w_034_2550, w_034_2551, w_034_2552, w_034_2553, w_034_2554, w_034_2557, w_034_2558, w_034_2560, w_034_2561, w_034_2562, w_034_2563, w_034_2564, w_034_2566, w_034_2567, w_034_2568, w_034_2569, w_034_2570, w_034_2571, w_034_2572, w_034_2573, w_034_2574, w_034_2575, w_034_2576, w_034_2577, w_034_2578, w_034_2579, w_034_2580, w_034_2582, w_034_2585, w_034_2586, w_034_2587, w_034_2588, w_034_2589, w_034_2591, w_034_2592, w_034_2593, w_034_2594, w_034_2595, w_034_2596, w_034_2598, w_034_2599, w_034_2601, w_034_2602, w_034_2603, w_034_2604, w_034_2605, w_034_2606, w_034_2607, w_034_2608, w_034_2609, w_034_2610, w_034_2611, w_034_2612, w_034_2613, w_034_2614, w_034_2615, w_034_2616, w_034_2617, w_034_2618, w_034_2619, w_034_2620, w_034_2621, w_034_2622, w_034_2623, w_034_2624, w_034_2625, w_034_2627, w_034_2628, w_034_2629, w_034_2630, w_034_2631, w_034_2632, w_034_2633, w_034_2634, w_034_2636, w_034_2637, w_034_2638, w_034_2639, w_034_2640, w_034_2641, w_034_2642, w_034_2644, w_034_2645, w_034_2647, w_034_2648, w_034_2649, w_034_2650, w_034_2651, w_034_2652, w_034_2653, w_034_2654, w_034_2655, w_034_2656, w_034_2658, w_034_2660, w_034_2663, w_034_2664, w_034_2665, w_034_2668, w_034_2669, w_034_2670, w_034_2671, w_034_2672, w_034_2673, w_034_2674, w_034_2675, w_034_2676, w_034_2677, w_034_2678, w_034_2679, w_034_2680, w_034_2682, w_034_2685, w_034_2686, w_034_2687, w_034_2688, w_034_2689, w_034_2690, w_034_2691, w_034_2692, w_034_2693, w_034_2694, w_034_2695, w_034_2697, w_034_2698, w_034_2699, w_034_2701, w_034_2702, w_034_2705, w_034_2708, w_034_2709, w_034_2710, w_034_2711, w_034_2713, w_034_2714, w_034_2715, w_034_2716, w_034_2717, w_034_2718, w_034_2719, w_034_2720, w_034_2721, w_034_2722, w_034_2726, w_034_2727, w_034_2729, w_034_2730, w_034_2731, w_034_2732, w_034_2733, w_034_2734, w_034_2735, w_034_2736, w_034_2737, w_034_2738, w_034_2739, w_034_2740, w_034_2742, w_034_2743, w_034_2744, w_034_2745, w_034_2746, w_034_2749, w_034_2750, w_034_2751, w_034_2752, w_034_2753, w_034_2754, w_034_2755, w_034_2757, w_034_2758, w_034_2759, w_034_2760, w_034_2761, w_034_2762, w_034_2763, w_034_2764, w_034_2766, w_034_2767, w_034_2768, w_034_2769, w_034_2770, w_034_2771, w_034_2773, w_034_2774, w_034_2775, w_034_2776, w_034_2777, w_034_2778, w_034_2781, w_034_2782, w_034_2783, w_034_2784, w_034_2785, w_034_2786, w_034_2787, w_034_2788, w_034_2789, w_034_2790, w_034_2791, w_034_2792, w_034_2793, w_034_2794, w_034_2795, w_034_2796, w_034_2797, w_034_2798, w_034_2799, w_034_2800, w_034_2801, w_034_2802, w_034_2803, w_034_2804, w_034_2805, w_034_2807, w_034_2808, w_034_2809, w_034_2810, w_034_2811, w_034_2812, w_034_2813, w_034_2814, w_034_2815, w_034_2816, w_034_2817, w_034_2818, w_034_2819, w_034_2820, w_034_2821, w_034_2822, w_034_2823, w_034_2825, w_034_2826, w_034_2827, w_034_2828, w_034_2829, w_034_2830, w_034_2831, w_034_2832, w_034_2833, w_034_2834, w_034_2835, w_034_2836, w_034_2837, w_034_2838, w_034_2839, w_034_2841, w_034_2842, w_034_2843, w_034_2845, w_034_2846, w_034_2847, w_034_2848, w_034_2850, w_034_2851, w_034_2854, w_034_2855, w_034_2857, w_034_2858, w_034_2859, w_034_2860, w_034_2861, w_034_2862, w_034_2863, w_034_2864, w_034_2865, w_034_2866, w_034_2868, w_034_2869, w_034_2870, w_034_2872, w_034_2874, w_034_2875, w_034_2878, w_034_2880, w_034_2881, w_034_2882, w_034_2884, w_034_2885, w_034_2886, w_034_2888, w_034_2889, w_034_2890, w_034_2891, w_034_2892, w_034_2893, w_034_2895, w_034_2896, w_034_2897, w_034_2898, w_034_2899, w_034_2900, w_034_2901, w_034_2903, w_034_2906, w_034_2907, w_034_2909, w_034_2910, w_034_2911, w_034_2913, w_034_2916, w_034_2917, w_034_2918, w_034_2920, w_034_2921, w_034_2923, w_034_2924, w_034_2925, w_034_2927, w_034_2928, w_034_2929, w_034_2930, w_034_2931, w_034_2932, w_034_2933, w_034_2934, w_034_2935, w_034_2937, w_034_2939, w_034_2941, w_034_2942, w_034_2943, w_034_2944, w_034_2945, w_034_2946, w_034_2947, w_034_2948, w_034_2949, w_034_2950, w_034_2951, w_034_2952, w_034_2953, w_034_2954, w_034_2955, w_034_2956, w_034_2959, w_034_2960, w_034_2963, w_034_2964, w_034_2965, w_034_2966, w_034_2968, w_034_2969, w_034_2970, w_034_2972, w_034_2974, w_034_2976, w_034_2980, w_034_2981, w_034_2982, w_034_2983, w_034_2984, w_034_2985, w_034_2987, w_034_2988, w_034_2990, w_034_2991, w_034_2992, w_034_2993, w_034_2994, w_034_2995, w_034_2996, w_034_2997, w_034_2998, w_034_2999, w_034_3000, w_034_3001, w_034_3003, w_034_3004, w_034_3005, w_034_3006, w_034_3007, w_034_3008, w_034_3010, w_034_3011, w_034_3012, w_034_3013, w_034_3014, w_034_3015, w_034_3016, w_034_3017, w_034_3018, w_034_3019, w_034_3020, w_034_3021, w_034_3023, w_034_3025, w_034_3026, w_034_3027, w_034_3030, w_034_3031, w_034_3033, w_034_3034, w_034_3036, w_034_3037, w_034_3038, w_034_3039, w_034_3040, w_034_3042, w_034_3043, w_034_3045, w_034_3046, w_034_3048, w_034_3049, w_034_3050, w_034_3051, w_034_3053, w_034_3054, w_034_3055, w_034_3058, w_034_3059, w_034_3061, w_034_3062, w_034_3063, w_034_3065, w_034_3067, w_034_3068, w_034_3069, w_034_3070, w_034_3074, w_034_3076, w_034_3077, w_034_3078, w_034_3079, w_034_3083, w_034_3085, w_034_3086, w_034_3087, w_034_3088, w_034_3089, w_034_3091, w_034_3092, w_034_3093, w_034_3094, w_034_3095, w_034_3096, w_034_3097, w_034_3098, w_034_3100, w_034_3101, w_034_3102, w_034_3103, w_034_3104, w_034_3105, w_034_3107, w_034_3108, w_034_3109, w_034_3110, w_034_3112, w_034_3113, w_034_3114, w_034_3115, w_034_3116, w_034_3119, w_034_3120, w_034_3121, w_034_3122, w_034_3123, w_034_3124, w_034_3125, w_034_3126, w_034_3132, w_034_3133, w_034_3134, w_034_3135, w_034_3136, w_034_3137, w_034_3140, w_034_3141, w_034_3142, w_034_3143, w_034_3144, w_034_3145, w_034_3146, w_034_3148, w_034_3149, w_034_3150, w_034_3152, w_034_3153, w_034_3154, w_034_3155, w_034_3156, w_034_3158, w_034_3159, w_034_3161, w_034_3162, w_034_3163, w_034_3165, w_034_3166, w_034_3167, w_034_3168, w_034_3169, w_034_3170, w_034_3171, w_034_3172, w_034_3173, w_034_3174, w_034_3175, w_034_3176, w_034_3178, w_034_3181, w_034_3182, w_034_3183, w_034_3184, w_034_3185, w_034_3186, w_034_3188, w_034_3189, w_034_3191, w_034_3192, w_034_3193, w_034_3194, w_034_3196, w_034_3197, w_034_3199, w_034_3200, w_034_3201, w_034_3202, w_034_3204, w_034_3205, w_034_3207, w_034_3208, w_034_3209, w_034_3210, w_034_3211, w_034_3213, w_034_3214, w_034_3215, w_034_3216, w_034_3217, w_034_3219, w_034_3222, w_034_3223, w_034_3225, w_034_3227, w_034_3228, w_034_3230, w_034_3231, w_034_3232, w_034_3233, w_034_3234, w_034_3235, w_034_3236, w_034_3237, w_034_3239, w_034_3240, w_034_3241, w_034_3242, w_034_3243, w_034_3244, w_034_3245, w_034_3246, w_034_3247, w_034_3248, w_034_3249, w_034_3250, w_034_3251, w_034_3254, w_034_3256, w_034_3257, w_034_3258, w_034_3259, w_034_3260, w_034_3261, w_034_3262, w_034_3263, w_034_3264, w_034_3265, w_034_3266, w_034_3267, w_034_3269, w_034_3270, w_034_3272, w_034_3274, w_034_3275, w_034_3276, w_034_3277, w_034_3278, w_034_3279, w_034_3280, w_034_3281, w_034_3282, w_034_3283, w_034_3284, w_034_3285, w_034_3286, w_034_3288, w_034_3289, w_034_3292, w_034_3293, w_034_3294, w_034_3295, w_034_3296, w_034_3297, w_034_3298, w_034_3300, w_034_3301, w_034_3302, w_034_3303, w_034_3304, w_034_3305, w_034_3308, w_034_3309, w_034_3312, w_034_3314, w_034_3315, w_034_3316, w_034_3317, w_034_3318, w_034_3319, w_034_3320, w_034_3321, w_034_3323, w_034_3324, w_034_3325, w_034_3326, w_034_3327, w_034_3329, w_034_3331, w_034_3333, w_034_3335, w_034_3336, w_034_3337, w_034_3338, w_034_3339, w_034_3340, w_034_3341, w_034_3342, w_034_3343, w_034_3344, w_034_3345, w_034_3346, w_034_3347, w_034_3348, w_034_3349, w_034_3351, w_034_3352, w_034_3353, w_034_3354, w_034_3356, w_034_3357, w_034_3358, w_034_3359, w_034_3360, w_034_3361, w_034_3362, w_034_3363, w_034_3364, w_034_3365, w_034_3366, w_034_3367, w_034_3368, w_034_3370, w_034_3371, w_034_3372, w_034_3374, w_034_3375, w_034_3376, w_034_3381, w_034_3382, w_034_3384, w_034_3386, w_034_3387, w_034_3388, w_034_3389, w_034_3390, w_034_3392, w_034_3394, w_034_3395, w_034_3396, w_034_3399, w_034_3401, w_034_3402, w_034_3403, w_034_3404, w_034_3406, w_034_3407, w_034_3410, w_034_3411, w_034_3413, w_034_3414, w_034_3422, w_034_3423, w_034_3424, w_034_3425, w_034_3426, w_034_3427, w_034_3429, w_034_3432, w_034_3433, w_034_3436, w_034_3437, w_034_3438, w_034_3439, w_034_3440, w_034_3441, w_034_3442, w_034_3443, w_034_3444, w_034_3445, w_034_3446, w_034_3447, w_034_3448, w_034_3449, w_034_3450, w_034_3452, w_034_3454, w_034_3455, w_034_3457, w_034_3458, w_034_3459, w_034_3460, w_034_3461, w_034_3462, w_034_3463, w_034_3464, w_034_3465, w_034_3466, w_034_3469, w_034_3471, w_034_3472, w_034_3473, w_034_3474, w_034_3475, w_034_3476, w_034_3477, w_034_3478, w_034_3479, w_034_3480, w_034_3481, w_034_3482, w_034_3483, w_034_3484, w_034_3485, w_034_3486, w_034_3487, w_034_3488, w_034_3490, w_034_3493, w_034_3494, w_034_3497, w_034_3498, w_034_3499, w_034_3500, w_034_3501, w_034_3502, w_034_3503, w_034_3505, w_034_3506, w_034_3508, w_034_3510, w_034_3511, w_034_3512, w_034_3513, w_034_3514, w_034_3515, w_034_3517, w_034_3518, w_034_3519, w_034_3520, w_034_3521, w_034_3522, w_034_3523, w_034_3524, w_034_3525, w_034_3526, w_034_3527, w_034_3528, w_034_3534, w_034_3535, w_034_3536, w_034_3539, w_034_3541, w_034_3542, w_034_3543, w_034_3547, w_034_3548, w_034_3549, w_034_3552, w_034_3553, w_034_3554, w_034_3555, w_034_3556, w_034_3557, w_034_3559, w_034_3560, w_034_3563, w_034_3567, w_034_3569, w_034_3570, w_034_3571, w_034_3572, w_034_3573, w_034_3576, w_034_3577, w_034_3578, w_034_3579, w_034_3582, w_034_3583, w_034_3584, w_034_3586, w_034_3587, w_034_3588, w_034_3589, w_034_3590, w_034_3591, w_034_3592, w_034_3594, w_034_3595, w_034_3596, w_034_3598, w_034_3599, w_034_3600, w_034_3601, w_034_3602, w_034_3603, w_034_3604, w_034_3605, w_034_3607, w_034_3608, w_034_3609, w_034_3610, w_034_3612, w_034_3613, w_034_3615, w_034_3617, w_034_3618, w_034_3619, w_034_3620, w_034_3621, w_034_3622, w_034_3623, w_034_3624, w_034_3625, w_034_3626, w_034_3629, w_034_3630, w_034_3631, w_034_3632, w_034_3633, w_034_3634, w_034_3635, w_034_3636, w_034_3637, w_034_3638, w_034_3639, w_034_3640, w_034_3641, w_034_3642, w_034_3643, w_034_3644, w_034_3645, w_034_3646, w_034_3647, w_034_3648, w_034_3649, w_034_3651, w_034_3652, w_034_3654, w_034_3655, w_034_3658, w_034_3659, w_034_3660, w_034_3661, w_034_3663, w_034_3664, w_034_3665, w_034_3666, w_034_3668, w_034_3669, w_034_3670, w_034_3671, w_034_3672, w_034_3673, w_034_3674, w_034_3675, w_034_3676, w_034_3677, w_034_3678, w_034_3679, w_034_3680, w_034_3682, w_034_3683, w_034_3684, w_034_3685, w_034_3686, w_034_3691, w_034_3692, w_034_3693, w_034_3694, w_034_3695, w_034_3697, w_034_3698, w_034_3699, w_034_3700, w_034_3701, w_034_3702, w_034_3703, w_034_3704, w_034_3707, w_034_3708, w_034_3710, w_034_3711, w_034_3712, w_034_3714, w_034_3716, w_034_3718, w_034_3720, w_034_3721, w_034_3722, w_034_3723, w_034_3724, w_034_3727, w_034_3728, w_034_3729, w_034_3730, w_034_3731, w_034_3733, w_034_3735, w_034_3736, w_034_3737, w_034_3739, w_034_3740, w_034_3742, w_034_3743, w_034_3744, w_034_3746, w_034_3747, w_034_3748, w_034_3749, w_034_3750, w_034_3752, w_034_3753, w_034_3754, w_034_3756, w_034_3758, w_034_3759, w_034_3760, w_034_3761, w_034_3762, w_034_3763, w_034_3764, w_034_3768, w_034_3769, w_034_3770, w_034_3773, w_034_3774, w_034_3775, w_034_3776, w_034_3777, w_034_3778, w_034_3780, w_034_3781, w_034_3782, w_034_3783, w_034_3784, w_034_3785, w_034_3787, w_034_3788, w_034_3789, w_034_3791, w_034_3792, w_034_3793, w_034_3794, w_034_3796, w_034_3797, w_034_3798, w_034_3799, w_034_3800, w_034_3801, w_034_3804, w_034_3806, w_034_3807, w_034_3808, w_034_3809, w_034_3811, w_034_3813, w_034_3814, w_034_3815, w_034_3817, w_034_3818, w_034_3821, w_034_3822, w_034_3823, w_034_3824, w_034_3825, w_034_3826, w_034_3828, w_034_3829, w_034_3830, w_034_3831, w_034_3832, w_034_3833, w_034_3835, w_034_3837, w_034_3838, w_034_3839, w_034_3841, w_034_3843, w_034_3844, w_034_3845, w_034_3846, w_034_3847, w_034_3848, w_034_3849, w_034_3850, w_034_3851, w_034_3852, w_034_3853, w_034_3854, w_034_3855, w_034_3856, w_034_3857, w_034_3858, w_034_3859, w_034_3862, w_034_3864, w_034_3866, w_034_3867, w_034_3868, w_034_3869, w_034_3870, w_034_3871, w_034_3872, w_034_3873, w_034_3875, w_034_3876, w_034_3877, w_034_3878, w_034_3879, w_034_3880, w_034_3881, w_034_3882, w_034_3883, w_034_3884, w_034_3885, w_034_3886, w_034_3887, w_034_3888, w_034_3889, w_034_3890, w_034_3891, w_034_3892, w_034_3895, w_034_3896, w_034_3897, w_034_3899, w_034_3900, w_034_3901, w_034_3902, w_034_3903, w_034_3904, w_034_3905, w_034_3907, w_034_3910, w_034_3911, w_034_3912, w_034_3913, w_034_3916, w_034_3919, w_034_3923, w_034_3924, w_034_3925, w_034_3926, w_034_3927, w_034_3929, w_034_3930, w_034_3931, w_034_3932, w_034_3934, w_034_3936, w_034_3937, w_034_3938, w_034_3939, w_034_3941, w_034_3942, w_034_3943, w_034_3945, w_034_3947, w_034_3949, w_034_3950, w_034_3952, w_034_3953, w_034_3954, w_034_3955, w_034_3956, w_034_3957, w_034_3958, w_034_3959, w_034_3960, w_034_3961, w_034_3962, w_034_3964, w_034_3967, w_034_3968, w_034_3969, w_034_3970, w_034_3971, w_034_3973, w_034_3975, w_034_3976, w_034_3978, w_034_3981, w_034_3983, w_034_3984, w_034_3985, w_034_3986, w_034_3988, w_034_3989, w_034_3990, w_034_3993, w_034_3994, w_034_3996, w_034_3997, w_034_4000, w_034_4003, w_034_4004, w_034_4005, w_034_4006, w_034_4007, w_034_4008, w_034_4009, w_034_4010, w_034_4011, w_034_4012, w_034_4013, w_034_4014, w_034_4015, w_034_4016, w_034_4017, w_034_4018, w_034_4019, w_034_4020, w_034_4021, w_034_4022, w_034_4023, w_034_4025, w_034_4027, w_034_4028, w_034_4029, w_034_4031, w_034_4032, w_034_4033, w_034_4034, w_034_4035, w_034_4036, w_034_4037, w_034_4038, w_034_4039, w_034_4040, w_034_4041, w_034_4042, w_034_4043, w_034_4044, w_034_4045, w_034_4046, w_034_4048, w_034_4049, w_034_4050, w_034_4051, w_034_4052, w_034_4053, w_034_4054, w_034_4055, w_034_4056, w_034_4057, w_034_4058, w_034_4059, w_034_4061, w_034_4062, w_034_4064, w_034_4065, w_034_4066, w_034_4067, w_034_4069, w_034_4071, w_034_4072, w_034_4073, w_034_4076, w_034_4078, w_034_4079, w_034_4080, w_034_4081, w_034_4083, w_034_4084, w_034_4085, w_034_4086, w_034_4087, w_034_4088, w_034_4089, w_034_4090, w_034_4091, w_034_4095, w_034_4097, w_034_4098, w_034_4099, w_034_4101, w_034_4103, w_034_4105, w_034_4106, w_034_4108, w_034_4109, w_034_4110, w_034_4111, w_034_4112, w_034_4113, w_034_4114, w_034_4115, w_034_4116, w_034_4118, w_034_4119, w_034_4120, w_034_4122, w_034_4123, w_034_4125, w_034_4126, w_034_4128, w_034_4129, w_034_4131, w_034_4132, w_034_4133, w_034_4135, w_034_4136, w_034_4137, w_034_4138, w_034_4139, w_034_4140, w_034_4143, w_034_4146, w_034_4148, w_034_4149, w_034_4150, w_034_4151, w_034_4152, w_034_4153, w_034_4154, w_034_4155, w_034_4156, w_034_4157, w_034_4158, w_034_4159, w_034_4160, w_034_4162, w_034_4163, w_034_4164, w_034_4165, w_034_4166, w_034_4167, w_034_4169, w_034_4170, w_034_4171, w_034_4173, w_034_4174, w_034_4175, w_034_4176, w_034_4177, w_034_4179, w_034_4180, w_034_4182, w_034_4183, w_034_4184, w_034_4186, w_034_4187, w_034_4188, w_034_4190, w_034_4191, w_034_4193, w_034_4194, w_034_4195, w_034_4196, w_034_4198, w_034_4199, w_034_4202, w_034_4204, w_034_4205, w_034_4206, w_034_4207, w_034_4208, w_034_4209, w_034_4211, w_034_4213, w_034_4214, w_034_4215, w_034_4216, w_034_4217, w_034_4218, w_034_4219, w_034_4220, w_034_4221, w_034_4223, w_034_4225, w_034_4226, w_034_4227, w_034_4228, w_034_4230, w_034_4231, w_034_4232, w_034_4233, w_034_4234, w_034_4235, w_034_4237, w_034_4238, w_034_4239, w_034_4241, w_034_4242, w_034_4243, w_034_4244, w_034_4245, w_034_4250, w_034_4251, w_034_4252, w_034_4253, w_034_4255, w_034_4256, w_034_4258, w_034_4259, w_034_4260, w_034_4261, w_034_4262, w_034_4265, w_034_4267, w_034_4269, w_034_4270, w_034_4271, w_034_4273, w_034_4274, w_034_4275, w_034_4276, w_034_4277, w_034_4280, w_034_4281, w_034_4282, w_034_4283, w_034_4285, w_034_4286, w_034_4287, w_034_4288, w_034_4289, w_034_4290, w_034_4291, w_034_4292, w_034_4293, w_034_4294, w_034_4295, w_034_4297, w_034_4298, w_034_4299, w_034_4300, w_034_4303, w_034_4304, w_034_4305, w_034_4306, w_034_4307, w_034_4308, w_034_4309, w_034_4310, w_034_4311, w_034_4315, w_034_4316, w_034_4317, w_034_4318, w_034_4320, w_034_4321, w_034_4323, w_034_4324, w_034_4326, w_034_4327, w_034_4328, w_034_4330, w_034_4331, w_034_4333, w_034_4334, w_034_4338, w_034_4339, w_034_4340, w_034_4341, w_034_4342, w_034_4343, w_034_4346, w_034_4347, w_034_4349, w_034_4351, w_034_4353, w_034_4354, w_034_4355, w_034_4356, w_034_4357, w_034_4358, w_034_4359, w_034_4360, w_034_4361, w_034_4362, w_034_4363, w_034_4364, w_034_4365, w_034_4366, w_034_4368, w_034_4369, w_034_4370, w_034_4371, w_034_4372, w_034_4374, w_034_4376, w_034_4377, w_034_4378, w_034_4379, w_034_4380, w_034_4382, w_034_4385, w_034_4386, w_034_4388, w_034_4389, w_034_4390, w_034_4391, w_034_4392, w_034_4393, w_034_4394, w_034_4396, w_034_4397, w_034_4398, w_034_4400, w_034_4401, w_034_4402, w_034_4404, w_034_4405, w_034_4406, w_034_4407, w_034_4408, w_034_4410, w_034_4412, w_034_4413, w_034_4414, w_034_4416, w_034_4418, w_034_4420, w_034_4422, w_034_4423, w_034_4424, w_034_4427, w_034_4428, w_034_4429, w_034_4430, w_034_4431, w_034_4432, w_034_4433, w_034_4434, w_034_4435, w_034_4437, w_034_4439, w_034_4440, w_034_4441, w_034_4442, w_034_4444, w_034_4445, w_034_4446, w_034_4447, w_034_4450, w_034_4451, w_034_4452, w_034_4453, w_034_4454, w_034_4455, w_034_4456, w_034_4457, w_034_4458, w_034_4459, w_034_4460, w_034_4461, w_034_4463, w_034_4464, w_034_4465, w_034_4468, w_034_4469, w_034_4470, w_034_4472, w_034_4474, w_034_4475, w_034_4476, w_034_4477, w_034_4479, w_034_4480, w_034_4482, w_034_4483, w_034_4484, w_034_4485, w_034_4486, w_034_4487, w_034_4488, w_034_4489, w_034_4490, w_034_4491, w_034_4492, w_034_4493, w_034_4494, w_034_4495, w_034_4496, w_034_4497, w_034_4498, w_034_4500, w_034_4501, w_034_4503, w_034_4506, w_034_4508, w_034_4509, w_034_4510, w_034_4511, w_034_4512, w_034_4513, w_034_4514, w_034_4515, w_034_4516, w_034_4517, w_034_4520, w_034_4521, w_034_4522, w_034_4523, w_034_4524, w_034_4525, w_034_4526, w_034_4527, w_034_4528, w_034_4529, w_034_4530, w_034_4531, w_034_4532, w_034_4533, w_034_4534, w_034_4535, w_034_4536, w_034_4537, w_034_4539, w_034_4540, w_034_4544, w_034_4545, w_034_4546, w_034_4548, w_034_4549, w_034_4550, w_034_4552, w_034_4553, w_034_4554, w_034_4557, w_034_4558, w_034_4559, w_034_4561, w_034_4563, w_034_4564, w_034_4565, w_034_4566, w_034_4568, w_034_4569, w_034_4571, w_034_4572, w_034_4573, w_034_4574, w_034_4575, w_034_4576, w_034_4577, w_034_4579, w_034_4580, w_034_4582, w_034_4585, w_034_4586, w_034_4587, w_034_4589, w_034_4590, w_034_4591, w_034_4592, w_034_4593, w_034_4594, w_034_4595, w_034_4596, w_034_4600, w_034_4601, w_034_4602, w_034_4603, w_034_4604, w_034_4605, w_034_4606, w_034_4607, w_034_4608, w_034_4609, w_034_4610, w_034_4612, w_034_4613, w_034_4614, w_034_4617, w_034_4618, w_034_4619, w_034_4620, w_034_4621, w_034_4623, w_034_4624, w_034_4626, w_034_4630, w_034_4632, w_034_4634, w_034_4636, w_034_4640, w_034_4641, w_034_4642, w_034_4644, w_034_4647, w_034_4653, w_034_4654, w_034_4657, w_034_4658, w_034_4659, w_034_4662, w_034_4663, w_034_4667, w_034_4671, w_034_4672, w_034_4673, w_034_4674, w_034_4675, w_034_4677, w_034_4679, w_034_4681, w_034_4683, w_034_4686, w_034_4687, w_034_4688, w_034_4693, w_034_4695, w_034_4696, w_034_4697, w_034_4702, w_034_4706, w_034_4708, w_034_4710, w_034_4713, w_034_4714, w_034_4717, w_034_4718, w_034_4719, w_034_4720, w_034_4722, w_034_4725, w_034_4727, w_034_4728, w_034_4729, w_034_4730, w_034_4731, w_034_4733, w_034_4734, w_034_4735, w_034_4738, w_034_4739, w_034_4740, w_034_4742, w_034_4743, w_034_4747, w_034_4748, w_034_4749, w_034_4751, w_034_4752, w_034_4754, w_034_4759, w_034_4760, w_034_4761, w_034_4762, w_034_4764, w_034_4765, w_034_4767, w_034_4774, w_034_4775, w_034_4779, w_034_4780, w_034_4781, w_034_4783, w_034_4784, w_034_4788, w_034_4793, w_034_4794, w_034_4795, w_034_4797, w_034_4798, w_034_4799, w_034_4800, w_034_4801, w_034_4802, w_034_4803, w_034_4805, w_034_4806, w_034_4807, w_034_4808, w_034_4809, w_034_4810, w_034_4811, w_034_4812, w_034_4813, w_034_4815, w_034_4816, w_034_4820, w_034_4823, w_034_4824, w_034_4826, w_034_4827, w_034_4829, w_034_4830, w_034_4832, w_034_4833, w_034_4834, w_034_4836, w_034_4838, w_034_4842, w_034_4843, w_034_4846, w_034_4847, w_034_4848, w_034_4851, w_034_4853, w_034_4854, w_034_4856, w_034_4857, w_034_4861, w_034_4862, w_034_4863, w_034_4866, w_034_4867, w_034_4868, w_034_4869, w_034_4872, w_034_4879, w_034_4884, w_034_4885, w_034_4888, w_034_4889, w_034_4890, w_034_4891, w_034_4892, w_034_4893, w_034_4895, w_034_4896, w_034_4897, w_034_4898, w_034_4900, w_034_4901, w_034_4903, w_034_4904, w_034_4905, w_034_4906, w_034_4908, w_034_4910, w_034_4912, w_034_4913, w_034_4915, w_034_4920, w_034_4923, w_034_4924, w_034_4925, w_034_4929, w_034_4932, w_034_4934, w_034_4935, w_034_4936, w_034_4939, w_034_4940, w_034_4941, w_034_4942, w_034_4944, w_034_4945, w_034_4946, w_034_4953, w_034_4955, w_034_4960, w_034_4964, w_034_4965, w_034_4967, w_034_4968, w_034_4973, w_034_4974, w_034_4975, w_034_4977, w_034_4980, w_034_4981, w_034_4983, w_034_4984, w_034_4985, w_034_4986, w_034_4989, w_034_4991, w_034_4992, w_034_4994, w_034_4995, w_034_4998, w_034_4999, w_034_5002, w_034_5005, w_034_5006, w_034_5007, w_034_5008, w_034_5009, w_034_5010, w_034_5014, w_034_5015, w_034_5018, w_034_5021, w_034_5025, w_034_5027, w_034_5029, w_034_5030, w_034_5031, w_034_5035, w_034_5036, w_034_5038, w_034_5039, w_034_5040, w_034_5041, w_034_5043, w_034_5046, w_034_5049, w_034_5051, w_034_5053, w_034_5054, w_034_5056, w_034_5059, w_034_5062, w_034_5064, w_034_5067, w_034_5068, w_034_5069, w_034_5071, w_034_5078, w_034_5079, w_034_5081, w_034_5082, w_034_5084, w_034_5085, w_034_5086, w_034_5089, w_034_5090, w_034_5094, w_034_5095, w_034_5096, w_034_5097, w_034_5098, w_034_5099, w_034_5101, w_034_5102, w_034_5105, w_034_5106, w_034_5109, w_034_5110, w_034_5112, w_034_5114, w_034_5115, w_034_5121, w_034_5123, w_034_5125, w_034_5126, w_034_5128, w_034_5130, w_034_5131, w_034_5132, w_034_5133, w_034_5135, w_034_5136, w_034_5139, w_034_5140, w_034_5144, w_034_5145, w_034_5147, w_034_5148, w_034_5149, w_034_5150, w_034_5152, w_034_5153, w_034_5154, w_034_5155, w_034_5158, w_034_5160, w_034_5162, w_034_5163, w_034_5168, w_034_5169, w_034_5170, w_034_5175, w_034_5176, w_034_5178, w_034_5182, w_034_5183, w_034_5185, w_034_5186, w_034_5187, w_034_5188, w_034_5190, w_034_5191, w_034_5192, w_034_5193, w_034_5203, w_034_5204, w_034_5206, w_034_5207, w_034_5208, w_034_5209, w_034_5211, w_034_5213, w_034_5214, w_034_5215, w_034_5217, w_034_5219, w_034_5223, w_034_5224, w_034_5226, w_034_5227, w_034_5228, w_034_5229, w_034_5230, w_034_5231, w_034_5232, w_034_5233, w_034_5237, w_034_5241, w_034_5242, w_034_5245, w_034_5247, w_034_5249, w_034_5250, w_034_5252, w_034_5253, w_034_5255, w_034_5261, w_034_5266, w_034_5267, w_034_5272, w_034_5274, w_034_5276, w_034_5277, w_034_5282, w_034_5283, w_034_5288, w_034_5289, w_034_5290, w_034_5291, w_034_5292, w_034_5293, w_034_5296, w_034_5301, w_034_5302, w_034_5308, w_034_5311, w_034_5312, w_034_5317, w_034_5318, w_034_5319, w_034_5321, w_034_5325, w_034_5327, w_034_5328, w_034_5332, w_034_5334, w_034_5335, w_034_5336, w_034_5337, w_034_5343, w_034_5345, w_034_5346, w_034_5347, w_034_5349, w_034_5350, w_034_5351, w_034_5353, w_034_5356, w_034_5359, w_034_5361, w_034_5365, w_034_5368, w_034_5369, w_034_5370, w_034_5371, w_034_5373, w_034_5374, w_034_5376, w_034_5377;
  wire w_035_001, w_035_004, w_035_006, w_035_009, w_035_010, w_035_011, w_035_012, w_035_013, w_035_014, w_035_016, w_035_017, w_035_018, w_035_020, w_035_021, w_035_022, w_035_024, w_035_025, w_035_026, w_035_027, w_035_029, w_035_030, w_035_031, w_035_032, w_035_033, w_035_034, w_035_035, w_035_036, w_035_037, w_035_038, w_035_039, w_035_040, w_035_042, w_035_044, w_035_045, w_035_046, w_035_048, w_035_051, w_035_052, w_035_053, w_035_054, w_035_055, w_035_060, w_035_062, w_035_063, w_035_064, w_035_065, w_035_066, w_035_067, w_035_068, w_035_071, w_035_072, w_035_074, w_035_076, w_035_077, w_035_078, w_035_079, w_035_080, w_035_081, w_035_084, w_035_085, w_035_086, w_035_087, w_035_089, w_035_090, w_035_091, w_035_092, w_035_093, w_035_094, w_035_096, w_035_098, w_035_099, w_035_100, w_035_101, w_035_102, w_035_103, w_035_105, w_035_107, w_035_108, w_035_109, w_035_110, w_035_112, w_035_114, w_035_115, w_035_116, w_035_117, w_035_118, w_035_119, w_035_120, w_035_121, w_035_122, w_035_123, w_035_126, w_035_127, w_035_128, w_035_129, w_035_130, w_035_131, w_035_132, w_035_133, w_035_134, w_035_135, w_035_136, w_035_138, w_035_139, w_035_141, w_035_145, w_035_146, w_035_148, w_035_150, w_035_151, w_035_153, w_035_154, w_035_155, w_035_156, w_035_158, w_035_159, w_035_160, w_035_161, w_035_162, w_035_163, w_035_166, w_035_167, w_035_168, w_035_169, w_035_170, w_035_171, w_035_173, w_035_175, w_035_176, w_035_180, w_035_181, w_035_182, w_035_184, w_035_185, w_035_186, w_035_187, w_035_188, w_035_189, w_035_190, w_035_191, w_035_192, w_035_193, w_035_194, w_035_197, w_035_199, w_035_200, w_035_202, w_035_203, w_035_204, w_035_205, w_035_206, w_035_207, w_035_208, w_035_209, w_035_210, w_035_211, w_035_212, w_035_213, w_035_215, w_035_216, w_035_217, w_035_218, w_035_219, w_035_223, w_035_224, w_035_225, w_035_227, w_035_229, w_035_230, w_035_231, w_035_232, w_035_235, w_035_238, w_035_240, w_035_241, w_035_242, w_035_243, w_035_245, w_035_246, w_035_247, w_035_248, w_035_249, w_035_250, w_035_254, w_035_256, w_035_258, w_035_259, w_035_260, w_035_262, w_035_264, w_035_265, w_035_267, w_035_269, w_035_271, w_035_272, w_035_273, w_035_275, w_035_276, w_035_277, w_035_279, w_035_280, w_035_281, w_035_283, w_035_284, w_035_288, w_035_290, w_035_291, w_035_292, w_035_293, w_035_294, w_035_295, w_035_296, w_035_297, w_035_301, w_035_302, w_035_303, w_035_305, w_035_306, w_035_307, w_035_309, w_035_310, w_035_312, w_035_313, w_035_314, w_035_315, w_035_316, w_035_317, w_035_318, w_035_319, w_035_320, w_035_321, w_035_323, w_035_324, w_035_326, w_035_327, w_035_328, w_035_331, w_035_332, w_035_333, w_035_334, w_035_335, w_035_337, w_035_338, w_035_343, w_035_344, w_035_345, w_035_346, w_035_347, w_035_350, w_035_351, w_035_354, w_035_356, w_035_357, w_035_358, w_035_360, w_035_362, w_035_363, w_035_364, w_035_365, w_035_366, w_035_367, w_035_369, w_035_370, w_035_371, w_035_372, w_035_373, w_035_375, w_035_378, w_035_379, w_035_380, w_035_382, w_035_383, w_035_384, w_035_385, w_035_386, w_035_387, w_035_388, w_035_390, w_035_392, w_035_393, w_035_394, w_035_395, w_035_396, w_035_397, w_035_398, w_035_399, w_035_400, w_035_401, w_035_403, w_035_405, w_035_406, w_035_407, w_035_410, w_035_411, w_035_416, w_035_418, w_035_421, w_035_422, w_035_424, w_035_425, w_035_426, w_035_427, w_035_428, w_035_429, w_035_430, w_035_431, w_035_434, w_035_437, w_035_438, w_035_439, w_035_440, w_035_441, w_035_442, w_035_443, w_035_444, w_035_445, w_035_446, w_035_447, w_035_449, w_035_450, w_035_452, w_035_453, w_035_454, w_035_455, w_035_456, w_035_457, w_035_458, w_035_459, w_035_460, w_035_461, w_035_462, w_035_463, w_035_466, w_035_467, w_035_468, w_035_471, w_035_472, w_035_473, w_035_474, w_035_475, w_035_476, w_035_477, w_035_479, w_035_481, w_035_485, w_035_486, w_035_487, w_035_489, w_035_490, w_035_491, w_035_492, w_035_493, w_035_496, w_035_497, w_035_499, w_035_501, w_035_502, w_035_503, w_035_504, w_035_505, w_035_506, w_035_508, w_035_509, w_035_510, w_035_512, w_035_514, w_035_515, w_035_516, w_035_517, w_035_518, w_035_519, w_035_520, w_035_522, w_035_523, w_035_524, w_035_525, w_035_526, w_035_527, w_035_528, w_035_529, w_035_530, w_035_531, w_035_533, w_035_534, w_035_536, w_035_537, w_035_538, w_035_539, w_035_540, w_035_541, w_035_542, w_035_543, w_035_545, w_035_546, w_035_547, w_035_549, w_035_551, w_035_552, w_035_553, w_035_555, w_035_556, w_035_557, w_035_558, w_035_559, w_035_561, w_035_562, w_035_563, w_035_564, w_035_568, w_035_569, w_035_570, w_035_571, w_035_572, w_035_573, w_035_574, w_035_575, w_035_576, w_035_577, w_035_580, w_035_582, w_035_583, w_035_585, w_035_586, w_035_587, w_035_588, w_035_589, w_035_591, w_035_592, w_035_593, w_035_594, w_035_596, w_035_597, w_035_598, w_035_601, w_035_602, w_035_604, w_035_605, w_035_606, w_035_607, w_035_608, w_035_609, w_035_611, w_035_612, w_035_613, w_035_614, w_035_615, w_035_616, w_035_617, w_035_618, w_035_619, w_035_620, w_035_621, w_035_622, w_035_623, w_035_624, w_035_625, w_035_626, w_035_627, w_035_629, w_035_630, w_035_632, w_035_633, w_035_634, w_035_637, w_035_639, w_035_640, w_035_644, w_035_645, w_035_647, w_035_648, w_035_652, w_035_653, w_035_654, w_035_656, w_035_658, w_035_659, w_035_660, w_035_661, w_035_662, w_035_663, w_035_664, w_035_665, w_035_666, w_035_668, w_035_671, w_035_672, w_035_673, w_035_674, w_035_675, w_035_676, w_035_677, w_035_679, w_035_680, w_035_681, w_035_682, w_035_683, w_035_684, w_035_685, w_035_686, w_035_689, w_035_690, w_035_692, w_035_693, w_035_694, w_035_695, w_035_696, w_035_698, w_035_699, w_035_700, w_035_701, w_035_704, w_035_705, w_035_707, w_035_709, w_035_710, w_035_711, w_035_712, w_035_713, w_035_714, w_035_715, w_035_717, w_035_718, w_035_719, w_035_720, w_035_721, w_035_723, w_035_724, w_035_725, w_035_728, w_035_729, w_035_731, w_035_733, w_035_734, w_035_735, w_035_738, w_035_739, w_035_740, w_035_744, w_035_746, w_035_747, w_035_748, w_035_749, w_035_750, w_035_751, w_035_752, w_035_753, w_035_755, w_035_756, w_035_758, w_035_759, w_035_760, w_035_761, w_035_762, w_035_763, w_035_764, w_035_765, w_035_766, w_035_767, w_035_768, w_035_769, w_035_772, w_035_774, w_035_775, w_035_776, w_035_779, w_035_780, w_035_784, w_035_785, w_035_786, w_035_788, w_035_791, w_035_792, w_035_794, w_035_797, w_035_798, w_035_800, w_035_801, w_035_802, w_035_805, w_035_806, w_035_807, w_035_809, w_035_813, w_035_814, w_035_815, w_035_816, w_035_817, w_035_818, w_035_819, w_035_821, w_035_822, w_035_824, w_035_825, w_035_826, w_035_830, w_035_831, w_035_833, w_035_834, w_035_835, w_035_837, w_035_838, w_035_840, w_035_841, w_035_842, w_035_843, w_035_844, w_035_845, w_035_847, w_035_849, w_035_850, w_035_851, w_035_852, w_035_854, w_035_855, w_035_856, w_035_857, w_035_858, w_035_860, w_035_862, w_035_865, w_035_867, w_035_868, w_035_869, w_035_871, w_035_872, w_035_873, w_035_875, w_035_876, w_035_877, w_035_878, w_035_879, w_035_880, w_035_882, w_035_883, w_035_884, w_035_885, w_035_886, w_035_888, w_035_889, w_035_890, w_035_891, w_035_892, w_035_893, w_035_895, w_035_897, w_035_898, w_035_900, w_035_903, w_035_904, w_035_905, w_035_906, w_035_907, w_035_908, w_035_909, w_035_910, w_035_911, w_035_912, w_035_913, w_035_914, w_035_916, w_035_918, w_035_919, w_035_920, w_035_921, w_035_923, w_035_924, w_035_925, w_035_927, w_035_928, w_035_929, w_035_930, w_035_931, w_035_932, w_035_934, w_035_935, w_035_936, w_035_938, w_035_939, w_035_940, w_035_941, w_035_942, w_035_943, w_035_946, w_035_947, w_035_949, w_035_950, w_035_952, w_035_953, w_035_956, w_035_958, w_035_960, w_035_961, w_035_962, w_035_966, w_035_967, w_035_968, w_035_970, w_035_971, w_035_972, w_035_973, w_035_974, w_035_975, w_035_976, w_035_978, w_035_980, w_035_982, w_035_984, w_035_985, w_035_987, w_035_988, w_035_989, w_035_990, w_035_991, w_035_992, w_035_993, w_035_994, w_035_995, w_035_997, w_035_998, w_035_999, w_035_1000, w_035_1003, w_035_1004, w_035_1005, w_035_1007, w_035_1008, w_035_1009, w_035_1010, w_035_1011, w_035_1012, w_035_1013, w_035_1014, w_035_1015, w_035_1016, w_035_1017, w_035_1018, w_035_1019, w_035_1020, w_035_1021, w_035_1023, w_035_1025, w_035_1026, w_035_1028, w_035_1029, w_035_1034, w_035_1036, w_035_1038, w_035_1039, w_035_1042, w_035_1045, w_035_1046, w_035_1047, w_035_1048, w_035_1049, w_035_1050, w_035_1051, w_035_1053, w_035_1055, w_035_1057, w_035_1058, w_035_1059, w_035_1062, w_035_1063, w_035_1066, w_035_1067, w_035_1068, w_035_1069, w_035_1070, w_035_1071, w_035_1072, w_035_1073, w_035_1075, w_035_1076, w_035_1078, w_035_1080, w_035_1082, w_035_1083, w_035_1084, w_035_1087, w_035_1088, w_035_1089, w_035_1090, w_035_1093, w_035_1094, w_035_1095, w_035_1096, w_035_1099, w_035_1100, w_035_1102, w_035_1104, w_035_1106, w_035_1107, w_035_1108, w_035_1110, w_035_1112, w_035_1114, w_035_1115, w_035_1116, w_035_1117, w_035_1118, w_035_1119, w_035_1120, w_035_1121, w_035_1122, w_035_1123, w_035_1126, w_035_1127, w_035_1128, w_035_1129, w_035_1130, w_035_1131, w_035_1132, w_035_1134, w_035_1135, w_035_1136, w_035_1137, w_035_1138, w_035_1141, w_035_1142, w_035_1144, w_035_1145, w_035_1146, w_035_1147, w_035_1149, w_035_1150, w_035_1151, w_035_1152, w_035_1153, w_035_1154, w_035_1155, w_035_1157, w_035_1158, w_035_1159, w_035_1160, w_035_1163, w_035_1165, w_035_1166, w_035_1168, w_035_1169, w_035_1170, w_035_1173, w_035_1174, w_035_1175, w_035_1176, w_035_1177, w_035_1179, w_035_1180, w_035_1183, w_035_1185, w_035_1188, w_035_1189, w_035_1190, w_035_1191, w_035_1192, w_035_1194, w_035_1196, w_035_1197, w_035_1199, w_035_1200, w_035_1201, w_035_1202, w_035_1203, w_035_1204, w_035_1205, w_035_1207, w_035_1208, w_035_1210, w_035_1212, w_035_1213, w_035_1214, w_035_1215, w_035_1217, w_035_1218, w_035_1219, w_035_1220, w_035_1221, w_035_1222, w_035_1223, w_035_1224, w_035_1225, w_035_1227, w_035_1228, w_035_1229, w_035_1230, w_035_1231, w_035_1232, w_035_1233, w_035_1234, w_035_1235, w_035_1236, w_035_1238, w_035_1240, w_035_1241, w_035_1242, w_035_1243, w_035_1244, w_035_1245, w_035_1247, w_035_1248, w_035_1249, w_035_1250, w_035_1251, w_035_1253, w_035_1254, w_035_1255, w_035_1256, w_035_1258, w_035_1259, w_035_1261, w_035_1262, w_035_1263, w_035_1265, w_035_1266, w_035_1267, w_035_1268, w_035_1269, w_035_1272, w_035_1273, w_035_1274, w_035_1275, w_035_1277, w_035_1278, w_035_1279, w_035_1280, w_035_1282, w_035_1283, w_035_1284, w_035_1285, w_035_1286, w_035_1287, w_035_1289, w_035_1290, w_035_1293, w_035_1294, w_035_1295, w_035_1296, w_035_1299, w_035_1300, w_035_1302, w_035_1303, w_035_1304, w_035_1305, w_035_1306, w_035_1307, w_035_1308, w_035_1309, w_035_1310, w_035_1311, w_035_1312, w_035_1313, w_035_1316, w_035_1317, w_035_1319, w_035_1320, w_035_1322, w_035_1323, w_035_1325, w_035_1326, w_035_1327, w_035_1328, w_035_1329, w_035_1330, w_035_1331, w_035_1332, w_035_1333, w_035_1334, w_035_1335, w_035_1336, w_035_1337, w_035_1340, w_035_1341, w_035_1342, w_035_1343, w_035_1344, w_035_1345, w_035_1346, w_035_1348, w_035_1349, w_035_1350, w_035_1352, w_035_1354, w_035_1357, w_035_1358, w_035_1359, w_035_1360, w_035_1361, w_035_1366, w_035_1367, w_035_1368, w_035_1370, w_035_1371, w_035_1372, w_035_1373, w_035_1374, w_035_1375, w_035_1376, w_035_1377, w_035_1378, w_035_1379, w_035_1380, w_035_1382, w_035_1383, w_035_1385, w_035_1386, w_035_1387, w_035_1390, w_035_1393, w_035_1394, w_035_1396, w_035_1397, w_035_1398, w_035_1400, w_035_1401, w_035_1402, w_035_1403, w_035_1404, w_035_1407, w_035_1408, w_035_1410, w_035_1411, w_035_1412, w_035_1413, w_035_1415, w_035_1417, w_035_1418, w_035_1419, w_035_1421, w_035_1423, w_035_1424, w_035_1426, w_035_1427, w_035_1428, w_035_1429, w_035_1430, w_035_1431, w_035_1432, w_035_1433, w_035_1434, w_035_1435, w_035_1436, w_035_1438, w_035_1439, w_035_1441, w_035_1443, w_035_1444, w_035_1445, w_035_1446, w_035_1447, w_035_1448, w_035_1449, w_035_1450, w_035_1451, w_035_1453, w_035_1454, w_035_1455, w_035_1457, w_035_1458, w_035_1460, w_035_1461, w_035_1462, w_035_1463, w_035_1464, w_035_1466, w_035_1467, w_035_1468, w_035_1469, w_035_1470, w_035_1471, w_035_1472, w_035_1474, w_035_1476, w_035_1477, w_035_1478, w_035_1479, w_035_1480, w_035_1481, w_035_1482, w_035_1483, w_035_1484, w_035_1485, w_035_1486, w_035_1487, w_035_1488, w_035_1489, w_035_1490, w_035_1491, w_035_1492, w_035_1494, w_035_1495, w_035_1496, w_035_1498, w_035_1499, w_035_1500, w_035_1501, w_035_1502, w_035_1505, w_035_1506, w_035_1507, w_035_1510, w_035_1511, w_035_1512, w_035_1513, w_035_1514, w_035_1515, w_035_1516, w_035_1517, w_035_1518, w_035_1519, w_035_1522, w_035_1524, w_035_1525, w_035_1526, w_035_1527, w_035_1528, w_035_1529, w_035_1531, w_035_1534, w_035_1535, w_035_1536, w_035_1537, w_035_1538, w_035_1539, w_035_1540, w_035_1541, w_035_1542, w_035_1543, w_035_1544, w_035_1545, w_035_1546, w_035_1547, w_035_1548, w_035_1550, w_035_1551, w_035_1552, w_035_1553, w_035_1555, w_035_1556, w_035_1557, w_035_1558, w_035_1559, w_035_1560, w_035_1561, w_035_1563, w_035_1564, w_035_1566, w_035_1567, w_035_1568, w_035_1569, w_035_1573, w_035_1575, w_035_1576, w_035_1577, w_035_1578, w_035_1579, w_035_1580, w_035_1581, w_035_1582, w_035_1584, w_035_1585, w_035_1586, w_035_1589, w_035_1590, w_035_1591, w_035_1592, w_035_1593, w_035_1594, w_035_1596, w_035_1598, w_035_1599, w_035_1600, w_035_1601, w_035_1602, w_035_1604, w_035_1605, w_035_1606, w_035_1608, w_035_1609, w_035_1611, w_035_1612, w_035_1613, w_035_1614, w_035_1616, w_035_1617, w_035_1618, w_035_1619, w_035_1620, w_035_1621, w_035_1622, w_035_1624, w_035_1625, w_035_1627, w_035_1628, w_035_1629, w_035_1630, w_035_1631, w_035_1633, w_035_1634, w_035_1635, w_035_1636, w_035_1637, w_035_1638, w_035_1639, w_035_1640, w_035_1641, w_035_1642, w_035_1643, w_035_1644, w_035_1646, w_035_1647, w_035_1649, w_035_1650, w_035_1652, w_035_1653, w_035_1654, w_035_1655, w_035_1656, w_035_1657, w_035_1658, w_035_1659, w_035_1661, w_035_1662, w_035_1663, w_035_1664, w_035_1665, w_035_1666, w_035_1667, w_035_1668, w_035_1670, w_035_1671, w_035_1672, w_035_1673, w_035_1674, w_035_1676, w_035_1678, w_035_1680, w_035_1681, w_035_1682, w_035_1684, w_035_1686, w_035_1687, w_035_1688, w_035_1690, w_035_1693, w_035_1694, w_035_1695, w_035_1696, w_035_1697, w_035_1698, w_035_1699, w_035_1700, w_035_1701, w_035_1702, w_035_1703, w_035_1704, w_035_1706, w_035_1707, w_035_1708, w_035_1709, w_035_1710, w_035_1711, w_035_1712, w_035_1713, w_035_1714, w_035_1716, w_035_1717, w_035_1718, w_035_1719, w_035_1720, w_035_1721, w_035_1722, w_035_1723, w_035_1725, w_035_1726, w_035_1727, w_035_1728, w_035_1729, w_035_1731, w_035_1732, w_035_1733, w_035_1735, w_035_1736, w_035_1737, w_035_1738, w_035_1739, w_035_1740, w_035_1741, w_035_1742, w_035_1743, w_035_1744, w_035_1745, w_035_1746, w_035_1747, w_035_1748, w_035_1750, w_035_1751, w_035_1752, w_035_1753, w_035_1754, w_035_1756, w_035_1757, w_035_1759, w_035_1760, w_035_1762, w_035_1763, w_035_1765, w_035_1766, w_035_1767, w_035_1768, w_035_1769, w_035_1770, w_035_1771, w_035_1773, w_035_1774, w_035_1775, w_035_1776, w_035_1778, w_035_1779, w_035_1780, w_035_1781, w_035_1782, w_035_1784, w_035_1785, w_035_1786, w_035_1787, w_035_1789, w_035_1790, w_035_1792, w_035_1793, w_035_1794, w_035_1799, w_035_1800, w_035_1801, w_035_1802, w_035_1803, w_035_1806, w_035_1807, w_035_1808, w_035_1809, w_035_1812, w_035_1815, w_035_1817, w_035_1820, w_035_1822, w_035_1823, w_035_1824, w_035_1825, w_035_1826, w_035_1827, w_035_1830, w_035_1831, w_035_1832, w_035_1834, w_035_1835, w_035_1837, w_035_1838, w_035_1839, w_035_1840, w_035_1841, w_035_1842, w_035_1843, w_035_1844, w_035_1845, w_035_1847, w_035_1848, w_035_1849, w_035_1851, w_035_1854, w_035_1855, w_035_1856, w_035_1857, w_035_1858, w_035_1860, w_035_1861, w_035_1862, w_035_1863, w_035_1864, w_035_1865, w_035_1867, w_035_1869, w_035_1871, w_035_1872, w_035_1874, w_035_1875, w_035_1878, w_035_1879, w_035_1881, w_035_1883, w_035_1884, w_035_1885, w_035_1886, w_035_1887, w_035_1889, w_035_1890, w_035_1891, w_035_1892, w_035_1893, w_035_1894, w_035_1895, w_035_1896, w_035_1899, w_035_1900, w_035_1901, w_035_1902, w_035_1903, w_035_1904, w_035_1905, w_035_1907, w_035_1909, w_035_1911, w_035_1913, w_035_1914, w_035_1915, w_035_1917, w_035_1921, w_035_1922, w_035_1923, w_035_1925, w_035_1926, w_035_1927, w_035_1928, w_035_1930, w_035_1931, w_035_1933, w_035_1934, w_035_1935, w_035_1936, w_035_1937, w_035_1938, w_035_1939, w_035_1940, w_035_1941, w_035_1942, w_035_1943, w_035_1945, w_035_1946, w_035_1947, w_035_1948, w_035_1949, w_035_1950, w_035_1951, w_035_1954, w_035_1955, w_035_1956, w_035_1957, w_035_1958, w_035_1959, w_035_1961, w_035_1963, w_035_1964, w_035_1965, w_035_1966, w_035_1967, w_035_1968, w_035_1969, w_035_1971, w_035_1972, w_035_1973, w_035_1974, w_035_1976, w_035_1977, w_035_1979, w_035_1980, w_035_1981, w_035_1983, w_035_1984, w_035_1985, w_035_1986, w_035_1987, w_035_1988, w_035_1989, w_035_1990, w_035_1991, w_035_1992, w_035_1993, w_035_1994, w_035_1995, w_035_1996, w_035_1997, w_035_1998, w_035_1999, w_035_2000, w_035_2002, w_035_2003, w_035_2004, w_035_2007, w_035_2008, w_035_2009, w_035_2011, w_035_2013, w_035_2014, w_035_2015, w_035_2016, w_035_2017, w_035_2018, w_035_2020, w_035_2021, w_035_2022, w_035_2023, w_035_2024, w_035_2025, w_035_2026, w_035_2027, w_035_2028, w_035_2029, w_035_2030, w_035_2031, w_035_2033, w_035_2035, w_035_2036, w_035_2037, w_035_2041, w_035_2042, w_035_2043, w_035_2044, w_035_2045, w_035_2048, w_035_2050, w_035_2051, w_035_2052, w_035_2053, w_035_2054, w_035_2055, w_035_2056, w_035_2057, w_035_2059, w_035_2060, w_035_2061, w_035_2063, w_035_2064, w_035_2065, w_035_2066, w_035_2067, w_035_2068, w_035_2069, w_035_2072, w_035_2073, w_035_2074, w_035_2075, w_035_2076, w_035_2077, w_035_2078, w_035_2080, w_035_2081, w_035_2083, w_035_2085, w_035_2087, w_035_2088, w_035_2089, w_035_2090, w_035_2091, w_035_2093, w_035_2095, w_035_2096, w_035_2098, w_035_2099, w_035_2102, w_035_2104, w_035_2106, w_035_2107, w_035_2108, w_035_2109, w_035_2110, w_035_2112, w_035_2114, w_035_2116, w_035_2117, w_035_2119, w_035_2120, w_035_2122, w_035_2123, w_035_2124, w_035_2125, w_035_2127, w_035_2128, w_035_2129, w_035_2132, w_035_2133, w_035_2136, w_035_2137, w_035_2138, w_035_2139, w_035_2141, w_035_2143, w_035_2144, w_035_2145, w_035_2146, w_035_2147, w_035_2149, w_035_2151, w_035_2152, w_035_2153, w_035_2156, w_035_2157, w_035_2158, w_035_2160, w_035_2161, w_035_2162, w_035_2163, w_035_2165, w_035_2166, w_035_2168, w_035_2171, w_035_2173, w_035_2174, w_035_2175, w_035_2176, w_035_2177, w_035_2179, w_035_2181, w_035_2182, w_035_2183, w_035_2186, w_035_2188, w_035_2189, w_035_2190, w_035_2191, w_035_2195, w_035_2199, w_035_2200, w_035_2202, w_035_2203, w_035_2205, w_035_2206, w_035_2207, w_035_2210, w_035_2211, w_035_2212, w_035_2213, w_035_2218, w_035_2219, w_035_2220, w_035_2222, w_035_2223, w_035_2224, w_035_2225, w_035_2226, w_035_2228, w_035_2230, w_035_2231, w_035_2232, w_035_2234, w_035_2235, w_035_2236, w_035_2240, w_035_2241, w_035_2242, w_035_2243, w_035_2244, w_035_2246, w_035_2247, w_035_2248, w_035_2249, w_035_2250, w_035_2252, w_035_2254, w_035_2255, w_035_2257, w_035_2258, w_035_2259, w_035_2260, w_035_2261, w_035_2262, w_035_2263, w_035_2264, w_035_2265, w_035_2268, w_035_2271, w_035_2273, w_035_2275, w_035_2276, w_035_2277, w_035_2278, w_035_2279, w_035_2280, w_035_2281, w_035_2284, w_035_2285, w_035_2287, w_035_2288, w_035_2289, w_035_2290, w_035_2291, w_035_2292, w_035_2293, w_035_2294, w_035_2295, w_035_2296, w_035_2297, w_035_2298, w_035_2299, w_035_2300, w_035_2303, w_035_2304, w_035_2305, w_035_2306, w_035_2308, w_035_2311, w_035_2313, w_035_2314, w_035_2316, w_035_2317, w_035_2318, w_035_2320, w_035_2321, w_035_2322, w_035_2323, w_035_2324, w_035_2325, w_035_2326, w_035_2329, w_035_2330, w_035_2332, w_035_2333, w_035_2334, w_035_2335, w_035_2337, w_035_2340, w_035_2341, w_035_2342, w_035_2343, w_035_2345, w_035_2347, w_035_2348, w_035_2349, w_035_2350, w_035_2351, w_035_2352, w_035_2353, w_035_2355, w_035_2357, w_035_2359, w_035_2360, w_035_2361, w_035_2362, w_035_2364, w_035_2365, w_035_2369, w_035_2370, w_035_2371, w_035_2373, w_035_2374, w_035_2376, w_035_2377, w_035_2378, w_035_2379, w_035_2380, w_035_2381, w_035_2382, w_035_2383, w_035_2384, w_035_2385, w_035_2386, w_035_2387, w_035_2388, w_035_2389, w_035_2390, w_035_2391, w_035_2392, w_035_2393, w_035_2394, w_035_2395, w_035_2396, w_035_2398, w_035_2399, w_035_2400, w_035_2401, w_035_2402, w_035_2403, w_035_2405, w_035_2406, w_035_2407, w_035_2408, w_035_2409, w_035_2410, w_035_2411, w_035_2412, w_035_2414, w_035_2416, w_035_2417, w_035_2419, w_035_2420, w_035_2422, w_035_2423, w_035_2424, w_035_2425, w_035_2426, w_035_2427, w_035_2428, w_035_2429, w_035_2430, w_035_2431, w_035_2432, w_035_2433, w_035_2434, w_035_2435, w_035_2436, w_035_2437, w_035_2438, w_035_2440, w_035_2441, w_035_2442, w_035_2443, w_035_2446, w_035_2447, w_035_2448, w_035_2452, w_035_2454, w_035_2456, w_035_2457, w_035_2458, w_035_2459, w_035_2462, w_035_2465, w_035_2468, w_035_2469, w_035_2470, w_035_2472, w_035_2473, w_035_2475, w_035_2476, w_035_2477, w_035_2478, w_035_2480, w_035_2481, w_035_2482, w_035_2483, w_035_2484, w_035_2486, w_035_2487, w_035_2488, w_035_2489, w_035_2490, w_035_2491, w_035_2494, w_035_2496, w_035_2497, w_035_2499, w_035_2500, w_035_2501, w_035_2504, w_035_2506, w_035_2509, w_035_2510, w_035_2511, w_035_2512, w_035_2515, w_035_2516, w_035_2517, w_035_2518, w_035_2519, w_035_2520, w_035_2522, w_035_2523, w_035_2524, w_035_2525, w_035_2526, w_035_2527, w_035_2528, w_035_2530, w_035_2531, w_035_2533, w_035_2534, w_035_2535, w_035_2536, w_035_2537, w_035_2538, w_035_2539, w_035_2540, w_035_2541, w_035_2542, w_035_2543, w_035_2544, w_035_2545, w_035_2546, w_035_2547, w_035_2548, w_035_2549, w_035_2550, w_035_2551, w_035_2552, w_035_2553, w_035_2555, w_035_2557, w_035_2558, w_035_2559, w_035_2560, w_035_2561, w_035_2562, w_035_2563, w_035_2564, w_035_2565, w_035_2566, w_035_2568, w_035_2569, w_035_2570, w_035_2572, w_035_2575, w_035_2577, w_035_2579, w_035_2582, w_035_2583, w_035_2584, w_035_2585, w_035_2586, w_035_2587, w_035_2588, w_035_2589, w_035_2591, w_035_2592, w_035_2593, w_035_2594, w_035_2596, w_035_2598, w_035_2599, w_035_2601, w_035_2602, w_035_2604, w_035_2605, w_035_2607, w_035_2608, w_035_2609, w_035_2610, w_035_2612, w_035_2613, w_035_2614, w_035_2616, w_035_2617, w_035_2618, w_035_2619, w_035_2620, w_035_2621, w_035_2623, w_035_2624, w_035_2625, w_035_2626, w_035_2628, w_035_2630, w_035_2631, w_035_2633, w_035_2634, w_035_2636, w_035_2638, w_035_2640, w_035_2641, w_035_2642, w_035_2644, w_035_2645, w_035_2646, w_035_2648, w_035_2649, w_035_2652, w_035_2653, w_035_2654, w_035_2655, w_035_2656, w_035_2658, w_035_2660, w_035_2661, w_035_2662, w_035_2663, w_035_2664, w_035_2665, w_035_2667, w_035_2668, w_035_2670, w_035_2671, w_035_2672, w_035_2673, w_035_2674, w_035_2675, w_035_2677, w_035_2678, w_035_2679, w_035_2680, w_035_2681, w_035_2682, w_035_2685, w_035_2686, w_035_2687, w_035_2688, w_035_2690, w_035_2691, w_035_2692, w_035_2694, w_035_2696, w_035_2697, w_035_2698, w_035_2699, w_035_2700, w_035_2701, w_035_2703, w_035_2704, w_035_2705, w_035_2706, w_035_2707, w_035_2709, w_035_2711, w_035_2712, w_035_2713, w_035_2714, w_035_2715, w_035_2716, w_035_2717, w_035_2718, w_035_2719, w_035_2720, w_035_2721, w_035_2722, w_035_2723, w_035_2724, w_035_2725, w_035_2726, w_035_2728, w_035_2729, w_035_2731, w_035_2732, w_035_2733, w_035_2734, w_035_2735, w_035_2736, w_035_2737, w_035_2738, w_035_2740, w_035_2741, w_035_2743, w_035_2744, w_035_2745, w_035_2746, w_035_2747, w_035_2748, w_035_2749, w_035_2750, w_035_2751, w_035_2752, w_035_2754, w_035_2755, w_035_2756, w_035_2757, w_035_2758, w_035_2759, w_035_2760, w_035_2761, w_035_2762, w_035_2766, w_035_2767, w_035_2768, w_035_2770, w_035_2771, w_035_2773, w_035_2774, w_035_2775, w_035_2777, w_035_2779, w_035_2780, w_035_2781, w_035_2782, w_035_2783, w_035_2784, w_035_2785, w_035_2786, w_035_2787, w_035_2788, w_035_2789, w_035_2791, w_035_2792, w_035_2794, w_035_2795, w_035_2796, w_035_2797, w_035_2798, w_035_2799, w_035_2800, w_035_2801, w_035_2802, w_035_2803, w_035_2804, w_035_2805, w_035_2806, w_035_2807, w_035_2809, w_035_2810, w_035_2811, w_035_2812, w_035_2813, w_035_2814, w_035_2816, w_035_2818, w_035_2819, w_035_2821, w_035_2822, w_035_2823, w_035_2824, w_035_2825, w_035_2826, w_035_2827, w_035_2828, w_035_2829, w_035_2830, w_035_2833, w_035_2835, w_035_2836, w_035_2838, w_035_2839, w_035_2840, w_035_2842, w_035_2843, w_035_2844, w_035_2845, w_035_2848, w_035_2849, w_035_2850, w_035_2851, w_035_2852, w_035_2853, w_035_2854, w_035_2855, w_035_2856, w_035_2857, w_035_2858, w_035_2859, w_035_2861, w_035_2862, w_035_2863, w_035_2864, w_035_2865, w_035_2866, w_035_2867, w_035_2868, w_035_2871, w_035_2872, w_035_2873, w_035_2875, w_035_2876, w_035_2877, w_035_2878, w_035_2879, w_035_2880, w_035_2882, w_035_2883, w_035_2884, w_035_2885, w_035_2886, w_035_2887, w_035_2889, w_035_2890, w_035_2891, w_035_2892, w_035_2893, w_035_2894, w_035_2895, w_035_2896, w_035_2898, w_035_2899, w_035_2901, w_035_2902, w_035_2903, w_035_2904, w_035_2905, w_035_2906, w_035_2907, w_035_2908, w_035_2911, w_035_2914, w_035_2916, w_035_2917, w_035_2918, w_035_2919, w_035_2920, w_035_2921, w_035_2923, w_035_2924, w_035_2926, w_035_2928, w_035_2929, w_035_2930, w_035_2931, w_035_2932, w_035_2933, w_035_2935, w_035_2936, w_035_2937, w_035_2938, w_035_2939, w_035_2940, w_035_2941, w_035_2943, w_035_2945, w_035_2946, w_035_2948, w_035_2949, w_035_2950, w_035_2951, w_035_2952, w_035_2953, w_035_2954, w_035_2955, w_035_2958, w_035_2960, w_035_2961, w_035_2963, w_035_2964, w_035_2965, w_035_2966, w_035_2967, w_035_2968, w_035_2969, w_035_2970, w_035_2971, w_035_2972, w_035_2973, w_035_2974, w_035_2977, w_035_2979, w_035_2980, w_035_2981, w_035_2982, w_035_2983, w_035_2984, w_035_2985, w_035_2986, w_035_2987, w_035_2988, w_035_2991, w_035_2992, w_035_2993, w_035_2994, w_035_2995, w_035_2996, w_035_2997, w_035_2998, w_035_2999, w_035_3000, w_035_3003, w_035_3004, w_035_3006, w_035_3007, w_035_3008, w_035_3010, w_035_3011, w_035_3012, w_035_3013, w_035_3014, w_035_3015, w_035_3022, w_035_3023, w_035_3024, w_035_3025, w_035_3026, w_035_3027, w_035_3029, w_035_3030, w_035_3032, w_035_3036, w_035_3037, w_035_3038, w_035_3039, w_035_3040, w_035_3041, w_035_3042, w_035_3044, w_035_3045, w_035_3046, w_035_3047, w_035_3051, w_035_3053, w_035_3054, w_035_3055, w_035_3056, w_035_3057, w_035_3058, w_035_3060, w_035_3062, w_035_3063, w_035_3066, w_035_3067, w_035_3068, w_035_3069, w_035_3070, w_035_3072, w_035_3073, w_035_3075, w_035_3076, w_035_3077, w_035_3078, w_035_3079, w_035_3080, w_035_3081, w_035_3082, w_035_3083, w_035_3084, w_035_3085, w_035_3087, w_035_3088, w_035_3092, w_035_3093, w_035_3094, w_035_3095, w_035_3098, w_035_3100, w_035_3101, w_035_3103, w_035_3104, w_035_3106, w_035_3107, w_035_3108, w_035_3109, w_035_3110, w_035_3111, w_035_3112, w_035_3113, w_035_3115, w_035_3116, w_035_3117, w_035_3119, w_035_3120, w_035_3121, w_035_3122, w_035_3123, w_035_3124, w_035_3125, w_035_3127, w_035_3128, w_035_3129, w_035_3130, w_035_3132, w_035_3133, w_035_3134, w_035_3135, w_035_3138, w_035_3140, w_035_3141, w_035_3142, w_035_3144, w_035_3145, w_035_3147, w_035_3149, w_035_3150, w_035_3151, w_035_3152, w_035_3153, w_035_3154, w_035_3155, w_035_3156, w_035_3157, w_035_3158, w_035_3159, w_035_3162, w_035_3166, w_035_3167, w_035_3168, w_035_3169, w_035_3170, w_035_3173, w_035_3174, w_035_3176, w_035_3177, w_035_3178, w_035_3181, w_035_3182, w_035_3183, w_035_3184, w_035_3185, w_035_3186, w_035_3187, w_035_3188, w_035_3193, w_035_3194, w_035_3195, w_035_3199, w_035_3200, w_035_3205, w_035_3206, w_035_3207, w_035_3208, w_035_3209, w_035_3210, w_035_3211, w_035_3212, w_035_3214, w_035_3215, w_035_3216, w_035_3218, w_035_3219, w_035_3224, w_035_3225, w_035_3227, w_035_3230, w_035_3232, w_035_3233, w_035_3234, w_035_3235, w_035_3237, w_035_3238, w_035_3239, w_035_3240, w_035_3242, w_035_3243, w_035_3244, w_035_3245, w_035_3248, w_035_3250, w_035_3253, w_035_3254, w_035_3255, w_035_3257, w_035_3258, w_035_3259, w_035_3260, w_035_3261, w_035_3262, w_035_3264, w_035_3265, w_035_3266, w_035_3268, w_035_3271, w_035_3272, w_035_3273, w_035_3274, w_035_3275, w_035_3276, w_035_3278, w_035_3279, w_035_3280, w_035_3282, w_035_3283, w_035_3285, w_035_3286, w_035_3287, w_035_3288, w_035_3289, w_035_3291, w_035_3293, w_035_3296, w_035_3297, w_035_3299, w_035_3300, w_035_3301, w_035_3302, w_035_3304, w_035_3305, w_035_3306, w_035_3307, w_035_3309, w_035_3310, w_035_3314, w_035_3315, w_035_3317, w_035_3318, w_035_3319, w_035_3321, w_035_3322, w_035_3323, w_035_3324, w_035_3325, w_035_3326, w_035_3328, w_035_3330, w_035_3332, w_035_3333, w_035_3334, w_035_3335, w_035_3336, w_035_3337, w_035_3338, w_035_3339, w_035_3340, w_035_3341, w_035_3343, w_035_3344, w_035_3348, w_035_3349, w_035_3350, w_035_3352, w_035_3353, w_035_3354, w_035_3355, w_035_3357, w_035_3359, w_035_3360, w_035_3363, w_035_3364, w_035_3365, w_035_3366, w_035_3367, w_035_3368, w_035_3369, w_035_3370, w_035_3372, w_035_3373, w_035_3374, w_035_3375, w_035_3376, w_035_3377, w_035_3378, w_035_3379, w_035_3380, w_035_3382, w_035_3384, w_035_3385, w_035_3386, w_035_3387, w_035_3388, w_035_3389, w_035_3390, w_035_3391, w_035_3392, w_035_3393, w_035_3395, w_035_3396, w_035_3397, w_035_3398, w_035_3400, w_035_3402, w_035_3403, w_035_3406, w_035_3407, w_035_3408, w_035_3409, w_035_3410, w_035_3412, w_035_3413, w_035_3414, w_035_3415, w_035_3416, w_035_3417, w_035_3418, w_035_3420, w_035_3422, w_035_3424, w_035_3426, w_035_3427, w_035_3430, w_035_3431, w_035_3433, w_035_3434, w_035_3435, w_035_3437, w_035_3438, w_035_3441, w_035_3442, w_035_3443, w_035_3444, w_035_3445, w_035_3446, w_035_3447, w_035_3448, w_035_3450, w_035_3451, w_035_3452, w_035_3453, w_035_3454, w_035_3455, w_035_3456, w_035_3458, w_035_3459, w_035_3462, w_035_3463, w_035_3464, w_035_3465, w_035_3467, w_035_3468, w_035_3469, w_035_3470, w_035_3471, w_035_3472, w_035_3473, w_035_3474, w_035_3475, w_035_3476, w_035_3478, w_035_3480, w_035_3481, w_035_3482, w_035_3483, w_035_3484, w_035_3485, w_035_3487, w_035_3488, w_035_3489, w_035_3490, w_035_3492, w_035_3493, w_035_3494, w_035_3495, w_035_3496, w_035_3498, w_035_3499, w_035_3500, w_035_3501, w_035_3502, w_035_3503, w_035_3505, w_035_3506, w_035_3507, w_035_3508, w_035_3510, w_035_3511, w_035_3513, w_035_3515, w_035_3516, w_035_3518, w_035_3519, w_035_3520, w_035_3521, w_035_3522, w_035_3524, w_035_3525, w_035_3527, w_035_3528, w_035_3529, w_035_3530, w_035_3531, w_035_3532, w_035_3534, w_035_3536, w_035_3537, w_035_3538, w_035_3539, w_035_3540, w_035_3541, w_035_3542, w_035_3543, w_035_3544, w_035_3546, w_035_3548, w_035_3549, w_035_3550, w_035_3552, w_035_3554, w_035_3556, w_035_3557, w_035_3559, w_035_3560, w_035_3561, w_035_3562, w_035_3563, w_035_3564, w_035_3565, w_035_3567, w_035_3568, w_035_3569, w_035_3570, w_035_3571, w_035_3572, w_035_3574, w_035_3575, w_035_3576, w_035_3578, w_035_3579, w_035_3580, w_035_3582, w_035_3583, w_035_3584, w_035_3585, w_035_3588, w_035_3589, w_035_3590, w_035_3591, w_035_3592, w_035_3593, w_035_3595, w_035_3597, w_035_3599, w_035_3600, w_035_3601, w_035_3602, w_035_3603, w_035_3604, w_035_3605, w_035_3606, w_035_3607, w_035_3608, w_035_3609, w_035_3611, w_035_3612, w_035_3616, w_035_3617, w_035_3618, w_035_3619, w_035_3620, w_035_3621, w_035_3622, w_035_3623, w_035_3624, w_035_3625, w_035_3626, w_035_3627, w_035_3628, w_035_3629, w_035_3630, w_035_3632, w_035_3633, w_035_3634, w_035_3636, w_035_3638, w_035_3639, w_035_3640, w_035_3641, w_035_3642, w_035_3643, w_035_3644, w_035_3645, w_035_3646, w_035_3647, w_035_3648, w_035_3649, w_035_3650, w_035_3652, w_035_3655, w_035_3656, w_035_3658, w_035_3660, w_035_3661, w_035_3662, w_035_3663, w_035_3664, w_035_3666, w_035_3667, w_035_3668, w_035_3669, w_035_3671, w_035_3672, w_035_3674, w_035_3675, w_035_3676, w_035_3677, w_035_3678, w_035_3679, w_035_3680, w_035_3681, w_035_3682, w_035_3683, w_035_3685, w_035_3686, w_035_3687, w_035_3689, w_035_3690, w_035_3691, w_035_3692, w_035_3694, w_035_3695, w_035_3696, w_035_3698, w_035_3699, w_035_3701, w_035_3702, w_035_3703, w_035_3704, w_035_3705, w_035_3706, w_035_3708, w_035_3709, w_035_3710, w_035_3711, w_035_3714, w_035_3715, w_035_3716, w_035_3717, w_035_3719, w_035_3720, w_035_3721, w_035_3723, w_035_3724, w_035_3725, w_035_3726, w_035_3727, w_035_3728, w_035_3729, w_035_3731, w_035_3732, w_035_3734, w_035_3735, w_035_3736, w_035_3737, w_035_3738, w_035_3740, w_035_3741, w_035_3745, w_035_3746, w_035_3747, w_035_3748, w_035_3749, w_035_3751, w_035_3753, w_035_3754, w_035_3755, w_035_3757, w_035_3758, w_035_3761, w_035_3763, w_035_3764, w_035_3765, w_035_3767, w_035_3768, w_035_3769, w_035_3770, w_035_3771, w_035_3772, w_035_3773, w_035_3774, w_035_3776, w_035_3778, w_035_3779, w_035_3780, w_035_3781, w_035_3782, w_035_3783, w_035_3784, w_035_3785, w_035_3786, w_035_3787, w_035_3788, w_035_3789, w_035_3790, w_035_3791, w_035_3792, w_035_3793, w_035_3795, w_035_3796, w_035_3798, w_035_3799, w_035_3800, w_035_3801, w_035_3802, w_035_3803, w_035_3804, w_035_3805, w_035_3806, w_035_3807, w_035_3808, w_035_3809, w_035_3811, w_035_3813, w_035_3815, w_035_3816, w_035_3818, w_035_3820, w_035_3821, w_035_3823, w_035_3824, w_035_3826, w_035_3827, w_035_3828, w_035_3829, w_035_3830, w_035_3831, w_035_3832, w_035_3835, w_035_3837, w_035_3839, w_035_3841, w_035_3842, w_035_3843, w_035_3844, w_035_3846, w_035_3847, w_035_3850, w_035_3851, w_035_3852, w_035_3853, w_035_3854, w_035_3858, w_035_3859, w_035_3860, w_035_3861, w_035_3862, w_035_3864, w_035_3869, w_035_3870, w_035_3871, w_035_3875, w_035_3876, w_035_3879, w_035_3880, w_035_3881, w_035_3882, w_035_3883, w_035_3884, w_035_3885, w_035_3886, w_035_3888, w_035_3889, w_035_3890, w_035_3891, w_035_3892, w_035_3893, w_035_3894, w_035_3895, w_035_3897, w_035_3899, w_035_3900, w_035_3901, w_035_3902, w_035_3903, w_035_3904, w_035_3905, w_035_3906, w_035_3907, w_035_3910, w_035_3911, w_035_3912, w_035_3914, w_035_3915, w_035_3916, w_035_3919, w_035_3920, w_035_3921, w_035_3922, w_035_3923, w_035_3924, w_035_3926, w_035_3929, w_035_3930, w_035_3932, w_035_3934, w_035_3935, w_035_3936, w_035_3937, w_035_3938, w_035_3939, w_035_3942, w_035_3943, w_035_3944, w_035_3946, w_035_3947, w_035_3949, w_035_3950, w_035_3953, w_035_3954, w_035_3956, w_035_3958, w_035_3959, w_035_3960, w_035_3962, w_035_3963, w_035_3964, w_035_3965, w_035_3966, w_035_3967, w_035_3970, w_035_3971, w_035_3973, w_035_3975, w_035_3976, w_035_3978, w_035_3979, w_035_3980, w_035_3981, w_035_3983, w_035_3984, w_035_3986, w_035_3987, w_035_3988, w_035_3990, w_035_3991, w_035_3992, w_035_3993, w_035_3995, w_035_3996, w_035_3997, w_035_3998, w_035_4000, w_035_4001, w_035_4002, w_035_4003, w_035_4004, w_035_4005, w_035_4007, w_035_4008, w_035_4009, w_035_4010, w_035_4011, w_035_4012, w_035_4013, w_035_4014, w_035_4015, w_035_4016, w_035_4017, w_035_4018, w_035_4019, w_035_4020, w_035_4021, w_035_4022, w_035_4023, w_035_4024, w_035_4025, w_035_4026, w_035_4027, w_035_4029, w_035_4030, w_035_4032, w_035_4033, w_035_4034, w_035_4035, w_035_4036, w_035_4040, w_035_4041, w_035_4043, w_035_4045, w_035_4046, w_035_4047, w_035_4049, w_035_4050, w_035_4051, w_035_4052, w_035_4053, w_035_4054, w_035_4055, w_035_4056, w_035_4057, w_035_4058, w_035_4060, w_035_4061, w_035_4062, w_035_4063, w_035_4064, w_035_4066, w_035_4067, w_035_4068, w_035_4069, w_035_4070, w_035_4071, w_035_4072, w_035_4074, w_035_4075, w_035_4078, w_035_4080, w_035_4081, w_035_4082, w_035_4083, w_035_4084, w_035_4085, w_035_4086, w_035_4088, w_035_4093, w_035_4094, w_035_4096, w_035_4097, w_035_4098, w_035_4099, w_035_4100, w_035_4101, w_035_4104, w_035_4105, w_035_4106, w_035_4107, w_035_4109, w_035_4111, w_035_4112, w_035_4113, w_035_4114, w_035_4117, w_035_4120, w_035_4121, w_035_4122, w_035_4124, w_035_4125, w_035_4127, w_035_4129, w_035_4130, w_035_4132, w_035_4134, w_035_4135, w_035_4136, w_035_4141, w_035_4142, w_035_4145, w_035_4147, w_035_4148, w_035_4149, w_035_4150, w_035_4153, w_035_4156, w_035_4159, w_035_4161, w_035_4162, w_035_4164, w_035_4165, w_035_4166, w_035_4167, w_035_4169, w_035_4170, w_035_4171, w_035_4173, w_035_4174, w_035_4176, w_035_4178, w_035_4179, w_035_4182, w_035_4183, w_035_4185, w_035_4187, w_035_4188, w_035_4189, w_035_4190, w_035_4191, w_035_4195, w_035_4196, w_035_4197, w_035_4199, w_035_4203, w_035_4204, w_035_4205, w_035_4206, w_035_4207, w_035_4208, w_035_4211, w_035_4214, w_035_4215, w_035_4216, w_035_4217, w_035_4219, w_035_4222, w_035_4223, w_035_4225, w_035_4227, w_035_4228, w_035_4231, w_035_4236, w_035_4238, w_035_4239, w_035_4242, w_035_4245, w_035_4249, w_035_4254, w_035_4255, w_035_4256, w_035_4257, w_035_4259, w_035_4261, w_035_4262, w_035_4266, w_035_4267, w_035_4268, w_035_4269, w_035_4270, w_035_4271, w_035_4272, w_035_4275, w_035_4276, w_035_4277, w_035_4279, w_035_4280, w_035_4281, w_035_4284, w_035_4285, w_035_4287, w_035_4288, w_035_4289, w_035_4290, w_035_4296, w_035_4297, w_035_4299, w_035_4302, w_035_4304, w_035_4305, w_035_4308, w_035_4309, w_035_4312, w_035_4313, w_035_4314, w_035_4315, w_035_4318, w_035_4320, w_035_4321, w_035_4322, w_035_4324, w_035_4325, w_035_4326, w_035_4328, w_035_4331, w_035_4335, w_035_4337, w_035_4338, w_035_4342, w_035_4343, w_035_4344, w_035_4345, w_035_4346, w_035_4348, w_035_4351, w_035_4352, w_035_4354, w_035_4356, w_035_4357, w_035_4359, w_035_4360, w_035_4361, w_035_4363, w_035_4365, w_035_4366, w_035_4369, w_035_4370, w_035_4375, w_035_4377, w_035_4378, w_035_4383, w_035_4384, w_035_4386, w_035_4387, w_035_4389, w_035_4390, w_035_4391, w_035_4392, w_035_4394, w_035_4395, w_035_4398, w_035_4399, w_035_4402, w_035_4403, w_035_4405, w_035_4409, w_035_4410, w_035_4411, w_035_4413, w_035_4415, w_035_4416, w_035_4417, w_035_4419, w_035_4421, w_035_4422, w_035_4423, w_035_4424, w_035_4425, w_035_4426, w_035_4427, w_035_4429, w_035_4432, w_035_4433, w_035_4434, w_035_4435, w_035_4440, w_035_4441, w_035_4443, w_035_4444, w_035_4445, w_035_4449, w_035_4450, w_035_4452, w_035_4453, w_035_4455, w_035_4457, w_035_4458, w_035_4465, w_035_4466, w_035_4467, w_035_4468, w_035_4470, w_035_4472, w_035_4476, w_035_4479, w_035_4480, w_035_4482, w_035_4483, w_035_4486, w_035_4487, w_035_4490, w_035_4491, w_035_4494, w_035_4495, w_035_4497, w_035_4498, w_035_4499, w_035_4501, w_035_4506, w_035_4507, w_035_4509, w_035_4512, w_035_4513, w_035_4515, w_035_4517, w_035_4518, w_035_4520, w_035_4522, w_035_4524, w_035_4525, w_035_4526, w_035_4527, w_035_4530, w_035_4532, w_035_4533, w_035_4535, w_035_4538, w_035_4539, w_035_4540, w_035_4542, w_035_4543, w_035_4545, w_035_4546, w_035_4547, w_035_4550, w_035_4551, w_035_4553, w_035_4556, w_035_4559, w_035_4560, w_035_4561, w_035_4562, w_035_4571, w_035_4573, w_035_4574, w_035_4576, w_035_4577, w_035_4578, w_035_4579, w_035_4580, w_035_4581, w_035_4585, w_035_4587, w_035_4588, w_035_4591, w_035_4592, w_035_4595, w_035_4596, w_035_4597, w_035_4599, w_035_4602, w_035_4603, w_035_4604, w_035_4606, w_035_4608, w_035_4612, w_035_4614, w_035_4615, w_035_4617, w_035_4621, w_035_4624, w_035_4626, w_035_4627, w_035_4629, w_035_4630, w_035_4631, w_035_4633, w_035_4634, w_035_4636, w_035_4637, w_035_4638, w_035_4639, w_035_4642, w_035_4643, w_035_4645, w_035_4646, w_035_4647, w_035_4648, w_035_4649, w_035_4650, w_035_4651, w_035_4652, w_035_4653, w_035_4658, w_035_4659, w_035_4661, w_035_4663, w_035_4666, w_035_4669, w_035_4671, w_035_4672, w_035_4676, w_035_4677, w_035_4678, w_035_4679, w_035_4681, w_035_4682, w_035_4683, w_035_4685, w_035_4686, w_035_4687, w_035_4690, w_035_4691, w_035_4693, w_035_4696, w_035_4697, w_035_4698, w_035_4699, w_035_4702, w_035_4703, w_035_4706, w_035_4707, w_035_4710, w_035_4711, w_035_4712, w_035_4713, w_035_4714, w_035_4715, w_035_4716, w_035_4717, w_035_4721, w_035_4724, w_035_4725, w_035_4726, w_035_4727, w_035_4728, w_035_4730, w_035_4731, w_035_4732, w_035_4734, w_035_4738, w_035_4739, w_035_4741, w_035_4742, w_035_4744, w_035_4746, w_035_4748, w_035_4750, w_035_4751, w_035_4754, w_035_4755, w_035_4762, w_035_4764, w_035_4765, w_035_4767, w_035_4771, w_035_4773, w_035_4775, w_035_4777, w_035_4779, w_035_4782, w_035_4784, w_035_4790, w_035_4793, w_035_4794, w_035_4795, w_035_4798, w_035_4800, w_035_4803, w_035_4805, w_035_4806, w_035_4807, w_035_4809, w_035_4810, w_035_4814, w_035_4815, w_035_4816, w_035_4817, w_035_4818, w_035_4819, w_035_4821, w_035_4824, w_035_4826, w_035_4828, w_035_4830, w_035_4833, w_035_4834, w_035_4837, w_035_4839, w_035_4840, w_035_4843, w_035_4847, w_035_4848, w_035_4852, w_035_4853, w_035_4855, w_035_4856, w_035_4857, w_035_4861, w_035_4863, w_035_4868, w_035_4869, w_035_4870, w_035_4871, w_035_4873, w_035_4874, w_035_4875, w_035_4876, w_035_4879, w_035_4880, w_035_4882, w_035_4884, w_035_4886, w_035_4887, w_035_4889, w_035_4893, w_035_4894, w_035_4895, w_035_4897, w_035_4898, w_035_4899, w_035_4904, w_035_4905, w_035_4909, w_035_4910, w_035_4911, w_035_4912, w_035_4913, w_035_4914, w_035_4916, w_035_4917, w_035_4919, w_035_4925, w_035_4926, w_035_4927, w_035_4929, w_035_4935, w_035_4938, w_035_4939, w_035_4940, w_035_4941, w_035_4944, w_035_4947, w_035_4948, w_035_4950, w_035_4952, w_035_4956, w_035_4957, w_035_4959, w_035_4962, w_035_4963, w_035_4965, w_035_4966, w_035_4968, w_035_4969, w_035_4971, w_035_4972, w_035_4973, w_035_4976, w_035_4978, w_035_4980, w_035_4982, w_035_4983, w_035_4985, w_035_4986, w_035_4987, w_035_4988, w_035_4990, w_035_4991, w_035_4992, w_035_4993, w_035_4994, w_035_4995, w_035_4996, w_035_4999, w_035_5002, w_035_5003, w_035_5004, w_035_5005, w_035_5010, w_035_5016, w_035_5017, w_035_5018, w_035_5019, w_035_5020, w_035_5021, w_035_5023, w_035_5024, w_035_5026, w_035_5028, w_035_5029, w_035_5030, w_035_5031, w_035_5033, w_035_5035, w_035_5036, w_035_5038, w_035_5039, w_035_5040, w_035_5043, w_035_5046, w_035_5050, w_035_5054, w_035_5057, w_035_5058, w_035_5059, w_035_5060, w_035_5061, w_035_5067, w_035_5068, w_035_5069, w_035_5072, w_035_5073, w_035_5076, w_035_5078, w_035_5082, w_035_5086, w_035_5088, w_035_5089, w_035_5090, w_035_5092, w_035_5093, w_035_5095, w_035_5098, w_035_5099, w_035_5104, w_035_5105, w_035_5106, w_035_5108, w_035_5109, w_035_5110, w_035_5112, w_035_5114, w_035_5115, w_035_5116, w_035_5117, w_035_5118, w_035_5119, w_035_5122, w_035_5123, w_035_5124, w_035_5125, w_035_5128, w_035_5129, w_035_5130, w_035_5133, w_035_5135, w_035_5137, w_035_5138, w_035_5139, w_035_5142, w_035_5147, w_035_5148, w_035_5149, w_035_5151, w_035_5153, w_035_5154, w_035_5158, w_035_5161, w_035_5164, w_035_5165, w_035_5166, w_035_5171, w_035_5172, w_035_5174, w_035_5176, w_035_5177, w_035_5178, w_035_5180, w_035_5181, w_035_5182, w_035_5183, w_035_5184, w_035_5185, w_035_5187, w_035_5189, w_035_5194, w_035_5195, w_035_5196, w_035_5197, w_035_5200, w_035_5201, w_035_5203, w_035_5205, w_035_5211, w_035_5215, w_035_5217, w_035_5218, w_035_5219, w_035_5220, w_035_5221, w_035_5223, w_035_5225, w_035_5229, w_035_5230, w_035_5234, w_035_5235, w_035_5238, w_035_5241, w_035_5242, w_035_5243, w_035_5244, w_035_5245, w_035_5246, w_035_5247, w_035_5251, w_035_5252, w_035_5253, w_035_5256, w_035_5259, w_035_5261, w_035_5263, w_035_5264, w_035_5265, w_035_5266, w_035_5267, w_035_5268, w_035_5269, w_035_5271, w_035_5274, w_035_5276, w_035_5277, w_035_5278, w_035_5283, w_035_5286, w_035_5288, w_035_5292, w_035_5298, w_035_5299, w_035_5300, w_035_5301, w_035_5302, w_035_5304, w_035_5310, w_035_5311, w_035_5312, w_035_5313, w_035_5314, w_035_5315, w_035_5317, w_035_5320, w_035_5321, w_035_5322, w_035_5324, w_035_5326, w_035_5327, w_035_5328, w_035_5329, w_035_5330, w_035_5331, w_035_5333, w_035_5336, w_035_5337, w_035_5338, w_035_5342, w_035_5344, w_035_5345, w_035_5347, w_035_5349, w_035_5350, w_035_5351, w_035_5352, w_035_5355, w_035_5360, w_035_5362, w_035_5365, w_035_5367, w_035_5368, w_035_5369, w_035_5371, w_035_5374, w_035_5376, w_035_5377, w_035_5378, w_035_5382, w_035_5383, w_035_5386, w_035_5387, w_035_5392, w_035_5395, w_035_5396, w_035_5397, w_035_5399, w_035_5400, w_035_5403, w_035_5404, w_035_5406, w_035_5408, w_035_5409, w_035_5410, w_035_5412, w_035_5416, w_035_5418, w_035_5419, w_035_5420, w_035_5422, w_035_5423, w_035_5430, w_035_5433, w_035_5436, w_035_5439, w_035_5441, w_035_5443, w_035_5444, w_035_5447, w_035_5449, w_035_5450, w_035_5451, w_035_5454, w_035_5455, w_035_5456, w_035_5457, w_035_5459, w_035_5460, w_035_5461, w_035_5462, w_035_5463, w_035_5467, w_035_5470, w_035_5471, w_035_5472, w_035_5475, w_035_5476, w_035_5479, w_035_5480, w_035_5484, w_035_5485, w_035_5486, w_035_5487, w_035_5492, w_035_5493, w_035_5494, w_035_5499, w_035_5500, w_035_5501, w_035_5502, w_035_5503, w_035_5504, w_035_5506, w_035_5508, w_035_5509, w_035_5511, w_035_5513, w_035_5514, w_035_5518, w_035_5520, w_035_5523, w_035_5525, w_035_5526, w_035_5528, w_035_5529, w_035_5531, w_035_5532, w_035_5533, w_035_5534, w_035_5536, w_035_5540, w_035_5541, w_035_5542, w_035_5544, w_035_5546, w_035_5547, w_035_5552, w_035_5554, w_035_5557, w_035_5558, w_035_5560, w_035_5562, w_035_5564, w_035_5573, w_035_5575, w_035_5576, w_035_5577, w_035_5579, w_035_5582, w_035_5584, w_035_5585, w_035_5586, w_035_5588, w_035_5589, w_035_5590, w_035_5591, w_035_5592, w_035_5597, w_035_5598, w_035_5600, w_035_5601, w_035_5602, w_035_5603, w_035_5607, w_035_5609, w_035_5611, w_035_5614, w_035_5617, w_035_5620, w_035_5621, w_035_5626, w_035_5627, w_035_5629, w_035_5630, w_035_5633, w_035_5634, w_035_5636, w_035_5638, w_035_5640, w_035_5642, w_035_5643, w_035_5644, w_035_5646, w_035_5647, w_035_5648, w_035_5651, w_035_5653, w_035_5657, w_035_5660, w_035_5661, w_035_5663, w_035_5666, w_035_5667, w_035_5670, w_035_5673, w_035_5674, w_035_5678, w_035_5683, w_035_5684, w_035_5687, w_035_5689, w_035_5690, w_035_5691, w_035_5692, w_035_5693, w_035_5695, w_035_5698, w_035_5699, w_035_5700, w_035_5701, w_035_5702, w_035_5710, w_035_5711, w_035_5712, w_035_5714, w_035_5719, w_035_5720, w_035_5721, w_035_5722, w_035_5723, w_035_5724, w_035_5725, w_035_5726, w_035_5727, w_035_5730, w_035_5732, w_035_5735, w_035_5736, w_035_5738, w_035_5739, w_035_5740, w_035_5741, w_035_5742, w_035_5743, w_035_5745, w_035_5748, w_035_5751, w_035_5755, w_035_5757, w_035_5761, w_035_5762, w_035_5763, w_035_5764, w_035_5770, w_035_5771, w_035_5774, w_035_5779, w_035_5780, w_035_5781, w_035_5783, w_035_5786, w_035_5787, w_035_5788, w_035_5789, w_035_5794, w_035_5796, w_035_5797, w_035_5798, w_035_5801, w_035_5802, w_035_5805, w_035_5808, w_035_5809, w_035_5810, w_035_5811, w_035_5813, w_035_5814, w_035_5816, w_035_5817, w_035_5819, w_035_5820, w_035_5821, w_035_5822, w_035_5825, w_035_5826, w_035_5827, w_035_5831, w_035_5833, w_035_5834, w_035_5835, w_035_5837, w_035_5838, w_035_5839, w_035_5840, w_035_5841, w_035_5844, w_035_5846, w_035_5847, w_035_5852, w_035_5856, w_035_5857, w_035_5860, w_035_5862, w_035_5863, w_035_5864, w_035_5865, w_035_5866;
  wire w_036_000, w_036_001, w_036_002, w_036_003, w_036_004, w_036_005, w_036_006, w_036_007, w_036_008, w_036_009, w_036_010, w_036_011, w_036_012, w_036_013, w_036_014, w_036_015, w_036_016, w_036_017, w_036_018, w_036_019, w_036_020, w_036_021, w_036_022, w_036_023, w_036_024, w_036_025, w_036_026, w_036_027, w_036_028, w_036_029, w_036_030, w_036_031, w_036_032, w_036_033, w_036_034, w_036_035, w_036_036, w_036_037, w_036_038, w_036_039, w_036_040, w_036_041, w_036_042, w_036_043, w_036_044, w_036_045, w_036_046, w_036_047, w_036_048, w_036_049, w_036_050, w_036_051, w_036_052, w_036_053, w_036_054, w_036_055, w_036_056, w_036_057, w_036_058, w_036_059, w_036_060, w_036_061, w_036_062, w_036_063, w_036_064, w_036_065, w_036_066, w_036_067, w_036_068, w_036_069, w_036_070, w_036_071, w_036_072, w_036_073, w_036_074, w_036_075, w_036_076, w_036_077, w_036_078, w_036_079, w_036_080, w_036_081, w_036_082, w_036_083, w_036_084, w_036_085, w_036_086, w_036_087, w_036_088, w_036_089, w_036_090, w_036_091, w_036_092, w_036_093, w_036_094, w_036_095, w_036_096, w_036_097, w_036_098, w_036_099, w_036_100, w_036_101, w_036_102, w_036_103, w_036_104, w_036_105, w_036_106, w_036_107, w_036_108, w_036_109, w_036_110, w_036_111, w_036_112, w_036_113, w_036_114, w_036_115, w_036_116, w_036_117, w_036_118, w_036_119, w_036_120, w_036_121, w_036_122, w_036_123, w_036_124, w_036_125, w_036_126, w_036_127, w_036_128, w_036_129, w_036_130, w_036_131, w_036_132, w_036_133, w_036_134, w_036_135, w_036_136, w_036_137, w_036_138, w_036_139, w_036_140, w_036_141, w_036_142, w_036_143, w_036_144, w_036_145, w_036_146, w_036_147, w_036_148, w_036_149, w_036_150, w_036_151, w_036_152, w_036_153, w_036_154, w_036_155, w_036_156, w_036_157, w_036_158, w_036_159, w_036_160, w_036_161, w_036_162, w_036_163, w_036_164, w_036_165, w_036_166, w_036_167, w_036_168, w_036_169, w_036_170, w_036_171, w_036_172, w_036_173, w_036_174, w_036_175, w_036_176, w_036_177, w_036_178, w_036_179, w_036_180, w_036_181, w_036_182, w_036_183, w_036_184, w_036_185, w_036_186, w_036_187, w_036_188, w_036_189, w_036_190, w_036_191, w_036_192, w_036_193, w_036_194, w_036_195, w_036_196, w_036_197, w_036_198, w_036_199, w_036_200, w_036_201, w_036_202, w_036_203, w_036_204, w_036_205, w_036_206, w_036_207, w_036_208, w_036_209, w_036_210, w_036_211, w_036_212, w_036_213, w_036_214, w_036_215, w_036_216, w_036_217, w_036_218, w_036_219, w_036_220, w_036_221, w_036_222, w_036_223, w_036_224, w_036_225, w_036_226, w_036_227, w_036_228, w_036_229, w_036_230, w_036_231, w_036_232, w_036_233, w_036_234, w_036_235, w_036_236, w_036_237, w_036_238, w_036_239, w_036_240, w_036_241, w_036_242, w_036_243, w_036_244, w_036_245, w_036_246, w_036_247, w_036_248, w_036_249, w_036_250, w_036_251, w_036_252, w_036_253, w_036_254, w_036_255, w_036_256, w_036_257, w_036_258, w_036_259, w_036_260, w_036_261, w_036_262, w_036_263, w_036_264, w_036_265, w_036_266, w_036_267, w_036_268, w_036_269, w_036_270, w_036_271, w_036_272, w_036_273, w_036_274, w_036_275, w_036_276, w_036_277, w_036_278, w_036_279, w_036_280, w_036_281, w_036_282, w_036_283, w_036_284, w_036_285, w_036_286, w_036_287, w_036_288, w_036_289, w_036_290, w_036_291, w_036_292, w_036_293, w_036_294, w_036_295, w_036_296, w_036_297, w_036_298, w_036_299, w_036_300, w_036_301, w_036_302, w_036_303, w_036_304, w_036_305, w_036_306, w_036_307, w_036_308, w_036_309, w_036_310, w_036_311, w_036_312, w_036_313, w_036_314, w_036_315, w_036_316, w_036_317, w_036_318, w_036_319, w_036_320, w_036_321, w_036_322, w_036_323, w_036_324, w_036_325, w_036_326, w_036_327, w_036_328, w_036_329, w_036_330, w_036_331, w_036_332, w_036_333, w_036_334, w_036_335, w_036_336, w_036_337, w_036_338, w_036_339, w_036_340, w_036_341, w_036_342, w_036_343, w_036_344, w_036_345, w_036_346, w_036_347, w_036_348, w_036_349, w_036_350, w_036_351, w_036_352, w_036_353, w_036_354, w_036_355, w_036_356, w_036_357, w_036_358, w_036_359, w_036_360, w_036_361, w_036_362, w_036_363, w_036_364, w_036_365, w_036_366, w_036_367, w_036_368, w_036_369, w_036_370, w_036_371, w_036_372, w_036_373, w_036_374, w_036_375, w_036_376, w_036_377, w_036_378, w_036_379, w_036_380, w_036_381, w_036_382, w_036_383, w_036_384, w_036_385, w_036_386, w_036_387, w_036_388, w_036_389, w_036_390, w_036_391, w_036_392, w_036_393, w_036_394, w_036_395, w_036_396, w_036_397, w_036_398, w_036_399, w_036_400, w_036_401, w_036_402, w_036_403, w_036_404, w_036_405, w_036_406, w_036_407, w_036_408, w_036_409, w_036_410, w_036_411, w_036_412, w_036_413, w_036_414, w_036_415, w_036_416, w_036_417, w_036_418, w_036_419, w_036_420, w_036_421, w_036_422, w_036_423, w_036_424, w_036_425, w_036_426, w_036_427, w_036_428, w_036_429, w_036_430, w_036_431, w_036_432, w_036_433, w_036_434, w_036_435, w_036_436, w_036_437, w_036_438, w_036_439, w_036_440, w_036_441, w_036_442, w_036_443, w_036_444, w_036_445, w_036_446, w_036_447, w_036_448, w_036_449, w_036_450, w_036_451, w_036_452, w_036_453, w_036_454, w_036_455, w_036_456, w_036_457, w_036_458, w_036_459, w_036_460, w_036_461, w_036_462, w_036_463, w_036_464, w_036_465, w_036_466, w_036_467, w_036_468, w_036_469, w_036_470, w_036_471, w_036_472, w_036_473, w_036_474, w_036_475, w_036_476, w_036_477, w_036_478, w_036_479, w_036_480, w_036_481, w_036_482, w_036_483, w_036_484, w_036_485, w_036_486, w_036_487, w_036_488, w_036_489, w_036_490, w_036_491, w_036_492, w_036_493, w_036_494, w_036_495, w_036_496, w_036_497, w_036_498, w_036_499, w_036_500, w_036_501, w_036_502, w_036_503, w_036_504, w_036_505, w_036_506, w_036_507, w_036_508, w_036_509, w_036_510, w_036_511, w_036_512, w_036_513, w_036_514, w_036_515, w_036_516, w_036_517, w_036_518, w_036_519, w_036_520, w_036_521, w_036_522, w_036_523, w_036_524, w_036_525, w_036_526, w_036_527, w_036_528, w_036_529, w_036_530, w_036_531, w_036_532, w_036_533, w_036_534, w_036_535, w_036_536, w_036_537, w_036_538, w_036_539, w_036_540, w_036_541, w_036_542, w_036_543, w_036_544, w_036_545, w_036_546, w_036_547, w_036_548, w_036_549, w_036_550, w_036_551, w_036_552, w_036_553, w_036_554, w_036_555, w_036_556, w_036_557, w_036_558, w_036_559, w_036_560, w_036_561, w_036_562, w_036_563, w_036_564, w_036_565, w_036_566, w_036_567, w_036_568, w_036_569, w_036_570, w_036_571, w_036_572, w_036_573, w_036_574, w_036_575, w_036_576, w_036_577, w_036_578, w_036_579, w_036_580, w_036_581, w_036_582, w_036_583, w_036_584, w_036_585, w_036_586, w_036_587, w_036_588, w_036_589, w_036_590, w_036_591, w_036_592, w_036_593, w_036_594, w_036_595, w_036_596, w_036_597, w_036_598, w_036_599, w_036_600, w_036_601, w_036_602, w_036_603, w_036_604, w_036_605, w_036_606, w_036_607, w_036_608, w_036_609, w_036_610, w_036_611, w_036_612, w_036_613, w_036_614, w_036_615, w_036_616, w_036_617, w_036_618, w_036_619, w_036_620, w_036_621, w_036_622, w_036_623, w_036_624, w_036_625, w_036_626, w_036_627, w_036_628, w_036_629, w_036_630, w_036_631, w_036_632, w_036_633, w_036_634, w_036_635, w_036_636, w_036_637, w_036_638, w_036_639, w_036_640, w_036_641, w_036_642, w_036_643, w_036_644, w_036_645, w_036_646, w_036_647, w_036_648, w_036_649, w_036_650, w_036_651, w_036_652, w_036_653, w_036_654, w_036_655, w_036_656, w_036_657, w_036_658, w_036_659, w_036_660, w_036_661, w_036_662, w_036_663, w_036_664, w_036_665, w_036_666, w_036_667, w_036_668, w_036_669, w_036_670, w_036_671, w_036_672, w_036_673, w_036_674, w_036_675, w_036_676, w_036_677, w_036_678, w_036_679, w_036_680, w_036_681, w_036_682, w_036_683, w_036_684, w_036_685, w_036_686, w_036_687, w_036_688, w_036_689, w_036_690, w_036_691, w_036_692, w_036_693, w_036_694, w_036_695, w_036_696, w_036_697, w_036_698, w_036_699, w_036_700, w_036_701, w_036_702, w_036_703, w_036_704, w_036_705, w_036_706, w_036_707, w_036_708, w_036_709, w_036_710, w_036_711, w_036_712;
  wire w_037_000, w_037_001, w_037_002, w_037_003, w_037_004, w_037_005, w_037_006, w_037_007, w_037_008, w_037_009, w_037_010, w_037_011, w_037_012, w_037_013, w_037_014, w_037_015, w_037_016, w_037_017, w_037_018, w_037_019, w_037_020, w_037_021, w_037_022, w_037_023, w_037_024, w_037_025, w_037_026, w_037_027, w_037_028, w_037_029, w_037_030, w_037_031, w_037_032, w_037_033, w_037_034, w_037_035, w_037_036, w_037_037, w_037_038, w_037_039, w_037_040, w_037_041, w_037_042, w_037_044, w_037_045, w_037_046, w_037_047, w_037_048, w_037_049, w_037_050, w_037_051, w_037_052, w_037_053, w_037_054, w_037_055, w_037_056, w_037_057, w_037_058, w_037_059, w_037_060, w_037_061, w_037_062, w_037_063, w_037_064, w_037_065, w_037_066, w_037_067, w_037_068, w_037_069, w_037_070, w_037_071, w_037_072, w_037_073, w_037_075, w_037_076, w_037_077, w_037_078, w_037_079, w_037_080, w_037_081, w_037_082, w_037_083, w_037_084, w_037_085, w_037_086, w_037_087, w_037_088, w_037_089, w_037_090, w_037_091, w_037_092, w_037_093, w_037_094, w_037_095, w_037_096, w_037_097, w_037_098, w_037_099, w_037_100, w_037_101, w_037_102, w_037_103, w_037_104, w_037_105, w_037_106, w_037_107, w_037_108, w_037_109, w_037_110, w_037_111, w_037_112, w_037_113, w_037_114, w_037_115, w_037_116, w_037_117, w_037_118, w_037_119, w_037_120, w_037_121, w_037_122, w_037_123, w_037_124, w_037_125, w_037_126, w_037_127, w_037_128, w_037_129, w_037_131, w_037_132, w_037_133, w_037_134, w_037_135, w_037_136, w_037_137, w_037_138, w_037_139, w_037_140, w_037_141, w_037_142, w_037_143, w_037_144, w_037_145, w_037_146, w_037_147, w_037_148, w_037_149, w_037_150, w_037_151, w_037_152, w_037_153, w_037_154, w_037_155, w_037_156, w_037_157, w_037_158, w_037_159, w_037_160, w_037_161, w_037_162, w_037_163, w_037_164, w_037_165, w_037_166, w_037_167, w_037_168, w_037_169, w_037_170, w_037_171, w_037_172, w_037_173, w_037_174, w_037_175, w_037_176, w_037_177, w_037_179, w_037_181, w_037_182, w_037_183, w_037_184, w_037_185, w_037_186, w_037_187, w_037_188, w_037_189, w_037_190, w_037_191, w_037_192, w_037_193, w_037_194, w_037_195, w_037_196, w_037_197, w_037_198, w_037_199, w_037_200, w_037_201, w_037_202, w_037_203, w_037_204, w_037_205, w_037_206, w_037_207, w_037_208, w_037_209, w_037_211, w_037_212, w_037_213, w_037_214, w_037_215, w_037_216, w_037_217, w_037_218, w_037_219, w_037_220, w_037_221, w_037_222, w_037_223, w_037_224, w_037_225, w_037_226, w_037_227, w_037_228, w_037_229, w_037_230, w_037_231, w_037_232, w_037_233, w_037_234, w_037_235, w_037_236, w_037_237, w_037_238, w_037_239, w_037_240, w_037_241, w_037_242, w_037_243, w_037_244, w_037_245, w_037_246, w_037_247, w_037_248, w_037_249, w_037_250, w_037_251, w_037_252, w_037_253, w_037_254, w_037_255, w_037_256, w_037_257, w_037_258, w_037_259, w_037_260, w_037_261, w_037_262, w_037_263, w_037_265, w_037_266, w_037_267, w_037_268, w_037_269, w_037_270, w_037_271, w_037_272, w_037_273, w_037_274, w_037_275, w_037_276, w_037_277, w_037_278, w_037_279, w_037_280, w_037_281, w_037_282, w_037_283, w_037_284, w_037_285, w_037_286, w_037_287, w_037_288, w_037_289, w_037_290, w_037_291, w_037_292, w_037_293, w_037_294, w_037_295, w_037_296, w_037_297, w_037_298, w_037_299, w_037_300, w_037_301, w_037_302, w_037_303, w_037_304, w_037_305, w_037_306, w_037_307, w_037_308, w_037_309, w_037_310, w_037_311, w_037_312, w_037_313, w_037_314, w_037_315, w_037_316, w_037_317, w_037_318, w_037_319, w_037_320, w_037_321, w_037_322, w_037_323, w_037_324, w_037_325, w_037_326, w_037_327, w_037_328, w_037_329, w_037_330, w_037_331, w_037_332, w_037_333, w_037_334, w_037_335, w_037_336, w_037_337, w_037_338, w_037_339, w_037_340, w_037_341, w_037_342, w_037_343, w_037_344, w_037_345, w_037_346, w_037_347, w_037_348, w_037_349, w_037_350, w_037_351, w_037_352, w_037_353, w_037_354, w_037_355, w_037_356, w_037_357, w_037_358, w_037_359, w_037_360, w_037_361, w_037_362, w_037_363, w_037_364, w_037_365, w_037_366, w_037_367, w_037_368, w_037_369, w_037_370, w_037_371, w_037_372, w_037_373, w_037_374, w_037_375, w_037_376, w_037_377, w_037_378, w_037_379, w_037_380, w_037_381, w_037_383, w_037_384, w_037_385, w_037_386, w_037_387, w_037_388, w_037_389, w_037_390, w_037_391, w_037_392, w_037_393, w_037_394, w_037_395, w_037_396, w_037_397, w_037_398, w_037_399, w_037_400, w_037_401, w_037_402, w_037_403, w_037_404, w_037_405, w_037_406, w_037_407, w_037_408, w_037_409, w_037_410, w_037_411, w_037_412, w_037_413, w_037_414, w_037_415, w_037_416, w_037_417, w_037_418, w_037_419, w_037_421, w_037_422, w_037_423, w_037_424, w_037_425, w_037_426, w_037_427, w_037_428, w_037_429, w_037_430, w_037_431, w_037_432, w_037_433, w_037_434, w_037_435, w_037_436, w_037_437, w_037_438, w_037_439, w_037_440, w_037_441, w_037_442, w_037_443, w_037_444, w_037_445, w_037_446, w_037_447, w_037_448, w_037_449, w_037_450, w_037_451, w_037_452, w_037_453, w_037_454, w_037_455, w_037_456, w_037_457, w_037_458, w_037_459, w_037_460, w_037_461, w_037_462, w_037_463, w_037_464, w_037_465, w_037_466, w_037_467, w_037_468, w_037_469, w_037_470, w_037_471, w_037_472, w_037_473, w_037_474, w_037_475, w_037_476, w_037_477, w_037_478, w_037_479, w_037_480, w_037_481, w_037_482, w_037_483, w_037_484, w_037_485, w_037_486, w_037_487, w_037_488, w_037_489, w_037_490, w_037_491, w_037_492, w_037_493, w_037_495, w_037_496, w_037_497, w_037_498, w_037_499, w_037_500, w_037_501, w_037_502, w_037_503, w_037_504, w_037_505, w_037_506, w_037_507, w_037_508, w_037_509, w_037_510, w_037_511, w_037_512, w_037_513, w_037_514, w_037_515, w_037_516, w_037_517, w_037_518, w_037_519, w_037_520, w_037_521, w_037_522, w_037_523, w_037_524, w_037_525, w_037_526, w_037_527, w_037_528, w_037_529, w_037_530, w_037_531, w_037_532, w_037_534, w_037_535, w_037_536, w_037_538, w_037_539, w_037_540, w_037_541, w_037_542, w_037_543, w_037_544, w_037_545, w_037_546, w_037_547, w_037_548, w_037_549, w_037_550, w_037_551, w_037_552, w_037_553, w_037_555, w_037_556, w_037_557, w_037_558, w_037_559, w_037_560, w_037_562, w_037_563, w_037_564, w_037_565, w_037_566, w_037_567, w_037_568, w_037_569, w_037_570, w_037_571, w_037_572, w_037_573, w_037_574, w_037_575, w_037_576, w_037_577, w_037_578, w_037_579, w_037_580, w_037_581, w_037_582, w_037_583, w_037_584, w_037_585, w_037_586, w_037_587, w_037_588, w_037_589, w_037_590, w_037_591, w_037_592, w_037_593, w_037_594, w_037_595, w_037_596, w_037_597, w_037_598, w_037_599, w_037_600, w_037_601, w_037_602, w_037_603, w_037_604, w_037_605, w_037_606, w_037_607, w_037_608, w_037_609, w_037_610, w_037_611, w_037_612, w_037_613, w_037_614, w_037_615, w_037_616, w_037_617, w_037_618, w_037_619, w_037_620, w_037_621, w_037_622, w_037_623, w_037_624, w_037_625, w_037_628, w_037_629, w_037_630, w_037_631, w_037_632, w_037_633, w_037_634, w_037_636, w_037_637, w_037_638, w_037_639, w_037_640, w_037_641, w_037_642, w_037_643, w_037_644, w_037_645, w_037_646, w_037_647, w_037_648, w_037_649, w_037_650, w_037_651, w_037_652, w_037_653, w_037_654, w_037_655, w_037_657, w_037_658, w_037_659, w_037_660, w_037_661, w_037_662, w_037_663, w_037_664, w_037_665, w_037_666, w_037_667, w_037_668, w_037_669, w_037_670, w_037_671, w_037_672, w_037_673, w_037_674, w_037_675, w_037_676, w_037_677, w_037_678, w_037_679, w_037_680, w_037_681, w_037_682, w_037_683, w_037_685, w_037_686, w_037_687, w_037_688, w_037_689, w_037_690, w_037_691, w_037_692, w_037_693, w_037_694, w_037_695, w_037_696, w_037_697, w_037_698, w_037_699, w_037_700, w_037_701, w_037_702, w_037_703, w_037_704, w_037_705, w_037_706, w_037_707, w_037_708, w_037_709, w_037_710, w_037_711, w_037_712, w_037_713, w_037_714, w_037_715, w_037_716, w_037_717, w_037_718, w_037_719, w_037_720, w_037_721, w_037_722, w_037_723, w_037_724, w_037_725, w_037_726, w_037_727, w_037_729, w_037_730, w_037_731, w_037_732, w_037_733, w_037_734, w_037_735, w_037_736, w_037_737, w_037_738, w_037_739, w_037_740, w_037_741, w_037_742, w_037_743, w_037_745, w_037_746, w_037_747, w_037_748, w_037_749, w_037_750, w_037_751, w_037_752, w_037_753, w_037_754, w_037_755, w_037_756, w_037_757, w_037_758, w_037_759, w_037_760, w_037_761, w_037_762, w_037_763, w_037_764, w_037_765, w_037_766, w_037_767, w_037_768, w_037_769, w_037_770, w_037_771, w_037_772, w_037_773, w_037_774, w_037_775, w_037_776, w_037_777, w_037_778, w_037_779, w_037_780, w_037_781, w_037_782, w_037_783, w_037_784, w_037_785, w_037_786, w_037_787, w_037_788, w_037_789, w_037_790, w_037_791, w_037_792, w_037_793, w_037_794, w_037_795, w_037_796, w_037_797, w_037_798, w_037_799, w_037_800, w_037_801, w_037_802, w_037_803, w_037_804, w_037_805, w_037_806, w_037_807, w_037_808, w_037_809, w_037_810, w_037_811, w_037_812, w_037_813, w_037_814, w_037_815, w_037_816, w_037_817, w_037_818, w_037_819, w_037_820, w_037_821, w_037_822, w_037_823, w_037_824, w_037_825, w_037_826, w_037_827, w_037_828, w_037_829, w_037_830, w_037_831, w_037_832, w_037_834, w_037_835, w_037_836, w_037_837, w_037_838, w_037_839, w_037_840, w_037_841, w_037_842, w_037_843, w_037_844, w_037_845, w_037_846, w_037_847, w_037_848, w_037_849, w_037_850, w_037_851, w_037_852, w_037_853, w_037_855, w_037_856, w_037_857, w_037_858, w_037_859, w_037_860, w_037_861, w_037_862, w_037_863, w_037_864, w_037_865, w_037_866, w_037_867, w_037_868, w_037_869, w_037_870, w_037_871, w_037_872, w_037_873, w_037_874, w_037_875, w_037_876, w_037_878, w_037_879, w_037_880, w_037_881, w_037_882, w_037_883, w_037_884, w_037_885, w_037_886, w_037_887, w_037_888, w_037_889, w_037_890, w_037_891, w_037_892, w_037_893, w_037_894, w_037_895, w_037_896, w_037_897, w_037_898, w_037_899, w_037_900, w_037_901, w_037_902, w_037_903, w_037_904, w_037_905, w_037_906, w_037_907, w_037_908, w_037_909, w_037_910, w_037_911, w_037_912, w_037_913, w_037_914, w_037_915, w_037_916, w_037_917, w_037_918, w_037_919, w_037_920, w_037_921, w_037_922, w_037_923, w_037_924, w_037_925, w_037_926, w_037_927, w_037_928, w_037_929, w_037_930, w_037_931, w_037_932, w_037_933, w_037_934, w_037_935, w_037_936, w_037_937, w_037_938, w_037_939, w_037_940, w_037_941, w_037_942, w_037_943, w_037_944, w_037_945, w_037_946, w_037_947, w_037_948, w_037_949, w_037_950, w_037_951, w_037_952, w_037_953, w_037_954, w_037_955, w_037_956, w_037_957, w_037_959, w_037_960, w_037_961, w_037_962, w_037_963, w_037_964, w_037_965, w_037_966, w_037_967, w_037_968, w_037_969, w_037_970, w_037_971, w_037_972, w_037_973, w_037_974, w_037_975, w_037_976, w_037_977, w_037_978, w_037_979, w_037_980, w_037_981, w_037_983, w_037_984, w_037_985, w_037_986, w_037_987, w_037_988, w_037_989, w_037_990, w_037_991, w_037_992, w_037_993, w_037_994, w_037_995, w_037_996, w_037_997, w_037_998, w_037_999, w_037_1000, w_037_1001, w_037_1002, w_037_1003, w_037_1004, w_037_1005, w_037_1006, w_037_1008, w_037_1009, w_037_1010, w_037_1011, w_037_1012, w_037_1013, w_037_1014, w_037_1015, w_037_1016, w_037_1017, w_037_1018, w_037_1019, w_037_1020, w_037_1021, w_037_1022, w_037_1023, w_037_1024, w_037_1025, w_037_1027, w_037_1028, w_037_1029, w_037_1030, w_037_1031, w_037_1032, w_037_1033, w_037_1034, w_037_1035, w_037_1036, w_037_1037, w_037_1038, w_037_1039, w_037_1040, w_037_1041, w_037_1042, w_037_1043, w_037_1044, w_037_1046, w_037_1048, w_037_1049, w_037_1050, w_037_1051, w_037_1052, w_037_1053, w_037_1054, w_037_1055, w_037_1056, w_037_1057, w_037_1058, w_037_1059, w_037_1060, w_037_1061, w_037_1062, w_037_1063, w_037_1064, w_037_1065, w_037_1066, w_037_1067, w_037_1068, w_037_1069, w_037_1070, w_037_1071, w_037_1072, w_037_1073, w_037_1074, w_037_1075, w_037_1076, w_037_1077, w_037_1078, w_037_1079, w_037_1081, w_037_1082, w_037_1083, w_037_1084, w_037_1086, w_037_1087, w_037_1088, w_037_1089, w_037_1090, w_037_1091, w_037_1092, w_037_1093, w_037_1094, w_037_1095, w_037_1096, w_037_1097, w_037_1098, w_037_1099, w_037_1100, w_037_1101, w_037_1102, w_037_1103, w_037_1104, w_037_1105, w_037_1106, w_037_1107, w_037_1108, w_037_1109, w_037_1110, w_037_1111, w_037_1112, w_037_1113, w_037_1114, w_037_1115, w_037_1116, w_037_1117, w_037_1118, w_037_1119, w_037_1120, w_037_1121, w_037_1122, w_037_1123, w_037_1124, w_037_1125, w_037_1126, w_037_1127, w_037_1128, w_037_1129, w_037_1130, w_037_1131, w_037_1132, w_037_1134, w_037_1135, w_037_1136, w_037_1137, w_037_1138, w_037_1139, w_037_1140, w_037_1141, w_037_1142, w_037_1143, w_037_1144, w_037_1145, w_037_1146, w_037_1147, w_037_1148, w_037_1149, w_037_1150, w_037_1151, w_037_1152, w_037_1153, w_037_1154, w_037_1155, w_037_1156, w_037_1157, w_037_1158, w_037_1160, w_037_1161, w_037_1162, w_037_1163, w_037_1164, w_037_1165, w_037_1166, w_037_1167, w_037_1168, w_037_1170, w_037_1171, w_037_1172, w_037_1173, w_037_1174, w_037_1175, w_037_1176, w_037_1177, w_037_1178, w_037_1179, w_037_1180, w_037_1181, w_037_1182, w_037_1183, w_037_1184, w_037_1185, w_037_1186, w_037_1187, w_037_1188, w_037_1189, w_037_1190, w_037_1191, w_037_1192, w_037_1193, w_037_1194, w_037_1195, w_037_1196, w_037_1197, w_037_1198, w_037_1199, w_037_1200, w_037_1201, w_037_1202, w_037_1203, w_037_1204, w_037_1205, w_037_1206, w_037_1207, w_037_1208, w_037_1209, w_037_1210, w_037_1211, w_037_1212, w_037_1213, w_037_1214, w_037_1215, w_037_1216, w_037_1217, w_037_1218, w_037_1219, w_037_1220, w_037_1221, w_037_1222, w_037_1223, w_037_1224, w_037_1225, w_037_1226, w_037_1228, w_037_1229, w_037_1230, w_037_1231, w_037_1232, w_037_1233, w_037_1234, w_037_1235, w_037_1236, w_037_1237, w_037_1238, w_037_1239, w_037_1240, w_037_1241, w_037_1242, w_037_1243, w_037_1244, w_037_1245, w_037_1246, w_037_1247, w_037_1248, w_037_1249, w_037_1250, w_037_1252, w_037_1253, w_037_1254, w_037_1255, w_037_1257, w_037_1258, w_037_1259, w_037_1260, w_037_1261, w_037_1262, w_037_1263, w_037_1264, w_037_1265, w_037_1266, w_037_1267, w_037_1268, w_037_1269, w_037_1270, w_037_1271, w_037_1272, w_037_1274, w_037_1275, w_037_1276, w_037_1277, w_037_1280, w_037_1281, w_037_1282, w_037_1283, w_037_1284, w_037_1285, w_037_1287, w_037_1288, w_037_1289, w_037_1290, w_037_1291, w_037_1292, w_037_1293, w_037_1294, w_037_1295, w_037_1296, w_037_1297, w_037_1298, w_037_1299, w_037_1300, w_037_1301, w_037_1302, w_037_1303, w_037_1304, w_037_1305, w_037_1306, w_037_1307, w_037_1308, w_037_1309, w_037_1310, w_037_1311, w_037_1312, w_037_1313, w_037_1314, w_037_1315, w_037_1316, w_037_1317, w_037_1318, w_037_1320, w_037_1321, w_037_1322, w_037_1323, w_037_1325, w_037_1326, w_037_1327, w_037_1328, w_037_1329, w_037_1330, w_037_1331, w_037_1332, w_037_1333, w_037_1334, w_037_1335, w_037_1336, w_037_1337, w_037_1338, w_037_1339, w_037_1340, w_037_1341, w_037_1342, w_037_1343, w_037_1344, w_037_1345, w_037_1346, w_037_1347, w_037_1348, w_037_1349, w_037_1350, w_037_1352, w_037_1353, w_037_1354, w_037_1355, w_037_1356, w_037_1357, w_037_1358, w_037_1359, w_037_1360, w_037_1361, w_037_1362, w_037_1363, w_037_1364, w_037_1366, w_037_1367, w_037_1368, w_037_1370, w_037_1371, w_037_1372, w_037_1373, w_037_1374, w_037_1375, w_037_1376, w_037_1377, w_037_1378, w_037_1379, w_037_1381, w_037_1383, w_037_1384, w_037_1385, w_037_1386, w_037_1387, w_037_1388, w_037_1389, w_037_1390, w_037_1391, w_037_1392, w_037_1393, w_037_1394, w_037_1395, w_037_1396, w_037_1397, w_037_1398, w_037_1399, w_037_1400, w_037_1401, w_037_1402, w_037_1403, w_037_1404, w_037_1406, w_037_1407, w_037_1408, w_037_1409, w_037_1410, w_037_1411, w_037_1412, w_037_1413, w_037_1414, w_037_1415, w_037_1416, w_037_1417, w_037_1418, w_037_1419, w_037_1420, w_037_1421, w_037_1422, w_037_1423, w_037_1424, w_037_1425, w_037_1426, w_037_1428, w_037_1429, w_037_1430, w_037_1431, w_037_1433, w_037_1435, w_037_1436, w_037_1437, w_037_1438, w_037_1439, w_037_1440, w_037_1441, w_037_1442, w_037_1443, w_037_1444, w_037_1445, w_037_1446, w_037_1447, w_037_1448, w_037_1449, w_037_1451, w_037_1452, w_037_1453, w_037_1454, w_037_1455, w_037_1457, w_037_1458, w_037_1459, w_037_1460, w_037_1461, w_037_1462, w_037_1463, w_037_1464, w_037_1465, w_037_1466, w_037_1467, w_037_1468, w_037_1469, w_037_1471, w_037_1472, w_037_1473, w_037_1474, w_037_1475, w_037_1476, w_037_1478, w_037_1479, w_037_1481, w_037_1482, w_037_1483, w_037_1484, w_037_1485, w_037_1486, w_037_1487, w_037_1488, w_037_1489, w_037_1490, w_037_1491, w_037_1492, w_037_1493, w_037_1494, w_037_1495, w_037_1496, w_037_1497, w_037_1498, w_037_1499, w_037_1500, w_037_1501, w_037_1502, w_037_1503, w_037_1504, w_037_1505, w_037_1506, w_037_1507, w_037_1508, w_037_1509, w_037_1510, w_037_1511, w_037_1512, w_037_1513, w_037_1514, w_037_1515, w_037_1516, w_037_1517, w_037_1518, w_037_1520, w_037_1521, w_037_1522, w_037_1523, w_037_1525, w_037_1526, w_037_1527, w_037_1528, w_037_1529, w_037_1530, w_037_1531, w_037_1532, w_037_1533, w_037_1534, w_037_1535, w_037_1536, w_037_1537, w_037_1538, w_037_1539, w_037_1540, w_037_1541, w_037_1542, w_037_1543, w_037_1544, w_037_1545, w_037_1546, w_037_1547, w_037_1548, w_037_1549, w_037_1551, w_037_1552, w_037_1553, w_037_1554, w_037_1555, w_037_1556, w_037_1557, w_037_1558, w_037_1559, w_037_1560, w_037_1561, w_037_1562, w_037_1563, w_037_1564, w_037_1565, w_037_1566, w_037_1567, w_037_1568, w_037_1569, w_037_1570, w_037_1571, w_037_1572, w_037_1573, w_037_1574, w_037_1575, w_037_1576, w_037_1577, w_037_1578, w_037_1579, w_037_1580, w_037_1581, w_037_1582, w_037_1583, w_037_1585, w_037_1586, w_037_1587, w_037_1588, w_037_1589, w_037_1590, w_037_1591, w_037_1592, w_037_1593, w_037_1594, w_037_1595, w_037_1596, w_037_1597, w_037_1598, w_037_1599, w_037_1600, w_037_1601, w_037_1602, w_037_1603, w_037_1604, w_037_1605, w_037_1607, w_037_1608, w_037_1609, w_037_1610, w_037_1611, w_037_1612, w_037_1613, w_037_1614, w_037_1615, w_037_1616, w_037_1617, w_037_1618, w_037_1619, w_037_1620, w_037_1621, w_037_1622, w_037_1623, w_037_1624, w_037_1625, w_037_1626, w_037_1627, w_037_1628, w_037_1629, w_037_1630, w_037_1631, w_037_1633, w_037_1634, w_037_1635, w_037_1636, w_037_1637, w_037_1638, w_037_1639, w_037_1640, w_037_1641, w_037_1642, w_037_1643, w_037_1644, w_037_1645, w_037_1646, w_037_1649, w_037_1650, w_037_1651, w_037_1652, w_037_1653, w_037_1654, w_037_1655, w_037_1656, w_037_1657, w_037_1658, w_037_1659, w_037_1661, w_037_1662, w_037_1663, w_037_1664, w_037_1665, w_037_1666, w_037_1667, w_037_1668, w_037_1669, w_037_1670, w_037_1671, w_037_1672, w_037_1673, w_037_1674, w_037_1675, w_037_1676, w_037_1677, w_037_1678, w_037_1679, w_037_1680, w_037_1681, w_037_1683, w_037_1684, w_037_1686, w_037_1687, w_037_1688, w_037_1689, w_037_1690, w_037_1691, w_037_1692, w_037_1694, w_037_1695, w_037_1696, w_037_1697, w_037_1698, w_037_1699, w_037_1700, w_037_1701, w_037_1703, w_037_1704, w_037_1705, w_037_1706, w_037_1707, w_037_1708, w_037_1709, w_037_1710, w_037_1711, w_037_1713, w_037_1714, w_037_1715, w_037_1716, w_037_1717, w_037_1718, w_037_1719, w_037_1720, w_037_1721, w_037_1722, w_037_1724, w_037_1725, w_037_1726, w_037_1727, w_037_1728, w_037_1730, w_037_1731, w_037_1732, w_037_1733, w_037_1734, w_037_1735, w_037_1736, w_037_1737, w_037_1738, w_037_1739, w_037_1740, w_037_1741, w_037_1742, w_037_1743, w_037_1744, w_037_1745, w_037_1746, w_037_1747, w_037_1748, w_037_1749, w_037_1750, w_037_1751, w_037_1752, w_037_1753, w_037_1754, w_037_1755, w_037_1756, w_037_1757, w_037_1758, w_037_1760, w_037_1761, w_037_1762, w_037_1763, w_037_1764, w_037_1767, w_037_1768, w_037_1769, w_037_1770, w_037_1771, w_037_1772, w_037_1773, w_037_1774, w_037_1775, w_037_1776, w_037_1777, w_037_1778, w_037_1779, w_037_1780, w_037_1781, w_037_1782, w_037_1783, w_037_1784, w_037_1785, w_037_1786, w_037_1787, w_037_1788, w_037_1789, w_037_1790, w_037_1791, w_037_1793, w_037_1794, w_037_1795, w_037_1797, w_037_1798, w_037_1799, w_037_1800, w_037_1801, w_037_1802, w_037_1803, w_037_1804, w_037_1805, w_037_1806, w_037_1807, w_037_1808, w_037_1809, w_037_1810, w_037_1811, w_037_1812, w_037_1813, w_037_1814, w_037_1815, w_037_1816, w_037_1817, w_037_1818, w_037_1819, w_037_1821, w_037_1822, w_037_1823, w_037_1824, w_037_1825, w_037_1827, w_037_1828, w_037_1829, w_037_1830, w_037_1831, w_037_1832, w_037_1833, w_037_1834, w_037_1835, w_037_1836, w_037_1837, w_037_1838, w_037_1839, w_037_1840, w_037_1841, w_037_1842, w_037_1844, w_037_1845, w_037_1846, w_037_1847, w_037_1848, w_037_1849, w_037_1850, w_037_1851, w_037_1852, w_037_1853, w_037_1854, w_037_1855, w_037_1856, w_037_1857, w_037_1859, w_037_1860, w_037_1861, w_037_1862, w_037_1863, w_037_1864, w_037_1865, w_037_1866, w_037_1867, w_037_1868, w_037_1869, w_037_1870, w_037_1871, w_037_1873, w_037_1874, w_037_1875, w_037_1876, w_037_1877, w_037_1878, w_037_1879, w_037_1880, w_037_1881, w_037_1883, w_037_1884, w_037_1885, w_037_1886, w_037_1887, w_037_1888, w_037_1889, w_037_1890, w_037_1892, w_037_1893, w_037_1894, w_037_1895, w_037_1896, w_037_1897, w_037_1898, w_037_1899, w_037_1900, w_037_1901, w_037_1902, w_037_1903, w_037_1904, w_037_1905, w_037_1908, w_037_1909, w_037_1910, w_037_1911, w_037_1912, w_037_1913, w_037_1914, w_037_1915, w_037_1916, w_037_1917, w_037_1918, w_037_1919, w_037_1920, w_037_1922, w_037_1924, w_037_1925, w_037_1926, w_037_1927, w_037_1928, w_037_1929, w_037_1930, w_037_1931, w_037_1932, w_037_1933, w_037_1935, w_037_1936, w_037_1937, w_037_1938, w_037_1939, w_037_1940, w_037_1941, w_037_1942, w_037_1943, w_037_1944, w_037_1945, w_037_1946, w_037_1947, w_037_1948, w_037_1949, w_037_1950, w_037_1951, w_037_1952, w_037_1953, w_037_1954, w_037_1955, w_037_1956, w_037_1957, w_037_1958, w_037_1959, w_037_1960, w_037_1961, w_037_1962, w_037_1963, w_037_1964, w_037_1965, w_037_1966, w_037_1967, w_037_1968, w_037_1969, w_037_1970, w_037_1971, w_037_1972, w_037_1973, w_037_1974, w_037_1975, w_037_1976, w_037_1977, w_037_1978, w_037_1979, w_037_1980, w_037_1981, w_037_1982, w_037_1983, w_037_1984, w_037_1986, w_037_1988, w_037_1989, w_037_1990, w_037_1991, w_037_1992, w_037_1993, w_037_1994, w_037_1995, w_037_1996, w_037_1997, w_037_1998, w_037_1999, w_037_2000, w_037_2001, w_037_2002, w_037_2003, w_037_2004, w_037_2005, w_037_2006, w_037_2007, w_037_2008, w_037_2009, w_037_2010, w_037_2011, w_037_2013, w_037_2014, w_037_2015, w_037_2016, w_037_2017, w_037_2018, w_037_2019, w_037_2020, w_037_2021, w_037_2022, w_037_2023, w_037_2024, w_037_2025, w_037_2026, w_037_2027, w_037_2028, w_037_2029, w_037_2030, w_037_2031, w_037_2032, w_037_2033, w_037_2034, w_037_2035, w_037_2036, w_037_2037, w_037_2038, w_037_2039, w_037_2040, w_037_2041, w_037_2042, w_037_2043, w_037_2044, w_037_2045, w_037_2046, w_037_2047, w_037_2048, w_037_2049, w_037_2051, w_037_2052, w_037_2053, w_037_2054, w_037_2055, w_037_2056, w_037_2057, w_037_2058, w_037_2059, w_037_2061, w_037_2062, w_037_2063, w_037_2064, w_037_2065, w_037_2066, w_037_2067, w_037_2069, w_037_2070, w_037_2071, w_037_2072, w_037_2073, w_037_2074, w_037_2075, w_037_2076, w_037_2077, w_037_2078, w_037_2079, w_037_2080, w_037_2081, w_037_2082, w_037_2084, w_037_2085, w_037_2086, w_037_2087, w_037_2089, w_037_2090, w_037_2091, w_037_2092, w_037_2093, w_037_2094, w_037_2095, w_037_2096, w_037_2097, w_037_2098, w_037_2099, w_037_2100, w_037_2101, w_037_2102, w_037_2103, w_037_2104, w_037_2105, w_037_2106, w_037_2107, w_037_2108, w_037_2109, w_037_2112, w_037_2113, w_037_2114, w_037_2115, w_037_2116, w_037_2117, w_037_2118, w_037_2119, w_037_2120, w_037_2121, w_037_2122, w_037_2123, w_037_2124, w_037_2125, w_037_2127, w_037_2128, w_037_2129, w_037_2130, w_037_2131, w_037_2132, w_037_2133, w_037_2134, w_037_2135, w_037_2136, w_037_2137, w_037_2138, w_037_2139, w_037_2140, w_037_2141, w_037_2142, w_037_2143, w_037_2144, w_037_2145, w_037_2146, w_037_2147, w_037_2148, w_037_2149, w_037_2150, w_037_2151, w_037_2152, w_037_2153, w_037_2154, w_037_2155, w_037_2157, w_037_2159, w_037_2160, w_037_2161, w_037_2162, w_037_2163, w_037_2164, w_037_2165, w_037_2166, w_037_2167, w_037_2168, w_037_2169, w_037_2170, w_037_2171, w_037_2172, w_037_2173, w_037_2174, w_037_2175, w_037_2176, w_037_2177, w_037_2178, w_037_2179, w_037_2180, w_037_2181, w_037_2182, w_037_2183, w_037_2184, w_037_2185, w_037_2186, w_037_2187, w_037_2188, w_037_2189, w_037_2190, w_037_2191, w_037_2192, w_037_2193, w_037_2194, w_037_2195, w_037_2196, w_037_2197, w_037_2198, w_037_2199, w_037_2200, w_037_2201, w_037_2202, w_037_2203, w_037_2204, w_037_2205, w_037_2206, w_037_2207, w_037_2208, w_037_2209, w_037_2210, w_037_2212, w_037_2213, w_037_2214, w_037_2215, w_037_2216, w_037_2217, w_037_2218, w_037_2219, w_037_2220, w_037_2221, w_037_2222, w_037_2223, w_037_2224, w_037_2225, w_037_2226, w_037_2227, w_037_2228, w_037_2229, w_037_2230, w_037_2231, w_037_2232, w_037_2233, w_037_2235, w_037_2236, w_037_2237, w_037_2238, w_037_2239, w_037_2240, w_037_2241, w_037_2242, w_037_2243, w_037_2244, w_037_2245, w_037_2246, w_037_2247, w_037_2248, w_037_2249, w_037_2250, w_037_2251, w_037_2252, w_037_2253, w_037_2254, w_037_2255, w_037_2256, w_037_2257, w_037_2258, w_037_2259, w_037_2260, w_037_2262, w_037_2263, w_037_2264, w_037_2266, w_037_2267, w_037_2268, w_037_2269, w_037_2270, w_037_2271, w_037_2272, w_037_2273, w_037_2274, w_037_2275, w_037_2276, w_037_2277, w_037_2278, w_037_2279, w_037_2280, w_037_2281, w_037_2282, w_037_2283, w_037_2284, w_037_2285;
  wire w_038_000, w_038_001, w_038_002, w_038_003, w_038_004, w_038_005, w_038_006, w_038_007, w_038_008, w_038_009, w_038_010, w_038_011, w_038_012, w_038_014, w_038_015, w_038_016, w_038_017, w_038_018, w_038_019, w_038_020, w_038_021, w_038_022, w_038_023, w_038_024, w_038_025, w_038_026, w_038_027, w_038_028, w_038_029, w_038_031, w_038_032, w_038_033, w_038_034, w_038_035, w_038_036, w_038_037, w_038_038, w_038_039, w_038_041, w_038_042, w_038_043, w_038_044, w_038_046, w_038_047, w_038_048, w_038_049, w_038_050, w_038_051, w_038_052, w_038_053, w_038_054, w_038_055, w_038_056, w_038_057, w_038_058, w_038_059, w_038_060, w_038_061, w_038_062, w_038_063, w_038_064, w_038_065, w_038_066, w_038_067, w_038_068, w_038_069, w_038_070, w_038_071, w_038_072, w_038_073, w_038_074, w_038_075, w_038_076, w_038_078, w_038_079, w_038_080, w_038_081, w_038_082, w_038_083, w_038_084, w_038_085, w_038_087, w_038_088, w_038_090, w_038_091, w_038_092, w_038_093, w_038_094, w_038_095, w_038_096, w_038_097, w_038_098, w_038_099, w_038_100, w_038_101, w_038_102, w_038_103, w_038_104, w_038_105, w_038_106, w_038_107, w_038_108, w_038_109, w_038_110, w_038_111, w_038_112, w_038_114, w_038_115, w_038_116, w_038_117, w_038_118, w_038_120, w_038_121, w_038_122, w_038_123, w_038_124, w_038_125, w_038_127, w_038_129, w_038_130, w_038_132, w_038_133, w_038_134, w_038_135, w_038_136, w_038_137, w_038_138, w_038_139, w_038_140, w_038_141, w_038_143, w_038_144, w_038_145, w_038_146, w_038_147, w_038_149, w_038_150, w_038_151, w_038_153, w_038_154, w_038_156, w_038_157, w_038_158, w_038_159, w_038_161, w_038_162, w_038_163, w_038_164, w_038_165, w_038_166, w_038_167, w_038_168, w_038_169, w_038_170, w_038_171, w_038_172, w_038_173, w_038_174, w_038_175, w_038_176, w_038_177, w_038_178, w_038_179, w_038_180, w_038_182, w_038_183, w_038_184, w_038_185, w_038_186, w_038_187, w_038_188, w_038_189, w_038_190, w_038_191, w_038_192, w_038_193, w_038_195, w_038_196, w_038_197, w_038_198, w_038_199, w_038_201, w_038_202, w_038_203, w_038_204, w_038_205, w_038_206, w_038_207, w_038_208, w_038_209, w_038_210, w_038_211, w_038_212, w_038_213, w_038_214, w_038_215, w_038_216, w_038_217, w_038_218, w_038_219, w_038_220, w_038_222, w_038_223, w_038_224, w_038_226, w_038_227, w_038_228, w_038_229, w_038_231, w_038_232, w_038_233, w_038_234, w_038_235, w_038_236, w_038_237, w_038_238, w_038_239, w_038_240, w_038_241, w_038_242, w_038_243, w_038_244, w_038_245, w_038_246, w_038_247, w_038_248, w_038_249, w_038_250, w_038_251, w_038_252, w_038_253, w_038_254, w_038_255, w_038_256, w_038_257, w_038_259, w_038_261, w_038_263, w_038_264, w_038_265, w_038_266, w_038_267, w_038_268, w_038_269, w_038_270, w_038_271, w_038_272, w_038_273, w_038_274, w_038_275, w_038_276, w_038_277, w_038_278, w_038_279, w_038_280, w_038_281, w_038_282, w_038_283, w_038_286, w_038_287, w_038_289, w_038_291, w_038_292, w_038_293, w_038_294, w_038_295, w_038_296, w_038_297, w_038_298, w_038_300, w_038_301, w_038_303, w_038_305, w_038_306, w_038_307, w_038_308, w_038_309, w_038_310, w_038_311, w_038_312, w_038_315, w_038_316, w_038_317, w_038_318, w_038_319, w_038_320, w_038_321, w_038_323, w_038_324, w_038_325, w_038_326, w_038_327, w_038_328, w_038_329, w_038_330, w_038_331, w_038_332, w_038_334, w_038_335, w_038_336, w_038_337, w_038_338, w_038_339, w_038_340, w_038_341, w_038_342, w_038_343, w_038_344, w_038_345, w_038_346, w_038_347, w_038_348, w_038_349, w_038_351, w_038_353, w_038_354, w_038_355, w_038_356, w_038_357, w_038_359, w_038_360, w_038_361, w_038_362, w_038_363, w_038_364, w_038_365, w_038_366, w_038_367, w_038_368, w_038_369, w_038_370, w_038_373, w_038_374, w_038_375, w_038_376, w_038_377, w_038_378, w_038_379, w_038_380, w_038_381, w_038_382, w_038_383, w_038_384, w_038_385, w_038_386, w_038_387, w_038_388, w_038_389, w_038_390, w_038_391, w_038_392, w_038_394, w_038_395, w_038_396, w_038_397, w_038_398, w_038_399, w_038_400, w_038_401, w_038_403, w_038_405, w_038_406, w_038_407, w_038_408, w_038_411, w_038_412, w_038_414, w_038_416, w_038_417, w_038_418, w_038_419, w_038_420, w_038_421, w_038_422, w_038_423, w_038_424, w_038_425, w_038_426, w_038_427, w_038_429, w_038_430, w_038_431, w_038_432, w_038_433, w_038_434, w_038_437, w_038_438, w_038_439, w_038_440, w_038_442, w_038_443, w_038_444, w_038_445, w_038_446, w_038_447, w_038_448, w_038_449, w_038_450, w_038_451, w_038_453, w_038_454, w_038_455, w_038_456, w_038_457, w_038_458, w_038_459, w_038_460, w_038_461, w_038_462, w_038_463, w_038_464, w_038_465, w_038_466, w_038_467, w_038_468, w_038_469, w_038_470, w_038_471, w_038_472, w_038_474, w_038_475, w_038_476, w_038_477, w_038_478, w_038_479, w_038_480, w_038_481, w_038_482, w_038_483, w_038_484, w_038_485, w_038_487, w_038_489, w_038_490, w_038_491, w_038_492, w_038_494, w_038_496, w_038_497, w_038_498, w_038_499, w_038_500, w_038_501, w_038_502, w_038_505, w_038_506, w_038_507, w_038_508, w_038_510, w_038_512, w_038_514, w_038_515, w_038_517, w_038_520, w_038_521, w_038_522, w_038_524, w_038_525, w_038_526, w_038_527, w_038_529, w_038_530, w_038_531, w_038_532, w_038_535, w_038_537, w_038_538, w_038_539, w_038_540, w_038_541, w_038_542, w_038_543, w_038_546, w_038_547, w_038_550, w_038_552, w_038_553, w_038_554, w_038_556, w_038_557, w_038_558, w_038_559, w_038_560, w_038_564, w_038_565, w_038_567, w_038_568, w_038_569, w_038_570, w_038_571, w_038_572, w_038_573, w_038_574, w_038_575, w_038_576, w_038_577, w_038_578, w_038_579, w_038_580, w_038_582, w_038_583, w_038_584, w_038_586, w_038_588, w_038_590, w_038_592, w_038_593, w_038_594, w_038_595, w_038_597, w_038_598, w_038_601, w_038_602, w_038_604, w_038_606, w_038_607, w_038_608, w_038_609, w_038_610, w_038_611, w_038_613, w_038_614, w_038_615, w_038_616, w_038_617, w_038_619, w_038_620, w_038_621, w_038_622, w_038_623, w_038_624, w_038_625, w_038_626, w_038_627, w_038_628, w_038_629, w_038_631, w_038_632, w_038_633, w_038_634, w_038_635, w_038_636, w_038_637, w_038_638, w_038_639, w_038_640, w_038_643, w_038_644, w_038_645, w_038_646, w_038_647, w_038_649, w_038_650, w_038_654, w_038_655, w_038_656, w_038_660, w_038_661, w_038_663, w_038_666, w_038_667, w_038_669, w_038_670, w_038_671, w_038_672, w_038_673, w_038_674, w_038_675, w_038_678, w_038_679, w_038_680, w_038_681, w_038_682, w_038_683, w_038_684, w_038_685, w_038_686, w_038_687, w_038_689, w_038_690, w_038_691, w_038_694, w_038_696, w_038_697, w_038_698, w_038_699, w_038_700, w_038_703, w_038_704, w_038_705, w_038_706, w_038_707, w_038_708, w_038_709, w_038_711, w_038_712, w_038_713, w_038_714, w_038_715, w_038_716, w_038_717, w_038_719, w_038_720, w_038_721, w_038_723, w_038_724, w_038_725, w_038_726, w_038_730, w_038_731, w_038_732, w_038_733, w_038_734, w_038_735, w_038_737, w_038_738, w_038_739, w_038_740, w_038_741, w_038_742, w_038_743, w_038_744, w_038_745, w_038_746, w_038_748, w_038_751, w_038_752, w_038_753, w_038_754, w_038_755, w_038_759, w_038_760, w_038_762, w_038_764, w_038_765, w_038_766, w_038_767, w_038_768, w_038_769, w_038_770, w_038_771, w_038_773, w_038_774, w_038_776, w_038_777, w_038_778, w_038_779, w_038_781, w_038_782, w_038_783, w_038_785, w_038_786, w_038_787, w_038_788, w_038_789, w_038_790, w_038_791, w_038_792, w_038_793, w_038_795, w_038_797, w_038_798, w_038_799, w_038_800, w_038_801, w_038_802, w_038_803, w_038_807, w_038_808, w_038_809, w_038_811, w_038_812, w_038_813, w_038_815, w_038_816, w_038_817, w_038_818, w_038_820, w_038_822, w_038_825, w_038_826, w_038_828, w_038_829, w_038_830, w_038_831, w_038_832, w_038_833, w_038_834, w_038_835, w_038_836, w_038_837, w_038_838, w_038_839, w_038_840, w_038_842, w_038_845, w_038_846, w_038_847, w_038_849, w_038_850, w_038_851, w_038_852, w_038_853, w_038_854, w_038_855, w_038_856, w_038_859, w_038_860, w_038_861, w_038_862, w_038_865, w_038_867, w_038_869, w_038_870, w_038_871, w_038_872, w_038_874, w_038_876, w_038_877, w_038_878, w_038_879, w_038_880, w_038_881, w_038_883, w_038_884, w_038_885, w_038_886, w_038_888, w_038_889, w_038_890, w_038_891, w_038_893, w_038_894, w_038_895, w_038_896, w_038_897, w_038_898, w_038_899, w_038_900, w_038_902, w_038_903, w_038_906, w_038_907, w_038_908, w_038_909, w_038_910, w_038_911, w_038_912, w_038_914, w_038_916, w_038_917, w_038_918, w_038_919, w_038_920, w_038_922, w_038_923, w_038_924, w_038_926, w_038_927, w_038_928, w_038_929, w_038_930, w_038_932, w_038_933, w_038_934, w_038_936, w_038_939, w_038_942, w_038_945, w_038_947, w_038_948, w_038_949, w_038_952, w_038_955, w_038_957, w_038_958, w_038_959, w_038_960, w_038_961, w_038_963, w_038_964, w_038_965, w_038_968, w_038_969, w_038_970, w_038_971, w_038_972, w_038_973, w_038_974, w_038_975, w_038_976, w_038_979, w_038_980, w_038_981, w_038_983, w_038_984, w_038_986, w_038_987, w_038_989, w_038_990, w_038_991, w_038_992, w_038_993, w_038_994, w_038_995, w_038_997, w_038_998, w_038_999, w_038_1000, w_038_1001, w_038_1003, w_038_1005, w_038_1006, w_038_1009, w_038_1010, w_038_1012, w_038_1013, w_038_1014, w_038_1015, w_038_1016, w_038_1017, w_038_1018, w_038_1019, w_038_1021, w_038_1022, w_038_1023, w_038_1024, w_038_1025, w_038_1026, w_038_1027, w_038_1028, w_038_1029, w_038_1031, w_038_1032, w_038_1033, w_038_1035, w_038_1036, w_038_1038, w_038_1039, w_038_1040, w_038_1041, w_038_1042, w_038_1043, w_038_1046, w_038_1047, w_038_1048, w_038_1049, w_038_1050, w_038_1051, w_038_1052, w_038_1054, w_038_1057, w_038_1058, w_038_1060, w_038_1061, w_038_1062, w_038_1063, w_038_1064, w_038_1065, w_038_1066, w_038_1067, w_038_1069, w_038_1072, w_038_1074, w_038_1075, w_038_1076, w_038_1078, w_038_1079, w_038_1080, w_038_1081, w_038_1082, w_038_1083, w_038_1084, w_038_1085, w_038_1087, w_038_1088, w_038_1089, w_038_1090, w_038_1091, w_038_1092, w_038_1094, w_038_1095, w_038_1098, w_038_1099, w_038_1100, w_038_1102, w_038_1103, w_038_1104, w_038_1105, w_038_1106, w_038_1107, w_038_1108, w_038_1109, w_038_1111, w_038_1112, w_038_1113, w_038_1114, w_038_1116, w_038_1117, w_038_1118, w_038_1119, w_038_1120, w_038_1121, w_038_1122, w_038_1123, w_038_1124, w_038_1126, w_038_1127, w_038_1128, w_038_1129, w_038_1130, w_038_1131, w_038_1132, w_038_1133, w_038_1134, w_038_1135, w_038_1136, w_038_1137, w_038_1138, w_038_1139, w_038_1140, w_038_1141, w_038_1142, w_038_1146, w_038_1147, w_038_1148, w_038_1149, w_038_1150, w_038_1151, w_038_1152, w_038_1155, w_038_1158, w_038_1159, w_038_1160, w_038_1161, w_038_1162, w_038_1163, w_038_1164, w_038_1165, w_038_1166, w_038_1167, w_038_1168, w_038_1169, w_038_1170, w_038_1172, w_038_1173, w_038_1174, w_038_1175, w_038_1176, w_038_1180, w_038_1181, w_038_1182, w_038_1184, w_038_1185, w_038_1186, w_038_1187, w_038_1188, w_038_1189, w_038_1192, w_038_1193, w_038_1194, w_038_1197, w_038_1198, w_038_1199, w_038_1202, w_038_1203, w_038_1204, w_038_1205, w_038_1206, w_038_1209, w_038_1210, w_038_1211, w_038_1212, w_038_1213, w_038_1214, w_038_1215, w_038_1218, w_038_1219, w_038_1220, w_038_1222, w_038_1224, w_038_1225, w_038_1228, w_038_1229, w_038_1231, w_038_1232, w_038_1234, w_038_1235, w_038_1236, w_038_1237, w_038_1241, w_038_1242, w_038_1243, w_038_1244, w_038_1247, w_038_1248, w_038_1250, w_038_1251, w_038_1252, w_038_1253, w_038_1254, w_038_1255, w_038_1257, w_038_1258, w_038_1259, w_038_1260, w_038_1261, w_038_1263, w_038_1264, w_038_1266, w_038_1267, w_038_1268, w_038_1269, w_038_1270, w_038_1273, w_038_1274, w_038_1275, w_038_1279, w_038_1281, w_038_1283, w_038_1284, w_038_1285, w_038_1287, w_038_1288, w_038_1289, w_038_1290, w_038_1291, w_038_1292, w_038_1293, w_038_1294, w_038_1295, w_038_1296, w_038_1297, w_038_1299, w_038_1300, w_038_1301, w_038_1302, w_038_1303, w_038_1304, w_038_1307, w_038_1311, w_038_1312, w_038_1313, w_038_1314, w_038_1317, w_038_1318, w_038_1319, w_038_1320, w_038_1321, w_038_1322, w_038_1323, w_038_1326, w_038_1327, w_038_1328, w_038_1330, w_038_1332, w_038_1333, w_038_1335, w_038_1336, w_038_1337, w_038_1338, w_038_1339, w_038_1341, w_038_1342, w_038_1343, w_038_1344, w_038_1345, w_038_1346, w_038_1347, w_038_1348, w_038_1349, w_038_1351, w_038_1352, w_038_1353, w_038_1354, w_038_1355, w_038_1356, w_038_1358, w_038_1359, w_038_1361, w_038_1362, w_038_1363, w_038_1364, w_038_1365, w_038_1367, w_038_1368, w_038_1369, w_038_1370, w_038_1371, w_038_1375, w_038_1378, w_038_1379, w_038_1380, w_038_1381, w_038_1382, w_038_1383, w_038_1384, w_038_1385, w_038_1386, w_038_1387, w_038_1390, w_038_1391, w_038_1393, w_038_1394, w_038_1396, w_038_1397, w_038_1400, w_038_1402, w_038_1403, w_038_1404, w_038_1406, w_038_1407, w_038_1408, w_038_1409, w_038_1410, w_038_1411, w_038_1412, w_038_1413, w_038_1415, w_038_1416, w_038_1417, w_038_1418, w_038_1419, w_038_1420, w_038_1424, w_038_1425, w_038_1426, w_038_1427, w_038_1428, w_038_1429, w_038_1430, w_038_1431, w_038_1432, w_038_1434, w_038_1436, w_038_1437, w_038_1438, w_038_1439, w_038_1440, w_038_1441, w_038_1442, w_038_1443, w_038_1445, w_038_1446, w_038_1448, w_038_1449, w_038_1450, w_038_1454, w_038_1456, w_038_1457, w_038_1458, w_038_1459, w_038_1460, w_038_1462, w_038_1463, w_038_1465, w_038_1468, w_038_1469, w_038_1470, w_038_1472, w_038_1473, w_038_1475, w_038_1477, w_038_1478, w_038_1480, w_038_1481, w_038_1483, w_038_1485, w_038_1486, w_038_1488, w_038_1489, w_038_1490, w_038_1491, w_038_1492, w_038_1493, w_038_1494, w_038_1495, w_038_1496, w_038_1497, w_038_1498, w_038_1499, w_038_1500, w_038_1501, w_038_1502, w_038_1503, w_038_1504, w_038_1506, w_038_1507, w_038_1508, w_038_1509, w_038_1510, w_038_1511, w_038_1512, w_038_1513, w_038_1515, w_038_1516, w_038_1517, w_038_1518, w_038_1519, w_038_1520, w_038_1523, w_038_1524, w_038_1525, w_038_1528, w_038_1529, w_038_1530, w_038_1532, w_038_1533, w_038_1536, w_038_1538, w_038_1539, w_038_1540, w_038_1541, w_038_1543, w_038_1548, w_038_1549, w_038_1550, w_038_1551, w_038_1552, w_038_1556, w_038_1557, w_038_1558, w_038_1559, w_038_1560, w_038_1562, w_038_1563, w_038_1564, w_038_1565, w_038_1566, w_038_1569, w_038_1570, w_038_1571, w_038_1573, w_038_1574, w_038_1576, w_038_1578, w_038_1579, w_038_1580, w_038_1581, w_038_1582, w_038_1583, w_038_1584, w_038_1589, w_038_1590, w_038_1591, w_038_1594, w_038_1595, w_038_1597, w_038_1598, w_038_1599, w_038_1600, w_038_1602, w_038_1603, w_038_1604, w_038_1605, w_038_1606, w_038_1608, w_038_1609, w_038_1610, w_038_1611, w_038_1613, w_038_1614, w_038_1616, w_038_1617, w_038_1618, w_038_1619, w_038_1621, w_038_1622, w_038_1623, w_038_1624, w_038_1626, w_038_1627, w_038_1628, w_038_1629, w_038_1630, w_038_1631, w_038_1632, w_038_1633, w_038_1634, w_038_1636, w_038_1638, w_038_1639, w_038_1641, w_038_1642, w_038_1647, w_038_1648, w_038_1649, w_038_1651, w_038_1654, w_038_1657, w_038_1658, w_038_1659, w_038_1660, w_038_1661, w_038_1662, w_038_1663, w_038_1664, w_038_1665, w_038_1666, w_038_1667, w_038_1668, w_038_1669, w_038_1670, w_038_1671, w_038_1673, w_038_1674, w_038_1675, w_038_1676, w_038_1679, w_038_1680, w_038_1681, w_038_1682, w_038_1683, w_038_1684, w_038_1685, w_038_1686, w_038_1687, w_038_1688, w_038_1690, w_038_1692, w_038_1693, w_038_1694, w_038_1695, w_038_1697, w_038_1698, w_038_1699, w_038_1700, w_038_1701, w_038_1703, w_038_1704, w_038_1705, w_038_1706, w_038_1707, w_038_1708, w_038_1709, w_038_1710, w_038_1711, w_038_1712, w_038_1713, w_038_1715, w_038_1716, w_038_1719, w_038_1720, w_038_1722, w_038_1724, w_038_1726, w_038_1727, w_038_1728, w_038_1729, w_038_1730, w_038_1734, w_038_1735, w_038_1736, w_038_1738, w_038_1739, w_038_1740, w_038_1741, w_038_1743, w_038_1744, w_038_1745, w_038_1746, w_038_1747, w_038_1748, w_038_1749, w_038_1751, w_038_1752, w_038_1754, w_038_1755, w_038_1756, w_038_1757, w_038_1758, w_038_1759, w_038_1762, w_038_1763, w_038_1765, w_038_1766, w_038_1767, w_038_1769, w_038_1770, w_038_1771, w_038_1772, w_038_1773, w_038_1774, w_038_1777, w_038_1780, w_038_1781, w_038_1782, w_038_1785, w_038_1787, w_038_1788, w_038_1789, w_038_1790, w_038_1791, w_038_1793, w_038_1795, w_038_1796, w_038_1797, w_038_1798, w_038_1799, w_038_1800, w_038_1801, w_038_1802, w_038_1803, w_038_1804, w_038_1806, w_038_1807, w_038_1809, w_038_1810, w_038_1812, w_038_1813, w_038_1815, w_038_1817, w_038_1818, w_038_1820, w_038_1821, w_038_1823, w_038_1825, w_038_1826, w_038_1828, w_038_1829, w_038_1830, w_038_1831, w_038_1832, w_038_1833, w_038_1834, w_038_1835, w_038_1836, w_038_1837, w_038_1840, w_038_1843, w_038_1844, w_038_1845, w_038_1848, w_038_1849, w_038_1850, w_038_1852, w_038_1853, w_038_1854, w_038_1855, w_038_1856, w_038_1857, w_038_1858, w_038_1860, w_038_1861, w_038_1862, w_038_1863, w_038_1864, w_038_1865, w_038_1866, w_038_1867, w_038_1868, w_038_1869, w_038_1870, w_038_1871, w_038_1872, w_038_1873, w_038_1874, w_038_1875, w_038_1876, w_038_1877, w_038_1878, w_038_1879, w_038_1880, w_038_1882, w_038_1883, w_038_1884, w_038_1885, w_038_1887, w_038_1889, w_038_1890, w_038_1891, w_038_1892, w_038_1894, w_038_1895, w_038_1896, w_038_1897, w_038_1899, w_038_1900, w_038_1902, w_038_1903, w_038_1906, w_038_1908, w_038_1910, w_038_1912, w_038_1914, w_038_1915, w_038_1916, w_038_1917, w_038_1918, w_038_1922, w_038_1924, w_038_1925, w_038_1927, w_038_1928, w_038_1929, w_038_1931, w_038_1933, w_038_1935, w_038_1936, w_038_1937, w_038_1938, w_038_1939, w_038_1940, w_038_1941, w_038_1942, w_038_1943, w_038_1945, w_038_1946, w_038_1947, w_038_1948, w_038_1949, w_038_1950, w_038_1952, w_038_1953, w_038_1954, w_038_1955, w_038_1956, w_038_1957, w_038_1958, w_038_1959, w_038_1960, w_038_1961, w_038_1963, w_038_1964, w_038_1965, w_038_1966, w_038_1967, w_038_1970, w_038_1971, w_038_1972, w_038_1973, w_038_1974, w_038_1976, w_038_1977, w_038_1979, w_038_1980, w_038_1981, w_038_1982, w_038_1983, w_038_1985, w_038_1986, w_038_1987, w_038_1988, w_038_1990, w_038_1991, w_038_1992, w_038_1993, w_038_1994, w_038_1995, w_038_1996, w_038_1998, w_038_1999, w_038_2000, w_038_2001, w_038_2003, w_038_2004, w_038_2005, w_038_2006, w_038_2007, w_038_2008, w_038_2009, w_038_2010, w_038_2011, w_038_2012, w_038_2014, w_038_2016, w_038_2020, w_038_2021, w_038_2022, w_038_2023, w_038_2024, w_038_2025, w_038_2027, w_038_2028, w_038_2029, w_038_2030, w_038_2031, w_038_2035, w_038_2036, w_038_2037, w_038_2039, w_038_2040, w_038_2042, w_038_2043, w_038_2047, w_038_2048, w_038_2050, w_038_2051, w_038_2052, w_038_2053, w_038_2054, w_038_2055, w_038_2056, w_038_2057, w_038_2058, w_038_2059, w_038_2060, w_038_2061, w_038_2063, w_038_2064, w_038_2066, w_038_2067, w_038_2069, w_038_2070, w_038_2071, w_038_2072, w_038_2074, w_038_2075, w_038_2078, w_038_2079, w_038_2080, w_038_2081, w_038_2082, w_038_2086, w_038_2088, w_038_2089, w_038_2090, w_038_2092, w_038_2094, w_038_2095, w_038_2096, w_038_2097, w_038_2098, w_038_2100, w_038_2101, w_038_2102, w_038_2105, w_038_2107, w_038_2108, w_038_2109, w_038_2110, w_038_2111, w_038_2112, w_038_2114, w_038_2116, w_038_2117, w_038_2118, w_038_2119, w_038_2120, w_038_2122, w_038_2123, w_038_2124, w_038_2125, w_038_2126, w_038_2127, w_038_2129, w_038_2130, w_038_2132, w_038_2133, w_038_2134, w_038_2136, w_038_2138, w_038_2139, w_038_2140, w_038_2141, w_038_2143, w_038_2144, w_038_2146, w_038_2147, w_038_2148, w_038_2149, w_038_2151, w_038_2152, w_038_2153, w_038_2156, w_038_2157, w_038_2159, w_038_2160, w_038_2162, w_038_2163, w_038_2164, w_038_2165, w_038_2166, w_038_2167, w_038_2168, w_038_2169, w_038_2170, w_038_2172, w_038_2173, w_038_2174, w_038_2175, w_038_2178, w_038_2179, w_038_2180, w_038_2181, w_038_2182, w_038_2183, w_038_2185, w_038_2186, w_038_2191, w_038_2192, w_038_2194, w_038_2195, w_038_2196, w_038_2200, w_038_2201, w_038_2202, w_038_2203, w_038_2204, w_038_2205, w_038_2206, w_038_2207, w_038_2208, w_038_2209, w_038_2210, w_038_2211, w_038_2212, w_038_2215, w_038_2216, w_038_2217, w_038_2220, w_038_2221, w_038_2222, w_038_2223, w_038_2224, w_038_2226, w_038_2227, w_038_2229, w_038_2230, w_038_2231, w_038_2232, w_038_2233, w_038_2235, w_038_2238, w_038_2239, w_038_2240, w_038_2242, w_038_2244, w_038_2245, w_038_2246, w_038_2247, w_038_2248, w_038_2249, w_038_2251, w_038_2252, w_038_2253, w_038_2254, w_038_2255, w_038_2256, w_038_2257, w_038_2259, w_038_2260, w_038_2261, w_038_2263, w_038_2264, w_038_2265, w_038_2266, w_038_2267, w_038_2271, w_038_2272, w_038_2274, w_038_2276, w_038_2277, w_038_2278, w_038_2279, w_038_2280, w_038_2282, w_038_2283, w_038_2284, w_038_2285, w_038_2287, w_038_2288, w_038_2289, w_038_2291, w_038_2292, w_038_2293, w_038_2295, w_038_2296, w_038_2297, w_038_2298, w_038_2301, w_038_2302, w_038_2304, w_038_2305, w_038_2308, w_038_2310, w_038_2311, w_038_2312, w_038_2313, w_038_2314, w_038_2315, w_038_2317, w_038_2318, w_038_2320, w_038_2321, w_038_2322, w_038_2323, w_038_2324, w_038_2325, w_038_2326, w_038_2328, w_038_2330, w_038_2331, w_038_2332, w_038_2333, w_038_2334, w_038_2335, w_038_2336, w_038_2337, w_038_2338, w_038_2339, w_038_2340, w_038_2341, w_038_2342, w_038_2343, w_038_2344, w_038_2346, w_038_2347, w_038_2348, w_038_2351, w_038_2352, w_038_2353, w_038_2354, w_038_2355, w_038_2356, w_038_2357, w_038_2359, w_038_2360, w_038_2361, w_038_2362, w_038_2363, w_038_2366, w_038_2367, w_038_2370, w_038_2371, w_038_2372, w_038_2374, w_038_2377, w_038_2379, w_038_2383, w_038_2384, w_038_2385, w_038_2386, w_038_2387, w_038_2388, w_038_2389, w_038_2390, w_038_2391, w_038_2393, w_038_2394, w_038_2396, w_038_2397, w_038_2398, w_038_2399, w_038_2400, w_038_2401, w_038_2403, w_038_2404, w_038_2406, w_038_2407, w_038_2408, w_038_2409, w_038_2410, w_038_2413, w_038_2414, w_038_2418, w_038_2419, w_038_2420, w_038_2422, w_038_2423, w_038_2424, w_038_2425, w_038_2426, w_038_2430, w_038_2431, w_038_2432, w_038_2435, w_038_2436, w_038_2437, w_038_2438, w_038_2439, w_038_2441, w_038_2442, w_038_2443, w_038_2444, w_038_2446, w_038_2447, w_038_2448, w_038_2449, w_038_2450, w_038_2451, w_038_2452, w_038_2453, w_038_2455, w_038_2457, w_038_2459, w_038_2460, w_038_2461, w_038_2462, w_038_2463, w_038_2464, w_038_2465, w_038_2466, w_038_2467, w_038_2468, w_038_2469, w_038_2471, w_038_2474, w_038_2475, w_038_2477, w_038_2478, w_038_2479, w_038_2481, w_038_2482, w_038_2484, w_038_2485, w_038_2486, w_038_2487, w_038_2488, w_038_2489, w_038_2490, w_038_2491, w_038_2492, w_038_2493, w_038_2494, w_038_2495, w_038_2496, w_038_2497, w_038_2498, w_038_2499, w_038_2501, w_038_2502, w_038_2503, w_038_2504, w_038_2505, w_038_2507, w_038_2508, w_038_2509, w_038_2510, w_038_2511, w_038_2512, w_038_2513, w_038_2515, w_038_2517, w_038_2518, w_038_2519, w_038_2521, w_038_2524, w_038_2526, w_038_2527, w_038_2528, w_038_2530, w_038_2531, w_038_2532, w_038_2533, w_038_2534, w_038_2535, w_038_2536, w_038_2537, w_038_2538, w_038_2540, w_038_2541, w_038_2542, w_038_2543, w_038_2544, w_038_2545, w_038_2546, w_038_2547, w_038_2548, w_038_2549, w_038_2550, w_038_2551, w_038_2553, w_038_2554, w_038_2555, w_038_2557, w_038_2558, w_038_2559, w_038_2560, w_038_2561, w_038_2562, w_038_2565, w_038_2566, w_038_2567, w_038_2568, w_038_2570, w_038_2572, w_038_2573, w_038_2574, w_038_2577, w_038_2579, w_038_2582, w_038_2583, w_038_2584, w_038_2585, w_038_2586, w_038_2587, w_038_2588, w_038_2590, w_038_2591, w_038_2592, w_038_2593, w_038_2594, w_038_2596, w_038_2597, w_038_2598, w_038_2600, w_038_2601, w_038_2602, w_038_2603, w_038_2604, w_038_2605, w_038_2608, w_038_2609, w_038_2613, w_038_2614, w_038_2616, w_038_2617, w_038_2618, w_038_2619, w_038_2620, w_038_2621, w_038_2622, w_038_2623, w_038_2624, w_038_2626, w_038_2627, w_038_2628, w_038_2629, w_038_2630, w_038_2631, w_038_2632, w_038_2633, w_038_2636, w_038_2638, w_038_2642, w_038_2643, w_038_2645, w_038_2646, w_038_2647, w_038_2648, w_038_2649, w_038_2651, w_038_2652, w_038_2653, w_038_2654, w_038_2655, w_038_2656, w_038_2657, w_038_2658, w_038_2659, w_038_2660, w_038_2661, w_038_2662, w_038_2663, w_038_2664, w_038_2665, w_038_2667, w_038_2668, w_038_2669, w_038_2670, w_038_2671, w_038_2672, w_038_2673, w_038_2674, w_038_2675, w_038_2677, w_038_2678, w_038_2679, w_038_2681, w_038_2683, w_038_2684, w_038_2685, w_038_2687, w_038_2689, w_038_2692, w_038_2693, w_038_2695, w_038_2696, w_038_2698, w_038_2699, w_038_2701, w_038_2702, w_038_2703, w_038_2704, w_038_2705, w_038_2706, w_038_2708, w_038_2709, w_038_2711, w_038_2712, w_038_2713, w_038_2714, w_038_2715, w_038_2717, w_038_2718, w_038_2719, w_038_2720, w_038_2722, w_038_2723, w_038_2724, w_038_2727, w_038_2729, w_038_2730, w_038_2733, w_038_2734, w_038_2736, w_038_2737, w_038_2738, w_038_2740, w_038_2741, w_038_2742, w_038_2744, w_038_2745, w_038_2746, w_038_2747, w_038_2749, w_038_2750, w_038_2752, w_038_2753, w_038_2754, w_038_2755, w_038_2757, w_038_2758, w_038_2759, w_038_2760, w_038_2761, w_038_2763, w_038_2765, w_038_2766, w_038_2768, w_038_2769, w_038_2771, w_038_2773, w_038_2774, w_038_2775, w_038_2776, w_038_2778, w_038_2779, w_038_2780, w_038_2781, w_038_2785, w_038_2786, w_038_2787, w_038_2789, w_038_2790, w_038_2791, w_038_2792, w_038_2793, w_038_2794, w_038_2796, w_038_2797, w_038_2798, w_038_2799, w_038_2802, w_038_2804, w_038_2805, w_038_2806, w_038_2810, w_038_2812, w_038_2813, w_038_2816, w_038_2817, w_038_2818, w_038_2819, w_038_2820, w_038_2821, w_038_2822, w_038_2823, w_038_2824, w_038_2825, w_038_2826, w_038_2829, w_038_2830, w_038_2831, w_038_2833, w_038_2834, w_038_2835, w_038_2836, w_038_2837, w_038_2838, w_038_2839, w_038_2840, w_038_2841, w_038_2842, w_038_2843, w_038_2844, w_038_2845, w_038_2846, w_038_2847, w_038_2848, w_038_2850, w_038_2851, w_038_2852, w_038_2853, w_038_2854, w_038_2855, w_038_2857, w_038_2858, w_038_2859, w_038_2860, w_038_2864, w_038_2865, w_038_2868, w_038_2869, w_038_2870, w_038_2871, w_038_2875, w_038_2876, w_038_2877, w_038_2879, w_038_2880, w_038_2881, w_038_2882, w_038_2884, w_038_2886, w_038_2887, w_038_2888, w_038_2889, w_038_2890, w_038_2891, w_038_2892, w_038_2893, w_038_2894, w_038_2895, w_038_2896, w_038_2897, w_038_2899, w_038_2901, w_038_2902, w_038_2903, w_038_2904, w_038_2905, w_038_2906, w_038_2907, w_038_2908, w_038_2909, w_038_2910, w_038_2913, w_038_2914, w_038_2915, w_038_2916, w_038_2918, w_038_2919, w_038_2921, w_038_2922, w_038_2924, w_038_2925, w_038_2926, w_038_2927, w_038_2928, w_038_2930, w_038_2932, w_038_2933, w_038_2934, w_038_2935, w_038_2936, w_038_2937, w_038_2939, w_038_2940, w_038_2941, w_038_2942, w_038_2943, w_038_2945, w_038_2947, w_038_2948, w_038_2949, w_038_2950, w_038_2951, w_038_2952, w_038_2953, w_038_2955, w_038_2956, w_038_2957, w_038_2958, w_038_2959, w_038_2960, w_038_2961, w_038_2963, w_038_2964, w_038_2965, w_038_2966, w_038_2968, w_038_2969, w_038_2970, w_038_2973, w_038_2974, w_038_2975, w_038_2978, w_038_2980, w_038_2981, w_038_2984, w_038_2985, w_038_2987, w_038_2988, w_038_2989, w_038_2990, w_038_2992, w_038_2994, w_038_2995, w_038_2996, w_038_2997, w_038_2999, w_038_3000, w_038_3002, w_038_3004, w_038_3005, w_038_3006, w_038_3007, w_038_3008, w_038_3010, w_038_3011, w_038_3012, w_038_3013, w_038_3014, w_038_3015, w_038_3017, w_038_3018, w_038_3019, w_038_3020, w_038_3021, w_038_3023, w_038_3025, w_038_3026, w_038_3027, w_038_3029, w_038_3030, w_038_3032, w_038_3033, w_038_3034, w_038_3035, w_038_3037, w_038_3038, w_038_3039, w_038_3040, w_038_3041, w_038_3042, w_038_3044, w_038_3045, w_038_3047, w_038_3048, w_038_3050, w_038_3051, w_038_3052, w_038_3053, w_038_3055, w_038_3056, w_038_3057, w_038_3058, w_038_3059, w_038_3060, w_038_3062, w_038_3063, w_038_3065, w_038_3066, w_038_3068, w_038_3069, w_038_3072, w_038_3073, w_038_3074, w_038_3075, w_038_3077, w_038_3078, w_038_3080, w_038_3081, w_038_3084, w_038_3085, w_038_3087, w_038_3088, w_038_3089, w_038_3090, w_038_3091, w_038_3092, w_038_3094, w_038_3095, w_038_3096, w_038_3097, w_038_3099, w_038_3100, w_038_3101, w_038_3102, w_038_3104, w_038_3105, w_038_3106, w_038_3107, w_038_3108, w_038_3109, w_038_3110, w_038_3111, w_038_3112, w_038_3113, w_038_3114, w_038_3115, w_038_3116, w_038_3117, w_038_3118, w_038_3119, w_038_3120, w_038_3121, w_038_3123, w_038_3124, w_038_3125, w_038_3126, w_038_3128, w_038_3130, w_038_3131, w_038_3132, w_038_3134, w_038_3135, w_038_3136, w_038_3137, w_038_3138, w_038_3139, w_038_3140, w_038_3142, w_038_3143, w_038_3146, w_038_3147, w_038_3149, w_038_3150, w_038_3153, w_038_3154, w_038_3155, w_038_3156, w_038_3159, w_038_3160, w_038_3162, w_038_3163, w_038_3165, w_038_3166, w_038_3167, w_038_3169, w_038_3172, w_038_3173, w_038_3174, w_038_3175, w_038_3176, w_038_3178, w_038_3179, w_038_3181, w_038_3183, w_038_3184, w_038_3186, w_038_3187, w_038_3188, w_038_3190, w_038_3191, w_038_3192, w_038_3194, w_038_3195, w_038_3197, w_038_3200, w_038_3201, w_038_3202, w_038_3203, w_038_3204, w_038_3205, w_038_3206, w_038_3208, w_038_3209, w_038_3211, w_038_3213, w_038_3216, w_038_3217, w_038_3218, w_038_3220, w_038_3221, w_038_3223, w_038_3224, w_038_3225, w_038_3227, w_038_3228, w_038_3230, w_038_3231, w_038_3233, w_038_3235, w_038_3236, w_038_3237, w_038_3240, w_038_3241, w_038_3243, w_038_3244, w_038_3245, w_038_3246, w_038_3247, w_038_3248, w_038_3249, w_038_3251, w_038_3252, w_038_3253, w_038_3254, w_038_3255, w_038_3256, w_038_3257, w_038_3259, w_038_3261, w_038_3262, w_038_3265, w_038_3267, w_038_3269, w_038_3271, w_038_3272, w_038_3273, w_038_3275, w_038_3276, w_038_3277, w_038_3278, w_038_3279, w_038_3280, w_038_3282, w_038_3283, w_038_3284, w_038_3286, w_038_3287, w_038_3288, w_038_3289, w_038_3290, w_038_3291, w_038_3292, w_038_3293, w_038_3294, w_038_3295, w_038_3296, w_038_3297, w_038_3298, w_038_3299, w_038_3300, w_038_3301, w_038_3303, w_038_3307, w_038_3309, w_038_3310, w_038_3311, w_038_3312, w_038_3314, w_038_3315, w_038_3316, w_038_3317, w_038_3318, w_038_3319, w_038_3320, w_038_3321, w_038_3322, w_038_3326, w_038_3328, w_038_3329, w_038_3330, w_038_3331, w_038_3334, w_038_3335, w_038_3336, w_038_3337, w_038_3339, w_038_3340, w_038_3344, w_038_3346, w_038_3347, w_038_3348, w_038_3350, w_038_3351, w_038_3352, w_038_3353, w_038_3354, w_038_3356, w_038_3357, w_038_3359, w_038_3364, w_038_3365, w_038_3366, w_038_3367, w_038_3369, w_038_3371, w_038_3373, w_038_3376, w_038_3377, w_038_3379, w_038_3380, w_038_3382, w_038_3384, w_038_3386, w_038_3387, w_038_3388, w_038_3390, w_038_3391, w_038_3392, w_038_3393, w_038_3395, w_038_3396, w_038_3397, w_038_3398, w_038_3399, w_038_3401, w_038_3402, w_038_3403, w_038_3407, w_038_3409, w_038_3410, w_038_3411, w_038_3413, w_038_3414, w_038_3415, w_038_3416, w_038_3417, w_038_3418, w_038_3419, w_038_3420, w_038_3421, w_038_3422, w_038_3423, w_038_3424, w_038_3425, w_038_3426, w_038_3427, w_038_3428, w_038_3431, w_038_3432, w_038_3434, w_038_3435, w_038_3437, w_038_3438, w_038_3440, w_038_3441, w_038_3442, w_038_3443, w_038_3444, w_038_3445, w_038_3446, w_038_3447, w_038_3449, w_038_3450, w_038_3452, w_038_3453, w_038_3455, w_038_3456, w_038_3457, w_038_3458, w_038_3459, w_038_3460, w_038_3461, w_038_3462, w_038_3463, w_038_3466, w_038_3467, w_038_3469, w_038_3470, w_038_3471, w_038_3473, w_038_3475, w_038_3476, w_038_3477, w_038_3478, w_038_3479, w_038_3480, w_038_3481, w_038_3484, w_038_3485, w_038_3486, w_038_3487, w_038_3488, w_038_3489, w_038_3492, w_038_3493, w_038_3495, w_038_3497, w_038_3498, w_038_3500, w_038_3503, w_038_3504, w_038_3505, w_038_3508, w_038_3510, w_038_3512, w_038_3514, w_038_3515, w_038_3516, w_038_3517, w_038_3519, w_038_3521, w_038_3522, w_038_3523, w_038_3524, w_038_3525, w_038_3526, w_038_3527, w_038_3528, w_038_3529, w_038_3531, w_038_3533, w_038_3534, w_038_3535, w_038_3538, w_038_3540, w_038_3541, w_038_3542, w_038_3544, w_038_3545, w_038_3546, w_038_3547, w_038_3548, w_038_3551, w_038_3552, w_038_3554, w_038_3555, w_038_3556, w_038_3557, w_038_3558, w_038_3559, w_038_3560, w_038_3561, w_038_3562, w_038_3563, w_038_3564, w_038_3566, w_038_3567, w_038_3568, w_038_3569, w_038_3570, w_038_3571, w_038_3576, w_038_3577, w_038_3578, w_038_3579, w_038_3581, w_038_3582, w_038_3583, w_038_3584, w_038_3585, w_038_3586, w_038_3587, w_038_3590, w_038_3592, w_038_3593, w_038_3596, w_038_3598, w_038_3599, w_038_3600, w_038_3601, w_038_3602, w_038_3603, w_038_3604, w_038_3606, w_038_3607, w_038_3608, w_038_3609, w_038_3610, w_038_3611, w_038_3612, w_038_3613, w_038_3617, w_038_3618, w_038_3619, w_038_3620, w_038_3622, w_038_3623, w_038_3626, w_038_3627, w_038_3628, w_038_3631, w_038_3632, w_038_3634, w_038_3635, w_038_3636, w_038_3638, w_038_3640, w_038_3641, w_038_3642, w_038_3644, w_038_3646, w_038_3648, w_038_3649, w_038_3651, w_038_3652, w_038_3653, w_038_3654, w_038_3656, w_038_3658, w_038_3659, w_038_3661, w_038_3662, w_038_3663, w_038_3667, w_038_3668, w_038_3669, w_038_3670, w_038_3671, w_038_3672, w_038_3673, w_038_3674, w_038_3675, w_038_3678, w_038_3680, w_038_3681, w_038_3683, w_038_3684, w_038_3685, w_038_3688, w_038_3689, w_038_3690, w_038_3691, w_038_3692, w_038_3694, w_038_3695, w_038_3696, w_038_3697, w_038_3698, w_038_3699, w_038_3700, w_038_3701, w_038_3702, w_038_3703, w_038_3706, w_038_3708, w_038_3709, w_038_3712, w_038_3713, w_038_3714, w_038_3716, w_038_3717, w_038_3718, w_038_3720, w_038_3721, w_038_3722, w_038_3723, w_038_3724, w_038_3725, w_038_3726, w_038_3727, w_038_3728, w_038_3730, w_038_3731, w_038_3732, w_038_3734, w_038_3736, w_038_3738, w_038_3740, w_038_3741, w_038_3742, w_038_3743, w_038_3745, w_038_3746, w_038_3747, w_038_3748, w_038_3750, w_038_3751, w_038_3752, w_038_3754, w_038_3755, w_038_3756, w_038_3757, w_038_3758, w_038_3759, w_038_3761, w_038_3766, w_038_3769, w_038_3770, w_038_3772, w_038_3774, w_038_3775, w_038_3777, w_038_3778, w_038_3779, w_038_3780, w_038_3782, w_038_3783, w_038_3784, w_038_3785, w_038_3786, w_038_3787, w_038_3788, w_038_3790, w_038_3791, w_038_3792, w_038_3793, w_038_3794, w_038_3795, w_038_3796, w_038_3797, w_038_3798, w_038_3799, w_038_3801, w_038_3802, w_038_3805, w_038_3806, w_038_3807, w_038_3808, w_038_3809, w_038_3810, w_038_3813, w_038_3814, w_038_3816, w_038_3817, w_038_3818, w_038_3819, w_038_3820, w_038_3821, w_038_3822, w_038_3823, w_038_3825, w_038_3826, w_038_3827, w_038_3828, w_038_3829, w_038_3830, w_038_3831, w_038_3832, w_038_3833, w_038_3834, w_038_3836, w_038_3838, w_038_3840, w_038_3841, w_038_3842, w_038_3843, w_038_3844, w_038_3845, w_038_3846, w_038_3847, w_038_3849, w_038_3850, w_038_3851, w_038_3853, w_038_3855, w_038_3856, w_038_3857, w_038_3858, w_038_3859, w_038_3860, w_038_3861, w_038_3862, w_038_3864, w_038_3866, w_038_3867, w_038_3868, w_038_3870, w_038_3872, w_038_3875, w_038_3876, w_038_3877, w_038_3880, w_038_3882, w_038_3884, w_038_3886, w_038_3887, w_038_3889, w_038_3890, w_038_3892, w_038_3893, w_038_3894, w_038_3895, w_038_3896, w_038_3898, w_038_3900, w_038_3901, w_038_3902, w_038_3904, w_038_3905, w_038_3906, w_038_3907, w_038_3908, w_038_3909, w_038_3910, w_038_3911, w_038_3912, w_038_3913, w_038_3914, w_038_3915, w_038_3916, w_038_3918, w_038_3919, w_038_3920, w_038_3922, w_038_3923, w_038_3926, w_038_3927, w_038_3928, w_038_3929, w_038_3930, w_038_3931, w_038_3932, w_038_3933, w_038_3934, w_038_3935, w_038_3936, w_038_3938, w_038_3939, w_038_3940, w_038_3941, w_038_3943, w_038_3944, w_038_3945, w_038_3946, w_038_3949, w_038_3950, w_038_3951, w_038_3952, w_038_3953, w_038_3954, w_038_3955, w_038_3956, w_038_3957, w_038_3958, w_038_3959, w_038_3962, w_038_3963, w_038_3964, w_038_3965, w_038_3966, w_038_3967, w_038_3968, w_038_3969, w_038_3971, w_038_3973, w_038_3974, w_038_3975, w_038_3976, w_038_3977, w_038_3978, w_038_3979, w_038_3980, w_038_3981, w_038_3982, w_038_3983, w_038_3984, w_038_3986, w_038_3987, w_038_3989, w_038_3990, w_038_3991, w_038_3992, w_038_3993, w_038_3995, w_038_3998, w_038_4000, w_038_4001, w_038_4002, w_038_4003, w_038_4004, w_038_4005, w_038_4007, w_038_4008, w_038_4009, w_038_4010, w_038_4011, w_038_4012, w_038_4013, w_038_4015, w_038_4016, w_038_4017, w_038_4018, w_038_4019, w_038_4020, w_038_4023, w_038_4027, w_038_4029, w_038_4031, w_038_4034, w_038_4035, w_038_4036, w_038_4037, w_038_4038, w_038_4039, w_038_4040, w_038_4041, w_038_4042, w_038_4043, w_038_4044, w_038_4046, w_038_4047, w_038_4048, w_038_4049, w_038_4050, w_038_4051, w_038_4054, w_038_4055, w_038_4056, w_038_4057, w_038_4058, w_038_4059, w_038_4060, w_038_4061, w_038_4062, w_038_4063, w_038_4065, w_038_4066, w_038_4068, w_038_4069, w_038_4071, w_038_4072, w_038_4073, w_038_4074, w_038_4075, w_038_4076, w_038_4078, w_038_4080, w_038_4082, w_038_4084, w_038_4085, w_038_4087, w_038_4088, w_038_4089, w_038_4092, w_038_4093, w_038_4094, w_038_4095, w_038_4096, w_038_4097, w_038_4099, w_038_4100, w_038_4101, w_038_4102, w_038_4104, w_038_4105, w_038_4106, w_038_4107, w_038_4108, w_038_4109, w_038_4110, w_038_4111, w_038_4112, w_038_4113, w_038_4115, w_038_4116, w_038_4117, w_038_4118, w_038_4119, w_038_4120, w_038_4121, w_038_4122, w_038_4123, w_038_4124, w_038_4125, w_038_4126, w_038_4127, w_038_4128, w_038_4129, w_038_4131, w_038_4132, w_038_4133, w_038_4134, w_038_4135, w_038_4137, w_038_4138, w_038_4139, w_038_4141, w_038_4142, w_038_4143, w_038_4144, w_038_4145, w_038_4146, w_038_4148, w_038_4149, w_038_4150, w_038_4151, w_038_4152, w_038_4153, w_038_4154, w_038_4155, w_038_4156, w_038_4157, w_038_4159, w_038_4160, w_038_4161, w_038_4162, w_038_4164, w_038_4165, w_038_4167, w_038_4170, w_038_4171, w_038_4173, w_038_4174, w_038_4176, w_038_4177, w_038_4178, w_038_4179, w_038_4180, w_038_4181, w_038_4182, w_038_4183, w_038_4184, w_038_4185, w_038_4186, w_038_4187, w_038_4188, w_038_4190, w_038_4191, w_038_4192, w_038_4193, w_038_4194, w_038_4195, w_038_4196, w_038_4197, w_038_4198, w_038_4199, w_038_4202, w_038_4204, w_038_4205, w_038_4206, w_038_4207, w_038_4208, w_038_4209, w_038_4210, w_038_4212, w_038_4213, w_038_4214, w_038_4215, w_038_4216, w_038_4217, w_038_4218, w_038_4219, w_038_4220, w_038_4222, w_038_4224, w_038_4225, w_038_4226, w_038_4227, w_038_4228, w_038_4229, w_038_4230, w_038_4231, w_038_4232, w_038_4233, w_038_4234, w_038_4239, w_038_4240, w_038_4241, w_038_4242, w_038_4243, w_038_4245, w_038_4246, w_038_4247, w_038_4248, w_038_4249, w_038_4250, w_038_4251, w_038_4253, w_038_4254, w_038_4255, w_038_4256, w_038_4258, w_038_4261, w_038_4263, w_038_4264, w_038_4265, w_038_4266, w_038_4267, w_038_4270, w_038_4271, w_038_4272, w_038_4273, w_038_4274, w_038_4276, w_038_4277, w_038_4278, w_038_4279, w_038_4281, w_038_4282, w_038_4283, w_038_4287, w_038_4288, w_038_4289, w_038_4292, w_038_4293, w_038_4294, w_038_4295, w_038_4297, w_038_4298, w_038_4299, w_038_4304, w_038_4307, w_038_4308, w_038_4309, w_038_4310, w_038_4311, w_038_4313, w_038_4314, w_038_4315, w_038_4316, w_038_4318, w_038_4319, w_038_4321, w_038_4322, w_038_4323, w_038_4324, w_038_4327, w_038_4328, w_038_4329, w_038_4330, w_038_4331, w_038_4332, w_038_4334, w_038_4335, w_038_4336, w_038_4337, w_038_4339, w_038_4340, w_038_4341, w_038_4342, w_038_4343, w_038_4344, w_038_4345, w_038_4346, w_038_4347, w_038_4348, w_038_4351, w_038_4352, w_038_4353, w_038_4354, w_038_4355, w_038_4356, w_038_4357, w_038_4358, w_038_4359, w_038_4360, w_038_4361, w_038_4362, w_038_4363, w_038_4365, w_038_4366, w_038_4367, w_038_4368, w_038_4369, w_038_4371, w_038_4372, w_038_4373, w_038_4375, w_038_4376, w_038_4377, w_038_4378, w_038_4379, w_038_4381, w_038_4382, w_038_4383, w_038_4387, w_038_4388, w_038_4391, w_038_4392, w_038_4393, w_038_4394, w_038_4395, w_038_4396, w_038_4397, w_038_4398, w_038_4399, w_038_4400, w_038_4401, w_038_4402, w_038_4403, w_038_4405, w_038_4406, w_038_4407, w_038_4408, w_038_4409, w_038_4410, w_038_4411, w_038_4412, w_038_4414, w_038_4415, w_038_4416, w_038_4417, w_038_4418, w_038_4419, w_038_4420, w_038_4421, w_038_4422, w_038_4425, w_038_4426, w_038_4427, w_038_4428, w_038_4429, w_038_4430, w_038_4431, w_038_4432, w_038_4433, w_038_4434, w_038_4435, w_038_4436, w_038_4439, w_038_4441, w_038_4444, w_038_4447, w_038_4448, w_038_4449, w_038_4450, w_038_4451, w_038_4452, w_038_4455, w_038_4456, w_038_4457, w_038_4458, w_038_4459, w_038_4460, w_038_4462, w_038_4463, w_038_4464, w_038_4465, w_038_4466, w_038_4467, w_038_4468, w_038_4469, w_038_4471, w_038_4472, w_038_4473, w_038_4475, w_038_4476, w_038_4477, w_038_4478, w_038_4479, w_038_4481, w_038_4482, w_038_4483, w_038_4484, w_038_4486, w_038_4487, w_038_4489, w_038_4491, w_038_4493, w_038_4494, w_038_4495, w_038_4496, w_038_4500, w_038_4501, w_038_4502, w_038_4503, w_038_4504, w_038_4505, w_038_4506, w_038_4508, w_038_4509, w_038_4510, w_038_4512, w_038_4513, w_038_4514, w_038_4515, w_038_4517, w_038_4518, w_038_4519, w_038_4520, w_038_4521, w_038_4522, w_038_4523, w_038_4524, w_038_4525, w_038_4526, w_038_4527, w_038_4528, w_038_4529, w_038_4530, w_038_4531, w_038_4532, w_038_4533, w_038_4534, w_038_4535, w_038_4536, w_038_4537, w_038_4538, w_038_4539, w_038_4540, w_038_4541, w_038_4549, w_038_4550, w_038_4551, w_038_4552, w_038_4553, w_038_4554, w_038_4555, w_038_4556, w_038_4560, w_038_4561, w_038_4562, w_038_4563, w_038_4565, w_038_4566, w_038_4567, w_038_4568, w_038_4569, w_038_4570, w_038_4572, w_038_4573, w_038_4574, w_038_4575, w_038_4576, w_038_4578, w_038_4579, w_038_4580, w_038_4583, w_038_4584, w_038_4585, w_038_4587, w_038_4589, w_038_4591, w_038_4594, w_038_4595, w_038_4598, w_038_4600, w_038_4601, w_038_4602, w_038_4603, w_038_4604, w_038_4605, w_038_4606, w_038_4607, w_038_4608, w_038_4610, w_038_4611, w_038_4613, w_038_4614, w_038_4615, w_038_4616, w_038_4618, w_038_4619, w_038_4620, w_038_4621, w_038_4622, w_038_4623, w_038_4624, w_038_4625, w_038_4626, w_038_4627, w_038_4628, w_038_4630, w_038_4631, w_038_4632, w_038_4633, w_038_4634, w_038_4635, w_038_4636, w_038_4637, w_038_4638, w_038_4639, w_038_4640, w_038_4641, w_038_4642, w_038_4643, w_038_4644, w_038_4646, w_038_4648, w_038_4650, w_038_4651, w_038_4652, w_038_4654, w_038_4655, w_038_4656, w_038_4657, w_038_4658, w_038_4660, w_038_4661, w_038_4663, w_038_4664, w_038_4665, w_038_4666, w_038_4669, w_038_4670, w_038_4671, w_038_4672, w_038_4673, w_038_4674, w_038_4675, w_038_4676, w_038_4677, w_038_4678, w_038_4680, w_038_4682, w_038_4683, w_038_4685, w_038_4686, w_038_4688, w_038_4689, w_038_4691, w_038_4692, w_038_4693, w_038_4694, w_038_4696, w_038_4699, w_038_4700, w_038_4701, w_038_4702, w_038_4703, w_038_4704, w_038_4705, w_038_4706, w_038_4707, w_038_4708, w_038_4709, w_038_4710, w_038_4711, w_038_4712, w_038_4714, w_038_4717, w_038_4718, w_038_4720, w_038_4721, w_038_4722, w_038_4724, w_038_4725, w_038_4726, w_038_4727, w_038_4728, w_038_4729, w_038_4732, w_038_4733, w_038_4734, w_038_4736, w_038_4739, w_038_4740, w_038_4741, w_038_4743, w_038_4744, w_038_4746, w_038_4749, w_038_4751, w_038_4752, w_038_4753, w_038_4754, w_038_4755;
  wire w_039_000, w_039_001, w_039_002, w_039_003, w_039_004, w_039_005, w_039_006, w_039_007, w_039_008, w_039_009, w_039_010, w_039_011, w_039_012, w_039_014, w_039_016, w_039_017, w_039_018, w_039_019, w_039_020, w_039_021, w_039_022, w_039_023, w_039_024, w_039_025, w_039_026, w_039_027, w_039_028, w_039_029, w_039_030, w_039_031, w_039_032, w_039_033, w_039_034, w_039_035, w_039_036, w_039_037, w_039_038, w_039_039, w_039_040, w_039_041, w_039_042, w_039_043, w_039_044, w_039_045, w_039_046, w_039_047, w_039_048, w_039_049, w_039_050, w_039_051, w_039_052, w_039_053, w_039_054, w_039_055, w_039_056, w_039_057, w_039_058, w_039_059, w_039_060, w_039_061, w_039_062, w_039_063, w_039_064, w_039_065, w_039_066, w_039_067, w_039_068, w_039_069, w_039_070, w_039_071, w_039_072, w_039_073, w_039_074, w_039_075, w_039_076, w_039_077, w_039_078, w_039_079, w_039_080, w_039_081, w_039_082, w_039_083, w_039_084, w_039_085, w_039_086, w_039_089, w_039_090, w_039_091, w_039_093, w_039_095, w_039_096, w_039_097, w_039_099, w_039_100, w_039_101, w_039_102, w_039_104, w_039_105, w_039_106, w_039_107, w_039_108, w_039_109, w_039_110, w_039_111, w_039_112, w_039_113, w_039_114, w_039_115, w_039_116, w_039_117, w_039_118, w_039_119, w_039_120, w_039_122, w_039_123, w_039_124, w_039_125, w_039_126, w_039_127, w_039_128, w_039_129, w_039_130, w_039_131, w_039_133, w_039_134, w_039_135, w_039_136, w_039_137, w_039_138, w_039_139, w_039_140, w_039_141, w_039_142, w_039_143, w_039_144, w_039_145, w_039_146, w_039_147, w_039_148, w_039_149, w_039_150, w_039_151, w_039_152, w_039_153, w_039_154, w_039_156, w_039_157, w_039_158, w_039_159, w_039_160, w_039_161, w_039_162, w_039_163, w_039_164, w_039_165, w_039_166, w_039_167, w_039_168, w_039_169, w_039_170, w_039_171, w_039_172, w_039_173, w_039_175, w_039_176, w_039_177, w_039_179, w_039_180, w_039_181, w_039_182, w_039_183, w_039_184, w_039_185, w_039_186, w_039_187, w_039_188, w_039_189, w_039_190, w_039_191, w_039_192, w_039_193, w_039_194, w_039_196, w_039_197, w_039_198, w_039_199, w_039_200, w_039_202, w_039_203, w_039_204, w_039_207, w_039_208, w_039_209, w_039_210, w_039_211, w_039_212, w_039_213, w_039_214, w_039_215, w_039_216, w_039_217, w_039_218, w_039_219, w_039_220, w_039_221, w_039_222, w_039_223, w_039_224, w_039_225, w_039_226, w_039_227, w_039_228, w_039_229, w_039_230, w_039_231, w_039_232, w_039_233, w_039_234, w_039_235, w_039_236, w_039_238, w_039_239, w_039_240, w_039_241, w_039_242, w_039_243, w_039_244, w_039_245, w_039_246, w_039_247, w_039_248, w_039_249, w_039_250, w_039_251, w_039_252, w_039_253, w_039_254, w_039_255, w_039_256, w_039_257, w_039_258, w_039_259, w_039_260, w_039_261, w_039_262, w_039_263, w_039_264, w_039_265, w_039_266, w_039_267, w_039_268, w_039_269, w_039_270, w_039_271, w_039_272, w_039_273, w_039_274, w_039_275, w_039_276, w_039_277, w_039_278, w_039_279, w_039_280, w_039_281, w_039_282, w_039_283, w_039_284, w_039_285, w_039_286, w_039_287, w_039_288, w_039_289, w_039_290, w_039_291, w_039_292, w_039_293, w_039_294, w_039_295, w_039_296, w_039_297, w_039_298, w_039_299, w_039_300, w_039_301, w_039_302, w_039_303, w_039_304, w_039_305, w_039_306, w_039_307, w_039_308, w_039_309, w_039_312, w_039_313, w_039_314, w_039_315, w_039_316, w_039_317, w_039_318, w_039_319, w_039_320, w_039_321, w_039_322, w_039_324, w_039_325, w_039_326, w_039_327, w_039_328, w_039_329, w_039_330, w_039_331, w_039_332, w_039_333, w_039_334, w_039_335, w_039_336, w_039_337, w_039_338, w_039_339, w_039_340, w_039_341, w_039_342, w_039_343, w_039_344, w_039_345, w_039_346, w_039_347, w_039_348, w_039_349, w_039_350, w_039_351, w_039_352, w_039_353, w_039_354, w_039_356, w_039_357, w_039_358, w_039_360, w_039_361, w_039_362, w_039_363, w_039_364, w_039_365, w_039_366, w_039_367, w_039_368, w_039_369, w_039_370, w_039_371, w_039_373, w_039_374, w_039_375, w_039_376, w_039_377, w_039_378, w_039_379, w_039_381, w_039_382, w_039_383, w_039_384, w_039_388, w_039_390, w_039_391, w_039_392, w_039_393, w_039_394, w_039_395, w_039_396, w_039_398, w_039_399, w_039_400, w_039_401, w_039_402, w_039_403, w_039_404, w_039_405, w_039_406, w_039_407, w_039_408, w_039_409, w_039_410, w_039_411, w_039_412, w_039_413, w_039_415, w_039_416, w_039_418, w_039_419, w_039_420, w_039_421, w_039_422, w_039_423, w_039_424, w_039_425, w_039_427, w_039_428, w_039_429, w_039_430, w_039_431, w_039_432, w_039_434, w_039_435, w_039_436, w_039_437, w_039_438, w_039_439, w_039_440, w_039_441, w_039_442, w_039_443, w_039_444, w_039_445, w_039_447, w_039_448, w_039_449, w_039_450, w_039_452, w_039_453, w_039_454, w_039_456, w_039_457, w_039_458, w_039_459, w_039_461, w_039_462, w_039_463, w_039_464, w_039_465, w_039_466, w_039_467, w_039_468, w_039_469, w_039_470, w_039_471, w_039_472, w_039_473, w_039_475, w_039_476, w_039_477, w_039_478, w_039_479, w_039_480, w_039_481, w_039_482, w_039_483, w_039_484, w_039_485, w_039_486, w_039_487, w_039_488, w_039_489, w_039_490, w_039_491, w_039_492, w_039_493, w_039_494, w_039_495, w_039_496, w_039_497, w_039_498, w_039_499, w_039_500, w_039_501, w_039_502, w_039_503, w_039_504, w_039_505, w_039_506, w_039_507, w_039_508, w_039_509, w_039_510, w_039_511, w_039_512, w_039_513, w_039_514, w_039_515, w_039_516, w_039_517, w_039_519, w_039_520, w_039_521, w_039_522, w_039_523, w_039_524, w_039_525, w_039_526, w_039_527, w_039_528, w_039_529, w_039_530, w_039_531, w_039_532, w_039_533, w_039_534, w_039_536, w_039_537, w_039_538, w_039_539, w_039_540, w_039_541, w_039_542, w_039_543, w_039_544, w_039_545, w_039_546, w_039_547, w_039_548, w_039_549, w_039_550, w_039_551, w_039_553, w_039_555, w_039_558, w_039_559, w_039_560, w_039_561, w_039_562, w_039_564, w_039_565, w_039_566, w_039_568, w_039_569, w_039_570, w_039_571, w_039_573, w_039_574, w_039_575, w_039_576, w_039_577, w_039_578, w_039_579, w_039_581, w_039_582, w_039_583, w_039_584, w_039_585, w_039_586, w_039_587, w_039_588, w_039_589, w_039_590, w_039_591, w_039_592, w_039_593, w_039_595, w_039_596, w_039_597, w_039_598, w_039_599, w_039_600, w_039_601, w_039_602, w_039_603, w_039_604, w_039_605, w_039_606, w_039_607, w_039_608, w_039_609, w_039_610, w_039_611, w_039_612, w_039_613, w_039_614, w_039_615, w_039_616, w_039_617, w_039_618, w_039_619, w_039_621, w_039_622, w_039_623, w_039_624, w_039_625, w_039_626, w_039_628, w_039_629, w_039_630, w_039_631, w_039_633, w_039_634, w_039_635, w_039_636, w_039_637, w_039_638, w_039_639, w_039_640, w_039_641, w_039_642, w_039_643, w_039_644, w_039_645, w_039_647, w_039_648, w_039_649, w_039_650, w_039_651, w_039_652, w_039_653, w_039_654, w_039_655, w_039_656, w_039_658, w_039_659, w_039_660, w_039_661, w_039_662, w_039_663, w_039_664, w_039_665, w_039_666, w_039_667, w_039_669, w_039_670, w_039_671, w_039_672, w_039_673, w_039_674, w_039_675, w_039_676, w_039_677, w_039_678, w_039_679, w_039_680, w_039_681, w_039_682, w_039_684, w_039_685, w_039_686, w_039_687, w_039_688, w_039_689, w_039_690, w_039_691, w_039_693, w_039_694, w_039_695, w_039_696, w_039_697, w_039_698, w_039_700, w_039_701, w_039_702, w_039_703, w_039_704, w_039_705, w_039_706, w_039_707, w_039_708, w_039_709, w_039_710, w_039_711, w_039_712, w_039_713, w_039_714, w_039_716, w_039_719, w_039_720, w_039_721, w_039_722, w_039_723, w_039_724, w_039_725, w_039_727, w_039_728, w_039_729, w_039_730, w_039_731, w_039_732, w_039_734, w_039_735, w_039_737, w_039_738, w_039_739, w_039_740, w_039_741, w_039_742, w_039_743, w_039_744, w_039_745, w_039_746, w_039_747, w_039_748, w_039_749, w_039_750, w_039_751, w_039_752, w_039_753, w_039_754, w_039_755, w_039_756, w_039_757, w_039_758, w_039_759, w_039_761, w_039_762, w_039_763, w_039_764, w_039_766, w_039_767, w_039_768, w_039_769, w_039_770, w_039_771, w_039_772, w_039_773, w_039_774, w_039_775, w_039_776, w_039_777, w_039_778, w_039_779, w_039_780, w_039_781, w_039_782, w_039_783, w_039_784, w_039_785, w_039_787, w_039_788, w_039_789, w_039_790, w_039_791, w_039_792, w_039_793, w_039_794, w_039_795, w_039_796, w_039_797, w_039_798, w_039_799, w_039_800, w_039_802, w_039_803, w_039_804, w_039_805, w_039_806, w_039_807, w_039_808, w_039_809, w_039_810, w_039_811, w_039_813, w_039_814, w_039_815, w_039_816, w_039_817, w_039_818, w_039_819, w_039_820, w_039_821, w_039_822, w_039_823, w_039_825, w_039_826, w_039_827, w_039_828, w_039_829, w_039_830, w_039_831, w_039_832, w_039_833, w_039_834, w_039_835, w_039_836, w_039_837, w_039_838, w_039_839, w_039_840, w_039_842, w_039_843, w_039_844, w_039_845, w_039_846, w_039_847, w_039_848, w_039_849, w_039_850, w_039_851, w_039_852, w_039_853, w_039_854, w_039_855, w_039_856, w_039_857, w_039_858, w_039_859, w_039_860, w_039_861, w_039_862, w_039_863, w_039_864, w_039_865, w_039_866, w_039_867, w_039_868, w_039_869, w_039_870, w_039_871, w_039_872, w_039_874, w_039_875, w_039_876, w_039_877, w_039_878, w_039_879, w_039_880, w_039_881, w_039_882, w_039_883, w_039_884, w_039_885, w_039_886, w_039_888, w_039_889, w_039_890, w_039_891, w_039_893, w_039_894, w_039_895, w_039_896, w_039_897, w_039_898, w_039_899, w_039_900, w_039_901, w_039_902, w_039_904, w_039_905, w_039_906, w_039_907, w_039_908, w_039_910, w_039_911, w_039_912, w_039_913, w_039_914, w_039_915, w_039_916, w_039_917, w_039_918, w_039_919, w_039_920, w_039_921, w_039_922, w_039_923, w_039_924, w_039_925, w_039_926, w_039_927, w_039_928, w_039_929, w_039_930, w_039_931, w_039_932, w_039_933, w_039_934, w_039_935, w_039_936, w_039_937, w_039_938, w_039_939, w_039_940, w_039_941, w_039_942, w_039_943, w_039_944, w_039_945, w_039_946, w_039_947, w_039_948, w_039_949, w_039_950, w_039_951, w_039_952, w_039_953, w_039_954, w_039_955, w_039_956, w_039_957, w_039_958, w_039_959, w_039_960, w_039_961, w_039_962, w_039_963, w_039_964, w_039_965, w_039_966, w_039_967, w_039_968, w_039_969, w_039_971, w_039_972, w_039_973, w_039_974, w_039_975, w_039_976, w_039_977, w_039_978, w_039_979, w_039_980, w_039_981, w_039_982, w_039_983, w_039_984, w_039_985, w_039_986, w_039_987, w_039_988, w_039_989, w_039_990, w_039_992, w_039_993, w_039_994, w_039_995, w_039_996, w_039_997, w_039_998, w_039_999, w_039_1000, w_039_1001, w_039_1002, w_039_1003, w_039_1004, w_039_1005, w_039_1006, w_039_1007, w_039_1008, w_039_1009, w_039_1010, w_039_1011, w_039_1012, w_039_1013, w_039_1014, w_039_1015, w_039_1016, w_039_1017, w_039_1018, w_039_1019, w_039_1020, w_039_1021, w_039_1022, w_039_1023, w_039_1024, w_039_1025, w_039_1026, w_039_1027, w_039_1029, w_039_1031, w_039_1032, w_039_1033, w_039_1034, w_039_1035, w_039_1036, w_039_1037, w_039_1038, w_039_1039, w_039_1040, w_039_1041, w_039_1042, w_039_1043, w_039_1044, w_039_1045, w_039_1046, w_039_1047, w_039_1048, w_039_1049, w_039_1050, w_039_1051, w_039_1052, w_039_1053, w_039_1054, w_039_1057, w_039_1058, w_039_1059, w_039_1060, w_039_1061, w_039_1062, w_039_1063, w_039_1064, w_039_1065, w_039_1066, w_039_1067, w_039_1069, w_039_1070, w_039_1071, w_039_1072, w_039_1073, w_039_1074, w_039_1075, w_039_1076, w_039_1077, w_039_1078, w_039_1079, w_039_1080, w_039_1081, w_039_1082, w_039_1083, w_039_1084, w_039_1085, w_039_1086, w_039_1087, w_039_1088, w_039_1089, w_039_1090, w_039_1091, w_039_1092, w_039_1093, w_039_1094, w_039_1095, w_039_1096, w_039_1097, w_039_1099, w_039_1100, w_039_1101, w_039_1103, w_039_1104, w_039_1105, w_039_1106, w_039_1107, w_039_1108, w_039_1109, w_039_1111, w_039_1112, w_039_1113, w_039_1114, w_039_1115, w_039_1116, w_039_1118, w_039_1119, w_039_1120, w_039_1121, w_039_1122, w_039_1123, w_039_1124, w_039_1125, w_039_1126, w_039_1127, w_039_1128, w_039_1129, w_039_1130, w_039_1131, w_039_1132, w_039_1133, w_039_1134, w_039_1135, w_039_1136, w_039_1137, w_039_1138, w_039_1139, w_039_1140, w_039_1141, w_039_1142, w_039_1143, w_039_1144, w_039_1145, w_039_1146, w_039_1148, w_039_1149, w_039_1150, w_039_1151, w_039_1152, w_039_1153, w_039_1154, w_039_1155, w_039_1156, w_039_1157, w_039_1158, w_039_1159, w_039_1160, w_039_1161, w_039_1162, w_039_1163, w_039_1164, w_039_1165, w_039_1166, w_039_1167, w_039_1168, w_039_1169, w_039_1170, w_039_1171, w_039_1172, w_039_1173, w_039_1175, w_039_1176, w_039_1177, w_039_1178, w_039_1179, w_039_1180, w_039_1181, w_039_1182, w_039_1183, w_039_1184, w_039_1185, w_039_1186, w_039_1188, w_039_1189, w_039_1190, w_039_1191, w_039_1192, w_039_1193, w_039_1194, w_039_1195, w_039_1196, w_039_1197, w_039_1198, w_039_1200, w_039_1201, w_039_1202, w_039_1203, w_039_1204, w_039_1205, w_039_1206, w_039_1207, w_039_1208, w_039_1209, w_039_1210, w_039_1211, w_039_1212, w_039_1214, w_039_1215, w_039_1216, w_039_1217, w_039_1218, w_039_1219, w_039_1220, w_039_1221, w_039_1222, w_039_1223, w_039_1224, w_039_1225, w_039_1226, w_039_1227, w_039_1228, w_039_1229, w_039_1230, w_039_1231, w_039_1232, w_039_1233, w_039_1234, w_039_1235, w_039_1236, w_039_1237, w_039_1238, w_039_1239, w_039_1240, w_039_1241, w_039_1242, w_039_1243, w_039_1244, w_039_1245, w_039_1246, w_039_1247, w_039_1248, w_039_1249, w_039_1250, w_039_1251, w_039_1252, w_039_1253, w_039_1254, w_039_1255, w_039_1256, w_039_1257, w_039_1258, w_039_1259, w_039_1260, w_039_1261, w_039_1262, w_039_1263, w_039_1264, w_039_1265, w_039_1266, w_039_1267, w_039_1268, w_039_1269, w_039_1270, w_039_1271, w_039_1272, w_039_1274, w_039_1275, w_039_1276, w_039_1277, w_039_1278, w_039_1279, w_039_1280, w_039_1281, w_039_1282, w_039_1283, w_039_1285, w_039_1286, w_039_1287, w_039_1288, w_039_1289, w_039_1290, w_039_1291, w_039_1292, w_039_1293, w_039_1294, w_039_1295, w_039_1296, w_039_1297, w_039_1298, w_039_1299, w_039_1300, w_039_1301, w_039_1302, w_039_1303, w_039_1304, w_039_1305, w_039_1306, w_039_1308, w_039_1309, w_039_1311, w_039_1312, w_039_1313, w_039_1314, w_039_1315, w_039_1316, w_039_1317, w_039_1318, w_039_1319, w_039_1320, w_039_1321, w_039_1322, w_039_1323, w_039_1324, w_039_1326, w_039_1327, w_039_1328, w_039_1329, w_039_1330, w_039_1331, w_039_1332, w_039_1333, w_039_1334, w_039_1335, w_039_1336, w_039_1338, w_039_1339, w_039_1340, w_039_1341, w_039_1342, w_039_1343, w_039_1344, w_039_1345, w_039_1346, w_039_1347, w_039_1348, w_039_1349, w_039_1350, w_039_1351, w_039_1352, w_039_1354, w_039_1355, w_039_1356, w_039_1357, w_039_1358, w_039_1359, w_039_1360, w_039_1361, w_039_1362, w_039_1363, w_039_1364, w_039_1365, w_039_1367, w_039_1368, w_039_1369, w_039_1370, w_039_1372, w_039_1373, w_039_1374, w_039_1375, w_039_1376, w_039_1377, w_039_1378, w_039_1380, w_039_1381, w_039_1382, w_039_1383, w_039_1384, w_039_1385, w_039_1386, w_039_1387, w_039_1389, w_039_1390, w_039_1391, w_039_1392, w_039_1393, w_039_1395, w_039_1396, w_039_1397, w_039_1398, w_039_1399, w_039_1401, w_039_1402, w_039_1403, w_039_1404, w_039_1405, w_039_1406, w_039_1408, w_039_1409, w_039_1410, w_039_1411, w_039_1412, w_039_1413, w_039_1414, w_039_1415, w_039_1416, w_039_1417, w_039_1418, w_039_1419, w_039_1420, w_039_1421, w_039_1422, w_039_1423, w_039_1424, w_039_1425, w_039_1426, w_039_1427, w_039_1428, w_039_1429, w_039_1430, w_039_1432, w_039_1433, w_039_1434, w_039_1435, w_039_1436, w_039_1437, w_039_1438, w_039_1439, w_039_1440, w_039_1442, w_039_1443, w_039_1444, w_039_1446, w_039_1447, w_039_1448, w_039_1449, w_039_1450, w_039_1451, w_039_1452, w_039_1453, w_039_1454, w_039_1455, w_039_1456, w_039_1457, w_039_1458, w_039_1459, w_039_1460, w_039_1461, w_039_1462, w_039_1463, w_039_1464, w_039_1465, w_039_1467, w_039_1468, w_039_1469, w_039_1470, w_039_1471, w_039_1472, w_039_1473, w_039_1475, w_039_1476, w_039_1477, w_039_1478, w_039_1479, w_039_1480, w_039_1481, w_039_1482, w_039_1483, w_039_1484, w_039_1485, w_039_1486, w_039_1487, w_039_1488, w_039_1489, w_039_1490, w_039_1491, w_039_1492, w_039_1494, w_039_1495, w_039_1497, w_039_1498, w_039_1499, w_039_1500, w_039_1501, w_039_1502, w_039_1503, w_039_1504, w_039_1505, w_039_1506, w_039_1507, w_039_1508, w_039_1509, w_039_1510, w_039_1511, w_039_1512, w_039_1514, w_039_1515, w_039_1516, w_039_1517, w_039_1518, w_039_1519, w_039_1520, w_039_1521, w_039_1522, w_039_1523, w_039_1524, w_039_1525, w_039_1526, w_039_1527, w_039_1528, w_039_1529, w_039_1530, w_039_1532, w_039_1533, w_039_1534, w_039_1535, w_039_1536, w_039_1537, w_039_1538, w_039_1539, w_039_1540, w_039_1541, w_039_1542, w_039_1543, w_039_1544, w_039_1545, w_039_1546, w_039_1547, w_039_1548, w_039_1549, w_039_1551, w_039_1552, w_039_1554, w_039_1555, w_039_1556, w_039_1557, w_039_1558, w_039_1559, w_039_1560, w_039_1561, w_039_1562, w_039_1563, w_039_1564, w_039_1565, w_039_1566, w_039_1567, w_039_1568, w_039_1569, w_039_1570, w_039_1572, w_039_1574, w_039_1575, w_039_1576, w_039_1577, w_039_1578, w_039_1579, w_039_1580, w_039_1581, w_039_1582, w_039_1583, w_039_1584, w_039_1585, w_039_1586, w_039_1587, w_039_1589, w_039_1591, w_039_1592, w_039_1593, w_039_1594, w_039_1596, w_039_1597, w_039_1598, w_039_1599, w_039_1600, w_039_1601, w_039_1602, w_039_1603, w_039_1604, w_039_1605, w_039_1606, w_039_1607, w_039_1608, w_039_1610, w_039_1611, w_039_1613, w_039_1614, w_039_1615, w_039_1616, w_039_1617, w_039_1618, w_039_1619, w_039_1620, w_039_1621, w_039_1623, w_039_1624, w_039_1625, w_039_1626, w_039_1627, w_039_1628, w_039_1629, w_039_1630, w_039_1631, w_039_1633, w_039_1634, w_039_1635, w_039_1636, w_039_1637, w_039_1638, w_039_1639, w_039_1640, w_039_1641, w_039_1642, w_039_1643, w_039_1644, w_039_1645, w_039_1646, w_039_1647, w_039_1648, w_039_1649, w_039_1651, w_039_1653, w_039_1654, w_039_1655, w_039_1656, w_039_1657, w_039_1658, w_039_1659, w_039_1660, w_039_1662, w_039_1663, w_039_1664, w_039_1665, w_039_1666, w_039_1667, w_039_1668, w_039_1669, w_039_1670, w_039_1671, w_039_1672, w_039_1674, w_039_1675, w_039_1676, w_039_1677, w_039_1678, w_039_1682, w_039_1683, w_039_1684, w_039_1686, w_039_1687, w_039_1688, w_039_1689, w_039_1690, w_039_1691, w_039_1693, w_039_1694, w_039_1695, w_039_1696, w_039_1698, w_039_1699, w_039_1700, w_039_1702, w_039_1703, w_039_1705, w_039_1706, w_039_1707, w_039_1708, w_039_1709, w_039_1710, w_039_1711, w_039_1712, w_039_1713, w_039_1714, w_039_1715, w_039_1716, w_039_1717, w_039_1718, w_039_1719, w_039_1720, w_039_1721, w_039_1722, w_039_1724, w_039_1725, w_039_1727, w_039_1728, w_039_1729, w_039_1730, w_039_1732, w_039_1733, w_039_1734, w_039_1736, w_039_1738, w_039_1739, w_039_1740, w_039_1741, w_039_1742, w_039_1743, w_039_1744, w_039_1745, w_039_1746, w_039_1748, w_039_1749, w_039_1754, w_039_1756, w_039_1757, w_039_1758, w_039_1759, w_039_1760, w_039_1761, w_039_1762, w_039_1763, w_039_1764, w_039_1765, w_039_1766, w_039_1767, w_039_1769, w_039_1770, w_039_1771, w_039_1772, w_039_1773, w_039_1774, w_039_1775, w_039_1776, w_039_1777, w_039_1778, w_039_1779, w_039_1780, w_039_1781, w_039_1782, w_039_1783, w_039_1784, w_039_1785, w_039_1786, w_039_1788, w_039_1789, w_039_1790, w_039_1791, w_039_1793, w_039_1794, w_039_1796, w_039_1798, w_039_1799, w_039_1800, w_039_1801, w_039_1802, w_039_1803, w_039_1804, w_039_1805, w_039_1806, w_039_1807, w_039_1808, w_039_1809, w_039_1810, w_039_1812, w_039_1813, w_039_1814, w_039_1815, w_039_1816, w_039_1817, w_039_1818, w_039_1819, w_039_1820, w_039_1821, w_039_1823, w_039_1824, w_039_1825, w_039_1826, w_039_1827, w_039_1828, w_039_1829, w_039_1830, w_039_1831, w_039_1832, w_039_1833, w_039_1834, w_039_1835, w_039_1837, w_039_1840, w_039_1841, w_039_1842, w_039_1844, w_039_1845, w_039_1846, w_039_1847, w_039_1848, w_039_1850, w_039_1851, w_039_1852, w_039_1853, w_039_1854, w_039_1855, w_039_1856, w_039_1857, w_039_1858, w_039_1859, w_039_1860, w_039_1861, w_039_1862, w_039_1863, w_039_1864, w_039_1865, w_039_1866, w_039_1867, w_039_1868, w_039_1869, w_039_1871, w_039_1872, w_039_1874, w_039_1875, w_039_1876, w_039_1877, w_039_1878, w_039_1879, w_039_1880, w_039_1882, w_039_1883, w_039_1884, w_039_1885, w_039_1886, w_039_1887, w_039_1889, w_039_1890, w_039_1891, w_039_1893, w_039_1894, w_039_1895, w_039_1896, w_039_1898, w_039_1899, w_039_1900, w_039_1901, w_039_1902, w_039_1903, w_039_1904, w_039_1905, w_039_1906, w_039_1908, w_039_1909, w_039_1911, w_039_1912, w_039_1913, w_039_1914, w_039_1915, w_039_1916, w_039_1918, w_039_1919, w_039_1920, w_039_1921, w_039_1922, w_039_1923, w_039_1924, w_039_1925, w_039_1926, w_039_1927, w_039_1928, w_039_1929, w_039_1930, w_039_1931, w_039_1932, w_039_1933, w_039_1934, w_039_1936, w_039_1937, w_039_1938, w_039_1939, w_039_1940, w_039_1943, w_039_1944, w_039_1946, w_039_1947, w_039_1948, w_039_1949, w_039_1951, w_039_1952, w_039_1953, w_039_1954, w_039_1955, w_039_1957, w_039_1958, w_039_1959, w_039_1960, w_039_1961, w_039_1962, w_039_1963, w_039_1964, w_039_1965, w_039_1966, w_039_1967, w_039_1968, w_039_1969, w_039_1970, w_039_1972, w_039_1973, w_039_1974, w_039_1975, w_039_1976, w_039_1977, w_039_1978, w_039_1979, w_039_1981, w_039_1982, w_039_1983, w_039_1984, w_039_1986, w_039_1987, w_039_1988, w_039_1989, w_039_1990, w_039_1991, w_039_1992, w_039_1993, w_039_1994, w_039_1995, w_039_1996, w_039_1997, w_039_1998, w_039_1999, w_039_2000, w_039_2001, w_039_2003, w_039_2004, w_039_2005, w_039_2006, w_039_2007, w_039_2008, w_039_2009, w_039_2010, w_039_2011, w_039_2012, w_039_2013, w_039_2014, w_039_2015, w_039_2016, w_039_2017, w_039_2019, w_039_2020, w_039_2021, w_039_2022, w_039_2023, w_039_2025, w_039_2026, w_039_2027, w_039_2028, w_039_2030, w_039_2031, w_039_2032, w_039_2033, w_039_2034, w_039_2035, w_039_2036, w_039_2037, w_039_2039, w_039_2040, w_039_2041, w_039_2042, w_039_2043, w_039_2044, w_039_2045, w_039_2046, w_039_2047, w_039_2048, w_039_2049, w_039_2050, w_039_2051, w_039_2052, w_039_2053, w_039_2055, w_039_2057, w_039_2058, w_039_2060, w_039_2061, w_039_2062, w_039_2064, w_039_2065, w_039_2066, w_039_2067, w_039_2068, w_039_2069, w_039_2070, w_039_2071, w_039_2072, w_039_2074, w_039_2076, w_039_2077, w_039_2078, w_039_2079, w_039_2080, w_039_2082, w_039_2083, w_039_2085, w_039_2086, w_039_2087, w_039_2089, w_039_2090, w_039_2091, w_039_2092, w_039_2093, w_039_2095, w_039_2096, w_039_2097, w_039_2098, w_039_2099, w_039_2101, w_039_2102, w_039_2103, w_039_2104, w_039_2105, w_039_2106, w_039_2108, w_039_2109, w_039_2110, w_039_2111, w_039_2112, w_039_2113, w_039_2114, w_039_2115, w_039_2116, w_039_2117, w_039_2118, w_039_2119, w_039_2121, w_039_2123, w_039_2124, w_039_2126, w_039_2127, w_039_2128, w_039_2129, w_039_2130, w_039_2131, w_039_2132, w_039_2133, w_039_2134, w_039_2135, w_039_2137, w_039_2138, w_039_2140, w_039_2141, w_039_2142, w_039_2143, w_039_2144, w_039_2145, w_039_2146, w_039_2147, w_039_2148, w_039_2150, w_039_2151, w_039_2152, w_039_2154, w_039_2155, w_039_2156, w_039_2158, w_039_2159, w_039_2160, w_039_2161, w_039_2163, w_039_2164, w_039_2165, w_039_2166, w_039_2167, w_039_2168, w_039_2169, w_039_2171, w_039_2172, w_039_2173, w_039_2174, w_039_2175, w_039_2176, w_039_2177, w_039_2178, w_039_2179, w_039_2180, w_039_2181, w_039_2182, w_039_2183, w_039_2184, w_039_2185, w_039_2186, w_039_2187, w_039_2188, w_039_2189, w_039_2191, w_039_2192, w_039_2193, w_039_2194, w_039_2195, w_039_2197, w_039_2198, w_039_2199, w_039_2200, w_039_2202, w_039_2204, w_039_2205, w_039_2206, w_039_2207, w_039_2208, w_039_2209, w_039_2210, w_039_2212, w_039_2213, w_039_2214, w_039_2216, w_039_2217, w_039_2219, w_039_2220, w_039_2221, w_039_2222, w_039_2223, w_039_2224, w_039_2225, w_039_2226, w_039_2228, w_039_2229, w_039_2230, w_039_2231, w_039_2232, w_039_2233, w_039_2234, w_039_2235, w_039_2236, w_039_2237, w_039_2238, w_039_2239, w_039_2240, w_039_2241, w_039_2242, w_039_2243, w_039_2244, w_039_2246, w_039_2247, w_039_2248, w_039_2249, w_039_2250, w_039_2251, w_039_2253, w_039_2254, w_039_2255, w_039_2256, w_039_2257, w_039_2258, w_039_2259, w_039_2260, w_039_2261, w_039_2262, w_039_2263, w_039_2264, w_039_2265, w_039_2266, w_039_2268, w_039_2270, w_039_2271, w_039_2273, w_039_2274, w_039_2275, w_039_2276, w_039_2277, w_039_2278, w_039_2279, w_039_2280, w_039_2281, w_039_2282, w_039_2283, w_039_2284, w_039_2285, w_039_2286, w_039_2287, w_039_2288, w_039_2289, w_039_2290, w_039_2291, w_039_2292, w_039_2293, w_039_2294, w_039_2295, w_039_2296, w_039_2297, w_039_2299, w_039_2300, w_039_2302, w_039_2303, w_039_2304, w_039_2305, w_039_2306, w_039_2307, w_039_2308, w_039_2309, w_039_2310, w_039_2311, w_039_2312, w_039_2313, w_039_2314, w_039_2315, w_039_2316, w_039_2317, w_039_2318, w_039_2319, w_039_2320, w_039_2321, w_039_2322, w_039_2323, w_039_2324, w_039_2325, w_039_2326, w_039_2327, w_039_2328, w_039_2329, w_039_2330, w_039_2331, w_039_2332, w_039_2333, w_039_2334, w_039_2335, w_039_2336, w_039_2337, w_039_2339, w_039_2340, w_039_2341, w_039_2342, w_039_2343, w_039_2345, w_039_2347, w_039_2348, w_039_2350, w_039_2351, w_039_2352, w_039_2353, w_039_2354, w_039_2355, w_039_2357, w_039_2358, w_039_2359, w_039_2360, w_039_2361, w_039_2362, w_039_2363, w_039_2364, w_039_2365, w_039_2366, w_039_2367, w_039_2368, w_039_2369, w_039_2370, w_039_2371, w_039_2372, w_039_2373, w_039_2374, w_039_2375, w_039_2376, w_039_2377, w_039_2378, w_039_2379, w_039_2380, w_039_2381, w_039_2382, w_039_2383, w_039_2384, w_039_2385, w_039_2386, w_039_2387, w_039_2388, w_039_2389, w_039_2390, w_039_2391, w_039_2392, w_039_2393, w_039_2395, w_039_2396, w_039_2397, w_039_2398, w_039_2399, w_039_2401, w_039_2402, w_039_2403, w_039_2405, w_039_2406, w_039_2407, w_039_2409, w_039_2410, w_039_2411, w_039_2412, w_039_2413, w_039_2414, w_039_2415, w_039_2416, w_039_2417, w_039_2418, w_039_2419, w_039_2420, w_039_2421, w_039_2423, w_039_2424, w_039_2425, w_039_2426, w_039_2427, w_039_2428, w_039_2429, w_039_2430, w_039_2431, w_039_2432, w_039_2434, w_039_2435, w_039_2436, w_039_2437, w_039_2438, w_039_2439, w_039_2440, w_039_2441, w_039_2442, w_039_2443, w_039_2444, w_039_2445, w_039_2446, w_039_2447, w_039_2448, w_039_2450, w_039_2451, w_039_2452, w_039_2453, w_039_2454, w_039_2455, w_039_2458, w_039_2459, w_039_2460, w_039_2462, w_039_2464, w_039_2465, w_039_2466, w_039_2467, w_039_2468, w_039_2469, w_039_2470, w_039_2471, w_039_2472, w_039_2475, w_039_2476, w_039_2477, w_039_2478, w_039_2479, w_039_2480, w_039_2481, w_039_2482, w_039_2483, w_039_2484, w_039_2485, w_039_2486, w_039_2488, w_039_2489, w_039_2490, w_039_2491, w_039_2492, w_039_2493, w_039_2494, w_039_2495, w_039_2496, w_039_2497, w_039_2498, w_039_2500, w_039_2501, w_039_2502, w_039_2504, w_039_2505, w_039_2506, w_039_2507, w_039_2509, w_039_2510, w_039_2511, w_039_2512, w_039_2513, w_039_2514, w_039_2515, w_039_2516, w_039_2518, w_039_2519, w_039_2520, w_039_2521, w_039_2522, w_039_2523, w_039_2525, w_039_2526, w_039_2527, w_039_2528, w_039_2529, w_039_2530, w_039_2531, w_039_2532, w_039_2533, w_039_2536, w_039_2537, w_039_2538, w_039_2539, w_039_2540, w_039_2541, w_039_2542, w_039_2543, w_039_2544, w_039_2545, w_039_2547, w_039_2548, w_039_2549, w_039_2550, w_039_2551, w_039_2553, w_039_2554, w_039_2557, w_039_2558, w_039_2559, w_039_2562, w_039_2563, w_039_2564, w_039_2565, w_039_2567, w_039_2569, w_039_2570, w_039_2571, w_039_2573, w_039_2575, w_039_2576, w_039_2577, w_039_2578, w_039_2579, w_039_2580, w_039_2581, w_039_2582, w_039_2583, w_039_2584, w_039_2585, w_039_2586, w_039_2587, w_039_2588, w_039_2589, w_039_2590, w_039_2591, w_039_2594, w_039_2595, w_039_2596, w_039_2597, w_039_2598, w_039_2599, w_039_2600, w_039_2601, w_039_2602, w_039_2603, w_039_2604, w_039_2605, w_039_2607, w_039_2608, w_039_2610, w_039_2612, w_039_2615, w_039_2616, w_039_2617, w_039_2619, w_039_2620, w_039_2621, w_039_2622, w_039_2623, w_039_2624, w_039_2626, w_039_2627, w_039_2628, w_039_2629, w_039_2630, w_039_2631, w_039_2632, w_039_2633, w_039_2634, w_039_2635, w_039_2638, w_039_2639, w_039_2641, w_039_2642, w_039_2644, w_039_2645, w_039_2646, w_039_2647, w_039_2648, w_039_2650, w_039_2652, w_039_2653, w_039_2654, w_039_2655, w_039_2657, w_039_2658, w_039_2659, w_039_2660, w_039_2661, w_039_2662, w_039_2663, w_039_2665, w_039_2666, w_039_2667, w_039_2668, w_039_2669, w_039_2670, w_039_2671, w_039_2672, w_039_2673, w_039_2674, w_039_2675, w_039_2676, w_039_2678, w_039_2679, w_039_2680, w_039_2681, w_039_2682, w_039_2684, w_039_2685, w_039_2687, w_039_2688, w_039_2689, w_039_2691, w_039_2693, w_039_2694, w_039_2695, w_039_2696, w_039_2698, w_039_2699, w_039_2700, w_039_2701, w_039_2703, w_039_2704, w_039_2705, w_039_2706, w_039_2708, w_039_2709, w_039_2710, w_039_2712, w_039_2713, w_039_2714, w_039_2715, w_039_2716, w_039_2717, w_039_2718, w_039_2719, w_039_2720, w_039_2721, w_039_2723, w_039_2724, w_039_2725, w_039_2726, w_039_2727, w_039_2728, w_039_2729, w_039_2730, w_039_2731, w_039_2732, w_039_2733, w_039_2734, w_039_2735, w_039_2736, w_039_2737, w_039_2738, w_039_2739, w_039_2740, w_039_2741, w_039_2742, w_039_2744, w_039_2745, w_039_2746, w_039_2747, w_039_2748, w_039_2749, w_039_2750, w_039_2751, w_039_2752, w_039_2753, w_039_2754, w_039_2755, w_039_2756, w_039_2757, w_039_2758, w_039_2759, w_039_2760, w_039_2761, w_039_2762, w_039_2763, w_039_2764, w_039_2765, w_039_2766, w_039_2767, w_039_2768, w_039_2771, w_039_2772, w_039_2773, w_039_2774, w_039_2775, w_039_2777, w_039_2778, w_039_2779, w_039_2780, w_039_2781, w_039_2782, w_039_2783, w_039_2784, w_039_2785, w_039_2786, w_039_2787, w_039_2788, w_039_2789, w_039_2790, w_039_2791, w_039_2792, w_039_2793, w_039_2795, w_039_2796, w_039_2797, w_039_2798, w_039_2800, w_039_2801, w_039_2802, w_039_2803, w_039_2804, w_039_2805, w_039_2806, w_039_2807, w_039_2809, w_039_2810, w_039_2812, w_039_2814, w_039_2815, w_039_2816, w_039_2817, w_039_2818;
  wire w_040_001, w_040_002, w_040_003, w_040_004, w_040_005, w_040_006, w_040_007, w_040_008, w_040_009, w_040_011, w_040_012, w_040_013, w_040_014, w_040_015, w_040_018, w_040_019, w_040_020, w_040_021, w_040_022, w_040_023, w_040_024, w_040_025, w_040_026, w_040_027, w_040_028, w_040_029, w_040_030, w_040_031, w_040_032, w_040_033, w_040_035, w_040_036, w_040_037, w_040_038, w_040_039, w_040_040, w_040_041, w_040_042, w_040_043, w_040_044, w_040_045, w_040_046, w_040_047, w_040_048, w_040_050, w_040_051, w_040_052, w_040_053, w_040_054, w_040_056, w_040_057, w_040_058, w_040_059, w_040_061, w_040_062, w_040_063, w_040_064, w_040_065, w_040_066, w_040_067, w_040_068, w_040_069, w_040_070, w_040_071, w_040_073, w_040_074, w_040_075, w_040_076, w_040_077, w_040_079, w_040_080, w_040_081, w_040_082, w_040_084, w_040_085, w_040_086, w_040_087, w_040_088, w_040_089, w_040_090, w_040_091, w_040_092, w_040_093, w_040_094, w_040_095, w_040_096, w_040_097, w_040_098, w_040_099, w_040_100, w_040_101, w_040_103, w_040_104, w_040_105, w_040_106, w_040_107, w_040_108, w_040_109, w_040_110, w_040_111, w_040_112, w_040_113, w_040_114, w_040_115, w_040_117, w_040_118, w_040_119, w_040_120, w_040_121, w_040_122, w_040_123, w_040_124, w_040_125, w_040_126, w_040_127, w_040_128, w_040_129, w_040_130, w_040_132, w_040_133, w_040_134, w_040_135, w_040_136, w_040_137, w_040_139, w_040_140, w_040_141, w_040_142, w_040_143, w_040_144, w_040_146, w_040_147, w_040_148, w_040_149, w_040_150, w_040_151, w_040_152, w_040_153, w_040_154, w_040_155, w_040_156, w_040_157, w_040_159, w_040_161, w_040_164, w_040_165, w_040_166, w_040_167, w_040_168, w_040_169, w_040_170, w_040_171, w_040_173, w_040_174, w_040_175, w_040_176, w_040_177, w_040_179, w_040_180, w_040_181, w_040_182, w_040_183, w_040_184, w_040_185, w_040_186, w_040_187, w_040_188, w_040_189, w_040_190, w_040_191, w_040_194, w_040_195, w_040_196, w_040_197, w_040_198, w_040_199, w_040_200, w_040_201, w_040_202, w_040_203, w_040_204, w_040_205, w_040_206, w_040_208, w_040_210, w_040_211, w_040_213, w_040_214, w_040_215, w_040_216, w_040_217, w_040_218, w_040_219, w_040_221, w_040_222, w_040_223, w_040_225, w_040_226, w_040_228, w_040_229, w_040_231, w_040_232, w_040_233, w_040_234, w_040_235, w_040_236, w_040_237, w_040_238, w_040_239, w_040_241, w_040_242, w_040_243, w_040_244, w_040_245, w_040_246, w_040_247, w_040_248, w_040_249, w_040_250, w_040_252, w_040_253, w_040_254, w_040_255, w_040_256, w_040_257, w_040_258, w_040_259, w_040_260, w_040_261, w_040_262, w_040_263, w_040_264, w_040_265, w_040_266, w_040_267, w_040_268, w_040_269, w_040_270, w_040_271, w_040_272, w_040_273, w_040_278, w_040_279, w_040_280, w_040_281, w_040_282, w_040_283, w_040_284, w_040_285, w_040_286, w_040_288, w_040_289, w_040_290, w_040_291, w_040_292, w_040_293, w_040_294, w_040_296, w_040_297, w_040_298, w_040_299, w_040_300, w_040_301, w_040_302, w_040_303, w_040_304, w_040_305, w_040_306, w_040_307, w_040_308, w_040_309, w_040_311, w_040_314, w_040_315, w_040_316, w_040_317, w_040_318, w_040_319, w_040_320, w_040_321, w_040_322, w_040_323, w_040_324, w_040_325, w_040_327, w_040_329, w_040_330, w_040_332, w_040_333, w_040_334, w_040_335, w_040_336, w_040_337, w_040_340, w_040_341, w_040_343, w_040_344, w_040_345, w_040_346, w_040_347, w_040_348, w_040_349, w_040_350, w_040_351, w_040_352, w_040_353, w_040_354, w_040_356, w_040_357, w_040_358, w_040_359, w_040_361, w_040_362, w_040_363, w_040_366, w_040_367, w_040_368, w_040_369, w_040_370, w_040_372, w_040_373, w_040_374, w_040_375, w_040_376, w_040_377, w_040_378, w_040_379, w_040_380, w_040_381, w_040_384, w_040_385, w_040_386, w_040_387, w_040_388, w_040_390, w_040_391, w_040_392, w_040_393, w_040_394, w_040_395, w_040_396, w_040_397, w_040_398, w_040_399, w_040_400, w_040_401, w_040_402, w_040_403, w_040_404, w_040_405, w_040_406, w_040_407, w_040_408, w_040_409, w_040_410, w_040_411, w_040_412, w_040_413, w_040_414, w_040_415, w_040_416, w_040_417, w_040_419, w_040_420, w_040_421, w_040_422, w_040_424, w_040_425, w_040_426, w_040_427, w_040_428, w_040_429, w_040_430, w_040_433, w_040_436, w_040_437, w_040_438, w_040_439, w_040_441, w_040_442, w_040_443, w_040_444, w_040_445, w_040_446, w_040_447, w_040_448, w_040_449, w_040_450, w_040_451, w_040_452, w_040_454, w_040_456, w_040_458, w_040_459, w_040_460, w_040_462, w_040_463, w_040_465, w_040_466, w_040_467, w_040_468, w_040_469, w_040_471, w_040_472, w_040_473, w_040_474, w_040_475, w_040_476, w_040_477, w_040_478, w_040_479, w_040_480, w_040_481, w_040_482, w_040_483, w_040_484, w_040_485, w_040_486, w_040_487, w_040_488, w_040_489, w_040_490, w_040_491, w_040_492, w_040_493, w_040_495, w_040_496, w_040_497, w_040_498, w_040_499, w_040_501, w_040_502, w_040_503, w_040_504, w_040_505, w_040_506, w_040_507, w_040_508, w_040_509, w_040_511, w_040_512, w_040_513, w_040_514, w_040_516, w_040_517, w_040_518, w_040_520, w_040_521, w_040_522, w_040_523, w_040_524, w_040_525, w_040_526, w_040_527, w_040_528, w_040_530, w_040_531, w_040_533, w_040_534, w_040_535, w_040_536, w_040_537, w_040_538, w_040_539, w_040_540, w_040_541, w_040_543, w_040_544, w_040_545, w_040_546, w_040_547, w_040_548, w_040_549, w_040_550, w_040_553, w_040_554, w_040_555, w_040_556, w_040_557, w_040_558, w_040_559, w_040_560, w_040_561, w_040_563, w_040_565, w_040_566, w_040_567, w_040_568, w_040_569, w_040_571, w_040_572, w_040_573, w_040_575, w_040_576, w_040_577, w_040_578, w_040_579, w_040_580, w_040_581, w_040_582, w_040_583, w_040_585, w_040_586, w_040_587, w_040_588, w_040_590, w_040_591, w_040_592, w_040_593, w_040_595, w_040_596, w_040_597, w_040_599, w_040_600, w_040_601, w_040_602, w_040_603, w_040_604, w_040_605, w_040_606, w_040_607, w_040_609, w_040_610, w_040_611, w_040_612, w_040_613, w_040_614, w_040_615, w_040_616, w_040_617, w_040_618, w_040_619, w_040_620, w_040_621, w_040_624, w_040_625, w_040_626, w_040_627, w_040_628, w_040_629, w_040_630, w_040_631, w_040_632, w_040_633, w_040_634, w_040_635, w_040_636, w_040_637, w_040_638, w_040_639, w_040_640, w_040_641, w_040_642, w_040_644, w_040_646, w_040_647, w_040_648, w_040_649, w_040_650, w_040_651, w_040_652, w_040_653, w_040_654, w_040_655, w_040_656, w_040_658, w_040_660, w_040_661, w_040_662, w_040_664, w_040_665, w_040_666, w_040_667, w_040_668, w_040_669, w_040_671, w_040_672, w_040_673, w_040_674, w_040_676, w_040_677, w_040_678, w_040_679, w_040_680, w_040_681, w_040_682, w_040_683, w_040_685, w_040_686, w_040_687, w_040_688, w_040_689, w_040_690, w_040_691, w_040_692, w_040_693, w_040_694, w_040_695, w_040_696, w_040_697, w_040_698, w_040_699, w_040_701, w_040_702, w_040_703, w_040_704, w_040_705, w_040_706, w_040_707, w_040_708, w_040_709, w_040_710, w_040_712, w_040_713, w_040_715, w_040_716, w_040_717, w_040_718, w_040_719, w_040_720, w_040_721, w_040_722, w_040_723, w_040_724, w_040_725, w_040_726, w_040_727, w_040_728, w_040_729, w_040_730, w_040_731, w_040_732, w_040_733, w_040_734, w_040_735, w_040_736, w_040_737, w_040_738, w_040_739, w_040_740, w_040_741, w_040_742, w_040_744, w_040_746, w_040_747, w_040_748, w_040_749, w_040_751, w_040_752, w_040_753, w_040_754, w_040_755, w_040_756, w_040_757, w_040_758, w_040_759, w_040_760, w_040_761, w_040_762, w_040_763, w_040_765, w_040_766, w_040_767, w_040_768, w_040_769, w_040_770, w_040_771, w_040_773, w_040_774, w_040_776, w_040_777, w_040_778, w_040_779, w_040_780, w_040_781, w_040_782, w_040_783, w_040_784, w_040_786, w_040_788, w_040_789, w_040_790, w_040_791, w_040_792, w_040_793, w_040_794, w_040_795, w_040_796, w_040_797, w_040_798, w_040_799, w_040_800, w_040_801, w_040_802, w_040_803, w_040_804, w_040_805, w_040_806, w_040_807, w_040_808, w_040_809, w_040_810, w_040_811, w_040_813, w_040_814, w_040_815, w_040_816, w_040_817, w_040_818, w_040_819, w_040_820, w_040_821, w_040_822, w_040_823, w_040_824, w_040_826, w_040_827, w_040_828, w_040_829, w_040_830, w_040_831, w_040_832, w_040_833, w_040_834, w_040_835, w_040_836, w_040_838, w_040_839, w_040_840, w_040_842, w_040_846, w_040_847, w_040_848, w_040_849, w_040_850, w_040_853, w_040_854, w_040_855, w_040_856, w_040_857, w_040_858, w_040_859, w_040_860, w_040_861, w_040_862, w_040_863, w_040_864, w_040_865, w_040_867, w_040_868, w_040_869, w_040_870, w_040_872, w_040_873, w_040_875, w_040_876, w_040_877, w_040_878, w_040_879, w_040_880, w_040_881, w_040_884, w_040_885, w_040_886, w_040_887, w_040_888, w_040_889, w_040_890, w_040_891, w_040_892, w_040_893, w_040_894, w_040_895, w_040_896, w_040_897, w_040_899, w_040_900, w_040_901, w_040_902, w_040_903, w_040_905, w_040_906, w_040_907, w_040_908, w_040_909, w_040_910, w_040_911, w_040_912, w_040_913, w_040_914, w_040_915, w_040_916, w_040_917, w_040_918, w_040_919, w_040_920, w_040_921, w_040_922, w_040_924, w_040_925, w_040_926, w_040_927, w_040_928, w_040_930, w_040_931, w_040_932, w_040_933, w_040_934, w_040_935, w_040_936, w_040_937, w_040_939, w_040_940, w_040_941, w_040_942, w_040_943, w_040_944, w_040_945, w_040_946, w_040_947, w_040_948, w_040_949, w_040_950, w_040_951, w_040_952, w_040_953, w_040_954, w_040_955, w_040_956, w_040_957, w_040_958, w_040_959, w_040_960, w_040_961, w_040_962, w_040_963, w_040_966, w_040_967, w_040_968, w_040_969, w_040_970, w_040_971, w_040_973, w_040_974, w_040_975, w_040_976, w_040_977, w_040_978, w_040_979, w_040_981, w_040_982, w_040_983, w_040_984, w_040_985, w_040_986, w_040_987, w_040_988, w_040_989, w_040_990, w_040_991, w_040_992, w_040_993, w_040_994, w_040_995, w_040_996, w_040_997, w_040_998, w_040_999, w_040_1000, w_040_1001, w_040_1002, w_040_1003, w_040_1004, w_040_1005, w_040_1006, w_040_1007, w_040_1008, w_040_1010, w_040_1011, w_040_1012, w_040_1013, w_040_1014, w_040_1015, w_040_1016, w_040_1018, w_040_1019, w_040_1020, w_040_1021, w_040_1022, w_040_1023, w_040_1024, w_040_1025, w_040_1026, w_040_1027, w_040_1028, w_040_1029, w_040_1031, w_040_1032, w_040_1033, w_040_1035, w_040_1036, w_040_1037, w_040_1038, w_040_1039, w_040_1040, w_040_1042, w_040_1043, w_040_1044, w_040_1045, w_040_1046, w_040_1048, w_040_1049, w_040_1051, w_040_1052, w_040_1053, w_040_1054, w_040_1055, w_040_1056, w_040_1057, w_040_1058, w_040_1059, w_040_1060, w_040_1061, w_040_1062, w_040_1063, w_040_1064, w_040_1065, w_040_1066, w_040_1067, w_040_1068, w_040_1069, w_040_1070, w_040_1071, w_040_1072, w_040_1073, w_040_1074, w_040_1077, w_040_1079, w_040_1080, w_040_1081, w_040_1083, w_040_1084, w_040_1085, w_040_1086, w_040_1087, w_040_1088, w_040_1090, w_040_1091, w_040_1092, w_040_1093, w_040_1094, w_040_1095, w_040_1096, w_040_1098, w_040_1099, w_040_1100, w_040_1101, w_040_1103, w_040_1104, w_040_1105, w_040_1106, w_040_1107, w_040_1108, w_040_1110, w_040_1111, w_040_1112, w_040_1113, w_040_1116, w_040_1117, w_040_1118, w_040_1119, w_040_1120, w_040_1121, w_040_1123, w_040_1125, w_040_1127, w_040_1128, w_040_1129, w_040_1130, w_040_1131, w_040_1132, w_040_1133, w_040_1134, w_040_1135, w_040_1137, w_040_1138, w_040_1139, w_040_1141, w_040_1142, w_040_1143, w_040_1144, w_040_1145, w_040_1146, w_040_1147, w_040_1148, w_040_1149, w_040_1150, w_040_1151, w_040_1152, w_040_1153, w_040_1154, w_040_1155, w_040_1156, w_040_1157, w_040_1158, w_040_1159, w_040_1160, w_040_1161, w_040_1162, w_040_1163, w_040_1164, w_040_1165, w_040_1166, w_040_1169, w_040_1170, w_040_1171, w_040_1172, w_040_1173, w_040_1174, w_040_1175, w_040_1176, w_040_1177, w_040_1178, w_040_1179, w_040_1180, w_040_1181, w_040_1182, w_040_1184, w_040_1185, w_040_1188, w_040_1189, w_040_1190, w_040_1191, w_040_1192, w_040_1193, w_040_1197, w_040_1199, w_040_1200, w_040_1201, w_040_1202, w_040_1203, w_040_1204, w_040_1205, w_040_1206, w_040_1207, w_040_1208, w_040_1209, w_040_1211, w_040_1212, w_040_1213, w_040_1214, w_040_1215, w_040_1216, w_040_1217, w_040_1218, w_040_1219, w_040_1220, w_040_1221, w_040_1222, w_040_1223, w_040_1224, w_040_1225, w_040_1226, w_040_1227, w_040_1228, w_040_1230, w_040_1231, w_040_1232, w_040_1233, w_040_1234, w_040_1235, w_040_1236, w_040_1237, w_040_1238, w_040_1239, w_040_1240, w_040_1241, w_040_1243, w_040_1245, w_040_1247, w_040_1248, w_040_1249, w_040_1250, w_040_1251, w_040_1252, w_040_1253, w_040_1255, w_040_1256, w_040_1258, w_040_1259, w_040_1260, w_040_1261, w_040_1262, w_040_1263, w_040_1264, w_040_1265, w_040_1267, w_040_1268, w_040_1269, w_040_1271, w_040_1272, w_040_1273, w_040_1274, w_040_1275, w_040_1276, w_040_1278, w_040_1279, w_040_1280, w_040_1282, w_040_1283, w_040_1284, w_040_1285, w_040_1286, w_040_1287, w_040_1288, w_040_1289, w_040_1291, w_040_1292, w_040_1293, w_040_1294, w_040_1295, w_040_1296, w_040_1297, w_040_1298, w_040_1299, w_040_1300, w_040_1301, w_040_1303, w_040_1304, w_040_1305, w_040_1306, w_040_1307, w_040_1308, w_040_1309, w_040_1310, w_040_1311, w_040_1312, w_040_1313, w_040_1314, w_040_1315, w_040_1316, w_040_1317, w_040_1318, w_040_1319, w_040_1320, w_040_1321, w_040_1322, w_040_1323, w_040_1324, w_040_1325, w_040_1326, w_040_1327, w_040_1328, w_040_1329, w_040_1330, w_040_1331, w_040_1332, w_040_1333, w_040_1335, w_040_1336, w_040_1337, w_040_1338, w_040_1339, w_040_1340, w_040_1341, w_040_1342, w_040_1345, w_040_1346, w_040_1348, w_040_1350, w_040_1351, w_040_1353, w_040_1354, w_040_1355, w_040_1356, w_040_1358, w_040_1360, w_040_1361, w_040_1362, w_040_1363, w_040_1364, w_040_1365, w_040_1366, w_040_1367, w_040_1368, w_040_1369, w_040_1370, w_040_1371, w_040_1372, w_040_1373, w_040_1374, w_040_1377, w_040_1378, w_040_1379, w_040_1380, w_040_1382, w_040_1384, w_040_1385, w_040_1386, w_040_1387, w_040_1388, w_040_1389, w_040_1390, w_040_1391, w_040_1392, w_040_1393, w_040_1394, w_040_1395, w_040_1396, w_040_1397, w_040_1398, w_040_1399, w_040_1400, w_040_1401, w_040_1402, w_040_1403, w_040_1404, w_040_1405, w_040_1406, w_040_1408, w_040_1409, w_040_1410, w_040_1411, w_040_1412, w_040_1414, w_040_1415, w_040_1416, w_040_1417, w_040_1418, w_040_1419, w_040_1420, w_040_1421, w_040_1422, w_040_1423, w_040_1425, w_040_1426, w_040_1427, w_040_1428, w_040_1429, w_040_1431, w_040_1432, w_040_1433, w_040_1434, w_040_1435, w_040_1436, w_040_1437, w_040_1438, w_040_1439, w_040_1440, w_040_1441, w_040_1442, w_040_1443, w_040_1444, w_040_1445, w_040_1447, w_040_1448, w_040_1450, w_040_1451, w_040_1452, w_040_1453, w_040_1454, w_040_1455, w_040_1456, w_040_1457, w_040_1458, w_040_1459, w_040_1460, w_040_1462, w_040_1463, w_040_1464, w_040_1465, w_040_1466, w_040_1467, w_040_1468, w_040_1469, w_040_1470, w_040_1472, w_040_1473, w_040_1474, w_040_1475, w_040_1476, w_040_1477, w_040_1479, w_040_1480, w_040_1481, w_040_1482, w_040_1483, w_040_1484, w_040_1485, w_040_1487, w_040_1488, w_040_1489, w_040_1490, w_040_1491, w_040_1492, w_040_1493, w_040_1494, w_040_1495, w_040_1496, w_040_1497, w_040_1498, w_040_1500, w_040_1501, w_040_1502, w_040_1503, w_040_1504, w_040_1505, w_040_1507, w_040_1508, w_040_1509, w_040_1511, w_040_1512, w_040_1513, w_040_1517, w_040_1518, w_040_1520, w_040_1521, w_040_1522, w_040_1523, w_040_1524, w_040_1525, w_040_1526, w_040_1527, w_040_1528, w_040_1530, w_040_1531, w_040_1532, w_040_1533, w_040_1534, w_040_1535, w_040_1536, w_040_1537, w_040_1538, w_040_1539, w_040_1541, w_040_1542, w_040_1543, w_040_1544, w_040_1546, w_040_1547, w_040_1548, w_040_1549, w_040_1550, w_040_1551, w_040_1552, w_040_1553, w_040_1555, w_040_1556, w_040_1557, w_040_1558, w_040_1559, w_040_1560, w_040_1562, w_040_1563, w_040_1564, w_040_1565, w_040_1566, w_040_1567, w_040_1568, w_040_1569, w_040_1571, w_040_1572, w_040_1573, w_040_1574, w_040_1575, w_040_1576, w_040_1577, w_040_1578, w_040_1579, w_040_1580, w_040_1581, w_040_1582, w_040_1583, w_040_1584, w_040_1587, w_040_1588, w_040_1589, w_040_1590, w_040_1591, w_040_1592, w_040_1593, w_040_1595, w_040_1596, w_040_1597, w_040_1598, w_040_1599, w_040_1600, w_040_1601, w_040_1602, w_040_1603, w_040_1604, w_040_1605, w_040_1606, w_040_1607, w_040_1608, w_040_1609, w_040_1612, w_040_1613, w_040_1615, w_040_1616, w_040_1617, w_040_1618, w_040_1619, w_040_1620, w_040_1621, w_040_1622, w_040_1623, w_040_1624, w_040_1625, w_040_1626, w_040_1627, w_040_1628, w_040_1631, w_040_1633, w_040_1634, w_040_1635, w_040_1636, w_040_1637, w_040_1638, w_040_1640, w_040_1641, w_040_1642, w_040_1643, w_040_1644, w_040_1645, w_040_1646, w_040_1647, w_040_1648, w_040_1649, w_040_1650, w_040_1652, w_040_1653, w_040_1654, w_040_1655, w_040_1656, w_040_1657, w_040_1658, w_040_1660, w_040_1661, w_040_1663, w_040_1664, w_040_1665, w_040_1666, w_040_1667, w_040_1668, w_040_1670, w_040_1671, w_040_1672, w_040_1673, w_040_1674, w_040_1675, w_040_1676, w_040_1677, w_040_1678, w_040_1679, w_040_1680, w_040_1681, w_040_1682, w_040_1685, w_040_1686, w_040_1687, w_040_1688, w_040_1689, w_040_1690, w_040_1691, w_040_1692, w_040_1693, w_040_1694, w_040_1695, w_040_1696, w_040_1698, w_040_1699, w_040_1701, w_040_1702, w_040_1703, w_040_1704, w_040_1706, w_040_1708, w_040_1709, w_040_1710, w_040_1711, w_040_1712, w_040_1713, w_040_1714, w_040_1715, w_040_1716, w_040_1717, w_040_1718, w_040_1719, w_040_1720, w_040_1722, w_040_1723, w_040_1724, w_040_1725, w_040_1726, w_040_1727, w_040_1728, w_040_1730, w_040_1731, w_040_1732, w_040_1734, w_040_1735, w_040_1736, w_040_1738, w_040_1740, w_040_1741, w_040_1742, w_040_1743, w_040_1744, w_040_1745, w_040_1746, w_040_1747, w_040_1748, w_040_1749, w_040_1751, w_040_1752, w_040_1753, w_040_1754, w_040_1755, w_040_1756, w_040_1757, w_040_1758, w_040_1760, w_040_1762, w_040_1764, w_040_1765, w_040_1766, w_040_1767, w_040_1768, w_040_1769, w_040_1770, w_040_1771, w_040_1772, w_040_1773, w_040_1774, w_040_1776, w_040_1778, w_040_1779, w_040_1780, w_040_1781, w_040_1782, w_040_1784, w_040_1786, w_040_1787, w_040_1789, w_040_1790, w_040_1791, w_040_1792, w_040_1793, w_040_1794, w_040_1795, w_040_1796, w_040_1799, w_040_1800, w_040_1801, w_040_1802, w_040_1804, w_040_1805, w_040_1806, w_040_1807, w_040_1809, w_040_1812, w_040_1814, w_040_1815, w_040_1816, w_040_1817, w_040_1818, w_040_1819, w_040_1820, w_040_1821, w_040_1822, w_040_1823, w_040_1824, w_040_1825, w_040_1826, w_040_1828, w_040_1829, w_040_1831, w_040_1832, w_040_1833, w_040_1834, w_040_1835, w_040_1836, w_040_1837, w_040_1838, w_040_1839, w_040_1840, w_040_1841, w_040_1842, w_040_1843, w_040_1844, w_040_1845, w_040_1846, w_040_1847, w_040_1848, w_040_1849, w_040_1850, w_040_1851, w_040_1852, w_040_1853, w_040_1854, w_040_1855, w_040_1856, w_040_1857, w_040_1858, w_040_1859, w_040_1860, w_040_1861, w_040_1863, w_040_1864, w_040_1865, w_040_1866, w_040_1867, w_040_1868, w_040_1869, w_040_1870, w_040_1872, w_040_1874, w_040_1875, w_040_1876, w_040_1877, w_040_1878, w_040_1879, w_040_1880, w_040_1881, w_040_1882, w_040_1883, w_040_1884, w_040_1885, w_040_1886, w_040_1887, w_040_1888, w_040_1889, w_040_1890, w_040_1891, w_040_1892, w_040_1893, w_040_1894, w_040_1895, w_040_1896, w_040_1897, w_040_1898, w_040_1900, w_040_1901, w_040_1903, w_040_1904, w_040_1905, w_040_1907, w_040_1910, w_040_1911, w_040_1913, w_040_1914, w_040_1916, w_040_1917, w_040_1918, w_040_1919, w_040_1920, w_040_1921, w_040_1922, w_040_1923, w_040_1924, w_040_1925, w_040_1926, w_040_1927, w_040_1928, w_040_1929, w_040_1932, w_040_1933, w_040_1934, w_040_1935, w_040_1936, w_040_1937, w_040_1939, w_040_1940, w_040_1941, w_040_1942, w_040_1943, w_040_1946, w_040_1947, w_040_1948, w_040_1949, w_040_1951, w_040_1952, w_040_1953, w_040_1954, w_040_1955, w_040_1956, w_040_1957, w_040_1958, w_040_1959, w_040_1960, w_040_1961, w_040_1962, w_040_1963, w_040_1964, w_040_1965, w_040_1966, w_040_1967, w_040_1968, w_040_1969, w_040_1970, w_040_1971, w_040_1972, w_040_1973, w_040_1975, w_040_1976, w_040_1977, w_040_1979, w_040_1980, w_040_1981, w_040_1982, w_040_1983, w_040_1984, w_040_1985, w_040_1987, w_040_1988, w_040_1989, w_040_1990, w_040_1991, w_040_1992, w_040_1993, w_040_1994, w_040_1995, w_040_1996, w_040_1997, w_040_1999, w_040_2001, w_040_2002, w_040_2003, w_040_2004, w_040_2005, w_040_2006, w_040_2008, w_040_2011, w_040_2012, w_040_2013, w_040_2014, w_040_2015, w_040_2016, w_040_2017, w_040_2018, w_040_2019, w_040_2020, w_040_2021, w_040_2022, w_040_2023, w_040_2024, w_040_2025, w_040_2026, w_040_2027, w_040_2028, w_040_2029, w_040_2030, w_040_2031, w_040_2033, w_040_2034, w_040_2035, w_040_2036, w_040_2038, w_040_2039, w_040_2040, w_040_2041, w_040_2043, w_040_2044, w_040_2045, w_040_2047, w_040_2048, w_040_2049, w_040_2050, w_040_2051, w_040_2053, w_040_2054, w_040_2056, w_040_2058, w_040_2060, w_040_2061, w_040_2063, w_040_2064, w_040_2065, w_040_2067, w_040_2068, w_040_2069, w_040_2070, w_040_2071, w_040_2073, w_040_2074, w_040_2075, w_040_2076, w_040_2077, w_040_2078, w_040_2079, w_040_2080, w_040_2081, w_040_2082, w_040_2083, w_040_2084, w_040_2085, w_040_2086, w_040_2087, w_040_2089, w_040_2090, w_040_2091, w_040_2093, w_040_2094, w_040_2095, w_040_2096, w_040_2099, w_040_2100, w_040_2102, w_040_2103, w_040_2104, w_040_2105, w_040_2106, w_040_2107, w_040_2110, w_040_2111, w_040_2112, w_040_2113, w_040_2114, w_040_2115, w_040_2116, w_040_2118, w_040_2119, w_040_2120, w_040_2121, w_040_2122, w_040_2123, w_040_2124, w_040_2125, w_040_2126, w_040_2127, w_040_2129, w_040_2130, w_040_2131, w_040_2132, w_040_2135, w_040_2137, w_040_2138, w_040_2140, w_040_2141, w_040_2143, w_040_2144, w_040_2145, w_040_2146, w_040_2147, w_040_2148, w_040_2149, w_040_2150, w_040_2153, w_040_2154, w_040_2155, w_040_2156, w_040_2158, w_040_2159, w_040_2160, w_040_2161, w_040_2162, w_040_2163, w_040_2165, w_040_2166, w_040_2167, w_040_2168, w_040_2169, w_040_2170, w_040_2171, w_040_2172, w_040_2173, w_040_2174, w_040_2175, w_040_2177, w_040_2178, w_040_2179, w_040_2181, w_040_2182, w_040_2183, w_040_2184, w_040_2187, w_040_2188, w_040_2189, w_040_2191, w_040_2192, w_040_2193, w_040_2195, w_040_2196, w_040_2197, w_040_2198, w_040_2199, w_040_2200, w_040_2201, w_040_2202, w_040_2203, w_040_2204, w_040_2205, w_040_2206, w_040_2207, w_040_2208, w_040_2209, w_040_2210, w_040_2211, w_040_2212, w_040_2213, w_040_2214, w_040_2215, w_040_2216, w_040_2217, w_040_2218, w_040_2219, w_040_2220, w_040_2221, w_040_2222, w_040_2223, w_040_2224, w_040_2225, w_040_2226, w_040_2227, w_040_2228, w_040_2229, w_040_2230, w_040_2231, w_040_2232, w_040_2233, w_040_2234, w_040_2235, w_040_2236, w_040_2237, w_040_2238, w_040_2240, w_040_2241, w_040_2242, w_040_2243, w_040_2245, w_040_2246, w_040_2247, w_040_2248, w_040_2249, w_040_2250, w_040_2251, w_040_2252, w_040_2254, w_040_2255, w_040_2256, w_040_2257, w_040_2258, w_040_2259, w_040_2261, w_040_2262, w_040_2263, w_040_2265, w_040_2267, w_040_2268, w_040_2269, w_040_2271, w_040_2273, w_040_2274, w_040_2275, w_040_2277, w_040_2278, w_040_2279, w_040_2280, w_040_2281, w_040_2282, w_040_2283, w_040_2284, w_040_2285, w_040_2286, w_040_2287, w_040_2289, w_040_2290, w_040_2291, w_040_2292, w_040_2293, w_040_2294, w_040_2295, w_040_2296, w_040_2297, w_040_2298, w_040_2299, w_040_2300, w_040_2301, w_040_2302, w_040_2303, w_040_2305, w_040_2306, w_040_2308, w_040_2309, w_040_2310, w_040_2311, w_040_2312, w_040_2313, w_040_2314, w_040_2316, w_040_2317, w_040_2318, w_040_2321, w_040_2323, w_040_2324, w_040_2325, w_040_2326, w_040_2327, w_040_2328, w_040_2329, w_040_2330, w_040_2331, w_040_2332, w_040_2333, w_040_2334, w_040_2335, w_040_2336, w_040_2337, w_040_2338, w_040_2339, w_040_2340, w_040_2341, w_040_2342, w_040_2343, w_040_2345, w_040_2346, w_040_2347, w_040_2349, w_040_2350, w_040_2351, w_040_2352, w_040_2353, w_040_2354, w_040_2355, w_040_2356, w_040_2357, w_040_2358, w_040_2359, w_040_2360, w_040_2364, w_040_2365, w_040_2366, w_040_2367, w_040_2368, w_040_2369, w_040_2370, w_040_2371, w_040_2373, w_040_2375, w_040_2376, w_040_2377, w_040_2378, w_040_2379, w_040_2380, w_040_2382, w_040_2383, w_040_2384, w_040_2385, w_040_2386, w_040_2387, w_040_2388, w_040_2389, w_040_2390, w_040_2391, w_040_2392, w_040_2393, w_040_2394, w_040_2395, w_040_2396, w_040_2397, w_040_2398, w_040_2401, w_040_2402, w_040_2403, w_040_2404, w_040_2405, w_040_2406, w_040_2407, w_040_2408, w_040_2409, w_040_2410, w_040_2412, w_040_2413, w_040_2414, w_040_2415, w_040_2416, w_040_2417, w_040_2418, w_040_2419, w_040_2420, w_040_2421, w_040_2422, w_040_2423, w_040_2424, w_040_2426, w_040_2427, w_040_2428, w_040_2429, w_040_2430, w_040_2431, w_040_2432, w_040_2434, w_040_2436, w_040_2438, w_040_2439, w_040_2440, w_040_2441, w_040_2442, w_040_2443, w_040_2444, w_040_2445, w_040_2446, w_040_2447, w_040_2448, w_040_2449, w_040_2450, w_040_2451, w_040_2452, w_040_2453, w_040_2456, w_040_2458, w_040_2459, w_040_2460, w_040_2461, w_040_2462, w_040_2464, w_040_2465, w_040_2466, w_040_2467, w_040_2468, w_040_2469, w_040_2470, w_040_2471, w_040_2472, w_040_2473, w_040_2474, w_040_2475, w_040_2478, w_040_2480, w_040_2481, w_040_2483, w_040_2485, w_040_2486, w_040_2487, w_040_2488, w_040_2489, w_040_2490, w_040_2491, w_040_2492, w_040_2493, w_040_2494, w_040_2495, w_040_2496, w_040_2498, w_040_2499, w_040_2500, w_040_2501, w_040_2502, w_040_2503, w_040_2504, w_040_2505, w_040_2506, w_040_2507, w_040_2508, w_040_2509, w_040_2513, w_040_2514, w_040_2515, w_040_2516, w_040_2517, w_040_2518, w_040_2519, w_040_2520, w_040_2521, w_040_2522, w_040_2523, w_040_2524, w_040_2526, w_040_2527, w_040_2528, w_040_2529, w_040_2530, w_040_2532, w_040_2533, w_040_2534, w_040_2535, w_040_2536, w_040_2537, w_040_2538, w_040_2539, w_040_2541, w_040_2542, w_040_2543, w_040_2544, w_040_2545, w_040_2546, w_040_2547, w_040_2548, w_040_2549, w_040_2550, w_040_2551, w_040_2552, w_040_2553, w_040_2554, w_040_2555, w_040_2556, w_040_2557, w_040_2559, w_040_2562, w_040_2563, w_040_2564, w_040_2565, w_040_2566, w_040_2567, w_040_2568, w_040_2569, w_040_2570, w_040_2571, w_040_2572, w_040_2573, w_040_2575, w_040_2576, w_040_2577, w_040_2578, w_040_2579, w_040_2580, w_040_2582, w_040_2583, w_040_2585, w_040_2586, w_040_2587, w_040_2588, w_040_2589, w_040_2590, w_040_2591, w_040_2592, w_040_2593, w_040_2594, w_040_2595, w_040_2596, w_040_2597, w_040_2601, w_040_2602, w_040_2603, w_040_2604, w_040_2606, w_040_2607, w_040_2608, w_040_2609, w_040_2610, w_040_2611, w_040_2612, w_040_2614, w_040_2615, w_040_2616, w_040_2619, w_040_2620, w_040_2621, w_040_2622, w_040_2624, w_040_2625, w_040_2626, w_040_2627, w_040_2628, w_040_2629, w_040_2630, w_040_2631, w_040_2632, w_040_2633, w_040_2634, w_040_2635, w_040_2637, w_040_2638, w_040_2639, w_040_2640, w_040_2641, w_040_2642, w_040_2643, w_040_2644, w_040_2645, w_040_2646, w_040_2647, w_040_2648, w_040_2649, w_040_2650, w_040_2652, w_040_2653, w_040_2654, w_040_2655, w_040_2656, w_040_2657, w_040_2658, w_040_2659, w_040_2661, w_040_2662, w_040_2663, w_040_2664, w_040_2667, w_040_2669, w_040_2670, w_040_2671, w_040_2672, w_040_2673, w_040_2674, w_040_2675, w_040_2676, w_040_2677, w_040_2678, w_040_2679, w_040_2680, w_040_2681, w_040_2682, w_040_2683, w_040_2684, w_040_2685, w_040_2686, w_040_2687, w_040_2688, w_040_2689, w_040_2690, w_040_2691, w_040_2693, w_040_2694, w_040_2695, w_040_2697, w_040_2698, w_040_2699, w_040_2701, w_040_2702, w_040_2704, w_040_2705, w_040_2706, w_040_2707, w_040_2708, w_040_2709, w_040_2710, w_040_2712, w_040_2713, w_040_2714, w_040_2715, w_040_2717, w_040_2718, w_040_2719, w_040_2720, w_040_2721, w_040_2722, w_040_2723, w_040_2724, w_040_2725, w_040_2726, w_040_2727, w_040_2728, w_040_2729, w_040_2731, w_040_2732, w_040_2733, w_040_2734, w_040_2736, w_040_2737, w_040_2738, w_040_2739, w_040_2740, w_040_2741, w_040_2742, w_040_2743, w_040_2744, w_040_2745, w_040_2746, w_040_2747, w_040_2748, w_040_2749, w_040_2750, w_040_2751, w_040_2753, w_040_2754, w_040_2755, w_040_2756, w_040_2758, w_040_2759, w_040_2761, w_040_2763, w_040_2764, w_040_2765, w_040_2766, w_040_2769, w_040_2770, w_040_2771, w_040_2772, w_040_2773, w_040_2775, w_040_2776, w_040_2777, w_040_2778, w_040_2780, w_040_2781, w_040_2782, w_040_2783, w_040_2784, w_040_2785, w_040_2786, w_040_2787, w_040_2788, w_040_2789, w_040_2790, w_040_2792, w_040_2793, w_040_2794, w_040_2795, w_040_2796, w_040_2797, w_040_2798, w_040_2799, w_040_2800, w_040_2801, w_040_2802, w_040_2803, w_040_2804, w_040_2805, w_040_2806, w_040_2808, w_040_2809, w_040_2810, w_040_2811, w_040_2812, w_040_2814, w_040_2815, w_040_2818, w_040_2819, w_040_2821, w_040_2822, w_040_2823, w_040_2825, w_040_2826, w_040_2827, w_040_2829, w_040_2830, w_040_2831, w_040_2832, w_040_2833, w_040_2834, w_040_2835, w_040_2837, w_040_2838, w_040_2840, w_040_2841, w_040_2842, w_040_2843, w_040_2844, w_040_2845, w_040_2846, w_040_2849, w_040_2851, w_040_2852, w_040_2853, w_040_2854, w_040_2855, w_040_2856, w_040_2857, w_040_2859, w_040_2861, w_040_2863, w_040_2864, w_040_2867, w_040_2868, w_040_2869, w_040_2872, w_040_2873, w_040_2875, w_040_2876, w_040_2877, w_040_2879, w_040_2880, w_040_2881, w_040_2882, w_040_2883, w_040_2884, w_040_2885, w_040_2886, w_040_2887, w_040_2888, w_040_2889, w_040_2890, w_040_2893, w_040_2894, w_040_2895, w_040_2896, w_040_2897, w_040_2898, w_040_2899, w_040_2901, w_040_2902, w_040_2903, w_040_2905, w_040_2906, w_040_2907, w_040_2909, w_040_2910, w_040_2911, w_040_2912, w_040_2913, w_040_2914, w_040_2915, w_040_2916, w_040_2917, w_040_2918, w_040_2920, w_040_2922, w_040_2923, w_040_2924, w_040_2926, w_040_2927, w_040_2928, w_040_2930, w_040_2931, w_040_2932, w_040_2933, w_040_2934, w_040_2936, w_040_2938, w_040_2939, w_040_2940, w_040_2941, w_040_2942, w_040_2943, w_040_2944, w_040_2946, w_040_2948, w_040_2949, w_040_2950, w_040_2951, w_040_2952, w_040_2953, w_040_2955, w_040_2957, w_040_2959, w_040_2960, w_040_2961, w_040_2962, w_040_2963, w_040_2964, w_040_2965, w_040_2966, w_040_2967, w_040_2972, w_040_2974, w_040_2975, w_040_2978, w_040_2979, w_040_2982, w_040_2983, w_040_2984, w_040_2985, w_040_2986, w_040_2988, w_040_2989, w_040_2990, w_040_2991, w_040_2992, w_040_2993, w_040_2995, w_040_2996, w_040_2997, w_040_2998, w_040_2999, w_040_3001, w_040_3002, w_040_3003, w_040_3004, w_040_3007, w_040_3008, w_040_3009, w_040_3010, w_040_3012, w_040_3013, w_040_3014, w_040_3016, w_040_3018, w_040_3019, w_040_3022, w_040_3023, w_040_3025, w_040_3026, w_040_3027, w_040_3029, w_040_3030, w_040_3031, w_040_3033, w_040_3035, w_040_3037, w_040_3039, w_040_3040, w_040_3041, w_040_3042, w_040_3045, w_040_3046, w_040_3047, w_040_3048, w_040_3049, w_040_3051, w_040_3052, w_040_3053, w_040_3054, w_040_3055, w_040_3056, w_040_3058, w_040_3059, w_040_3060, w_040_3061, w_040_3062, w_040_3063, w_040_3065, w_040_3071, w_040_3073, w_040_3074, w_040_3075, w_040_3077, w_040_3079, w_040_3080, w_040_3081, w_040_3082, w_040_3084, w_040_3086, w_040_3087, w_040_3088, w_040_3092, w_040_3093, w_040_3094, w_040_3095, w_040_3097, w_040_3099, w_040_3100, w_040_3102, w_040_3104, w_040_3105, w_040_3106, w_040_3107, w_040_3108, w_040_3109, w_040_3110, w_040_3111, w_040_3112, w_040_3118, w_040_3119, w_040_3120, w_040_3121, w_040_3122, w_040_3123, w_040_3124, w_040_3125, w_040_3127, w_040_3128, w_040_3129, w_040_3131, w_040_3132, w_040_3133, w_040_3135, w_040_3136, w_040_3137, w_040_3139, w_040_3140, w_040_3141, w_040_3144, w_040_3145, w_040_3146, w_040_3148, w_040_3149, w_040_3150, w_040_3151, w_040_3152, w_040_3154, w_040_3155, w_040_3156, w_040_3157, w_040_3159, w_040_3160, w_040_3161, w_040_3162, w_040_3165, w_040_3166, w_040_3167, w_040_3168, w_040_3170, w_040_3171, w_040_3174, w_040_3175, w_040_3176, w_040_3177, w_040_3178, w_040_3181, w_040_3182, w_040_3183, w_040_3184, w_040_3186, w_040_3190, w_040_3191, w_040_3193, w_040_3195, w_040_3196, w_040_3197, w_040_3198, w_040_3199, w_040_3200, w_040_3201, w_040_3203, w_040_3204, w_040_3205, w_040_3206, w_040_3207, w_040_3208, w_040_3210, w_040_3211, w_040_3213, w_040_3215, w_040_3216, w_040_3218, w_040_3219, w_040_3220, w_040_3221, w_040_3222, w_040_3224, w_040_3225, w_040_3226, w_040_3227, w_040_3228, w_040_3229, w_040_3230, w_040_3233, w_040_3234, w_040_3236, w_040_3237, w_040_3239, w_040_3240, w_040_3241, w_040_3243, w_040_3244, w_040_3245, w_040_3246, w_040_3248, w_040_3251, w_040_3252, w_040_3254, w_040_3255, w_040_3256, w_040_3257, w_040_3259, w_040_3260, w_040_3261, w_040_3262, w_040_3263, w_040_3264, w_040_3265, w_040_3267, w_040_3268, w_040_3269, w_040_3270, w_040_3271, w_040_3272, w_040_3273, w_040_3274, w_040_3275, w_040_3278, w_040_3279, w_040_3282, w_040_3285, w_040_3287, w_040_3289, w_040_3291, w_040_3292, w_040_3293, w_040_3294, w_040_3296, w_040_3298, w_040_3299, w_040_3300, w_040_3301, w_040_3302, w_040_3303, w_040_3304, w_040_3305, w_040_3306, w_040_3307, w_040_3308, w_040_3309, w_040_3310, w_040_3312, w_040_3313, w_040_3314, w_040_3318, w_040_3319, w_040_3320, w_040_3321, w_040_3322, w_040_3323, w_040_3324, w_040_3325, w_040_3326, w_040_3327, w_040_3328, w_040_3329, w_040_3330, w_040_3332, w_040_3333, w_040_3334, w_040_3335, w_040_3336, w_040_3337, w_040_3338, w_040_3339, w_040_3340, w_040_3341, w_040_3342, w_040_3343, w_040_3344, w_040_3346, w_040_3347, w_040_3348, w_040_3349, w_040_3350, w_040_3351, w_040_3352, w_040_3353, w_040_3354, w_040_3355, w_040_3356, w_040_3358, w_040_3359, w_040_3361, w_040_3362, w_040_3363, w_040_3365, w_040_3366, w_040_3367, w_040_3370, w_040_3371, w_040_3372, w_040_3373, w_040_3375, w_040_3376, w_040_3377, w_040_3378, w_040_3381, w_040_3382, w_040_3383, w_040_3385, w_040_3386, w_040_3387, w_040_3388, w_040_3389, w_040_3390, w_040_3391, w_040_3392, w_040_3395, w_040_3397, w_040_3399, w_040_3400, w_040_3401, w_040_3402, w_040_3404, w_040_3407, w_040_3409, w_040_3410, w_040_3415, w_040_3416, w_040_3417, w_040_3419, w_040_3420, w_040_3421, w_040_3422, w_040_3424, w_040_3425, w_040_3426, w_040_3427, w_040_3428, w_040_3429, w_040_3430, w_040_3432, w_040_3433, w_040_3435, w_040_3437, w_040_3439, w_040_3442, w_040_3443, w_040_3446, w_040_3447, w_040_3449, w_040_3450, w_040_3452, w_040_3454, w_040_3456, w_040_3457, w_040_3458, w_040_3459, w_040_3460, w_040_3461, w_040_3464, w_040_3465, w_040_3466, w_040_3467, w_040_3468, w_040_3469, w_040_3470, w_040_3471, w_040_3472, w_040_3473, w_040_3474, w_040_3476, w_040_3478, w_040_3479, w_040_3480, w_040_3482, w_040_3487, w_040_3488, w_040_3489, w_040_3491, w_040_3492, w_040_3494, w_040_3496, w_040_3498, w_040_3500, w_040_3502, w_040_3504, w_040_3506, w_040_3507, w_040_3508, w_040_3510, w_040_3512, w_040_3513, w_040_3515, w_040_3516, w_040_3518, w_040_3520, w_040_3521, w_040_3522, w_040_3523, w_040_3524, w_040_3525, w_040_3526, w_040_3527, w_040_3528, w_040_3529, w_040_3530, w_040_3531, w_040_3533, w_040_3534, w_040_3535, w_040_3536, w_040_3538, w_040_3539, w_040_3540, w_040_3541, w_040_3542, w_040_3543, w_040_3545, w_040_3546, w_040_3547, w_040_3548, w_040_3549, w_040_3550, w_040_3553, w_040_3554, w_040_3556, w_040_3557, w_040_3558, w_040_3561, w_040_3563, w_040_3564, w_040_3565, w_040_3566, w_040_3567, w_040_3568, w_040_3570, w_040_3571, w_040_3572, w_040_3573, w_040_3574, w_040_3575, w_040_3577, w_040_3578, w_040_3579, w_040_3580, w_040_3581, w_040_3582, w_040_3583, w_040_3585, w_040_3586, w_040_3588, w_040_3589, w_040_3590, w_040_3591, w_040_3593, w_040_3594, w_040_3596;
  wire w_041_001, w_041_002, w_041_003, w_041_004, w_041_005, w_041_006, w_041_007, w_041_008, w_041_009, w_041_010, w_041_012, w_041_013, w_041_014, w_041_015, w_041_016, w_041_018, w_041_019, w_041_020, w_041_021, w_041_022, w_041_023, w_041_024, w_041_025, w_041_027, w_041_028, w_041_029, w_041_031, w_041_032, w_041_033, w_041_036, w_041_037, w_041_038, w_041_039, w_041_040, w_041_041, w_041_042, w_041_043, w_041_044, w_041_045, w_041_046, w_041_047, w_041_049, w_041_051, w_041_052, w_041_053, w_041_055, w_041_056, w_041_057, w_041_058, w_041_059, w_041_060, w_041_061, w_041_062, w_041_063, w_041_064, w_041_065, w_041_066, w_041_067, w_041_068, w_041_069, w_041_070, w_041_071, w_041_072, w_041_073, w_041_074, w_041_077, w_041_078, w_041_080, w_041_081, w_041_082, w_041_083, w_041_084, w_041_085, w_041_086, w_041_087, w_041_088, w_041_089, w_041_090, w_041_091, w_041_092, w_041_094, w_041_095, w_041_096, w_041_097, w_041_098, w_041_099, w_041_100, w_041_104, w_041_105, w_041_106, w_041_107, w_041_108, w_041_110, w_041_111, w_041_113, w_041_114, w_041_115, w_041_116, w_041_117, w_041_118, w_041_119, w_041_120, w_041_121, w_041_122, w_041_123, w_041_124, w_041_125, w_041_126, w_041_127, w_041_128, w_041_129, w_041_130, w_041_131, w_041_132, w_041_133, w_041_134, w_041_135, w_041_136, w_041_137, w_041_139, w_041_140, w_041_141, w_041_142, w_041_143, w_041_144, w_041_146, w_041_147, w_041_148, w_041_149, w_041_150, w_041_152, w_041_153, w_041_154, w_041_155, w_041_156, w_041_157, w_041_158, w_041_159, w_041_160, w_041_162, w_041_163, w_041_164, w_041_165, w_041_166, w_041_168, w_041_169, w_041_170, w_041_171, w_041_172, w_041_176, w_041_177, w_041_178, w_041_179, w_041_180, w_041_182, w_041_183, w_041_184, w_041_185, w_041_186, w_041_187, w_041_188, w_041_189, w_041_190, w_041_191, w_041_192, w_041_195, w_041_196, w_041_197, w_041_198, w_041_199, w_041_200, w_041_202, w_041_203, w_041_204, w_041_205, w_041_206, w_041_208, w_041_210, w_041_213, w_041_214, w_041_215, w_041_218, w_041_219, w_041_220, w_041_221, w_041_223, w_041_224, w_041_225, w_041_226, w_041_227, w_041_228, w_041_229, w_041_231, w_041_232, w_041_233, w_041_235, w_041_236, w_041_237, w_041_238, w_041_239, w_041_240, w_041_242, w_041_243, w_041_244, w_041_245, w_041_246, w_041_247, w_041_248, w_041_249, w_041_250, w_041_251, w_041_253, w_041_254, w_041_255, w_041_256, w_041_257, w_041_258, w_041_259, w_041_260, w_041_261, w_041_262, w_041_264, w_041_265, w_041_266, w_041_267, w_041_268, w_041_269, w_041_271, w_041_273, w_041_274, w_041_275, w_041_276, w_041_277, w_041_278, w_041_279, w_041_280, w_041_281, w_041_283, w_041_284, w_041_285, w_041_286, w_041_287, w_041_288, w_041_289, w_041_290, w_041_291, w_041_292, w_041_293, w_041_294, w_041_295, w_041_296, w_041_297, w_041_298, w_041_299, w_041_300, w_041_301, w_041_302, w_041_303, w_041_304, w_041_305, w_041_306, w_041_307, w_041_308, w_041_309, w_041_310, w_041_312, w_041_313, w_041_316, w_041_317, w_041_318, w_041_319, w_041_321, w_041_324, w_041_325, w_041_326, w_041_327, w_041_328, w_041_330, w_041_331, w_041_332, w_041_333, w_041_334, w_041_335, w_041_336, w_041_337, w_041_338, w_041_339, w_041_340, w_041_341, w_041_342, w_041_343, w_041_345, w_041_348, w_041_349, w_041_350, w_041_351, w_041_352, w_041_354, w_041_355, w_041_356, w_041_357, w_041_358, w_041_359, w_041_360, w_041_361, w_041_363, w_041_364, w_041_365, w_041_366, w_041_367, w_041_368, w_041_369, w_041_370, w_041_372, w_041_373, w_041_376, w_041_379, w_041_380, w_041_381, w_041_383, w_041_384, w_041_385, w_041_386, w_041_387, w_041_388, w_041_389, w_041_390, w_041_391, w_041_393, w_041_394, w_041_395, w_041_396, w_041_397, w_041_398, w_041_399, w_041_400, w_041_401, w_041_402, w_041_403, w_041_404, w_041_405, w_041_406, w_041_407, w_041_408, w_041_409, w_041_410, w_041_411, w_041_412, w_041_413, w_041_414, w_041_415, w_041_416, w_041_417, w_041_418, w_041_419, w_041_420, w_041_421, w_041_422, w_041_423, w_041_424, w_041_425, w_041_426, w_041_427, w_041_428, w_041_429, w_041_430, w_041_431, w_041_432, w_041_433, w_041_434, w_041_435, w_041_436, w_041_438, w_041_440, w_041_442, w_041_443, w_041_444, w_041_445, w_041_446, w_041_447, w_041_449, w_041_450, w_041_452, w_041_453, w_041_454, w_041_455, w_041_456, w_041_457, w_041_458, w_041_459, w_041_460, w_041_461, w_041_462, w_041_463, w_041_464, w_041_465, w_041_466, w_041_467, w_041_469, w_041_471, w_041_472, w_041_473, w_041_474, w_041_475, w_041_476, w_041_479, w_041_480, w_041_481, w_041_482, w_041_483, w_041_484, w_041_485, w_041_486, w_041_487, w_041_488, w_041_489, w_041_490, w_041_491, w_041_492, w_041_493, w_041_494, w_041_495, w_041_496, w_041_497, w_041_498, w_041_499, w_041_501, w_041_503, w_041_504, w_041_505, w_041_507, w_041_508, w_041_510, w_041_511, w_041_514, w_041_515, w_041_516, w_041_517, w_041_518, w_041_519, w_041_520, w_041_521, w_041_522, w_041_523, w_041_524, w_041_525, w_041_526, w_041_527, w_041_529, w_041_530, w_041_531, w_041_532, w_041_533, w_041_534, w_041_535, w_041_536, w_041_537, w_041_539, w_041_540, w_041_541, w_041_544, w_041_546, w_041_547, w_041_548, w_041_549, w_041_550, w_041_552, w_041_553, w_041_554, w_041_556, w_041_558, w_041_559, w_041_560, w_041_561, w_041_562, w_041_563, w_041_564, w_041_565, w_041_567, w_041_568, w_041_569, w_041_570, w_041_572, w_041_573, w_041_574, w_041_575, w_041_576, w_041_577, w_041_578, w_041_579, w_041_580, w_041_581, w_041_582, w_041_585, w_041_586, w_041_588, w_041_589, w_041_590, w_041_591, w_041_592, w_041_593, w_041_594, w_041_595, w_041_596, w_041_597, w_041_598, w_041_600, w_041_601, w_041_602, w_041_603, w_041_604, w_041_606, w_041_608, w_041_609, w_041_610, w_041_611, w_041_612, w_041_613, w_041_615, w_041_616, w_041_617, w_041_618, w_041_619, w_041_620, w_041_621, w_041_622, w_041_623, w_041_625, w_041_626, w_041_627, w_041_628, w_041_629, w_041_630, w_041_631, w_041_632, w_041_633, w_041_634, w_041_635, w_041_636, w_041_637, w_041_638, w_041_639, w_041_640, w_041_641, w_041_642, w_041_643, w_041_644, w_041_645, w_041_646, w_041_647, w_041_648, w_041_649, w_041_650, w_041_651, w_041_652, w_041_653, w_041_654, w_041_655, w_041_656, w_041_657, w_041_658, w_041_659, w_041_660, w_041_661, w_041_663, w_041_664, w_041_665, w_041_667, w_041_668, w_041_669, w_041_670, w_041_671, w_041_672, w_041_673, w_041_674, w_041_675, w_041_676, w_041_677, w_041_678, w_041_679, w_041_680, w_041_681, w_041_682, w_041_683, w_041_684, w_041_685, w_041_686, w_041_687, w_041_688, w_041_689, w_041_690, w_041_691, w_041_692, w_041_693, w_041_694, w_041_695, w_041_696, w_041_697, w_041_698, w_041_699, w_041_700, w_041_701, w_041_702, w_041_703, w_041_705, w_041_708, w_041_709, w_041_710, w_041_711, w_041_712, w_041_713, w_041_714, w_041_716, w_041_720, w_041_721, w_041_722, w_041_723, w_041_724, w_041_725, w_041_726, w_041_727, w_041_728, w_041_730, w_041_731, w_041_732, w_041_733, w_041_734, w_041_735, w_041_736, w_041_737, w_041_738, w_041_741, w_041_742, w_041_743, w_041_744, w_041_746, w_041_748, w_041_749, w_041_750, w_041_752, w_041_753, w_041_754, w_041_756, w_041_757, w_041_758, w_041_759, w_041_760, w_041_761, w_041_762, w_041_763, w_041_764, w_041_765, w_041_766, w_041_767, w_041_768, w_041_769, w_041_773, w_041_774, w_041_775, w_041_776, w_041_777, w_041_778, w_041_779, w_041_780, w_041_781, w_041_783, w_041_784, w_041_785, w_041_787, w_041_788, w_041_789, w_041_790, w_041_791, w_041_793, w_041_796, w_041_797, w_041_798, w_041_799, w_041_800, w_041_801, w_041_802, w_041_803, w_041_804, w_041_805, w_041_806, w_041_807, w_041_808, w_041_810, w_041_811, w_041_812, w_041_813, w_041_815, w_041_816, w_041_817, w_041_818, w_041_819, w_041_820, w_041_821, w_041_823, w_041_824, w_041_825, w_041_826, w_041_827, w_041_828, w_041_829, w_041_830, w_041_831, w_041_832, w_041_833, w_041_834, w_041_836, w_041_838, w_041_839, w_041_840, w_041_841, w_041_842, w_041_843, w_041_844, w_041_845, w_041_846, w_041_847, w_041_850, w_041_852, w_041_853, w_041_854, w_041_855, w_041_856, w_041_857, w_041_858, w_041_859, w_041_861, w_041_862, w_041_863, w_041_864, w_041_865, w_041_867, w_041_868, w_041_869, w_041_870, w_041_871, w_041_872, w_041_874, w_041_875, w_041_877, w_041_878, w_041_879, w_041_880, w_041_881, w_041_883, w_041_884, w_041_885, w_041_886, w_041_887, w_041_889, w_041_891, w_041_892, w_041_893, w_041_894, w_041_895, w_041_896, w_041_897, w_041_898, w_041_899, w_041_901, w_041_902, w_041_903, w_041_904, w_041_905, w_041_910, w_041_911, w_041_912, w_041_913, w_041_914, w_041_915, w_041_916, w_041_917, w_041_918, w_041_920, w_041_921, w_041_922, w_041_923, w_041_926, w_041_927, w_041_928, w_041_929, w_041_930, w_041_931, w_041_932, w_041_933, w_041_934, w_041_935, w_041_936, w_041_937, w_041_938, w_041_939, w_041_940, w_041_944, w_041_945, w_041_946, w_041_947, w_041_948, w_041_949, w_041_951, w_041_952, w_041_953, w_041_954, w_041_955, w_041_956, w_041_957, w_041_958, w_041_959, w_041_960, w_041_961, w_041_962, w_041_963, w_041_964, w_041_965, w_041_966, w_041_967, w_041_968, w_041_969, w_041_970, w_041_971, w_041_972, w_041_973, w_041_974, w_041_975, w_041_976, w_041_977, w_041_978, w_041_979, w_041_980, w_041_981, w_041_983, w_041_985, w_041_986, w_041_987, w_041_988, w_041_989, w_041_990, w_041_992, w_041_993, w_041_994, w_041_995, w_041_996, w_041_997, w_041_1000, w_041_1001, w_041_1002, w_041_1003, w_041_1004, w_041_1005, w_041_1006, w_041_1007, w_041_1008, w_041_1009, w_041_1010, w_041_1011, w_041_1012, w_041_1013, w_041_1014, w_041_1015, w_041_1016, w_041_1017, w_041_1019, w_041_1020, w_041_1021, w_041_1022, w_041_1023, w_041_1024, w_041_1025, w_041_1026, w_041_1027, w_041_1028, w_041_1031, w_041_1032, w_041_1033, w_041_1034, w_041_1035, w_041_1036, w_041_1037, w_041_1038, w_041_1039, w_041_1040, w_041_1041, w_041_1042, w_041_1043, w_041_1044, w_041_1045, w_041_1046, w_041_1048, w_041_1049, w_041_1051, w_041_1052, w_041_1053, w_041_1054, w_041_1055, w_041_1056, w_041_1057, w_041_1058, w_041_1059, w_041_1060, w_041_1061, w_041_1062, w_041_1063, w_041_1064, w_041_1066, w_041_1067, w_041_1069, w_041_1070, w_041_1071, w_041_1072, w_041_1073, w_041_1074, w_041_1075, w_041_1076, w_041_1077, w_041_1078, w_041_1080, w_041_1082, w_041_1083, w_041_1084, w_041_1085, w_041_1086, w_041_1087, w_041_1088, w_041_1092, w_041_1093, w_041_1094, w_041_1095, w_041_1096, w_041_1097, w_041_1098, w_041_1099, w_041_1100, w_041_1101, w_041_1102, w_041_1103, w_041_1104, w_041_1105, w_041_1106, w_041_1107, w_041_1109, w_041_1110, w_041_1111, w_041_1112, w_041_1113, w_041_1114, w_041_1115, w_041_1116, w_041_1117, w_041_1119, w_041_1120, w_041_1121, w_041_1122, w_041_1123, w_041_1124, w_041_1125, w_041_1126, w_041_1127, w_041_1128, w_041_1129, w_041_1132, w_041_1133, w_041_1134, w_041_1136, w_041_1137, w_041_1138, w_041_1140, w_041_1141, w_041_1142, w_041_1143, w_041_1144, w_041_1145, w_041_1146, w_041_1147, w_041_1148, w_041_1149, w_041_1150, w_041_1151, w_041_1152, w_041_1153, w_041_1154, w_041_1155, w_041_1156, w_041_1157, w_041_1158, w_041_1159, w_041_1160, w_041_1161, w_041_1162, w_041_1163, w_041_1164, w_041_1165, w_041_1166, w_041_1167, w_041_1168, w_041_1170, w_041_1171, w_041_1173, w_041_1174, w_041_1175, w_041_1176, w_041_1177, w_041_1178, w_041_1179, w_041_1180, w_041_1181, w_041_1182, w_041_1183, w_041_1184, w_041_1187, w_041_1188, w_041_1189, w_041_1190, w_041_1192, w_041_1193, w_041_1194, w_041_1196, w_041_1198, w_041_1199, w_041_1200, w_041_1201, w_041_1202, w_041_1203, w_041_1204, w_041_1205, w_041_1206, w_041_1208, w_041_1209, w_041_1210, w_041_1211, w_041_1212, w_041_1213, w_041_1214, w_041_1215, w_041_1216, w_041_1217, w_041_1218, w_041_1219, w_041_1220, w_041_1221, w_041_1222, w_041_1223, w_041_1224, w_041_1226, w_041_1227, w_041_1228, w_041_1230, w_041_1231, w_041_1233, w_041_1234, w_041_1236, w_041_1237, w_041_1238, w_041_1239, w_041_1240, w_041_1241, w_041_1242, w_041_1243, w_041_1245, w_041_1247, w_041_1248, w_041_1249, w_041_1250, w_041_1251, w_041_1252, w_041_1253, w_041_1254, w_041_1255, w_041_1257, w_041_1258, w_041_1259, w_041_1261, w_041_1262, w_041_1263, w_041_1265, w_041_1266, w_041_1267, w_041_1268, w_041_1269, w_041_1270, w_041_1271, w_041_1272, w_041_1273, w_041_1274, w_041_1275, w_041_1276, w_041_1279, w_041_1280, w_041_1281, w_041_1282, w_041_1283, w_041_1284, w_041_1285, w_041_1286, w_041_1287, w_041_1288, w_041_1289, w_041_1290, w_041_1292, w_041_1293, w_041_1294, w_041_1295, w_041_1296, w_041_1297, w_041_1298, w_041_1299, w_041_1300, w_041_1301, w_041_1302, w_041_1303, w_041_1304, w_041_1305, w_041_1306, w_041_1307, w_041_1308, w_041_1309, w_041_1310, w_041_1311, w_041_1312, w_041_1314, w_041_1315, w_041_1316, w_041_1317, w_041_1320, w_041_1321, w_041_1322, w_041_1323, w_041_1324, w_041_1325, w_041_1326, w_041_1327, w_041_1328, w_041_1329, w_041_1330, w_041_1331, w_041_1332, w_041_1333, w_041_1334, w_041_1336, w_041_1337, w_041_1338, w_041_1339, w_041_1340, w_041_1341, w_041_1342, w_041_1343, w_041_1344, w_041_1345, w_041_1349, w_041_1350, w_041_1351, w_041_1353, w_041_1354, w_041_1355, w_041_1356, w_041_1358, w_041_1359, w_041_1360, w_041_1361, w_041_1363, w_041_1364, w_041_1365, w_041_1366, w_041_1367, w_041_1368, w_041_1369, w_041_1370, w_041_1371, w_041_1372, w_041_1373, w_041_1374, w_041_1375, w_041_1377, w_041_1379, w_041_1380, w_041_1384, w_041_1385, w_041_1386, w_041_1387, w_041_1388, w_041_1389, w_041_1390, w_041_1391, w_041_1392, w_041_1393, w_041_1394, w_041_1395, w_041_1396, w_041_1397, w_041_1398, w_041_1399, w_041_1400, w_041_1401, w_041_1402, w_041_1403, w_041_1405, w_041_1406, w_041_1407, w_041_1408, w_041_1409, w_041_1410, w_041_1411, w_041_1412, w_041_1413, w_041_1414, w_041_1416, w_041_1417, w_041_1419, w_041_1420, w_041_1421, w_041_1422, w_041_1423, w_041_1424, w_041_1425, w_041_1426, w_041_1427, w_041_1428, w_041_1429, w_041_1430, w_041_1431, w_041_1432, w_041_1433, w_041_1434, w_041_1436, w_041_1437, w_041_1438, w_041_1440, w_041_1441, w_041_1442, w_041_1443, w_041_1445, w_041_1446, w_041_1448, w_041_1449, w_041_1450, w_041_1451, w_041_1453, w_041_1454, w_041_1455, w_041_1457, w_041_1458, w_041_1459, w_041_1460, w_041_1461, w_041_1462, w_041_1463, w_041_1464, w_041_1465, w_041_1466, w_041_1467, w_041_1468, w_041_1469, w_041_1470, w_041_1471, w_041_1472, w_041_1473, w_041_1474, w_041_1476, w_041_1479, w_041_1480, w_041_1481, w_041_1482, w_041_1483, w_041_1484, w_041_1485, w_041_1486, w_041_1487, w_041_1488, w_041_1489, w_041_1490, w_041_1491, w_041_1493, w_041_1494, w_041_1496, w_041_1498, w_041_1499, w_041_1500, w_041_1501, w_041_1502, w_041_1503, w_041_1504, w_041_1505, w_041_1506, w_041_1507, w_041_1509, w_041_1510, w_041_1511, w_041_1512, w_041_1513, w_041_1514, w_041_1515, w_041_1518, w_041_1520, w_041_1521, w_041_1522, w_041_1523, w_041_1524, w_041_1525, w_041_1526, w_041_1527, w_041_1528, w_041_1529, w_041_1530, w_041_1531, w_041_1533, w_041_1534, w_041_1536, w_041_1537, w_041_1538, w_041_1539, w_041_1540, w_041_1541, w_041_1542, w_041_1543, w_041_1544, w_041_1545, w_041_1547, w_041_1549, w_041_1551, w_041_1552, w_041_1553, w_041_1554, w_041_1555, w_041_1556, w_041_1557, w_041_1558, w_041_1559, w_041_1562, w_041_1563, w_041_1564, w_041_1565, w_041_1566, w_041_1567, w_041_1569, w_041_1570, w_041_1571, w_041_1572, w_041_1573, w_041_1574, w_041_1575, w_041_1576, w_041_1578, w_041_1579, w_041_1580, w_041_1581, w_041_1582, w_041_1583, w_041_1584, w_041_1585, w_041_1587, w_041_1588, w_041_1590, w_041_1591, w_041_1592, w_041_1593, w_041_1594, w_041_1595, w_041_1596, w_041_1597, w_041_1598, w_041_1599, w_041_1600, w_041_1601, w_041_1602, w_041_1603, w_041_1604, w_041_1605, w_041_1607, w_041_1608, w_041_1610, w_041_1611, w_041_1612, w_041_1613, w_041_1614, w_041_1615, w_041_1616, w_041_1617, w_041_1618, w_041_1619, w_041_1620, w_041_1621, w_041_1622, w_041_1623, w_041_1624, w_041_1625, w_041_1626, w_041_1627, w_041_1629, w_041_1630, w_041_1631, w_041_1632, w_041_1633, w_041_1634, w_041_1635, w_041_1636, w_041_1637, w_041_1638, w_041_1639, w_041_1640, w_041_1641, w_041_1642, w_041_1643, w_041_1644, w_041_1645, w_041_1647, w_041_1649, w_041_1650, w_041_1651, w_041_1652, w_041_1654, w_041_1655, w_041_1657, w_041_1658, w_041_1659, w_041_1660, w_041_1661, w_041_1664, w_041_1665, w_041_1666, w_041_1667, w_041_1668, w_041_1669, w_041_1670, w_041_1671, w_041_1672, w_041_1673, w_041_1674, w_041_1675, w_041_1677, w_041_1678, w_041_1679, w_041_1680, w_041_1681, w_041_1682, w_041_1684, w_041_1685, w_041_1687, w_041_1688, w_041_1689, w_041_1690, w_041_1691, w_041_1693, w_041_1694, w_041_1695, w_041_1696, w_041_1698, w_041_1700, w_041_1701, w_041_1702, w_041_1704, w_041_1705, w_041_1707, w_041_1708, w_041_1709, w_041_1711, w_041_1712, w_041_1713, w_041_1714, w_041_1715, w_041_1716, w_041_1717, w_041_1718, w_041_1719, w_041_1720, w_041_1721, w_041_1722, w_041_1723, w_041_1724, w_041_1726, w_041_1727, w_041_1728, w_041_1730, w_041_1731, w_041_1732, w_041_1733, w_041_1734, w_041_1735, w_041_1736, w_041_1737, w_041_1738, w_041_1739, w_041_1741, w_041_1742, w_041_1743, w_041_1744, w_041_1745, w_041_1746, w_041_1747, w_041_1748, w_041_1749, w_041_1750, w_041_1751, w_041_1752, w_041_1753, w_041_1754, w_041_1755, w_041_1756, w_041_1757, w_041_1758, w_041_1761, w_041_1762, w_041_1763, w_041_1764, w_041_1765, w_041_1766, w_041_1768, w_041_1770, w_041_1771, w_041_1772, w_041_1773, w_041_1774, w_041_1776, w_041_1778, w_041_1779, w_041_1781, w_041_1782, w_041_1784, w_041_1785, w_041_1786, w_041_1787, w_041_1788, w_041_1789, w_041_1790, w_041_1791, w_041_1792, w_041_1793, w_041_1794, w_041_1795, w_041_1796, w_041_1798, w_041_1799, w_041_1801, w_041_1802, w_041_1803, w_041_1804, w_041_1806, w_041_1809, w_041_1810, w_041_1811, w_041_1812, w_041_1813, w_041_1814, w_041_1816, w_041_1817, w_041_1818, w_041_1820, w_041_1823, w_041_1824, w_041_1825, w_041_1826, w_041_1827, w_041_1828, w_041_1830, w_041_1831, w_041_1832, w_041_1834, w_041_1836, w_041_1837, w_041_1838, w_041_1839, w_041_1840, w_041_1841, w_041_1842, w_041_1843, w_041_1845, w_041_1846, w_041_1847, w_041_1849, w_041_1850, w_041_1851, w_041_1852, w_041_1853, w_041_1855, w_041_1856, w_041_1857, w_041_1858, w_041_1859, w_041_1860, w_041_1861, w_041_1863, w_041_1864, w_041_1865, w_041_1866, w_041_1867, w_041_1868, w_041_1869, w_041_1871, w_041_1872, w_041_1873, w_041_1874, w_041_1875, w_041_1876, w_041_1877, w_041_1878, w_041_1879, w_041_1880, w_041_1881, w_041_1882, w_041_1883, w_041_1884, w_041_1885, w_041_1886, w_041_1887, w_041_1888, w_041_1889, w_041_1891, w_041_1893, w_041_1894, w_041_1895, w_041_1896, w_041_1897, w_041_1898, w_041_1899, w_041_1900, w_041_1901, w_041_1903, w_041_1904, w_041_1905, w_041_1906, w_041_1908, w_041_1910, w_041_1911, w_041_1913, w_041_1915, w_041_1916, w_041_1917, w_041_1920, w_041_1922, w_041_1923, w_041_1924, w_041_1925, w_041_1927, w_041_1928, w_041_1929, w_041_1930, w_041_1931, w_041_1932, w_041_1933, w_041_1935, w_041_1936, w_041_1937, w_041_1938, w_041_1939, w_041_1940, w_041_1941, w_041_1942, w_041_1944, w_041_1945, w_041_1946, w_041_1947, w_041_1948, w_041_1949, w_041_1950, w_041_1953, w_041_1954, w_041_1955, w_041_1956, w_041_1958, w_041_1959, w_041_1960, w_041_1961, w_041_1962, w_041_1963, w_041_1964, w_041_1965, w_041_1966, w_041_1967, w_041_1968, w_041_1969, w_041_1970, w_041_1971, w_041_1972, w_041_1973, w_041_1974, w_041_1975, w_041_1976, w_041_1977, w_041_1978, w_041_1979, w_041_1980, w_041_1981, w_041_1982, w_041_1983, w_041_1984, w_041_1985, w_041_1987, w_041_1988, w_041_1989, w_041_1992, w_041_1993, w_041_1995, w_041_1997, w_041_1998, w_041_2000, w_041_2001, w_041_2002, w_041_2003, w_041_2004, w_041_2005, w_041_2007, w_041_2008, w_041_2009, w_041_2010, w_041_2012, w_041_2014, w_041_2015, w_041_2016, w_041_2017, w_041_2018, w_041_2019, w_041_2020, w_041_2023, w_041_2024, w_041_2026, w_041_2027, w_041_2028, w_041_2029, w_041_2030, w_041_2031, w_041_2032, w_041_2033, w_041_2034, w_041_2035, w_041_2036, w_041_2037, w_041_2038, w_041_2039, w_041_2040, w_041_2041, w_041_2042, w_041_2044, w_041_2046, w_041_2047, w_041_2048, w_041_2049, w_041_2050, w_041_2051, w_041_2052, w_041_2053, w_041_2054, w_041_2055, w_041_2056, w_041_2058, w_041_2059, w_041_2061, w_041_2062, w_041_2063, w_041_2064, w_041_2065, w_041_2066, w_041_2067, w_041_2069, w_041_2071, w_041_2072, w_041_2073, w_041_2074, w_041_2076, w_041_2077, w_041_2079, w_041_2080, w_041_2081, w_041_2082, w_041_2083, w_041_2084, w_041_2085, w_041_2086, w_041_2087, w_041_2089, w_041_2090, w_041_2091, w_041_2092, w_041_2093, w_041_2094, w_041_2095, w_041_2096, w_041_2097, w_041_2099, w_041_2100, w_041_2101, w_041_2102, w_041_2104, w_041_2105, w_041_2106, w_041_2107, w_041_2108, w_041_2111, w_041_2113, w_041_2114, w_041_2115, w_041_2116, w_041_2117, w_041_2120, w_041_2121, w_041_2123, w_041_2124, w_041_2125, w_041_2126, w_041_2127, w_041_2130, w_041_2133, w_041_2134, w_041_2136, w_041_2137, w_041_2138, w_041_2139, w_041_2140, w_041_2141, w_041_2142, w_041_2143, w_041_2144, w_041_2146, w_041_2148, w_041_2149, w_041_2151, w_041_2152, w_041_2153, w_041_2154, w_041_2155, w_041_2156, w_041_2157, w_041_2158, w_041_2159, w_041_2161, w_041_2162, w_041_2163, w_041_2165, w_041_2166, w_041_2167, w_041_2169, w_041_2170, w_041_2171, w_041_2173, w_041_2176, w_041_2178, w_041_2179, w_041_2180, w_041_2181, w_041_2182, w_041_2183, w_041_2186, w_041_2190, w_041_2192, w_041_2193, w_041_2194, w_041_2195, w_041_2196, w_041_2197, w_041_2198, w_041_2200, w_041_2201, w_041_2202, w_041_2203, w_041_2204, w_041_2205, w_041_2206, w_041_2207, w_041_2208, w_041_2211, w_041_2213, w_041_2214, w_041_2215, w_041_2216, w_041_2217, w_041_2218, w_041_2220, w_041_2221, w_041_2223, w_041_2224, w_041_2225, w_041_2226, w_041_2227, w_041_2228, w_041_2229, w_041_2230, w_041_2231, w_041_2232, w_041_2234, w_041_2235, w_041_2236, w_041_2237, w_041_2238, w_041_2239, w_041_2240, w_041_2241, w_041_2242, w_041_2243, w_041_2244, w_041_2245, w_041_2246, w_041_2247, w_041_2249, w_041_2250, w_041_2251, w_041_2253, w_041_2254, w_041_2255, w_041_2257, w_041_2258, w_041_2261, w_041_2266, w_041_2267, w_041_2268, w_041_2270, w_041_2272, w_041_2273, w_041_2274, w_041_2275, w_041_2276, w_041_2277, w_041_2278, w_041_2279, w_041_2281, w_041_2283, w_041_2285, w_041_2286, w_041_2287, w_041_2288, w_041_2290, w_041_2292, w_041_2293, w_041_2294, w_041_2295, w_041_2296, w_041_2300, w_041_2301, w_041_2303, w_041_2307, w_041_2308, w_041_2309, w_041_2310, w_041_2313, w_041_2314, w_041_2315, w_041_2316, w_041_2317, w_041_2318, w_041_2319, w_041_2320, w_041_2321, w_041_2322, w_041_2323, w_041_2324, w_041_2325, w_041_2326, w_041_2327, w_041_2329, w_041_2331, w_041_2332, w_041_2333, w_041_2336, w_041_2338, w_041_2339, w_041_2340, w_041_2341, w_041_2342, w_041_2343, w_041_2344, w_041_2345, w_041_2346, w_041_2347, w_041_2348, w_041_2351, w_041_2352, w_041_2353, w_041_2354, w_041_2355, w_041_2357, w_041_2358, w_041_2360, w_041_2362, w_041_2363, w_041_2364, w_041_2365, w_041_2366, w_041_2367, w_041_2368, w_041_2369, w_041_2373, w_041_2375, w_041_2376, w_041_2377, w_041_2382, w_041_2383, w_041_2384, w_041_2385, w_041_2386, w_041_2387, w_041_2388, w_041_2390, w_041_2391, w_041_2394, w_041_2395, w_041_2396, w_041_2397, w_041_2398, w_041_2399, w_041_2400, w_041_2401, w_041_2402, w_041_2404, w_041_2405, w_041_2406, w_041_2407, w_041_2409, w_041_2412, w_041_2413, w_041_2414, w_041_2415, w_041_2416, w_041_2417, w_041_2418, w_041_2420, w_041_2421, w_041_2425, w_041_2427, w_041_2428, w_041_2429, w_041_2432, w_041_2433, w_041_2434, w_041_2435, w_041_2436, w_041_2437, w_041_2439, w_041_2440, w_041_2441, w_041_2442, w_041_2443, w_041_2444, w_041_2446, w_041_2447, w_041_2448, w_041_2451, w_041_2452, w_041_2454, w_041_2455, w_041_2456, w_041_2457, w_041_2459, w_041_2460, w_041_2461, w_041_2462, w_041_2463, w_041_2464, w_041_2466, w_041_2468, w_041_2469, w_041_2470, w_041_2472, w_041_2474, w_041_2475, w_041_2476, w_041_2477, w_041_2478, w_041_2480, w_041_2481, w_041_2482, w_041_2483, w_041_2484, w_041_2486, w_041_2488, w_041_2489, w_041_2491, w_041_2492, w_041_2494, w_041_2496, w_041_2497, w_041_2498, w_041_2499, w_041_2500, w_041_2501, w_041_2503, w_041_2504, w_041_2505, w_041_2506, w_041_2508, w_041_2509, w_041_2512, w_041_2514, w_041_2515, w_041_2516, w_041_2517, w_041_2518, w_041_2520, w_041_2521, w_041_2522, w_041_2523, w_041_2524, w_041_2525, w_041_2526, w_041_2527, w_041_2528, w_041_2530, w_041_2531, w_041_2535, w_041_2536, w_041_2538, w_041_2539, w_041_2540, w_041_2541, w_041_2543, w_041_2544, w_041_2546, w_041_2547, w_041_2548, w_041_2549, w_041_2550, w_041_2552, w_041_2553, w_041_2554, w_041_2558, w_041_2559, w_041_2560, w_041_2561, w_041_2562, w_041_2563, w_041_2566, w_041_2567, w_041_2568, w_041_2569, w_041_2570, w_041_2571, w_041_2573, w_041_2574, w_041_2575, w_041_2577, w_041_2578, w_041_2579, w_041_2580, w_041_2583, w_041_2584, w_041_2585, w_041_2587, w_041_2590, w_041_2592, w_041_2593, w_041_2597, w_041_2598, w_041_2601, w_041_2602, w_041_2603, w_041_2606, w_041_2608, w_041_2609, w_041_2610, w_041_2611, w_041_2612, w_041_2613, w_041_2614, w_041_2615, w_041_2617, w_041_2618, w_041_2619, w_041_2620, w_041_2622, w_041_2623, w_041_2624, w_041_2625, w_041_2626, w_041_2628, w_041_2629, w_041_2630, w_041_2632, w_041_2634, w_041_2635, w_041_2637, w_041_2639, w_041_2640, w_041_2642, w_041_2643, w_041_2645, w_041_2646, w_041_2647, w_041_2648, w_041_2649, w_041_2650, w_041_2651, w_041_2652, w_041_2653, w_041_2654, w_041_2655, w_041_2656, w_041_2657, w_041_2658, w_041_2659, w_041_2661, w_041_2663, w_041_2664, w_041_2665, w_041_2666, w_041_2667, w_041_2668, w_041_2671, w_041_2674, w_041_2675, w_041_2676, w_041_2677, w_041_2678, w_041_2682, w_041_2683, w_041_2684, w_041_2685, w_041_2686, w_041_2687, w_041_2689, w_041_2690, w_041_2692, w_041_2693, w_041_2694, w_041_2695, w_041_2696, w_041_2697, w_041_2698, w_041_2699, w_041_2700, w_041_2701, w_041_2703, w_041_2705, w_041_2706, w_041_2711, w_041_2714, w_041_2715, w_041_2716, w_041_2718, w_041_2720, w_041_2722, w_041_2723, w_041_2724, w_041_2727, w_041_2728, w_041_2729, w_041_2730, w_041_2732, w_041_2733, w_041_2735, w_041_2736, w_041_2737, w_041_2739, w_041_2741, w_041_2742, w_041_2743, w_041_2744, w_041_2745, w_041_2746, w_041_2747, w_041_2749, w_041_2750, w_041_2751, w_041_2752, w_041_2754, w_041_2755, w_041_2756, w_041_2759, w_041_2761, w_041_2762, w_041_2764, w_041_2765, w_041_2766, w_041_2767, w_041_2769, w_041_2770, w_041_2775, w_041_2776, w_041_2778, w_041_2779, w_041_2780, w_041_2782, w_041_2783, w_041_2784, w_041_2786, w_041_2787, w_041_2788, w_041_2789, w_041_2791, w_041_2792, w_041_2794, w_041_2795, w_041_2796, w_041_2797, w_041_2798, w_041_2799, w_041_2800, w_041_2801, w_041_2802, w_041_2805, w_041_2806, w_041_2807, w_041_2811, w_041_2812, w_041_2815, w_041_2816, w_041_2819, w_041_2820, w_041_2821, w_041_2822, w_041_2824, w_041_2825, w_041_2827, w_041_2828, w_041_2830, w_041_2832, w_041_2833, w_041_2834, w_041_2836, w_041_2837, w_041_2838, w_041_2839, w_041_2840, w_041_2841, w_041_2844, w_041_2847, w_041_2849, w_041_2853, w_041_2854, w_041_2855, w_041_2857, w_041_2859, w_041_2860, w_041_2861, w_041_2862, w_041_2863, w_041_2864, w_041_2865, w_041_2866, w_041_2870, w_041_2871, w_041_2873, w_041_2874, w_041_2875, w_041_2876, w_041_2877, w_041_2878, w_041_2880, w_041_2881, w_041_2882, w_041_2883, w_041_2884, w_041_2886, w_041_2890, w_041_2891, w_041_2892, w_041_2893, w_041_2894, w_041_2895, w_041_2896, w_041_2899, w_041_2900, w_041_2901, w_041_2903, w_041_2904, w_041_2905, w_041_2907, w_041_2908, w_041_2909, w_041_2911, w_041_2913, w_041_2914, w_041_2915, w_041_2916, w_041_2917, w_041_2918, w_041_2919, w_041_2920, w_041_2921, w_041_2922, w_041_2923, w_041_2924, w_041_2925, w_041_2926, w_041_2927, w_041_2928, w_041_2929, w_041_2931, w_041_2935, w_041_2936, w_041_2937, w_041_2938, w_041_2939, w_041_2941, w_041_2945, w_041_2946, w_041_2949, w_041_2950, w_041_2952, w_041_2953, w_041_2954, w_041_2955, w_041_2957, w_041_2958, w_041_2959, w_041_2960, w_041_2961, w_041_2962, w_041_2965, w_041_2966, w_041_2967, w_041_2968, w_041_2970, w_041_2972, w_041_2973, w_041_2974, w_041_2975, w_041_2976, w_041_2977, w_041_2979, w_041_2980, w_041_2983, w_041_2986, w_041_2988, w_041_2989, w_041_2992, w_041_2993, w_041_2994, w_041_2995, w_041_2996, w_041_2997, w_041_2998, w_041_2999, w_041_3002, w_041_3004, w_041_3005, w_041_3006, w_041_3008, w_041_3010, w_041_3011, w_041_3012, w_041_3015, w_041_3018, w_041_3019, w_041_3022, w_041_3023, w_041_3025, w_041_3028, w_041_3030, w_041_3031, w_041_3032, w_041_3033, w_041_3034, w_041_3035, w_041_3038, w_041_3039, w_041_3040, w_041_3041, w_041_3043, w_041_3044, w_041_3045, w_041_3046, w_041_3047, w_041_3048, w_041_3049, w_041_3053, w_041_3054, w_041_3055, w_041_3056, w_041_3059, w_041_3060, w_041_3061, w_041_3062, w_041_3063, w_041_3064, w_041_3066, w_041_3067, w_041_3069, w_041_3071, w_041_3072, w_041_3073, w_041_3075, w_041_3076, w_041_3077, w_041_3078, w_041_3080, w_041_3082, w_041_3083, w_041_3084, w_041_3085, w_041_3089, w_041_3090, w_041_3091, w_041_3093, w_041_3095, w_041_3096, w_041_3097, w_041_3098, w_041_3099, w_041_3100, w_041_3101, w_041_3103, w_041_3104, w_041_3106, w_041_3107, w_041_3110, w_041_3111, w_041_3112, w_041_3114, w_041_3116, w_041_3117, w_041_3118, w_041_3120, w_041_3121, w_041_3122, w_041_3123, w_041_3124, w_041_3125, w_041_3126, w_041_3127, w_041_3129, w_041_3132, w_041_3134, w_041_3136, w_041_3138, w_041_3139, w_041_3140, w_041_3141, w_041_3142, w_041_3146, w_041_3147, w_041_3148, w_041_3149, w_041_3150, w_041_3151, w_041_3152, w_041_3153, w_041_3156, w_041_3157, w_041_3158, w_041_3159, w_041_3160, w_041_3161, w_041_3162, w_041_3163, w_041_3165, w_041_3170, w_041_3171, w_041_3172, w_041_3173, w_041_3174, w_041_3175, w_041_3176, w_041_3177, w_041_3178, w_041_3179, w_041_3180, w_041_3181, w_041_3186, w_041_3188, w_041_3189, w_041_3191, w_041_3193, w_041_3194, w_041_3196, w_041_3197, w_041_3199, w_041_3200, w_041_3201, w_041_3202, w_041_3204, w_041_3206, w_041_3207, w_041_3208, w_041_3209, w_041_3210, w_041_3211, w_041_3212, w_041_3213, w_041_3214, w_041_3215, w_041_3216, w_041_3217, w_041_3218, w_041_3219, w_041_3220, w_041_3221, w_041_3222, w_041_3223, w_041_3224, w_041_3225, w_041_3226, w_041_3228, w_041_3229, w_041_3230, w_041_3231, w_041_3232, w_041_3233, w_041_3234, w_041_3235, w_041_3236, w_041_3237, w_041_3238, w_041_3239, w_041_3240, w_041_3241, w_041_3242, w_041_3245, w_041_3246, w_041_3247, w_041_3248, w_041_3249, w_041_3250, w_041_3252, w_041_3253, w_041_3254, w_041_3256, w_041_3258, w_041_3259, w_041_3260, w_041_3261, w_041_3263, w_041_3265, w_041_3266, w_041_3267, w_041_3268, w_041_3269, w_041_3270, w_041_3271, w_041_3272, w_041_3273, w_041_3275, w_041_3276, w_041_3277, w_041_3278, w_041_3279, w_041_3280, w_041_3281, w_041_3283, w_041_3284, w_041_3287, w_041_3288, w_041_3289, w_041_3290, w_041_3292, w_041_3293, w_041_3294, w_041_3295, w_041_3296, w_041_3298, w_041_3301, w_041_3303, w_041_3304, w_041_3306, w_041_3307, w_041_3308, w_041_3309, w_041_3310, w_041_3311, w_041_3312, w_041_3313, w_041_3314, w_041_3315, w_041_3316, w_041_3320, w_041_3321, w_041_3327, w_041_3328, w_041_3329, w_041_3330, w_041_3331, w_041_3333, w_041_3334, w_041_3335, w_041_3336, w_041_3337, w_041_3338, w_041_3339, w_041_3341, w_041_3343, w_041_3344, w_041_3345, w_041_3346, w_041_3347, w_041_3348, w_041_3349, w_041_3350, w_041_3352, w_041_3354, w_041_3355, w_041_3356, w_041_3360, w_041_3361, w_041_3362, w_041_3363, w_041_3365, w_041_3366, w_041_3367, w_041_3368, w_041_3369, w_041_3370, w_041_3371, w_041_3372, w_041_3373, w_041_3374, w_041_3377, w_041_3378, w_041_3379, w_041_3380, w_041_3381, w_041_3382, w_041_3383, w_041_3384, w_041_3385, w_041_3386, w_041_3387, w_041_3389, w_041_3390, w_041_3392, w_041_3393, w_041_3394, w_041_3396, w_041_3397, w_041_3398, w_041_3400, w_041_3401, w_041_3404, w_041_3405, w_041_3406, w_041_3407, w_041_3409, w_041_3410, w_041_3411, w_041_3413, w_041_3414, w_041_3415, w_041_3416, w_041_3418, w_041_3419, w_041_3422, w_041_3423, w_041_3424, w_041_3426, w_041_3427, w_041_3429, w_041_3431, w_041_3432, w_041_3433, w_041_3434, w_041_3435, w_041_3436, w_041_3437, w_041_3438, w_041_3439, w_041_3440, w_041_3441, w_041_3442, w_041_3443, w_041_3444, w_041_3446, w_041_3447, w_041_3448, w_041_3450, w_041_3451, w_041_3453, w_041_3454, w_041_3455, w_041_3457, w_041_3458, w_041_3460, w_041_3461, w_041_3462, w_041_3464, w_041_3465, w_041_3466, w_041_3467, w_041_3468, w_041_3469, w_041_3470, w_041_3471, w_041_3473, w_041_3474, w_041_3476, w_041_3479, w_041_3480, w_041_3481, w_041_3482, w_041_3483, w_041_3484, w_041_3485, w_041_3486, w_041_3488, w_041_3489, w_041_3490, w_041_3491, w_041_3492, w_041_3493, w_041_3494, w_041_3495, w_041_3498, w_041_3500, w_041_3501, w_041_3502, w_041_3503, w_041_3505, w_041_3506, w_041_3507, w_041_3508, w_041_3512, w_041_3513, w_041_3514, w_041_3515, w_041_3516, w_041_3517, w_041_3518, w_041_3519, w_041_3520, w_041_3521, w_041_3523, w_041_3525, w_041_3526, w_041_3527, w_041_3528, w_041_3529, w_041_3530, w_041_3531, w_041_3532, w_041_3534, w_041_3535, w_041_3536, w_041_3538, w_041_3539, w_041_3540, w_041_3541, w_041_3542, w_041_3544, w_041_3545, w_041_3546, w_041_3548, w_041_3550, w_041_3552, w_041_3553, w_041_3556, w_041_3557, w_041_3558, w_041_3560, w_041_3563, w_041_3564, w_041_3565, w_041_3567, w_041_3569, w_041_3570, w_041_3571, w_041_3572, w_041_3573, w_041_3574, w_041_3575, w_041_3576, w_041_3577, w_041_3578, w_041_3580, w_041_3581, w_041_3582, w_041_3583, w_041_3584, w_041_3585, w_041_3586, w_041_3587, w_041_3589, w_041_3590, w_041_3591, w_041_3592, w_041_3593, w_041_3594, w_041_3595, w_041_3596, w_041_3597, w_041_3598, w_041_3599, w_041_3600, w_041_3601, w_041_3602, w_041_3604, w_041_3605, w_041_3607, w_041_3608, w_041_3609, w_041_3610, w_041_3611, w_041_3612, w_041_3613, w_041_3616, w_041_3617, w_041_3618, w_041_3619, w_041_3620, w_041_3621, w_041_3622, w_041_3624, w_041_3625, w_041_3626, w_041_3627, w_041_3628, w_041_3629, w_041_3630, w_041_3631, w_041_3632, w_041_3633, w_041_3636, w_041_3637, w_041_3640, w_041_3642, w_041_3644, w_041_3645, w_041_3647, w_041_3648, w_041_3649, w_041_3651, w_041_3652, w_041_3655, w_041_3657, w_041_3659, w_041_3660, w_041_3663, w_041_3664, w_041_3665, w_041_3666, w_041_3667, w_041_3668, w_041_3669, w_041_3670, w_041_3673, w_041_3674, w_041_3675, w_041_3676, w_041_3678, w_041_3680, w_041_3681, w_041_3682, w_041_3684, w_041_3685, w_041_3686, w_041_3687, w_041_3689, w_041_3690, w_041_3691, w_041_3692, w_041_3695, w_041_3696, w_041_3697, w_041_3698, w_041_3702, w_041_3703, w_041_3706, w_041_3708, w_041_3710, w_041_3711, w_041_3712, w_041_3713, w_041_3714, w_041_3716, w_041_3717, w_041_3720, w_041_3721, w_041_3723, w_041_3724, w_041_3725, w_041_3727, w_041_3728, w_041_3729, w_041_3730, w_041_3731, w_041_3732, w_041_3733, w_041_3734, w_041_3735, w_041_3736, w_041_3738, w_041_3740, w_041_3741, w_041_3742, w_041_3743, w_041_3744, w_041_3746, w_041_3747, w_041_3750, w_041_3753, w_041_3754, w_041_3755, w_041_3757, w_041_3758, w_041_3760, w_041_3762, w_041_3763, w_041_3766, w_041_3767, w_041_3768, w_041_3769, w_041_3770, w_041_3771, w_041_3772, w_041_3773, w_041_3774, w_041_3775, w_041_3777, w_041_3780, w_041_3782, w_041_3783, w_041_3785, w_041_3786, w_041_3787, w_041_3788, w_041_3789, w_041_3791, w_041_3792, w_041_3793, w_041_3794, w_041_3796, w_041_3798, w_041_3799, w_041_3801, w_041_3802, w_041_3803, w_041_3804, w_041_3805, w_041_3806, w_041_3807, w_041_3809, w_041_3812, w_041_3814, w_041_3816, w_041_3817, w_041_3818, w_041_3819, w_041_3820, w_041_3821, w_041_3822, w_041_3824, w_041_3825, w_041_3826, w_041_3827, w_041_3830, w_041_3831, w_041_3834, w_041_3836, w_041_3837, w_041_3838, w_041_3839, w_041_3840, w_041_3842, w_041_3845, w_041_3847, w_041_3848, w_041_3850, w_041_3851, w_041_3852, w_041_3853, w_041_3855, w_041_3856, w_041_3857, w_041_3861, w_041_3862, w_041_3864, w_041_3866, w_041_3867, w_041_3868, w_041_3869, w_041_3870, w_041_3871, w_041_3872, w_041_3874, w_041_3876, w_041_3877, w_041_3880, w_041_3882, w_041_3883, w_041_3884, w_041_3885, w_041_3886, w_041_3887, w_041_3889, w_041_3890, w_041_3892, w_041_3893, w_041_3894, w_041_3895, w_041_3896, w_041_3898, w_041_3899, w_041_3901, w_041_3902, w_041_3903, w_041_3904, w_041_3905, w_041_3907, w_041_3909, w_041_3910, w_041_3911, w_041_3912, w_041_3913, w_041_3916, w_041_3917, w_041_3918, w_041_3919, w_041_3920, w_041_3922, w_041_3923, w_041_3924, w_041_3925, w_041_3926, w_041_3928, w_041_3929, w_041_3930, w_041_3931, w_041_3932, w_041_3935;
  wire w_042_000, w_042_001, w_042_002, w_042_003, w_042_004, w_042_005, w_042_006, w_042_007, w_042_008, w_042_009, w_042_010, w_042_011, w_042_012, w_042_013, w_042_014, w_042_015, w_042_016, w_042_017, w_042_018, w_042_019, w_042_020, w_042_021, w_042_022, w_042_023, w_042_024, w_042_025, w_042_026, w_042_027, w_042_028, w_042_029, w_042_030, w_042_031, w_042_032, w_042_033, w_042_034, w_042_035, w_042_036, w_042_037, w_042_038, w_042_039, w_042_040, w_042_041, w_042_042, w_042_043, w_042_044, w_042_045, w_042_046, w_042_047, w_042_048, w_042_049, w_042_050, w_042_051, w_042_052, w_042_053, w_042_054, w_042_056, w_042_057, w_042_058, w_042_059, w_042_060, w_042_061, w_042_062, w_042_063, w_042_064, w_042_065, w_042_066, w_042_067, w_042_068, w_042_069, w_042_070, w_042_071, w_042_072, w_042_073, w_042_074, w_042_075, w_042_076, w_042_077, w_042_078, w_042_079, w_042_080, w_042_081, w_042_082, w_042_083, w_042_084, w_042_085, w_042_086, w_042_087, w_042_088, w_042_089, w_042_090, w_042_091, w_042_092, w_042_093, w_042_094, w_042_095, w_042_096, w_042_097, w_042_098, w_042_099, w_042_100, w_042_101, w_042_102, w_042_103, w_042_104, w_042_105, w_042_106, w_042_107, w_042_108, w_042_109, w_042_110, w_042_111, w_042_112, w_042_113, w_042_114, w_042_115, w_042_116, w_042_117, w_042_118, w_042_119, w_042_120, w_042_121, w_042_122, w_042_123, w_042_124, w_042_125, w_042_126, w_042_127, w_042_128, w_042_129, w_042_130, w_042_131, w_042_132, w_042_133, w_042_134, w_042_136, w_042_137, w_042_138, w_042_139, w_042_140, w_042_141, w_042_142, w_042_143, w_042_144, w_042_145, w_042_146, w_042_147, w_042_148, w_042_149, w_042_150, w_042_151, w_042_152, w_042_153, w_042_154, w_042_155, w_042_156, w_042_157, w_042_158, w_042_159, w_042_160, w_042_161, w_042_162, w_042_163, w_042_164, w_042_165, w_042_166, w_042_167, w_042_168, w_042_169, w_042_170, w_042_171, w_042_172, w_042_173, w_042_174, w_042_175, w_042_176, w_042_177, w_042_178, w_042_179, w_042_180, w_042_181, w_042_182, w_042_183, w_042_184, w_042_185, w_042_186, w_042_187, w_042_188, w_042_189, w_042_190, w_042_191, w_042_192, w_042_193, w_042_194, w_042_195, w_042_196, w_042_197, w_042_198, w_042_199, w_042_200, w_042_201, w_042_202, w_042_203, w_042_204, w_042_205, w_042_206, w_042_207, w_042_208, w_042_209, w_042_210, w_042_211, w_042_212, w_042_213, w_042_214, w_042_215, w_042_216, w_042_217, w_042_218, w_042_219, w_042_220, w_042_221, w_042_222, w_042_223, w_042_224, w_042_225, w_042_226, w_042_227, w_042_228, w_042_229, w_042_230, w_042_231, w_042_232, w_042_233, w_042_234, w_042_235, w_042_236, w_042_237, w_042_238, w_042_239, w_042_240, w_042_241, w_042_242, w_042_243, w_042_244, w_042_245, w_042_246, w_042_247, w_042_248, w_042_249, w_042_250, w_042_251, w_042_252, w_042_253, w_042_255, w_042_256, w_042_257, w_042_258, w_042_259, w_042_260, w_042_261, w_042_262, w_042_263, w_042_264, w_042_265, w_042_266, w_042_267, w_042_268, w_042_269, w_042_270, w_042_271, w_042_272, w_042_273, w_042_274, w_042_275, w_042_276, w_042_277, w_042_278, w_042_279, w_042_280, w_042_281, w_042_282, w_042_283, w_042_284, w_042_285, w_042_286, w_042_287, w_042_288, w_042_290, w_042_291, w_042_292, w_042_293, w_042_294, w_042_295, w_042_296, w_042_297, w_042_298, w_042_299, w_042_300, w_042_301, w_042_302, w_042_303, w_042_304, w_042_305, w_042_306, w_042_307, w_042_308, w_042_309, w_042_310, w_042_311, w_042_312, w_042_313, w_042_314, w_042_315, w_042_316, w_042_317, w_042_318, w_042_319, w_042_320, w_042_321, w_042_322, w_042_323, w_042_324, w_042_325, w_042_326, w_042_327, w_042_328, w_042_329, w_042_331, w_042_332, w_042_333, w_042_334, w_042_335, w_042_337, w_042_338, w_042_339, w_042_340, w_042_341, w_042_342, w_042_343, w_042_344, w_042_345, w_042_346, w_042_347, w_042_348, w_042_349, w_042_350, w_042_351, w_042_352, w_042_353, w_042_354, w_042_355, w_042_356, w_042_357, w_042_358, w_042_360, w_042_361, w_042_362, w_042_363, w_042_364, w_042_365, w_042_366, w_042_367, w_042_369, w_042_370, w_042_371, w_042_372, w_042_373, w_042_374, w_042_375, w_042_376, w_042_377, w_042_378, w_042_379, w_042_380, w_042_381, w_042_382, w_042_383, w_042_384, w_042_385, w_042_386, w_042_387, w_042_388, w_042_389, w_042_390, w_042_391, w_042_392, w_042_393, w_042_395, w_042_396, w_042_397, w_042_398, w_042_399, w_042_400, w_042_401, w_042_402, w_042_403, w_042_405, w_042_406, w_042_407, w_042_408, w_042_409, w_042_410, w_042_411, w_042_412, w_042_413, w_042_414, w_042_415, w_042_416, w_042_417, w_042_418, w_042_419, w_042_420, w_042_421, w_042_422, w_042_423, w_042_424, w_042_425, w_042_426, w_042_427, w_042_428, w_042_429, w_042_430, w_042_431, w_042_432, w_042_433, w_042_434, w_042_435, w_042_436, w_042_437, w_042_438, w_042_439, w_042_440, w_042_441, w_042_442, w_042_443, w_042_444, w_042_445, w_042_446, w_042_447, w_042_448, w_042_449, w_042_450, w_042_451, w_042_452, w_042_453, w_042_454, w_042_455, w_042_457, w_042_458, w_042_459, w_042_460, w_042_461, w_042_462, w_042_463, w_042_464, w_042_465, w_042_466, w_042_467, w_042_468, w_042_469, w_042_470, w_042_471, w_042_472, w_042_473, w_042_474, w_042_477, w_042_478, w_042_479, w_042_480, w_042_481, w_042_482, w_042_483, w_042_484, w_042_485, w_042_486, w_042_487, w_042_488, w_042_490, w_042_491, w_042_492, w_042_493, w_042_494, w_042_495, w_042_496, w_042_497, w_042_498, w_042_499, w_042_500, w_042_501, w_042_502, w_042_503, w_042_504, w_042_505, w_042_506, w_042_507, w_042_508, w_042_509, w_042_510, w_042_511, w_042_512, w_042_513, w_042_514, w_042_515, w_042_516, w_042_518, w_042_519, w_042_520, w_042_521, w_042_522, w_042_523, w_042_524, w_042_525, w_042_526, w_042_527, w_042_528, w_042_529, w_042_530, w_042_531, w_042_532, w_042_533, w_042_534, w_042_535, w_042_536, w_042_537, w_042_538, w_042_539, w_042_540, w_042_541, w_042_542, w_042_543, w_042_544, w_042_545, w_042_546, w_042_547, w_042_548, w_042_549, w_042_550, w_042_551, w_042_552, w_042_553, w_042_554, w_042_555, w_042_556, w_042_557, w_042_559, w_042_560, w_042_561, w_042_562, w_042_563, w_042_564, w_042_565, w_042_566, w_042_567, w_042_568, w_042_569, w_042_570, w_042_571, w_042_573, w_042_574, w_042_575, w_042_576, w_042_577, w_042_578, w_042_579, w_042_580, w_042_581, w_042_582, w_042_583, w_042_584, w_042_585, w_042_586, w_042_587, w_042_588, w_042_589, w_042_590, w_042_591, w_042_592, w_042_593, w_042_594, w_042_595, w_042_596, w_042_597, w_042_598, w_042_599, w_042_600, w_042_601, w_042_602, w_042_603, w_042_604, w_042_605, w_042_606, w_042_607, w_042_608, w_042_610, w_042_612, w_042_613, w_042_614, w_042_615, w_042_616, w_042_617, w_042_618, w_042_619, w_042_620, w_042_621, w_042_622, w_042_623, w_042_624, w_042_625, w_042_626, w_042_627, w_042_628, w_042_629, w_042_630, w_042_631, w_042_632, w_042_633, w_042_634, w_042_635, w_042_636, w_042_637, w_042_638, w_042_639, w_042_640, w_042_641, w_042_642, w_042_643, w_042_644, w_042_645, w_042_646, w_042_647, w_042_648, w_042_649, w_042_650, w_042_651, w_042_652, w_042_653, w_042_654, w_042_655, w_042_656, w_042_657, w_042_658, w_042_659, w_042_660, w_042_661, w_042_662, w_042_663, w_042_664, w_042_665, w_042_666, w_042_667, w_042_668, w_042_669, w_042_670, w_042_671, w_042_672, w_042_673, w_042_674, w_042_675, w_042_676, w_042_677, w_042_678, w_042_679, w_042_680, w_042_681, w_042_682, w_042_683, w_042_684, w_042_686, w_042_687, w_042_688, w_042_689, w_042_690, w_042_691, w_042_692, w_042_693, w_042_694, w_042_695, w_042_696, w_042_697, w_042_698, w_042_699, w_042_700, w_042_701, w_042_702, w_042_703, w_042_704, w_042_705, w_042_706, w_042_707, w_042_708, w_042_709, w_042_710, w_042_711, w_042_712, w_042_713, w_042_714, w_042_715, w_042_716, w_042_718, w_042_719, w_042_720, w_042_721, w_042_722, w_042_723, w_042_724, w_042_725, w_042_726, w_042_727, w_042_728, w_042_729, w_042_730, w_042_731, w_042_732, w_042_733, w_042_734, w_042_735, w_042_736, w_042_737, w_042_738, w_042_739, w_042_740, w_042_741, w_042_742, w_042_743, w_042_744, w_042_745, w_042_746, w_042_747, w_042_748, w_042_749, w_042_750, w_042_752, w_042_753, w_042_754, w_042_755, w_042_756, w_042_757, w_042_758, w_042_759, w_042_760, w_042_761, w_042_762, w_042_764, w_042_765, w_042_766, w_042_767, w_042_768, w_042_769, w_042_770, w_042_771, w_042_772, w_042_773, w_042_774, w_042_775, w_042_776, w_042_777, w_042_778, w_042_779, w_042_780, w_042_781, w_042_782, w_042_783, w_042_784, w_042_785, w_042_786, w_042_787, w_042_789, w_042_790, w_042_791, w_042_792, w_042_793, w_042_794, w_042_795, w_042_796, w_042_797, w_042_798, w_042_799, w_042_800, w_042_801, w_042_802, w_042_803, w_042_805, w_042_806, w_042_807, w_042_808, w_042_809, w_042_810, w_042_811, w_042_812, w_042_813, w_042_814, w_042_815, w_042_816, w_042_817, w_042_818, w_042_819, w_042_820, w_042_821, w_042_822, w_042_823, w_042_824, w_042_825, w_042_826, w_042_827, w_042_828, w_042_829, w_042_830, w_042_831, w_042_832, w_042_833, w_042_834, w_042_835, w_042_836, w_042_837, w_042_838, w_042_839, w_042_840, w_042_841, w_042_842, w_042_843, w_042_844, w_042_845, w_042_846, w_042_847, w_042_848, w_042_849, w_042_850, w_042_851, w_042_852, w_042_853, w_042_854, w_042_855, w_042_856, w_042_857, w_042_858, w_042_859, w_042_860, w_042_863, w_042_864, w_042_865, w_042_866, w_042_867, w_042_868, w_042_869, w_042_871, w_042_872, w_042_873, w_042_874, w_042_875, w_042_876, w_042_877, w_042_878, w_042_879, w_042_880, w_042_881, w_042_882, w_042_883, w_042_884, w_042_885, w_042_886, w_042_887, w_042_888, w_042_889, w_042_890, w_042_891, w_042_892, w_042_893, w_042_894, w_042_895, w_042_896, w_042_897, w_042_898, w_042_900, w_042_902, w_042_903, w_042_904, w_042_905, w_042_906, w_042_907, w_042_908, w_042_909, w_042_910, w_042_911, w_042_913, w_042_914, w_042_915, w_042_916, w_042_917, w_042_918, w_042_919, w_042_920, w_042_921, w_042_922, w_042_923, w_042_925, w_042_926, w_042_928, w_042_929, w_042_930, w_042_931, w_042_932, w_042_933, w_042_934, w_042_935, w_042_936, w_042_937, w_042_938, w_042_939, w_042_941, w_042_942, w_042_943, w_042_944, w_042_945, w_042_946, w_042_947, w_042_948, w_042_949, w_042_950, w_042_951, w_042_952, w_042_953, w_042_954, w_042_955, w_042_956, w_042_957, w_042_958, w_042_960, w_042_961, w_042_962, w_042_963, w_042_964, w_042_965, w_042_966, w_042_967, w_042_968, w_042_969, w_042_970, w_042_971, w_042_972, w_042_973, w_042_974, w_042_975, w_042_976, w_042_977, w_042_978, w_042_979, w_042_980, w_042_981, w_042_982, w_042_984, w_042_985, w_042_986, w_042_987, w_042_988, w_042_989, w_042_990, w_042_991, w_042_992, w_042_993, w_042_994, w_042_995, w_042_996, w_042_997, w_042_998, w_042_999, w_042_1000, w_042_1001, w_042_1002, w_042_1003, w_042_1004, w_042_1005, w_042_1006, w_042_1007, w_042_1009, w_042_1010, w_042_1011, w_042_1012, w_042_1013, w_042_1014, w_042_1015, w_042_1016, w_042_1017, w_042_1018, w_042_1019, w_042_1020, w_042_1021, w_042_1023, w_042_1024, w_042_1025, w_042_1026, w_042_1027, w_042_1028, w_042_1029, w_042_1031, w_042_1032, w_042_1033, w_042_1034, w_042_1036, w_042_1037, w_042_1038, w_042_1039, w_042_1040, w_042_1041, w_042_1042, w_042_1043, w_042_1044, w_042_1045, w_042_1046, w_042_1047, w_042_1048, w_042_1049, w_042_1050, w_042_1051, w_042_1052, w_042_1053, w_042_1054, w_042_1055, w_042_1056, w_042_1057, w_042_1058, w_042_1059, w_042_1060, w_042_1061, w_042_1062, w_042_1063, w_042_1064, w_042_1065, w_042_1066, w_042_1067, w_042_1068, w_042_1069, w_042_1070, w_042_1071, w_042_1072, w_042_1073, w_042_1074, w_042_1075, w_042_1076, w_042_1077, w_042_1078, w_042_1079, w_042_1080, w_042_1081, w_042_1082, w_042_1083, w_042_1084, w_042_1085, w_042_1086, w_042_1087, w_042_1088, w_042_1089, w_042_1090, w_042_1091, w_042_1092, w_042_1093, w_042_1094, w_042_1095, w_042_1096, w_042_1097, w_042_1098, w_042_1099, w_042_1100, w_042_1101, w_042_1102, w_042_1103, w_042_1104, w_042_1105, w_042_1106, w_042_1107, w_042_1108, w_042_1109, w_042_1111, w_042_1112, w_042_1114, w_042_1115, w_042_1116, w_042_1117, w_042_1118, w_042_1119, w_042_1120, w_042_1121, w_042_1122, w_042_1123, w_042_1126, w_042_1127, w_042_1128, w_042_1129, w_042_1130, w_042_1131, w_042_1132, w_042_1133, w_042_1134, w_042_1135, w_042_1136, w_042_1137, w_042_1138, w_042_1139, w_042_1140, w_042_1141, w_042_1142, w_042_1144, w_042_1145, w_042_1146, w_042_1147, w_042_1148, w_042_1149, w_042_1150, w_042_1151, w_042_1152, w_042_1153, w_042_1154, w_042_1155, w_042_1156, w_042_1157, w_042_1158, w_042_1159, w_042_1160, w_042_1161, w_042_1162, w_042_1163, w_042_1164, w_042_1165, w_042_1166, w_042_1167, w_042_1168, w_042_1169, w_042_1170, w_042_1171, w_042_1172, w_042_1173, w_042_1174, w_042_1175, w_042_1176, w_042_1177, w_042_1178, w_042_1179, w_042_1180, w_042_1181, w_042_1182, w_042_1183, w_042_1184, w_042_1185, w_042_1186, w_042_1187, w_042_1188, w_042_1189, w_042_1190, w_042_1191, w_042_1192, w_042_1193, w_042_1194, w_042_1195, w_042_1196, w_042_1197, w_042_1198, w_042_1199, w_042_1200, w_042_1201, w_042_1202, w_042_1203, w_042_1204, w_042_1205, w_042_1208, w_042_1209, w_042_1210, w_042_1211, w_042_1212, w_042_1213, w_042_1214, w_042_1215, w_042_1216, w_042_1217, w_042_1218, w_042_1220, w_042_1221, w_042_1222, w_042_1223, w_042_1224, w_042_1225, w_042_1226, w_042_1227, w_042_1228, w_042_1229, w_042_1230, w_042_1231, w_042_1232, w_042_1233, w_042_1234, w_042_1235, w_042_1236, w_042_1237, w_042_1238, w_042_1239, w_042_1240, w_042_1242, w_042_1243, w_042_1244, w_042_1245, w_042_1246, w_042_1247, w_042_1248, w_042_1249, w_042_1251, w_042_1252, w_042_1254, w_042_1255, w_042_1256, w_042_1257, w_042_1258, w_042_1259, w_042_1260, w_042_1261, w_042_1262, w_042_1263, w_042_1264, w_042_1265, w_042_1266, w_042_1267, w_042_1268, w_042_1269, w_042_1270, w_042_1272, w_042_1274, w_042_1275, w_042_1276, w_042_1277, w_042_1278, w_042_1279, w_042_1280, w_042_1281, w_042_1282, w_042_1283, w_042_1284, w_042_1285, w_042_1286, w_042_1287, w_042_1288, w_042_1289, w_042_1290, w_042_1291, w_042_1292, w_042_1293, w_042_1294, w_042_1295, w_042_1296, w_042_1297, w_042_1298, w_042_1299, w_042_1300, w_042_1301, w_042_1302, w_042_1303, w_042_1305, w_042_1306, w_042_1307, w_042_1309, w_042_1310, w_042_1311, w_042_1312, w_042_1313, w_042_1314, w_042_1315, w_042_1316, w_042_1317, w_042_1318, w_042_1319, w_042_1320, w_042_1321, w_042_1322, w_042_1323, w_042_1324, w_042_1325, w_042_1326, w_042_1327, w_042_1328, w_042_1329, w_042_1330, w_042_1331, w_042_1332, w_042_1333, w_042_1334, w_042_1335, w_042_1336, w_042_1337, w_042_1338, w_042_1339, w_042_1341, w_042_1342, w_042_1343, w_042_1344, w_042_1345, w_042_1346, w_042_1347, w_042_1348, w_042_1349, w_042_1350, w_042_1351, w_042_1352, w_042_1353, w_042_1354, w_042_1355, w_042_1356, w_042_1357, w_042_1358, w_042_1359, w_042_1360, w_042_1361, w_042_1362, w_042_1363, w_042_1364, w_042_1365, w_042_1366, w_042_1367, w_042_1368, w_042_1369, w_042_1370, w_042_1371, w_042_1372, w_042_1373, w_042_1374, w_042_1375, w_042_1376, w_042_1377, w_042_1378, w_042_1379, w_042_1380, w_042_1381, w_042_1382, w_042_1383, w_042_1384, w_042_1385, w_042_1386, w_042_1387, w_042_1388, w_042_1389, w_042_1390, w_042_1391, w_042_1392, w_042_1393, w_042_1394, w_042_1395, w_042_1396, w_042_1397, w_042_1398, w_042_1399, w_042_1400, w_042_1401, w_042_1402, w_042_1403, w_042_1404, w_042_1405, w_042_1406, w_042_1407, w_042_1408, w_042_1409, w_042_1410, w_042_1411, w_042_1412, w_042_1413, w_042_1414, w_042_1416, w_042_1417, w_042_1418, w_042_1419, w_042_1420, w_042_1421, w_042_1422, w_042_1423, w_042_1424, w_042_1425, w_042_1426, w_042_1427, w_042_1428, w_042_1429, w_042_1430, w_042_1431, w_042_1432, w_042_1433, w_042_1434, w_042_1435, w_042_1436, w_042_1437, w_042_1438, w_042_1439, w_042_1440, w_042_1441, w_042_1442, w_042_1443, w_042_1444, w_042_1445, w_042_1446, w_042_1447, w_042_1448, w_042_1449, w_042_1450, w_042_1451, w_042_1452, w_042_1453, w_042_1454, w_042_1455, w_042_1456, w_042_1457, w_042_1458, w_042_1459, w_042_1460, w_042_1461, w_042_1463, w_042_1464, w_042_1465, w_042_1466, w_042_1467, w_042_1468, w_042_1469, w_042_1470, w_042_1471, w_042_1473, w_042_1474, w_042_1475, w_042_1476, w_042_1477, w_042_1479, w_042_1480, w_042_1481, w_042_1482, w_042_1483, w_042_1484, w_042_1485, w_042_1486, w_042_1487, w_042_1488, w_042_1489, w_042_1490, w_042_1491, w_042_1492, w_042_1493, w_042_1494, w_042_1495, w_042_1496, w_042_1497, w_042_1498, w_042_1499, w_042_1500, w_042_1501, w_042_1502, w_042_1503, w_042_1504, w_042_1505, w_042_1506, w_042_1507, w_042_1508, w_042_1509, w_042_1510, w_042_1511, w_042_1512, w_042_1514, w_042_1515, w_042_1516, w_042_1517, w_042_1518, w_042_1519, w_042_1520, w_042_1521, w_042_1522, w_042_1523, w_042_1524, w_042_1525, w_042_1526, w_042_1527, w_042_1528, w_042_1529, w_042_1530, w_042_1531, w_042_1532, w_042_1533, w_042_1534, w_042_1535, w_042_1536, w_042_1537, w_042_1538, w_042_1539, w_042_1540, w_042_1541, w_042_1542, w_042_1543, w_042_1545, w_042_1546, w_042_1547, w_042_1548, w_042_1549, w_042_1550, w_042_1551, w_042_1552, w_042_1553, w_042_1554, w_042_1555, w_042_1556, w_042_1557, w_042_1558, w_042_1559, w_042_1560, w_042_1561, w_042_1562, w_042_1563, w_042_1564, w_042_1565, w_042_1566, w_042_1567, w_042_1568, w_042_1569, w_042_1570, w_042_1571, w_042_1572, w_042_1573, w_042_1574, w_042_1575, w_042_1576, w_042_1577, w_042_1578, w_042_1579, w_042_1580, w_042_1581, w_042_1582, w_042_1584, w_042_1585, w_042_1586, w_042_1587, w_042_1588, w_042_1589, w_042_1590, w_042_1591, w_042_1592, w_042_1593, w_042_1594, w_042_1595, w_042_1596, w_042_1597, w_042_1598, w_042_1599, w_042_1600, w_042_1601, w_042_1602, w_042_1603, w_042_1604, w_042_1605, w_042_1606, w_042_1607, w_042_1608, w_042_1609, w_042_1610, w_042_1611, w_042_1612, w_042_1613, w_042_1614, w_042_1615, w_042_1617, w_042_1619, w_042_1620, w_042_1621, w_042_1622, w_042_1623, w_042_1624, w_042_1625, w_042_1626, w_042_1627, w_042_1628, w_042_1629, w_042_1630, w_042_1631, w_042_1632, w_042_1633, w_042_1634, w_042_1635, w_042_1636, w_042_1637, w_042_1638, w_042_1639, w_042_1640, w_042_1641, w_042_1642, w_042_1643, w_042_1644, w_042_1645, w_042_1646, w_042_1647, w_042_1648, w_042_1649, w_042_1650, w_042_1651, w_042_1652, w_042_1653, w_042_1654, w_042_1655, w_042_1656, w_042_1657, w_042_1658, w_042_1659, w_042_1660, w_042_1661, w_042_1662, w_042_1663, w_042_1664, w_042_1665, w_042_1666, w_042_1667, w_042_1668, w_042_1669, w_042_1670, w_042_1671, w_042_1672, w_042_1673, w_042_1675, w_042_1676, w_042_1677, w_042_1678, w_042_1679, w_042_1680, w_042_1681, w_042_1682, w_042_1683, w_042_1684, w_042_1685, w_042_1687, w_042_1688, w_042_1689, w_042_1690, w_042_1691, w_042_1692, w_042_1693, w_042_1694, w_042_1695, w_042_1696, w_042_1697, w_042_1698, w_042_1699, w_042_1700, w_042_1701, w_042_1702, w_042_1703, w_042_1704, w_042_1705, w_042_1706, w_042_1707, w_042_1708, w_042_1709, w_042_1710, w_042_1711, w_042_1712, w_042_1714, w_042_1715, w_042_1716, w_042_1717, w_042_1718, w_042_1719, w_042_1720, w_042_1721, w_042_1722, w_042_1723, w_042_1724, w_042_1725, w_042_1726, w_042_1727, w_042_1728, w_042_1729, w_042_1730, w_042_1731, w_042_1732, w_042_1733, w_042_1734, w_042_1735, w_042_1736, w_042_1737, w_042_1738, w_042_1739, w_042_1740, w_042_1741, w_042_1742, w_042_1743, w_042_1744, w_042_1745, w_042_1746, w_042_1747, w_042_1748, w_042_1749, w_042_1750, w_042_1751, w_042_1753, w_042_1754, w_042_1755, w_042_1756, w_042_1757, w_042_1759, w_042_1760, w_042_1761, w_042_1762, w_042_1763, w_042_1764, w_042_1765, w_042_1766, w_042_1767, w_042_1769, w_042_1770, w_042_1771, w_042_1772, w_042_1773, w_042_1774, w_042_1775, w_042_1776, w_042_1777, w_042_1778, w_042_1779, w_042_1780, w_042_1781, w_042_1782, w_042_1783, w_042_1784, w_042_1785, w_042_1786, w_042_1787, w_042_1788, w_042_1789, w_042_1790, w_042_1791, w_042_1792, w_042_1793, w_042_1794, w_042_1795, w_042_1796, w_042_1797, w_042_1798, w_042_1799, w_042_1800, w_042_1801, w_042_1802, w_042_1803, w_042_1804, w_042_1805, w_042_1806, w_042_1807, w_042_1808, w_042_1809, w_042_1810, w_042_1811, w_042_1812, w_042_1814, w_042_1815, w_042_1816, w_042_1817, w_042_1818, w_042_1819, w_042_1820, w_042_1821, w_042_1822, w_042_1823, w_042_1824, w_042_1825, w_042_1826, w_042_1827, w_042_1828, w_042_1829, w_042_1830, w_042_1831, w_042_1832, w_042_1833, w_042_1834, w_042_1835, w_042_1836, w_042_1837, w_042_1838, w_042_1839, w_042_1840, w_042_1841, w_042_1842, w_042_1843, w_042_1845, w_042_1847, w_042_1848, w_042_1849, w_042_1850, w_042_1851, w_042_1852, w_042_1853, w_042_1854, w_042_1855, w_042_1856, w_042_1857, w_042_1858, w_042_1859, w_042_1860, w_042_1861, w_042_1862, w_042_1863, w_042_1864, w_042_1866, w_042_1867, w_042_1868, w_042_1869, w_042_1870, w_042_1871, w_042_1872, w_042_1873, w_042_1874, w_042_1875, w_042_1876, w_042_1877, w_042_1878, w_042_1879, w_042_1880, w_042_1881, w_042_1882, w_042_1883, w_042_1884, w_042_1885, w_042_1886, w_042_1887, w_042_1888, w_042_1889, w_042_1890, w_042_1891, w_042_1892, w_042_1893, w_042_1894, w_042_1895, w_042_1896, w_042_1897, w_042_1898, w_042_1899, w_042_1900, w_042_1901, w_042_1902, w_042_1903, w_042_1904, w_042_1905, w_042_1906, w_042_1907, w_042_1908, w_042_1909, w_042_1910, w_042_1911, w_042_1912, w_042_1913, w_042_1914, w_042_1915, w_042_1916, w_042_1917, w_042_1918, w_042_1919, w_042_1920, w_042_1921, w_042_1922, w_042_1923, w_042_1924, w_042_1925, w_042_1926, w_042_1927, w_042_1928, w_042_1929, w_042_1930, w_042_1931, w_042_1932, w_042_1933, w_042_1934, w_042_1935, w_042_1936, w_042_1937, w_042_1938, w_042_1939, w_042_1940, w_042_1941, w_042_1942, w_042_1943, w_042_1944, w_042_1945, w_042_1946, w_042_1947, w_042_1948, w_042_1949, w_042_1950, w_042_1951, w_042_1952, w_042_1953;
  wire w_043_000, w_043_003, w_043_004, w_043_006, w_043_007, w_043_011, w_043_012, w_043_014, w_043_015, w_043_016, w_043_017, w_043_018, w_043_020, w_043_021, w_043_022, w_043_024, w_043_026, w_043_029, w_043_031, w_043_036, w_043_037, w_043_038, w_043_039, w_043_040, w_043_044, w_043_045, w_043_047, w_043_049, w_043_050, w_043_051, w_043_052, w_043_053, w_043_055, w_043_056, w_043_057, w_043_058, w_043_060, w_043_061, w_043_063, w_043_065, w_043_067, w_043_069, w_043_070, w_043_073, w_043_075, w_043_078, w_043_079, w_043_080, w_043_083, w_043_084, w_043_085, w_043_086, w_043_087, w_043_088, w_043_089, w_043_090, w_043_091, w_043_093, w_043_094, w_043_095, w_043_096, w_043_097, w_043_098, w_043_099, w_043_100, w_043_103, w_043_104, w_043_105, w_043_107, w_043_108, w_043_112, w_043_113, w_043_114, w_043_116, w_043_118, w_043_120, w_043_121, w_043_122, w_043_124, w_043_125, w_043_126, w_043_128, w_043_129, w_043_130, w_043_131, w_043_132, w_043_133, w_043_136, w_043_137, w_043_139, w_043_140, w_043_141, w_043_142, w_043_144, w_043_145, w_043_146, w_043_150, w_043_151, w_043_152, w_043_153, w_043_154, w_043_156, w_043_157, w_043_159, w_043_161, w_043_163, w_043_164, w_043_165, w_043_166, w_043_167, w_043_168, w_043_172, w_043_173, w_043_175, w_043_176, w_043_177, w_043_178, w_043_179, w_043_184, w_043_185, w_043_188, w_043_189, w_043_191, w_043_193, w_043_196, w_043_197, w_043_198, w_043_200, w_043_202, w_043_203, w_043_204, w_043_205, w_043_206, w_043_207, w_043_209, w_043_211, w_043_212, w_043_213, w_043_214, w_043_215, w_043_216, w_043_217, w_043_218, w_043_220, w_043_221, w_043_222, w_043_223, w_043_226, w_043_227, w_043_228, w_043_229, w_043_230, w_043_232, w_043_233, w_043_234, w_043_237, w_043_238, w_043_239, w_043_240, w_043_242, w_043_243, w_043_246, w_043_247, w_043_248, w_043_250, w_043_251, w_043_252, w_043_253, w_043_254, w_043_255, w_043_256, w_043_261, w_043_262, w_043_263, w_043_264, w_043_265, w_043_266, w_043_267, w_043_268, w_043_269, w_043_270, w_043_271, w_043_272, w_043_273, w_043_276, w_043_278, w_043_279, w_043_280, w_043_281, w_043_282, w_043_284, w_043_285, w_043_286, w_043_287, w_043_290, w_043_291, w_043_293, w_043_295, w_043_296, w_043_297, w_043_298, w_043_299, w_043_302, w_043_305, w_043_306, w_043_307, w_043_308, w_043_309, w_043_310, w_043_312, w_043_313, w_043_315, w_043_316, w_043_317, w_043_318, w_043_319, w_043_320, w_043_321, w_043_322, w_043_324, w_043_325, w_043_326, w_043_327, w_043_328, w_043_330, w_043_331, w_043_333, w_043_335, w_043_336, w_043_339, w_043_340, w_043_342, w_043_344, w_043_345, w_043_347, w_043_349, w_043_350, w_043_354, w_043_355, w_043_356, w_043_357, w_043_358, w_043_359, w_043_360, w_043_361, w_043_362, w_043_365, w_043_366, w_043_367, w_043_369, w_043_370, w_043_371, w_043_372, w_043_375, w_043_376, w_043_377, w_043_378, w_043_380, w_043_381, w_043_382, w_043_383, w_043_384, w_043_388, w_043_390, w_043_391, w_043_392, w_043_393, w_043_394, w_043_395, w_043_396, w_043_397, w_043_398, w_043_399, w_043_401, w_043_402, w_043_403, w_043_405, w_043_407, w_043_408, w_043_409, w_043_411, w_043_413, w_043_414, w_043_415, w_043_416, w_043_417, w_043_418, w_043_419, w_043_420, w_043_422, w_043_423, w_043_426, w_043_427, w_043_428, w_043_431, w_043_432, w_043_433, w_043_434, w_043_435, w_043_438, w_043_439, w_043_440, w_043_441, w_043_442, w_043_446, w_043_447, w_043_448, w_043_449, w_043_451, w_043_452, w_043_454, w_043_458, w_043_459, w_043_461, w_043_463, w_043_464, w_043_465, w_043_466, w_043_470, w_043_471, w_043_472, w_043_474, w_043_476, w_043_477, w_043_479, w_043_480, w_043_481, w_043_482, w_043_483, w_043_485, w_043_486, w_043_487, w_043_488, w_043_489, w_043_493, w_043_495, w_043_499, w_043_500, w_043_502, w_043_504, w_043_505, w_043_510, w_043_512, w_043_513, w_043_514, w_043_515, w_043_517, w_043_518, w_043_519, w_043_521, w_043_522, w_043_523, w_043_524, w_043_525, w_043_526, w_043_527, w_043_528, w_043_529, w_043_530, w_043_531, w_043_533, w_043_536, w_043_537, w_043_538, w_043_539, w_043_542, w_043_544, w_043_545, w_043_546, w_043_548, w_043_549, w_043_550, w_043_551, w_043_552, w_043_553, w_043_556, w_043_557, w_043_563, w_043_564, w_043_565, w_043_566, w_043_570, w_043_571, w_043_574, w_043_575, w_043_576, w_043_578, w_043_580, w_043_582, w_043_583, w_043_584, w_043_585, w_043_586, w_043_588, w_043_589, w_043_590, w_043_591, w_043_592, w_043_593, w_043_596, w_043_597, w_043_599, w_043_605, w_043_608, w_043_609, w_043_611, w_043_613, w_043_615, w_043_616, w_043_617, w_043_618, w_043_619, w_043_620, w_043_621, w_043_625, w_043_627, w_043_628, w_043_629, w_043_630, w_043_632, w_043_634, w_043_635, w_043_636, w_043_637, w_043_638, w_043_643, w_043_644, w_043_645, w_043_646, w_043_647, w_043_648, w_043_650, w_043_651, w_043_652, w_043_653, w_043_655, w_043_657, w_043_658, w_043_659, w_043_660, w_043_661, w_043_662, w_043_663, w_043_665, w_043_666, w_043_667, w_043_668, w_043_669, w_043_670, w_043_671, w_043_672, w_043_673, w_043_674, w_043_675, w_043_676, w_043_677, w_043_678, w_043_679, w_043_680, w_043_681, w_043_682, w_043_684, w_043_685, w_043_686, w_043_687, w_043_692, w_043_693, w_043_694, w_043_695, w_043_696, w_043_697, w_043_700, w_043_705, w_043_706, w_043_707, w_043_708, w_043_709, w_043_710, w_043_711, w_043_712, w_043_713, w_043_714, w_043_715, w_043_716, w_043_717, w_043_719, w_043_720, w_043_721, w_043_722, w_043_723, w_043_724, w_043_726, w_043_728, w_043_729, w_043_730, w_043_731, w_043_732, w_043_733, w_043_734, w_043_736, w_043_737, w_043_738, w_043_739, w_043_740, w_043_741, w_043_742, w_043_744, w_043_745, w_043_746, w_043_749, w_043_752, w_043_754, w_043_755, w_043_756, w_043_757, w_043_758, w_043_759, w_043_761, w_043_762, w_043_765, w_043_766, w_043_767, w_043_768, w_043_772, w_043_773, w_043_774, w_043_775, w_043_776, w_043_780, w_043_782, w_043_783, w_043_784, w_043_786, w_043_787, w_043_791, w_043_792, w_043_794, w_043_796, w_043_798, w_043_800, w_043_801, w_043_802, w_043_803, w_043_806, w_043_807, w_043_808, w_043_809, w_043_811, w_043_812, w_043_813, w_043_814, w_043_815, w_043_817, w_043_823, w_043_825, w_043_827, w_043_828, w_043_830, w_043_831, w_043_832, w_043_833, w_043_834, w_043_837, w_043_839, w_043_841, w_043_842, w_043_843, w_043_845, w_043_846, w_043_847, w_043_848, w_043_849, w_043_850, w_043_851, w_043_853, w_043_855, w_043_857, w_043_858, w_043_860, w_043_861, w_043_863, w_043_864, w_043_865, w_043_866, w_043_870, w_043_871, w_043_872, w_043_873, w_043_874, w_043_877, w_043_878, w_043_879, w_043_882, w_043_883, w_043_884, w_043_885, w_043_886, w_043_887, w_043_890, w_043_891, w_043_892, w_043_893, w_043_894, w_043_897, w_043_898, w_043_899, w_043_900, w_043_901, w_043_902, w_043_906, w_043_907, w_043_908, w_043_913, w_043_914, w_043_915, w_043_916, w_043_920, w_043_921, w_043_922, w_043_924, w_043_926, w_043_927, w_043_928, w_043_932, w_043_933, w_043_935, w_043_936, w_043_939, w_043_940, w_043_941, w_043_942, w_043_943, w_043_944, w_043_945, w_043_946, w_043_947, w_043_948, w_043_949, w_043_950, w_043_952, w_043_953, w_043_954, w_043_956, w_043_958, w_043_963, w_043_964, w_043_966, w_043_967, w_043_968, w_043_970, w_043_971, w_043_972, w_043_973, w_043_975, w_043_976, w_043_977, w_043_978, w_043_979, w_043_981, w_043_982, w_043_983, w_043_984, w_043_986, w_043_987, w_043_989, w_043_990, w_043_991, w_043_992, w_043_994, w_043_995, w_043_996, w_043_997, w_043_998, w_043_1000, w_043_1001, w_043_1002, w_043_1003, w_043_1004, w_043_1005, w_043_1006, w_043_1008, w_043_1009, w_043_1010, w_043_1011, w_043_1013, w_043_1015, w_043_1016, w_043_1017, w_043_1018, w_043_1019, w_043_1020, w_043_1021, w_043_1022, w_043_1023, w_043_1025, w_043_1026, w_043_1028, w_043_1030, w_043_1032, w_043_1034, w_043_1035, w_043_1036, w_043_1037, w_043_1038, w_043_1039, w_043_1040, w_043_1041, w_043_1043, w_043_1044, w_043_1046, w_043_1047, w_043_1048, w_043_1050, w_043_1051, w_043_1052, w_043_1055, w_043_1056, w_043_1057, w_043_1058, w_043_1062, w_043_1065, w_043_1066, w_043_1067, w_043_1068, w_043_1069, w_043_1070, w_043_1071, w_043_1073, w_043_1077, w_043_1078, w_043_1079, w_043_1080, w_043_1081, w_043_1082, w_043_1083, w_043_1084, w_043_1086, w_043_1087, w_043_1088, w_043_1090, w_043_1091, w_043_1092, w_043_1093, w_043_1094, w_043_1095, w_043_1096, w_043_1097, w_043_1098, w_043_1099, w_043_1100, w_043_1101, w_043_1102, w_043_1103, w_043_1105, w_043_1106, w_043_1107, w_043_1109, w_043_1111, w_043_1112, w_043_1115, w_043_1116, w_043_1119, w_043_1120, w_043_1122, w_043_1126, w_043_1127, w_043_1128, w_043_1129, w_043_1131, w_043_1132, w_043_1133, w_043_1134, w_043_1135, w_043_1136, w_043_1137, w_043_1138, w_043_1139, w_043_1140, w_043_1141, w_043_1144, w_043_1145, w_043_1148, w_043_1149, w_043_1152, w_043_1153, w_043_1155, w_043_1157, w_043_1158, w_043_1160, w_043_1161, w_043_1162, w_043_1163, w_043_1164, w_043_1165, w_043_1166, w_043_1167, w_043_1168, w_043_1169, w_043_1170, w_043_1171, w_043_1172, w_043_1176, w_043_1178, w_043_1180, w_043_1183, w_043_1184, w_043_1185, w_043_1187, w_043_1188, w_043_1189, w_043_1190, w_043_1191, w_043_1192, w_043_1193, w_043_1195, w_043_1196, w_043_1197, w_043_1198, w_043_1199, w_043_1200, w_043_1201, w_043_1203, w_043_1204, w_043_1205, w_043_1206, w_043_1207, w_043_1208, w_043_1209, w_043_1211, w_043_1214, w_043_1215, w_043_1216, w_043_1219, w_043_1221, w_043_1222, w_043_1223, w_043_1224, w_043_1225, w_043_1227, w_043_1228, w_043_1230, w_043_1231, w_043_1232, w_043_1233, w_043_1235, w_043_1236, w_043_1237, w_043_1238, w_043_1240, w_043_1242, w_043_1244, w_043_1245, w_043_1246, w_043_1247, w_043_1249, w_043_1250, w_043_1251, w_043_1252, w_043_1253, w_043_1254, w_043_1255, w_043_1257, w_043_1258, w_043_1259, w_043_1261, w_043_1263, w_043_1264, w_043_1265, w_043_1267, w_043_1268, w_043_1270, w_043_1271, w_043_1272, w_043_1273, w_043_1275, w_043_1276, w_043_1277, w_043_1278, w_043_1279, w_043_1280, w_043_1283, w_043_1284, w_043_1285, w_043_1288, w_043_1289, w_043_1290, w_043_1292, w_043_1293, w_043_1296, w_043_1298, w_043_1300, w_043_1302, w_043_1303, w_043_1305, w_043_1306, w_043_1307, w_043_1309, w_043_1311, w_043_1312, w_043_1313, w_043_1315, w_043_1317, w_043_1318, w_043_1319, w_043_1320, w_043_1322, w_043_1323, w_043_1324, w_043_1326, w_043_1327, w_043_1328, w_043_1330, w_043_1331, w_043_1332, w_043_1333, w_043_1335, w_043_1336, w_043_1337, w_043_1338, w_043_1339, w_043_1340, w_043_1341, w_043_1346, w_043_1347, w_043_1349, w_043_1350, w_043_1351, w_043_1352, w_043_1354, w_043_1355, w_043_1357, w_043_1359, w_043_1360, w_043_1361, w_043_1362, w_043_1363, w_043_1364, w_043_1365, w_043_1366, w_043_1367, w_043_1368, w_043_1369, w_043_1371, w_043_1373, w_043_1374, w_043_1375, w_043_1376, w_043_1377, w_043_1378, w_043_1379, w_043_1380, w_043_1381, w_043_1382, w_043_1383, w_043_1384, w_043_1385, w_043_1388, w_043_1390, w_043_1391, w_043_1392, w_043_1393, w_043_1394, w_043_1395, w_043_1396, w_043_1397, w_043_1399, w_043_1402, w_043_1404, w_043_1408, w_043_1410, w_043_1411, w_043_1412, w_043_1414, w_043_1416, w_043_1418, w_043_1419, w_043_1420, w_043_1421, w_043_1422, w_043_1423, w_043_1424, w_043_1425, w_043_1427, w_043_1428, w_043_1429, w_043_1431, w_043_1433, w_043_1434, w_043_1436, w_043_1437, w_043_1438, w_043_1439, w_043_1440, w_043_1441, w_043_1442, w_043_1443, w_043_1444, w_043_1445, w_043_1446, w_043_1447, w_043_1448, w_043_1450, w_043_1451, w_043_1452, w_043_1454, w_043_1455, w_043_1456, w_043_1457, w_043_1458, w_043_1459, w_043_1460, w_043_1461, w_043_1462, w_043_1463, w_043_1464, w_043_1465, w_043_1466, w_043_1467, w_043_1470, w_043_1471, w_043_1472, w_043_1474, w_043_1476, w_043_1477, w_043_1478, w_043_1479, w_043_1480, w_043_1482, w_043_1483, w_043_1484, w_043_1487, w_043_1488, w_043_1491, w_043_1492, w_043_1493, w_043_1494, w_043_1496, w_043_1497, w_043_1498, w_043_1499, w_043_1500, w_043_1502, w_043_1503, w_043_1504, w_043_1505, w_043_1506, w_043_1507, w_043_1508, w_043_1510, w_043_1512, w_043_1513, w_043_1514, w_043_1515, w_043_1517, w_043_1518, w_043_1520, w_043_1522, w_043_1523, w_043_1524, w_043_1525, w_043_1527, w_043_1528, w_043_1529, w_043_1530, w_043_1531, w_043_1535, w_043_1536, w_043_1537, w_043_1538, w_043_1539, w_043_1540, w_043_1541, w_043_1544, w_043_1545, w_043_1547, w_043_1548, w_043_1549, w_043_1550, w_043_1552, w_043_1553, w_043_1554, w_043_1556, w_043_1558, w_043_1559, w_043_1561, w_043_1562, w_043_1563, w_043_1564, w_043_1565, w_043_1566, w_043_1567, w_043_1569, w_043_1571, w_043_1573, w_043_1574, w_043_1576, w_043_1577, w_043_1578, w_043_1579, w_043_1580, w_043_1581, w_043_1585, w_043_1586, w_043_1587, w_043_1591, w_043_1592, w_043_1593, w_043_1595, w_043_1596, w_043_1599, w_043_1600, w_043_1603, w_043_1604, w_043_1605, w_043_1606, w_043_1608, w_043_1610, w_043_1611, w_043_1612, w_043_1614, w_043_1615, w_043_1617, w_043_1618, w_043_1619, w_043_1620, w_043_1621, w_043_1622, w_043_1623, w_043_1626, w_043_1627, w_043_1628, w_043_1629, w_043_1630, w_043_1631, w_043_1635, w_043_1637, w_043_1638, w_043_1641, w_043_1642, w_043_1643, w_043_1644, w_043_1648, w_043_1649, w_043_1651, w_043_1652, w_043_1653, w_043_1654, w_043_1655, w_043_1656, w_043_1657, w_043_1658, w_043_1659, w_043_1660, w_043_1663, w_043_1664, w_043_1665, w_043_1666, w_043_1668, w_043_1670, w_043_1671, w_043_1672, w_043_1673, w_043_1675, w_043_1676, w_043_1677, w_043_1678, w_043_1679, w_043_1680, w_043_1681, w_043_1682, w_043_1683, w_043_1686, w_043_1687, w_043_1688, w_043_1689, w_043_1690, w_043_1691, w_043_1692, w_043_1693, w_043_1694, w_043_1696, w_043_1699, w_043_1700, w_043_1701, w_043_1702, w_043_1704, w_043_1705, w_043_1706, w_043_1707, w_043_1708, w_043_1709, w_043_1710, w_043_1711, w_043_1712, w_043_1713, w_043_1714, w_043_1715, w_043_1716, w_043_1718, w_043_1719, w_043_1720, w_043_1722, w_043_1723, w_043_1724, w_043_1725, w_043_1726, w_043_1727, w_043_1728, w_043_1729, w_043_1731, w_043_1732, w_043_1734, w_043_1736, w_043_1737, w_043_1738, w_043_1740, w_043_1742, w_043_1744, w_043_1745, w_043_1746, w_043_1747, w_043_1748, w_043_1749, w_043_1750, w_043_1751, w_043_1752, w_043_1753, w_043_1754, w_043_1755, w_043_1757, w_043_1759, w_043_1760, w_043_1761, w_043_1762, w_043_1763, w_043_1764, w_043_1765, w_043_1766, w_043_1767, w_043_1768, w_043_1769, w_043_1770, w_043_1771, w_043_1774, w_043_1775, w_043_1777, w_043_1778, w_043_1781, w_043_1783, w_043_1784, w_043_1785, w_043_1786, w_043_1787, w_043_1788, w_043_1789, w_043_1791, w_043_1793, w_043_1794, w_043_1795, w_043_1796, w_043_1797, w_043_1798, w_043_1799, w_043_1800, w_043_1801, w_043_1803, w_043_1804, w_043_1805, w_043_1806, w_043_1807, w_043_1808, w_043_1809, w_043_1810, w_043_1811, w_043_1813, w_043_1814, w_043_1815, w_043_1816, w_043_1817, w_043_1818, w_043_1819, w_043_1820, w_043_1826, w_043_1827, w_043_1828, w_043_1829, w_043_1833, w_043_1834, w_043_1835, w_043_1836, w_043_1837, w_043_1838, w_043_1842, w_043_1843, w_043_1844, w_043_1846, w_043_1848, w_043_1850, w_043_1851, w_043_1852, w_043_1853, w_043_1854, w_043_1855, w_043_1856, w_043_1858, w_043_1859, w_043_1860, w_043_1861, w_043_1863, w_043_1864, w_043_1865, w_043_1869, w_043_1870, w_043_1871, w_043_1872, w_043_1873, w_043_1874, w_043_1875, w_043_1876, w_043_1880, w_043_1881, w_043_1882, w_043_1885, w_043_1886, w_043_1887, w_043_1889, w_043_1890, w_043_1891, w_043_1892, w_043_1893, w_043_1894, w_043_1896, w_043_1897, w_043_1899, w_043_1901, w_043_1902, w_043_1903, w_043_1904, w_043_1905, w_043_1906, w_043_1907, w_043_1908, w_043_1911, w_043_1912, w_043_1913, w_043_1914, w_043_1915, w_043_1916, w_043_1917, w_043_1920, w_043_1921, w_043_1922, w_043_1923, w_043_1925, w_043_1928, w_043_1929, w_043_1930, w_043_1931, w_043_1933, w_043_1934, w_043_1937, w_043_1938, w_043_1939, w_043_1940, w_043_1941, w_043_1942, w_043_1943, w_043_1944, w_043_1946, w_043_1947, w_043_1948, w_043_1953, w_043_1954, w_043_1955, w_043_1956, w_043_1957, w_043_1959, w_043_1960, w_043_1961, w_043_1962, w_043_1963, w_043_1964, w_043_1965, w_043_1966, w_043_1967, w_043_1968, w_043_1969, w_043_1971, w_043_1972, w_043_1973, w_043_1974, w_043_1976, w_043_1978, w_043_1979, w_043_1980, w_043_1981, w_043_1982, w_043_1983, w_043_1985, w_043_1987, w_043_1988, w_043_1990, w_043_1991, w_043_1992, w_043_1994, w_043_1995, w_043_1996, w_043_1997, w_043_1998, w_043_1999, w_043_2000, w_043_2001, w_043_2003, w_043_2004, w_043_2005, w_043_2006, w_043_2007, w_043_2010, w_043_2012, w_043_2013, w_043_2015, w_043_2016, w_043_2017, w_043_2018, w_043_2019, w_043_2021, w_043_2022, w_043_2024, w_043_2025, w_043_2026, w_043_2027, w_043_2029, w_043_2030, w_043_2032, w_043_2034, w_043_2035, w_043_2036, w_043_2037, w_043_2038, w_043_2040, w_043_2041, w_043_2042, w_043_2043, w_043_2045, w_043_2047, w_043_2049, w_043_2051, w_043_2052, w_043_2053, w_043_2054, w_043_2056, w_043_2057, w_043_2058, w_043_2059, w_043_2060, w_043_2061, w_043_2062, w_043_2063, w_043_2064, w_043_2066, w_043_2068, w_043_2069, w_043_2070, w_043_2071, w_043_2072, w_043_2073, w_043_2074, w_043_2075, w_043_2076, w_043_2078, w_043_2079, w_043_2080, w_043_2082, w_043_2083, w_043_2084, w_043_2085, w_043_2086, w_043_2087, w_043_2088, w_043_2089, w_043_2091, w_043_2093, w_043_2094, w_043_2096, w_043_2098, w_043_2099, w_043_2100, w_043_2101, w_043_2102, w_043_2103, w_043_2104, w_043_2105, w_043_2106, w_043_2107, w_043_2109, w_043_2110, w_043_2111, w_043_2112, w_043_2113, w_043_2114, w_043_2115, w_043_2118, w_043_2119, w_043_2120, w_043_2121, w_043_2122, w_043_2123, w_043_2125, w_043_2126, w_043_2128, w_043_2129, w_043_2130, w_043_2131, w_043_2132, w_043_2133, w_043_2134, w_043_2135, w_043_2136, w_043_2138, w_043_2139, w_043_2140, w_043_2141, w_043_2142, w_043_2143, w_043_2144, w_043_2145, w_043_2146, w_043_2147, w_043_2148, w_043_2149, w_043_2150, w_043_2152, w_043_2153, w_043_2154, w_043_2155, w_043_2156, w_043_2157, w_043_2158, w_043_2161, w_043_2163, w_043_2165, w_043_2166, w_043_2167, w_043_2169, w_043_2171, w_043_2173, w_043_2174, w_043_2176, w_043_2178, w_043_2179, w_043_2180, w_043_2181, w_043_2182, w_043_2183, w_043_2184, w_043_2185, w_043_2186, w_043_2187, w_043_2188, w_043_2189, w_043_2190, w_043_2191, w_043_2192, w_043_2194, w_043_2195, w_043_2197, w_043_2198, w_043_2199, w_043_2200, w_043_2201, w_043_2202, w_043_2203, w_043_2204, w_043_2205, w_043_2207, w_043_2208, w_043_2209, w_043_2210, w_043_2213, w_043_2214, w_043_2215, w_043_2216, w_043_2217, w_043_2218, w_043_2219, w_043_2220, w_043_2221, w_043_2222, w_043_2223, w_043_2225, w_043_2227, w_043_2229, w_043_2230, w_043_2231, w_043_2232, w_043_2233, w_043_2235, w_043_2238, w_043_2239, w_043_2240, w_043_2242, w_043_2243, w_043_2244, w_043_2247, w_043_2248, w_043_2249, w_043_2250, w_043_2252, w_043_2253, w_043_2254, w_043_2255, w_043_2256, w_043_2258, w_043_2259, w_043_2260, w_043_2262, w_043_2264, w_043_2265, w_043_2267, w_043_2270, w_043_2272, w_043_2273, w_043_2274, w_043_2275, w_043_2276, w_043_2277, w_043_2278, w_043_2279, w_043_2280, w_043_2281, w_043_2283, w_043_2285, w_043_2286, w_043_2287, w_043_2289, w_043_2292, w_043_2293, w_043_2295, w_043_2297, w_043_2298, w_043_2300, w_043_2301, w_043_2302, w_043_2303, w_043_2304, w_043_2305, w_043_2306, w_043_2308, w_043_2309, w_043_2310, w_043_2311, w_043_2312, w_043_2313, w_043_2314, w_043_2315, w_043_2316, w_043_2317, w_043_2318, w_043_2320, w_043_2321, w_043_2322, w_043_2323, w_043_2324, w_043_2325, w_043_2326, w_043_2327, w_043_2328, w_043_2334, w_043_2335, w_043_2336, w_043_2338, w_043_2339, w_043_2340, w_043_2341, w_043_2342, w_043_2343, w_043_2344, w_043_2345, w_043_2346, w_043_2347, w_043_2348, w_043_2349, w_043_2350, w_043_2352, w_043_2353, w_043_2354, w_043_2356, w_043_2357, w_043_2358, w_043_2359, w_043_2360, w_043_2361, w_043_2362, w_043_2363, w_043_2364, w_043_2365, w_043_2366, w_043_2367, w_043_2368, w_043_2369, w_043_2370, w_043_2373, w_043_2377, w_043_2378, w_043_2379, w_043_2380, w_043_2381, w_043_2382, w_043_2384, w_043_2385, w_043_2391, w_043_2392, w_043_2394, w_043_2395, w_043_2396, w_043_2397, w_043_2398, w_043_2400, w_043_2401, w_043_2403, w_043_2405, w_043_2406, w_043_2407, w_043_2408, w_043_2409, w_043_2410, w_043_2411, w_043_2412, w_043_2413, w_043_2415, w_043_2418, w_043_2420, w_043_2421, w_043_2423, w_043_2424, w_043_2425, w_043_2426, w_043_2427, w_043_2428, w_043_2429, w_043_2430, w_043_2431, w_043_2432, w_043_2433, w_043_2434, w_043_2435, w_043_2437, w_043_2438, w_043_2439, w_043_2440, w_043_2441, w_043_2442, w_043_2443, w_043_2446, w_043_2447, w_043_2448, w_043_2450, w_043_2451, w_043_2452, w_043_2454, w_043_2455, w_043_2456, w_043_2457, w_043_2459, w_043_2460, w_043_2461, w_043_2462, w_043_2464, w_043_2466, w_043_2468, w_043_2469, w_043_2470, w_043_2471, w_043_2472, w_043_2473, w_043_2475, w_043_2476, w_043_2477, w_043_2479, w_043_2480, w_043_2481, w_043_2482, w_043_2483, w_043_2485, w_043_2486, w_043_2487, w_043_2488, w_043_2489, w_043_2491, w_043_2492, w_043_2493, w_043_2495, w_043_2496, w_043_2498, w_043_2501, w_043_2504, w_043_2506, w_043_2507, w_043_2509, w_043_2513, w_043_2514, w_043_2515, w_043_2516, w_043_2520, w_043_2521, w_043_2523, w_043_2524, w_043_2525, w_043_2526, w_043_2528, w_043_2529, w_043_2530, w_043_2531, w_043_2532, w_043_2533, w_043_2535, w_043_2536, w_043_2538, w_043_2539, w_043_2540, w_043_2543, w_043_2545, w_043_2546, w_043_2547, w_043_2550, w_043_2551, w_043_2552, w_043_2553, w_043_2554, w_043_2555, w_043_2556, w_043_2557, w_043_2558, w_043_2559, w_043_2561, w_043_2562, w_043_2565, w_043_2566, w_043_2568, w_043_2569, w_043_2571, w_043_2574, w_043_2575, w_043_2576, w_043_2577, w_043_2579, w_043_2580, w_043_2581, w_043_2582, w_043_2583, w_043_2584, w_043_2585, w_043_2588, w_043_2589, w_043_2591, w_043_2592, w_043_2593, w_043_2594, w_043_2595, w_043_2597, w_043_2598, w_043_2599, w_043_2601, w_043_2602, w_043_2603, w_043_2604, w_043_2606, w_043_2607, w_043_2608, w_043_2609, w_043_2610, w_043_2611, w_043_2612, w_043_2613, w_043_2614, w_043_2615, w_043_2617, w_043_2618, w_043_2619, w_043_2622, w_043_2623, w_043_2624, w_043_2625, w_043_2626, w_043_2627, w_043_2629, w_043_2630, w_043_2631, w_043_2633, w_043_2634, w_043_2636, w_043_2637, w_043_2638, w_043_2639, w_043_2641, w_043_2644, w_043_2645, w_043_2646, w_043_2648, w_043_2649, w_043_2650, w_043_2651, w_043_2652, w_043_2654, w_043_2655, w_043_2656, w_043_2657, w_043_2658, w_043_2660, w_043_2661, w_043_2662, w_043_2663, w_043_2664, w_043_2665, w_043_2666, w_043_2667, w_043_2668, w_043_2670, w_043_2671, w_043_2672, w_043_2673, w_043_2676, w_043_2677, w_043_2678, w_043_2682, w_043_2685, w_043_2686, w_043_2688, w_043_2690, w_043_2691, w_043_2692, w_043_2693, w_043_2695, w_043_2697, w_043_2698, w_043_2699, w_043_2700, w_043_2701, w_043_2703, w_043_2704, w_043_2705, w_043_2706, w_043_2709, w_043_2710, w_043_2711, w_043_2712, w_043_2713, w_043_2716, w_043_2717, w_043_2718, w_043_2720, w_043_2721, w_043_2723, w_043_2724, w_043_2725, w_043_2726, w_043_2727, w_043_2728, w_043_2729, w_043_2730, w_043_2731, w_043_2734, w_043_2735, w_043_2736, w_043_2737, w_043_2738, w_043_2739, w_043_2741, w_043_2742, w_043_2743, w_043_2744, w_043_2745, w_043_2746, w_043_2747, w_043_2749, w_043_2750, w_043_2751, w_043_2752, w_043_2754, w_043_2755, w_043_2756, w_043_2758, w_043_2760, w_043_2762, w_043_2763, w_043_2765, w_043_2766, w_043_2767, w_043_2768, w_043_2769, w_043_2770, w_043_2772, w_043_2773, w_043_2774, w_043_2775, w_043_2776, w_043_2777, w_043_2778, w_043_2779, w_043_2781, w_043_2782, w_043_2783, w_043_2785, w_043_2786, w_043_2787, w_043_2789, w_043_2790, w_043_2791, w_043_2792, w_043_2793, w_043_2794, w_043_2796, w_043_2799, w_043_2800, w_043_2801, w_043_2802, w_043_2804, w_043_2805, w_043_2811, w_043_2812, w_043_2814, w_043_2817, w_043_2818, w_043_2819, w_043_2820, w_043_2821, w_043_2822, w_043_2824, w_043_2825, w_043_2828, w_043_2829, w_043_2830, w_043_2831, w_043_2832, w_043_2833, w_043_2834, w_043_2836, w_043_2837, w_043_2838, w_043_2839, w_043_2840, w_043_2841, w_043_2842, w_043_2843, w_043_2844, w_043_2845, w_043_2846, w_043_2847, w_043_2849, w_043_2850, w_043_2851, w_043_2852, w_043_2853, w_043_2854, w_043_2856, w_043_2857, w_043_2858, w_043_2859, w_043_2860, w_043_2862, w_043_2863, w_043_2865, w_043_2867, w_043_2868, w_043_2869, w_043_2870, w_043_2872, w_043_2873, w_043_2874, w_043_2876, w_043_2878, w_043_2879, w_043_2881, w_043_2882, w_043_2884, w_043_2885, w_043_2886, w_043_2888, w_043_2889, w_043_2890, w_043_2891, w_043_2892, w_043_2893, w_043_2894, w_043_2895, w_043_2896, w_043_2897, w_043_2898, w_043_2899, w_043_2900, w_043_2901, w_043_2903, w_043_2904, w_043_2907, w_043_2908, w_043_2909, w_043_2910, w_043_2911, w_043_2913, w_043_2914, w_043_2915, w_043_2916, w_043_2917, w_043_2918, w_043_2920, w_043_2922, w_043_2924, w_043_2925, w_043_2927, w_043_2928, w_043_2929, w_043_2930, w_043_2932, w_043_2933, w_043_2935, w_043_2936, w_043_2937, w_043_2938, w_043_2939, w_043_2940, w_043_2941, w_043_2942, w_043_2944, w_043_2945, w_043_2946, w_043_2947, w_043_2948, w_043_2949, w_043_2950, w_043_2951, w_043_2952, w_043_2953, w_043_2954, w_043_2957, w_043_2958, w_043_2959, w_043_2960, w_043_2961, w_043_2963, w_043_2965, w_043_2966, w_043_2967, w_043_2969, w_043_2971, w_043_2972, w_043_2973, w_043_2974, w_043_2975, w_043_2976, w_043_2977, w_043_2978, w_043_2979, w_043_2980, w_043_2981, w_043_2983, w_043_2985, w_043_2986, w_043_2988, w_043_2989, w_043_2990, w_043_2992, w_043_2994, w_043_2995, w_043_3001, w_043_3002, w_043_3003, w_043_3004, w_043_3005, w_043_3006, w_043_3007, w_043_3008, w_043_3009, w_043_3011, w_043_3012, w_043_3014, w_043_3015, w_043_3017, w_043_3019, w_043_3022, w_043_3024, w_043_3026, w_043_3027, w_043_3028, w_043_3029, w_043_3030, w_043_3031, w_043_3032, w_043_3033, w_043_3034, w_043_3035, w_043_3036, w_043_3037, w_043_3038, w_043_3040, w_043_3041, w_043_3042, w_043_3043, w_043_3044, w_043_3046, w_043_3047, w_043_3048, w_043_3050, w_043_3051, w_043_3054, w_043_3057, w_043_3058, w_043_3059, w_043_3061, w_043_3062, w_043_3063, w_043_3064, w_043_3066, w_043_3067, w_043_3068, w_043_3070, w_043_3071, w_043_3072, w_043_3074, w_043_3075, w_043_3076, w_043_3077, w_043_3078, w_043_3079, w_043_3084, w_043_3086, w_043_3087, w_043_3089, w_043_3090, w_043_3091, w_043_3092, w_043_3094, w_043_3096, w_043_3097, w_043_3098, w_043_3099, w_043_3101, w_043_3102, w_043_3104, w_043_3108, w_043_3109, w_043_3110, w_043_3111, w_043_3117, w_043_3118, w_043_3119, w_043_3120, w_043_3121, w_043_3122, w_043_3123, w_043_3124, w_043_3125, w_043_3126, w_043_3127, w_043_3129, w_043_3130, w_043_3131, w_043_3132, w_043_3133, w_043_3134, w_043_3136, w_043_3137, w_043_3138, w_043_3140, w_043_3141, w_043_3142, w_043_3145, w_043_3146, w_043_3148, w_043_3149, w_043_3150, w_043_3151, w_043_3152, w_043_3154, w_043_3155, w_043_3158, w_043_3159, w_043_3160, w_043_3161, w_043_3165, w_043_3166, w_043_3167, w_043_3169, w_043_3170, w_043_3171, w_043_3172, w_043_3173, w_043_3174, w_043_3175, w_043_3176, w_043_3177, w_043_3178, w_043_3179, w_043_3181, w_043_3182, w_043_3183, w_043_3185, w_043_3187, w_043_3188, w_043_3189, w_043_3190, w_043_3191, w_043_3192, w_043_3193, w_043_3195, w_043_3196, w_043_3197, w_043_3198, w_043_3199, w_043_3200, w_043_3201, w_043_3205, w_043_3206, w_043_3207, w_043_3208, w_043_3212, w_043_3213, w_043_3216, w_043_3218, w_043_3220, w_043_3221, w_043_3224, w_043_3225, w_043_3226, w_043_3227, w_043_3228, w_043_3229, w_043_3230, w_043_3231, w_043_3232, w_043_3233, w_043_3234, w_043_3235, w_043_3237, w_043_3239, w_043_3241, w_043_3242, w_043_3244, w_043_3245, w_043_3247, w_043_3249, w_043_3250, w_043_3252, w_043_3253, w_043_3254, w_043_3255, w_043_3256, w_043_3257, w_043_3258, w_043_3259, w_043_3260, w_043_3261, w_043_3262, w_043_3263, w_043_3265, w_043_3266, w_043_3268, w_043_3269, w_043_3271, w_043_3272, w_043_3273, w_043_3274, w_043_3275, w_043_3276, w_043_3277, w_043_3278, w_043_3279, w_043_3282, w_043_3283, w_043_3285, w_043_3286, w_043_3287, w_043_3289, w_043_3291, w_043_3293, w_043_3294, w_043_3296, w_043_3297, w_043_3298, w_043_3299, w_043_3300, w_043_3301, w_043_3302, w_043_3303, w_043_3304, w_043_3306, w_043_3308, w_043_3309, w_043_3310, w_043_3311, w_043_3312, w_043_3314, w_043_3315, w_043_3316, w_043_3318, w_043_3319, w_043_3320, w_043_3322, w_043_3323, w_043_3325, w_043_3326, w_043_3328, w_043_3329, w_043_3331, w_043_3332, w_043_3333, w_043_3335, w_043_3336, w_043_3337, w_043_3340, w_043_3341, w_043_3343, w_043_3345, w_043_3346, w_043_3347, w_043_3348, w_043_3351, w_043_3352, w_043_3353, w_043_3354, w_043_3355, w_043_3357, w_043_3360, w_043_3361, w_043_3363, w_043_3365, w_043_3366, w_043_3367, w_043_3368, w_043_3369, w_043_3371, w_043_3373, w_043_3374, w_043_3375, w_043_3376, w_043_3378, w_043_3379, w_043_3380, w_043_3381, w_043_3382, w_043_3384, w_043_3386, w_043_3387, w_043_3388, w_043_3389, w_043_3390, w_043_3391, w_043_3392, w_043_3393, w_043_3395, w_043_3396, w_043_3397, w_043_3399, w_043_3401, w_043_3405, w_043_3406, w_043_3407, w_043_3408, w_043_3409, w_043_3410, w_043_3411, w_043_3412, w_043_3415, w_043_3417, w_043_3418, w_043_3420, w_043_3422, w_043_3423, w_043_3424, w_043_3425, w_043_3426, w_043_3427, w_043_3428, w_043_3430, w_043_3431, w_043_3432, w_043_3434, w_043_3435, w_043_3436, w_043_3437, w_043_3438, w_043_3439, w_043_3440, w_043_3441, w_043_3442, w_043_3443, w_043_3445, w_043_3446, w_043_3447, w_043_3448, w_043_3450, w_043_3451, w_043_3452, w_043_3453, w_043_3454, w_043_3455, w_043_3456, w_043_3457, w_043_3458, w_043_3459, w_043_3460, w_043_3463, w_043_3464, w_043_3465, w_043_3467, w_043_3469, w_043_3470, w_043_3471, w_043_3472, w_043_3473, w_043_3474, w_043_3475, w_043_3476, w_043_3477, w_043_3478, w_043_3479, w_043_3480, w_043_3483, w_043_3486, w_043_3487, w_043_3488, w_043_3489, w_043_3490, w_043_3492, w_043_3493, w_043_3495, w_043_3496, w_043_3497, w_043_3499, w_043_3500, w_043_3501, w_043_3504, w_043_3506, w_043_3508, w_043_3509, w_043_3510, w_043_3511, w_043_3513, w_043_3514, w_043_3515, w_043_3516, w_043_3518, w_043_3519, w_043_3520, w_043_3521, w_043_3522, w_043_3523, w_043_3525, w_043_3526, w_043_3528, w_043_3529, w_043_3530, w_043_3531, w_043_3532, w_043_3533, w_043_3534, w_043_3535, w_043_3536, w_043_3537, w_043_3538, w_043_3539, w_043_3541, w_043_3543, w_043_3544, w_043_3546, w_043_3547, w_043_3549, w_043_3550, w_043_3551, w_043_3552, w_043_3553, w_043_3554, w_043_3555, w_043_3556, w_043_3557, w_043_3559, w_043_3560, w_043_3562, w_043_3563, w_043_3564, w_043_3565, w_043_3568, w_043_3569, w_043_3571, w_043_3573, w_043_3574, w_043_3575, w_043_3576, w_043_3577, w_043_3578, w_043_3579, w_043_3582, w_043_3583, w_043_3584, w_043_3586, w_043_3587, w_043_3588, w_043_3591, w_043_3592, w_043_3593, w_043_3594, w_043_3595, w_043_3596, w_043_3598, w_043_3599, w_043_3600, w_043_3601, w_043_3603, w_043_3605, w_043_3606, w_043_3607, w_043_3608, w_043_3609, w_043_3610, w_043_3611, w_043_3612, w_043_3614, w_043_3615, w_043_3616, w_043_3617, w_043_3619, w_043_3620, w_043_3621, w_043_3625, w_043_3626, w_043_3627, w_043_3628, w_043_3629, w_043_3630, w_043_3632, w_043_3633, w_043_3634, w_043_3635, w_043_3636, w_043_3638, w_043_3639, w_043_3640, w_043_3641, w_043_3642, w_043_3643, w_043_3644, w_043_3645, w_043_3646, w_043_3647, w_043_3648, w_043_3650, w_043_3651, w_043_3656, w_043_3657, w_043_3658, w_043_3659, w_043_3660, w_043_3662, w_043_3663, w_043_3664, w_043_3667, w_043_3670, w_043_3671, w_043_3672, w_043_3674, w_043_3675, w_043_3678, w_043_3679, w_043_3680, w_043_3681, w_043_3682, w_043_3683, w_043_3684, w_043_3685, w_043_3686, w_043_3687, w_043_3690, w_043_3691, w_043_3692, w_043_3693, w_043_3695, w_043_3697, w_043_3699, w_043_3700, w_043_3701, w_043_3703, w_043_3704, w_043_3705, w_043_3706, w_043_3707, w_043_3708, w_043_3709, w_043_3713, w_043_3714, w_043_3716, w_043_3717, w_043_3718, w_043_3719, w_043_3720, w_043_3721, w_043_3722, w_043_3723, w_043_3724, w_043_3727, w_043_3728, w_043_3729, w_043_3730, w_043_3732, w_043_3733, w_043_3734, w_043_3735, w_043_3736, w_043_3737, w_043_3738, w_043_3739, w_043_3740, w_043_3741, w_043_3742, w_043_3743, w_043_3745, w_043_3746, w_043_3747, w_043_3749, w_043_3750, w_043_3751, w_043_3753, w_043_3756, w_043_3760, w_043_3761, w_043_3763, w_043_3767, w_043_3768, w_043_3769, w_043_3770, w_043_3771, w_043_3772, w_043_3774, w_043_3775, w_043_3776, w_043_3777, w_043_3779, w_043_3780, w_043_3781, w_043_3782, w_043_3783, w_043_3785, w_043_3786, w_043_3788, w_043_3789, w_043_3792, w_043_3793, w_043_3794, w_043_3796, w_043_3797, w_043_3798, w_043_3799, w_043_3800, w_043_3801, w_043_3806, w_043_3807, w_043_3809, w_043_3811, w_043_3813, w_043_3814, w_043_3815, w_043_3816, w_043_3817, w_043_3818, w_043_3819, w_043_3821, w_043_3822, w_043_3823, w_043_3824, w_043_3825, w_043_3827, w_043_3828, w_043_3830, w_043_3831, w_043_3832, w_043_3833, w_043_3834, w_043_3835, w_043_3836, w_043_3837, w_043_3839, w_043_3841, w_043_3842, w_043_3845, w_043_3846, w_043_3847, w_043_3848, w_043_3849, w_043_3850, w_043_3852, w_043_3853, w_043_3854, w_043_3855, w_043_3856, w_043_3858, w_043_3859, w_043_3860, w_043_3862, w_043_3863, w_043_3864, w_043_3866, w_043_3868, w_043_3869, w_043_3871, w_043_3872, w_043_3874, w_043_3875, w_043_3876, w_043_3877, w_043_3878, w_043_3880, w_043_3881, w_043_3883, w_043_3885, w_043_3886, w_043_3891, w_043_3893, w_043_3894, w_043_3896, w_043_3897, w_043_3898, w_043_3903, w_043_3904, w_043_3905, w_043_3906, w_043_3907, w_043_3908, w_043_3909, w_043_3910, w_043_3911, w_043_3916, w_043_3919, w_043_3921, w_043_3922, w_043_3923, w_043_3924, w_043_3925, w_043_3926, w_043_3928, w_043_3929, w_043_3935, w_043_3938, w_043_3939, w_043_3940, w_043_3941, w_043_3946, w_043_3949, w_043_3951, w_043_3954, w_043_3958, w_043_3962, w_043_3964, w_043_3968, w_043_3973, w_043_3975, w_043_3976, w_043_3977, w_043_3981, w_043_3983, w_043_3985, w_043_3988, w_043_3989, w_043_3991, w_043_3992, w_043_3995, w_043_3996, w_043_3998, w_043_4002, w_043_4006, w_043_4007, w_043_4008, w_043_4010, w_043_4012, w_043_4014, w_043_4015, w_043_4018, w_043_4020, w_043_4025, w_043_4026, w_043_4027, w_043_4030, w_043_4031, w_043_4036, w_043_4038, w_043_4039, w_043_4041, w_043_4044, w_043_4045, w_043_4050, w_043_4051, w_043_4055, w_043_4059, w_043_4060, w_043_4065, w_043_4067, w_043_4068, w_043_4071, w_043_4072, w_043_4073, w_043_4077, w_043_4081, w_043_4083, w_043_4084, w_043_4088, w_043_4090, w_043_4091, w_043_4094, w_043_4095, w_043_4096, w_043_4098, w_043_4099, w_043_4100, w_043_4102, w_043_4104, w_043_4107, w_043_4109, w_043_4110, w_043_4111, w_043_4113, w_043_4114, w_043_4115, w_043_4120, w_043_4122, w_043_4123, w_043_4124, w_043_4126, w_043_4127, w_043_4128, w_043_4130, w_043_4134, w_043_4139, w_043_4141, w_043_4142, w_043_4145, w_043_4147, w_043_4150, w_043_4151, w_043_4154, w_043_4155, w_043_4157, w_043_4160, w_043_4164, w_043_4167, w_043_4168, w_043_4169, w_043_4171, w_043_4175, w_043_4177, w_043_4178, w_043_4179, w_043_4184, w_043_4186, w_043_4187, w_043_4194, w_043_4198, w_043_4199, w_043_4201, w_043_4209, w_043_4211, w_043_4213, w_043_4215, w_043_4217, w_043_4218, w_043_4219, w_043_4222, w_043_4223, w_043_4227, w_043_4228, w_043_4234, w_043_4235, w_043_4241, w_043_4242, w_043_4244, w_043_4246, w_043_4250, w_043_4252, w_043_4257, w_043_4258, w_043_4261, w_043_4273, w_043_4276, w_043_4282, w_043_4283, w_043_4284, w_043_4285, w_043_4287, w_043_4289, w_043_4290, w_043_4292, w_043_4293, w_043_4294, w_043_4296, w_043_4297, w_043_4298, w_043_4299, w_043_4303, w_043_4304, w_043_4309, w_043_4310, w_043_4312, w_043_4314, w_043_4315, w_043_4316, w_043_4318, w_043_4320, w_043_4324, w_043_4330, w_043_4332, w_043_4333, w_043_4335, w_043_4337, w_043_4339, w_043_4341, w_043_4344, w_043_4346, w_043_4348, w_043_4349, w_043_4350, w_043_4353, w_043_4355, w_043_4359, w_043_4362, w_043_4366, w_043_4367, w_043_4368, w_043_4370, w_043_4372, w_043_4374, w_043_4375, w_043_4377, w_043_4378, w_043_4379, w_043_4384, w_043_4388, w_043_4389, w_043_4393, w_043_4394, w_043_4396, w_043_4399, w_043_4400, w_043_4401, w_043_4404, w_043_4407, w_043_4408, w_043_4411, w_043_4412, w_043_4417, w_043_4418, w_043_4419, w_043_4423, w_043_4425, w_043_4426, w_043_4434, w_043_4436, w_043_4437, w_043_4444, w_043_4450, w_043_4451, w_043_4452, w_043_4454, w_043_4456, w_043_4458, w_043_4460, w_043_4463, w_043_4464, w_043_4466, w_043_4467, w_043_4471, w_043_4472, w_043_4473, w_043_4475, w_043_4476, w_043_4479, w_043_4480, w_043_4484, w_043_4485, w_043_4486, w_043_4488, w_043_4489, w_043_4490, w_043_4497, w_043_4499, w_043_4502, w_043_4506, w_043_4508, w_043_4510, w_043_4512, w_043_4513, w_043_4514, w_043_4517, w_043_4518, w_043_4520, w_043_4523, w_043_4524, w_043_4526, w_043_4527, w_043_4530, w_043_4531, w_043_4532, w_043_4534, w_043_4535, w_043_4538, w_043_4540, w_043_4542, w_043_4543, w_043_4544, w_043_4545, w_043_4546, w_043_4549, w_043_4550, w_043_4551, w_043_4553, w_043_4555, w_043_4556, w_043_4557, w_043_4558, w_043_4559, w_043_4560, w_043_4561, w_043_4562, w_043_4564, w_043_4565, w_043_4566, w_043_4570, w_043_4572, w_043_4576, w_043_4579, w_043_4580, w_043_4581, w_043_4582, w_043_4584, w_043_4585, w_043_4586, w_043_4588, w_043_4591, w_043_4594, w_043_4595, w_043_4597, w_043_4598, w_043_4600, w_043_4604, w_043_4605, w_043_4606, w_043_4607, w_043_4608, w_043_4611, w_043_4614, w_043_4616, w_043_4617, w_043_4619, w_043_4620, w_043_4623, w_043_4624, w_043_4628, w_043_4630, w_043_4634, w_043_4635, w_043_4636, w_043_4638, w_043_4639, w_043_4642, w_043_4644, w_043_4645, w_043_4646, w_043_4647, w_043_4650, w_043_4653, w_043_4655, w_043_4658, w_043_4663, w_043_4665, w_043_4666, w_043_4669, w_043_4671, w_043_4672, w_043_4673, w_043_4677, w_043_4678, w_043_4682, w_043_4683, w_043_4685, w_043_4687, w_043_4692, w_043_4694, w_043_4695, w_043_4697, w_043_4698, w_043_4699, w_043_4700, w_043_4701, w_043_4702, w_043_4703, w_043_4704, w_043_4706, w_043_4707, w_043_4708, w_043_4710, w_043_4712, w_043_4715, w_043_4717, w_043_4724, w_043_4725, w_043_4727, w_043_4730, w_043_4732, w_043_4737, w_043_4738, w_043_4739, w_043_4743, w_043_4744, w_043_4745, w_043_4747, w_043_4753, w_043_4755, w_043_4757, w_043_4759, w_043_4762, w_043_4765, w_043_4766, w_043_4767, w_043_4768, w_043_4770, w_043_4773, w_043_4774, w_043_4779, w_043_4780, w_043_4781, w_043_4784, w_043_4785, w_043_4786, w_043_4798, w_043_4802, w_043_4803, w_043_4806, w_043_4808, w_043_4811, w_043_4812, w_043_4814, w_043_4815, w_043_4816, w_043_4821, w_043_4823, w_043_4825, w_043_4826, w_043_4828, w_043_4834, w_043_4838, w_043_4839, w_043_4848, w_043_4851, w_043_4852, w_043_4853, w_043_4854, w_043_4855, w_043_4856, w_043_4857, w_043_4861, w_043_4862, w_043_4863, w_043_4864, w_043_4865, w_043_4866, w_043_4867, w_043_4868, w_043_4871, w_043_4875, w_043_4880, w_043_4882, w_043_4883, w_043_4884, w_043_4887, w_043_4889, w_043_4890, w_043_4891, w_043_4894, w_043_4895, w_043_4899, w_043_4903, w_043_4908, w_043_4909, w_043_4911, w_043_4913, w_043_4914, w_043_4916, w_043_4920, w_043_4921, w_043_4922, w_043_4923, w_043_4924, w_043_4925, w_043_4927, w_043_4928, w_043_4929, w_043_4935, w_043_4937, w_043_4941, w_043_4942, w_043_4944, w_043_4949, w_043_4954, w_043_4955, w_043_4956, w_043_4958, w_043_4959, w_043_4963, w_043_4964, w_043_4967, w_043_4971, w_043_4973, w_043_4979, w_043_4982, w_043_4983, w_043_4985, w_043_4987, w_043_4989, w_043_4991, w_043_4992, w_043_4993, w_043_4994, w_043_4996, w_043_4997, w_043_4998, w_043_4999, w_043_5000, w_043_5004, w_043_5005, w_043_5009, w_043_5012, w_043_5013, w_043_5014, w_043_5016, w_043_5017, w_043_5019, w_043_5021, w_043_5025, w_043_5026, w_043_5027, w_043_5033, w_043_5034, w_043_5035, w_043_5038, w_043_5039, w_043_5045, w_043_5047, w_043_5048, w_043_5049, w_043_5051, w_043_5052, w_043_5053, w_043_5054, w_043_5059, w_043_5061, w_043_5066, w_043_5072, w_043_5073, w_043_5074, w_043_5075, w_043_5076, w_043_5077, w_043_5079, w_043_5085, w_043_5086, w_043_5087, w_043_5089, w_043_5090, w_043_5092, w_043_5094, w_043_5095, w_043_5097, w_043_5098, w_043_5100, w_043_5102, w_043_5104, w_043_5105, w_043_5108, w_043_5109, w_043_5111, w_043_5112, w_043_5113, w_043_5115, w_043_5117, w_043_5121, w_043_5123, w_043_5124, w_043_5126, w_043_5127, w_043_5128, w_043_5129, w_043_5130, w_043_5131, w_043_5135, w_043_5136, w_043_5137, w_043_5138, w_043_5139, w_043_5141, w_043_5142, w_043_5143, w_043_5145, w_043_5146, w_043_5150, w_043_5151, w_043_5156, w_043_5158, w_043_5161, w_043_5162, w_043_5164, w_043_5168, w_043_5169, w_043_5171, w_043_5173, w_043_5174, w_043_5176, w_043_5177, w_043_5178, w_043_5180, w_043_5183, w_043_5185, w_043_5192, w_043_5193, w_043_5194, w_043_5200, w_043_5202, w_043_5204, w_043_5205, w_043_5208, w_043_5212, w_043_5213, w_043_5214, w_043_5217, w_043_5218, w_043_5219, w_043_5222, w_043_5225, w_043_5227, w_043_5229, w_043_5231, w_043_5236, w_043_5238, w_043_5239, w_043_5240, w_043_5242, w_043_5243, w_043_5244, w_043_5246, w_043_5248, w_043_5251, w_043_5253, w_043_5254, w_043_5255, w_043_5256, w_043_5260, w_043_5263, w_043_5265, w_043_5266, w_043_5269, w_043_5275, w_043_5276, w_043_5280, w_043_5285, w_043_5290, w_043_5291, w_043_5294, w_043_5296, w_043_5297, w_043_5302, w_043_5305, w_043_5307, w_043_5308, w_043_5310, w_043_5313, w_043_5318, w_043_5321, w_043_5323, w_043_5324, w_043_5325, w_043_5326, w_043_5329, w_043_5330, w_043_5332, w_043_5343, w_043_5345, w_043_5351, w_043_5352, w_043_5353, w_043_5357, w_043_5358, w_043_5359, w_043_5362, w_043_5365, w_043_5366, w_043_5371, w_043_5372, w_043_5373, w_043_5375, w_043_5376, w_043_5377, w_043_5379, w_043_5384, w_043_5387, w_043_5388, w_043_5390, w_043_5391, w_043_5393, w_043_5394, w_043_5395, w_043_5396, w_043_5398, w_043_5399, w_043_5400, w_043_5402, w_043_5405, w_043_5406, w_043_5407, w_043_5411, w_043_5413, w_043_5414, w_043_5416, w_043_5417, w_043_5418, w_043_5419, w_043_5421, w_043_5423, w_043_5424, w_043_5426, w_043_5427, w_043_5438, w_043_5440, w_043_5445, w_043_5446, w_043_5449, w_043_5453, w_043_5454, w_043_5457, w_043_5460, w_043_5461, w_043_5462, w_043_5463, w_043_5465, w_043_5466, w_043_5468, w_043_5470, w_043_5472, w_043_5476, w_043_5478, w_043_5481, w_043_5486, w_043_5489, w_043_5496, w_043_5497, w_043_5498, w_043_5499, w_043_5500, w_043_5501, w_043_5503, w_043_5504, w_043_5505, w_043_5506, w_043_5507, w_043_5508, w_043_5513, w_043_5514, w_043_5516, w_043_5519, w_043_5520, w_043_5521, w_043_5524, w_043_5525, w_043_5533, w_043_5534, w_043_5535, w_043_5538, w_043_5539, w_043_5541, w_043_5544, w_043_5550, w_043_5551, w_043_5552, w_043_5553, w_043_5555, w_043_5559, w_043_5562, w_043_5565, w_043_5568, w_043_5579, w_043_5580, w_043_5581, w_043_5587, w_043_5589, w_043_5591, w_043_5594, w_043_5595, w_043_5598, w_043_5599, w_043_5601, w_043_5602, w_043_5603, w_043_5604, w_043_5605, w_043_5607, w_043_5610, w_043_5611, w_043_5613, w_043_5616, w_043_5618, w_043_5619, w_043_5621, w_043_5622, w_043_5624, w_043_5625, w_043_5626, w_043_5627, w_043_5628, w_043_5630, w_043_5631, w_043_5633, w_043_5636, w_043_5638, w_043_5640, w_043_5642, w_043_5643, w_043_5646, w_043_5647, w_043_5649, w_043_5650, w_043_5652, w_043_5654, w_043_5655, w_043_5656, w_043_5659, w_043_5660, w_043_5662, w_043_5663, w_043_5664, w_043_5666, w_043_5667, w_043_5668, w_043_5669, w_043_5670, w_043_5672, w_043_5674, w_043_5676, w_043_5680, w_043_5681, w_043_5682, w_043_5685, w_043_5686, w_043_5687, w_043_5691, w_043_5695, w_043_5703, w_043_5704, w_043_5708, w_043_5710, w_043_5713, w_043_5717, w_043_5721, w_043_5727, w_043_5734, w_043_5736, w_043_5738, w_043_5740, w_043_5741, w_043_5742, w_043_5744, w_043_5746, w_043_5749, w_043_5750, w_043_5753, w_043_5759, w_043_5761, w_043_5763, w_043_5765, w_043_5766, w_043_5769, w_043_5770, w_043_5771, w_043_5772, w_043_5773, w_043_5774, w_043_5778, w_043_5779, w_043_5781, w_043_5784, w_043_5785, w_043_5788, w_043_5789, w_043_5796, w_043_5798, w_043_5799, w_043_5800, w_043_5802, w_043_5803, w_043_5805, w_043_5806, w_043_5810, w_043_5811, w_043_5816, w_043_5819, w_043_5825, w_043_5826, w_043_5827, w_043_5828, w_043_5829, w_043_5831, w_043_5832, w_043_5836, w_043_5843, w_043_5844, w_043_5845, w_043_5847, w_043_5848, w_043_5849, w_043_5853, w_043_5854, w_043_5856, w_043_5857, w_043_5859, w_043_5860, w_043_5863, w_043_5864, w_043_5868, w_043_5869, w_043_5871, w_043_5872, w_043_5873, w_043_5879, w_043_5880, w_043_5881, w_043_5882, w_043_5886, w_043_5887, w_043_5891, w_043_5894, w_043_5895, w_043_5896, w_043_5899, w_043_5902, w_043_5905, w_043_5907, w_043_5910, w_043_5912, w_043_5917, w_043_5922, w_043_5923, w_043_5924, w_043_5928, w_043_5929, w_043_5931, w_043_5934, w_043_5936, w_043_5938, w_043_5941, w_043_5943, w_043_5947, w_043_5950, w_043_5953, w_043_5954, w_043_5955, w_043_5956, w_043_5957, w_043_5960, w_043_5961, w_043_5962, w_043_5963, w_043_5966, w_043_5967, w_043_5969, w_043_5972, w_043_5973, w_043_5978, w_043_5979, w_043_5984, w_043_5986, w_043_5987, w_043_5988, w_043_5990, w_043_5993, w_043_5994, w_043_5995, w_043_5998, w_043_5999, w_043_6002, w_043_6005, w_043_6013, w_043_6014, w_043_6016, w_043_6017, w_043_6018, w_043_6019, w_043_6020, w_043_6023, w_043_6024, w_043_6026, w_043_6029, w_043_6031, w_043_6033, w_043_6034, w_043_6035, w_043_6038, w_043_6039, w_043_6041, w_043_6042, w_043_6043, w_043_6044, w_043_6045, w_043_6048, w_043_6050, w_043_6054, w_043_6055, w_043_6058, w_043_6062, w_043_6065, w_043_6066, w_043_6069, w_043_6070, w_043_6071, w_043_6072, w_043_6073, w_043_6075, w_043_6076, w_043_6082, w_043_6084;
  wire w_044_000, w_044_001, w_044_002, w_044_003, w_044_004, w_044_006, w_044_008, w_044_011, w_044_013, w_044_014, w_044_015, w_044_017, w_044_018, w_044_020, w_044_021, w_044_022, w_044_023, w_044_024, w_044_025, w_044_026, w_044_027, w_044_029, w_044_032, w_044_034, w_044_035, w_044_037, w_044_038, w_044_040, w_044_043, w_044_044, w_044_045, w_044_046, w_044_047, w_044_048, w_044_052, w_044_054, w_044_055, w_044_056, w_044_057, w_044_058, w_044_059, w_044_060, w_044_061, w_044_063, w_044_065, w_044_066, w_044_067, w_044_068, w_044_070, w_044_072, w_044_074, w_044_075, w_044_077, w_044_078, w_044_080, w_044_081, w_044_082, w_044_083, w_044_084, w_044_085, w_044_086, w_044_087, w_044_089, w_044_091, w_044_093, w_044_094, w_044_100, w_044_101, w_044_102, w_044_104, w_044_105, w_044_106, w_044_108, w_044_109, w_044_110, w_044_111, w_044_112, w_044_113, w_044_114, w_044_115, w_044_118, w_044_122, w_044_123, w_044_124, w_044_125, w_044_126, w_044_127, w_044_128, w_044_129, w_044_130, w_044_131, w_044_132, w_044_133, w_044_135, w_044_137, w_044_138, w_044_140, w_044_142, w_044_143, w_044_144, w_044_145, w_044_146, w_044_148, w_044_149, w_044_150, w_044_151, w_044_152, w_044_154, w_044_155, w_044_157, w_044_158, w_044_159, w_044_162, w_044_163, w_044_164, w_044_166, w_044_167, w_044_168, w_044_170, w_044_171, w_044_172, w_044_173, w_044_174, w_044_175, w_044_176, w_044_177, w_044_178, w_044_181, w_044_182, w_044_183, w_044_184, w_044_187, w_044_188, w_044_190, w_044_191, w_044_193, w_044_195, w_044_196, w_044_198, w_044_201, w_044_202, w_044_207, w_044_208, w_044_209, w_044_211, w_044_213, w_044_214, w_044_215, w_044_216, w_044_217, w_044_218, w_044_219, w_044_220, w_044_221, w_044_222, w_044_226, w_044_227, w_044_229, w_044_230, w_044_231, w_044_232, w_044_233, w_044_234, w_044_235, w_044_236, w_044_237, w_044_238, w_044_239, w_044_240, w_044_241, w_044_242, w_044_244, w_044_245, w_044_248, w_044_249, w_044_250, w_044_252, w_044_253, w_044_254, w_044_255, w_044_258, w_044_259, w_044_260, w_044_261, w_044_262, w_044_263, w_044_264, w_044_265, w_044_266, w_044_267, w_044_268, w_044_269, w_044_271, w_044_272, w_044_273, w_044_276, w_044_277, w_044_279, w_044_280, w_044_281, w_044_284, w_044_285, w_044_286, w_044_287, w_044_288, w_044_290, w_044_291, w_044_293, w_044_294, w_044_295, w_044_296, w_044_297, w_044_298, w_044_300, w_044_302, w_044_303, w_044_305, w_044_306, w_044_308, w_044_310, w_044_311, w_044_312, w_044_313, w_044_314, w_044_315, w_044_316, w_044_317, w_044_319, w_044_321, w_044_324, w_044_326, w_044_327, w_044_330, w_044_331, w_044_334, w_044_336, w_044_337, w_044_338, w_044_339, w_044_340, w_044_341, w_044_344, w_044_345, w_044_346, w_044_348, w_044_349, w_044_351, w_044_353, w_044_354, w_044_355, w_044_356, w_044_358, w_044_359, w_044_360, w_044_361, w_044_362, w_044_363, w_044_365, w_044_367, w_044_368, w_044_373, w_044_374, w_044_375, w_044_376, w_044_378, w_044_379, w_044_381, w_044_385, w_044_386, w_044_388, w_044_391, w_044_393, w_044_394, w_044_395, w_044_397, w_044_398, w_044_400, w_044_402, w_044_403, w_044_406, w_044_408, w_044_411, w_044_413, w_044_416, w_044_417, w_044_418, w_044_419, w_044_420, w_044_421, w_044_424, w_044_425, w_044_426, w_044_427, w_044_429, w_044_430, w_044_431, w_044_432, w_044_433, w_044_436, w_044_437, w_044_438, w_044_440, w_044_441, w_044_442, w_044_443, w_044_446, w_044_449, w_044_452, w_044_454, w_044_455, w_044_456, w_044_459, w_044_460, w_044_461, w_044_462, w_044_463, w_044_464, w_044_467, w_044_468, w_044_469, w_044_470, w_044_471, w_044_475, w_044_476, w_044_477, w_044_478, w_044_479, w_044_482, w_044_483, w_044_484, w_044_486, w_044_487, w_044_488, w_044_489, w_044_490, w_044_491, w_044_492, w_044_494, w_044_496, w_044_498, w_044_502, w_044_503, w_044_505, w_044_508, w_044_509, w_044_510, w_044_511, w_044_512, w_044_513, w_044_514, w_044_517, w_044_518, w_044_521, w_044_523, w_044_524, w_044_525, w_044_526, w_044_528, w_044_529, w_044_530, w_044_531, w_044_532, w_044_533, w_044_535, w_044_536, w_044_537, w_044_539, w_044_540, w_044_541, w_044_543, w_044_544, w_044_545, w_044_547, w_044_548, w_044_549, w_044_550, w_044_551, w_044_552, w_044_553, w_044_554, w_044_555, w_044_556, w_044_558, w_044_559, w_044_560, w_044_561, w_044_562, w_044_563, w_044_569, w_044_570, w_044_571, w_044_572, w_044_574, w_044_575, w_044_577, w_044_578, w_044_579, w_044_580, w_044_581, w_044_582, w_044_583, w_044_584, w_044_585, w_044_587, w_044_588, w_044_589, w_044_590, w_044_591, w_044_593, w_044_596, w_044_598, w_044_599, w_044_600, w_044_602, w_044_603, w_044_604, w_044_606, w_044_607, w_044_609, w_044_610, w_044_613, w_044_614, w_044_615, w_044_616, w_044_617, w_044_618, w_044_620, w_044_621, w_044_623, w_044_626, w_044_629, w_044_630, w_044_632, w_044_633, w_044_637, w_044_638, w_044_640, w_044_643, w_044_645, w_044_646, w_044_647, w_044_649, w_044_651, w_044_652, w_044_653, w_044_654, w_044_656, w_044_657, w_044_658, w_044_659, w_044_660, w_044_661, w_044_666, w_044_667, w_044_668, w_044_669, w_044_670, w_044_675, w_044_676, w_044_677, w_044_678, w_044_679, w_044_680, w_044_681, w_044_682, w_044_683, w_044_684, w_044_688, w_044_692, w_044_693, w_044_694, w_044_696, w_044_697, w_044_699, w_044_701, w_044_703, w_044_704, w_044_705, w_044_706, w_044_710, w_044_711, w_044_712, w_044_713, w_044_714, w_044_716, w_044_717, w_044_718, w_044_719, w_044_721, w_044_722, w_044_723, w_044_729, w_044_730, w_044_731, w_044_733, w_044_734, w_044_735, w_044_736, w_044_737, w_044_739, w_044_740, w_044_741, w_044_742, w_044_743, w_044_744, w_044_748, w_044_749, w_044_751, w_044_754, w_044_756, w_044_761, w_044_762, w_044_763, w_044_764, w_044_765, w_044_766, w_044_767, w_044_769, w_044_772, w_044_775, w_044_777, w_044_779, w_044_780, w_044_784, w_044_785, w_044_787, w_044_789, w_044_790, w_044_791, w_044_792, w_044_793, w_044_794, w_044_795, w_044_796, w_044_797, w_044_798, w_044_799, w_044_801, w_044_803, w_044_804, w_044_805, w_044_806, w_044_807, w_044_809, w_044_810, w_044_811, w_044_814, w_044_815, w_044_817, w_044_819, w_044_825, w_044_826, w_044_828, w_044_829, w_044_831, w_044_832, w_044_833, w_044_836, w_044_837, w_044_838, w_044_839, w_044_840, w_044_841, w_044_844, w_044_847, w_044_848, w_044_849, w_044_853, w_044_854, w_044_857, w_044_858, w_044_859, w_044_860, w_044_861, w_044_864, w_044_866, w_044_867, w_044_868, w_044_869, w_044_870, w_044_872, w_044_873, w_044_876, w_044_878, w_044_879, w_044_880, w_044_882, w_044_884, w_044_888, w_044_889, w_044_891, w_044_893, w_044_894, w_044_897, w_044_899, w_044_900, w_044_901, w_044_902, w_044_903, w_044_904, w_044_905, w_044_906, w_044_909, w_044_910, w_044_911, w_044_913, w_044_914, w_044_915, w_044_916, w_044_918, w_044_919, w_044_921, w_044_922, w_044_924, w_044_925, w_044_926, w_044_927, w_044_928, w_044_929, w_044_930, w_044_931, w_044_935, w_044_937, w_044_938, w_044_939, w_044_940, w_044_941, w_044_942, w_044_944, w_044_945, w_044_946, w_044_947, w_044_948, w_044_950, w_044_951, w_044_953, w_044_954, w_044_955, w_044_958, w_044_959, w_044_961, w_044_962, w_044_966, w_044_967, w_044_968, w_044_969, w_044_970, w_044_972, w_044_973, w_044_978, w_044_979, w_044_982, w_044_985, w_044_986, w_044_987, w_044_988, w_044_989, w_044_990, w_044_991, w_044_993, w_044_994, w_044_995, w_044_1001, w_044_1002, w_044_1003, w_044_1004, w_044_1006, w_044_1007, w_044_1008, w_044_1009, w_044_1010, w_044_1011, w_044_1012, w_044_1013, w_044_1014, w_044_1016, w_044_1017, w_044_1018, w_044_1019, w_044_1020, w_044_1023, w_044_1027, w_044_1028, w_044_1030, w_044_1032, w_044_1033, w_044_1034, w_044_1035, w_044_1036, w_044_1038, w_044_1039, w_044_1042, w_044_1043, w_044_1044, w_044_1045, w_044_1046, w_044_1047, w_044_1048, w_044_1049, w_044_1052, w_044_1054, w_044_1055, w_044_1056, w_044_1057, w_044_1060, w_044_1062, w_044_1063, w_044_1064, w_044_1065, w_044_1066, w_044_1067, w_044_1068, w_044_1069, w_044_1070, w_044_1071, w_044_1072, w_044_1073, w_044_1075, w_044_1076, w_044_1077, w_044_1080, w_044_1081, w_044_1083, w_044_1084, w_044_1085, w_044_1086, w_044_1087, w_044_1090, w_044_1091, w_044_1092, w_044_1093, w_044_1094, w_044_1095, w_044_1099, w_044_1100, w_044_1101, w_044_1102, w_044_1103, w_044_1105, w_044_1106, w_044_1107, w_044_1108, w_044_1109, w_044_1110, w_044_1111, w_044_1113, w_044_1114, w_044_1116, w_044_1117, w_044_1118, w_044_1119, w_044_1123, w_044_1127, w_044_1128, w_044_1129, w_044_1130, w_044_1131, w_044_1132, w_044_1133, w_044_1134, w_044_1135, w_044_1136, w_044_1137, w_044_1138, w_044_1140, w_044_1142, w_044_1143, w_044_1144, w_044_1145, w_044_1146, w_044_1147, w_044_1149, w_044_1150, w_044_1151, w_044_1152, w_044_1153, w_044_1154, w_044_1157, w_044_1158, w_044_1159, w_044_1160, w_044_1162, w_044_1163, w_044_1164, w_044_1166, w_044_1167, w_044_1168, w_044_1169, w_044_1170, w_044_1171, w_044_1172, w_044_1173, w_044_1174, w_044_1175, w_044_1176, w_044_1177, w_044_1180, w_044_1181, w_044_1185, w_044_1186, w_044_1187, w_044_1188, w_044_1189, w_044_1195, w_044_1196, w_044_1197, w_044_1198, w_044_1199, w_044_1201, w_044_1202, w_044_1203, w_044_1204, w_044_1206, w_044_1208, w_044_1209, w_044_1213, w_044_1214, w_044_1215, w_044_1216, w_044_1217, w_044_1220, w_044_1221, w_044_1222, w_044_1223, w_044_1224, w_044_1229, w_044_1230, w_044_1232, w_044_1233, w_044_1238, w_044_1239, w_044_1240, w_044_1241, w_044_1245, w_044_1248, w_044_1250, w_044_1251, w_044_1253, w_044_1257, w_044_1258, w_044_1260, w_044_1261, w_044_1262, w_044_1263, w_044_1264, w_044_1266, w_044_1267, w_044_1269, w_044_1270, w_044_1271, w_044_1272, w_044_1273, w_044_1274, w_044_1275, w_044_1276, w_044_1277, w_044_1278, w_044_1280, w_044_1281, w_044_1282, w_044_1283, w_044_1284, w_044_1285, w_044_1286, w_044_1287, w_044_1291, w_044_1292, w_044_1293, w_044_1295, w_044_1296, w_044_1297, w_044_1298, w_044_1300, w_044_1304, w_044_1306, w_044_1307, w_044_1311, w_044_1313, w_044_1314, w_044_1316, w_044_1317, w_044_1318, w_044_1319, w_044_1321, w_044_1322, w_044_1324, w_044_1325, w_044_1326, w_044_1328, w_044_1330, w_044_1332, w_044_1335, w_044_1336, w_044_1337, w_044_1339, w_044_1340, w_044_1342, w_044_1343, w_044_1344, w_044_1345, w_044_1346, w_044_1347, w_044_1348, w_044_1352, w_044_1353, w_044_1354, w_044_1360, w_044_1361, w_044_1363, w_044_1364, w_044_1365, w_044_1366, w_044_1367, w_044_1368, w_044_1369, w_044_1370, w_044_1372, w_044_1373, w_044_1375, w_044_1376, w_044_1378, w_044_1380, w_044_1381, w_044_1382, w_044_1383, w_044_1384, w_044_1385, w_044_1386, w_044_1388, w_044_1391, w_044_1393, w_044_1394, w_044_1395, w_044_1396, w_044_1397, w_044_1398, w_044_1399, w_044_1401, w_044_1402, w_044_1403, w_044_1404, w_044_1405, w_044_1407, w_044_1409, w_044_1410, w_044_1412, w_044_1413, w_044_1414, w_044_1416, w_044_1418, w_044_1419, w_044_1420, w_044_1423, w_044_1427, w_044_1430, w_044_1431, w_044_1435, w_044_1437, w_044_1438, w_044_1439, w_044_1440, w_044_1441, w_044_1442, w_044_1444, w_044_1445, w_044_1447, w_044_1448, w_044_1451, w_044_1452, w_044_1453, w_044_1454, w_044_1457, w_044_1461, w_044_1462, w_044_1463, w_044_1464, w_044_1465, w_044_1466, w_044_1467, w_044_1469, w_044_1470, w_044_1473, w_044_1474, w_044_1475, w_044_1476, w_044_1477, w_044_1478, w_044_1479, w_044_1480, w_044_1481, w_044_1482, w_044_1488, w_044_1489, w_044_1490, w_044_1491, w_044_1492, w_044_1494, w_044_1495, w_044_1496, w_044_1497, w_044_1498, w_044_1499, w_044_1500, w_044_1501, w_044_1502, w_044_1505, w_044_1506, w_044_1509, w_044_1510, w_044_1511, w_044_1514, w_044_1516, w_044_1517, w_044_1518, w_044_1521, w_044_1522, w_044_1524, w_044_1525, w_044_1526, w_044_1527, w_044_1528, w_044_1529, w_044_1534, w_044_1535, w_044_1536, w_044_1537, w_044_1539, w_044_1541, w_044_1542, w_044_1543, w_044_1544, w_044_1545, w_044_1546, w_044_1547, w_044_1549, w_044_1551, w_044_1553, w_044_1554, w_044_1555, w_044_1556, w_044_1559, w_044_1560, w_044_1561, w_044_1563, w_044_1564, w_044_1565, w_044_1566, w_044_1567, w_044_1569, w_044_1571, w_044_1572, w_044_1573, w_044_1574, w_044_1575, w_044_1579, w_044_1582, w_044_1583, w_044_1584, w_044_1585, w_044_1586, w_044_1587, w_044_1588, w_044_1589, w_044_1590, w_044_1591, w_044_1593, w_044_1594, w_044_1595, w_044_1596, w_044_1597, w_044_1598, w_044_1600, w_044_1601, w_044_1602, w_044_1603, w_044_1605, w_044_1606, w_044_1607, w_044_1608, w_044_1609, w_044_1611, w_044_1612, w_044_1613, w_044_1616, w_044_1617, w_044_1618, w_044_1619, w_044_1620, w_044_1621, w_044_1622, w_044_1623, w_044_1624, w_044_1625, w_044_1626, w_044_1627, w_044_1629, w_044_1630, w_044_1632, w_044_1633, w_044_1634, w_044_1635, w_044_1636, w_044_1637, w_044_1638, w_044_1639, w_044_1640, w_044_1641, w_044_1642, w_044_1644, w_044_1645, w_044_1647, w_044_1649, w_044_1650, w_044_1651, w_044_1652, w_044_1653, w_044_1654, w_044_1655, w_044_1656, w_044_1657, w_044_1658, w_044_1659, w_044_1661, w_044_1662, w_044_1664, w_044_1667, w_044_1669, w_044_1670, w_044_1672, w_044_1674, w_044_1675, w_044_1676, w_044_1677, w_044_1678, w_044_1680, w_044_1682, w_044_1683, w_044_1686, w_044_1687, w_044_1689, w_044_1690, w_044_1692, w_044_1693, w_044_1694, w_044_1697, w_044_1698, w_044_1699, w_044_1700, w_044_1701, w_044_1702, w_044_1703, w_044_1705, w_044_1706, w_044_1707, w_044_1709, w_044_1710, w_044_1711, w_044_1712, w_044_1713, w_044_1716, w_044_1717, w_044_1720, w_044_1721, w_044_1722, w_044_1723, w_044_1724, w_044_1725, w_044_1726, w_044_1727, w_044_1730, w_044_1732, w_044_1733, w_044_1734, w_044_1735, w_044_1736, w_044_1737, w_044_1738, w_044_1739, w_044_1740, w_044_1741, w_044_1744, w_044_1745, w_044_1746, w_044_1747, w_044_1748, w_044_1749, w_044_1750, w_044_1751, w_044_1752, w_044_1753, w_044_1754, w_044_1756, w_044_1757, w_044_1758, w_044_1760, w_044_1761, w_044_1763, w_044_1764, w_044_1765, w_044_1766, w_044_1767, w_044_1770, w_044_1771, w_044_1772, w_044_1775, w_044_1776, w_044_1777, w_044_1778, w_044_1779, w_044_1781, w_044_1782, w_044_1784, w_044_1785, w_044_1787, w_044_1788, w_044_1789, w_044_1790, w_044_1791, w_044_1794, w_044_1795, w_044_1796, w_044_1798, w_044_1799, w_044_1801, w_044_1802, w_044_1803, w_044_1805, w_044_1806, w_044_1807, w_044_1809, w_044_1810, w_044_1811, w_044_1812, w_044_1813, w_044_1815, w_044_1816, w_044_1817, w_044_1818, w_044_1819, w_044_1822, w_044_1823, w_044_1824, w_044_1825, w_044_1826, w_044_1829, w_044_1830, w_044_1832, w_044_1833, w_044_1834, w_044_1835, w_044_1836, w_044_1837, w_044_1838, w_044_1839, w_044_1841, w_044_1842, w_044_1843, w_044_1845, w_044_1846, w_044_1847, w_044_1848, w_044_1849, w_044_1850, w_044_1852, w_044_1853, w_044_1854, w_044_1855, w_044_1856, w_044_1857, w_044_1858, w_044_1859, w_044_1860, w_044_1861, w_044_1862, w_044_1863, w_044_1865, w_044_1866, w_044_1867, w_044_1868, w_044_1870, w_044_1871, w_044_1872, w_044_1873, w_044_1875, w_044_1876, w_044_1877, w_044_1878, w_044_1880, w_044_1882, w_044_1883, w_044_1885, w_044_1886, w_044_1887, w_044_1889, w_044_1890, w_044_1891, w_044_1893, w_044_1896, w_044_1897, w_044_1898, w_044_1899, w_044_1900, w_044_1903, w_044_1904, w_044_1905, w_044_1907, w_044_1908, w_044_1911, w_044_1912, w_044_1913, w_044_1914, w_044_1915, w_044_1917, w_044_1918, w_044_1919, w_044_1920, w_044_1921, w_044_1922, w_044_1924, w_044_1926, w_044_1927, w_044_1928, w_044_1929, w_044_1930, w_044_1931, w_044_1932, w_044_1933, w_044_1934, w_044_1935, w_044_1937, w_044_1939, w_044_1941, w_044_1943, w_044_1944, w_044_1945, w_044_1946, w_044_1947, w_044_1948, w_044_1949, w_044_1952, w_044_1953, w_044_1954, w_044_1956, w_044_1957, w_044_1959, w_044_1960, w_044_1961, w_044_1963, w_044_1964, w_044_1965, w_044_1967, w_044_1969, w_044_1970, w_044_1971, w_044_1972, w_044_1973, w_044_1974, w_044_1976, w_044_1977, w_044_1978, w_044_1979, w_044_1980, w_044_1982, w_044_1983, w_044_1984, w_044_1987, w_044_1988, w_044_1989, w_044_1990, w_044_1991, w_044_1992, w_044_1994, w_044_1995, w_044_1996, w_044_1997, w_044_1998, w_044_2000, w_044_2001, w_044_2002, w_044_2003, w_044_2004, w_044_2005, w_044_2006, w_044_2007, w_044_2009, w_044_2010, w_044_2011, w_044_2012, w_044_2015, w_044_2016, w_044_2017, w_044_2018, w_044_2019, w_044_2020, w_044_2024, w_044_2027, w_044_2030, w_044_2031, w_044_2032, w_044_2033, w_044_2034, w_044_2036, w_044_2037, w_044_2041, w_044_2044, w_044_2045, w_044_2047, w_044_2048, w_044_2050, w_044_2051, w_044_2052, w_044_2053, w_044_2054, w_044_2055, w_044_2056, w_044_2057, w_044_2058, w_044_2060, w_044_2061, w_044_2063, w_044_2064, w_044_2065, w_044_2066, w_044_2069, w_044_2070, w_044_2072, w_044_2073, w_044_2074, w_044_2075, w_044_2076, w_044_2077, w_044_2078, w_044_2080, w_044_2082, w_044_2083, w_044_2084, w_044_2085, w_044_2086, w_044_2087, w_044_2088, w_044_2089, w_044_2092, w_044_2093, w_044_2097, w_044_2100, w_044_2102, w_044_2103, w_044_2104, w_044_2105, w_044_2106, w_044_2107, w_044_2109, w_044_2110, w_044_2111, w_044_2112, w_044_2113, w_044_2115, w_044_2116, w_044_2118, w_044_2119, w_044_2121, w_044_2123, w_044_2125, w_044_2126, w_044_2127, w_044_2128, w_044_2129, w_044_2130, w_044_2131, w_044_2132, w_044_2133, w_044_2134, w_044_2135, w_044_2137, w_044_2138, w_044_2139, w_044_2140, w_044_2141, w_044_2145, w_044_2146, w_044_2147, w_044_2149, w_044_2150, w_044_2151, w_044_2154, w_044_2157, w_044_2158, w_044_2159, w_044_2160, w_044_2161, w_044_2162, w_044_2163, w_044_2164, w_044_2165, w_044_2167, w_044_2169, w_044_2170, w_044_2171, w_044_2172, w_044_2173, w_044_2176, w_044_2177, w_044_2180, w_044_2181, w_044_2183, w_044_2184, w_044_2186, w_044_2187, w_044_2188, w_044_2189, w_044_2190, w_044_2192, w_044_2193, w_044_2195, w_044_2196, w_044_2197, w_044_2200, w_044_2201, w_044_2203, w_044_2204, w_044_2205, w_044_2206, w_044_2207, w_044_2208, w_044_2213, w_044_2215, w_044_2216, w_044_2217, w_044_2218, w_044_2219, w_044_2220, w_044_2221, w_044_2222, w_044_2223, w_044_2224, w_044_2225, w_044_2226, w_044_2227, w_044_2228, w_044_2229, w_044_2230, w_044_2231, w_044_2233, w_044_2234, w_044_2235, w_044_2236, w_044_2237, w_044_2241, w_044_2243, w_044_2246, w_044_2247, w_044_2248, w_044_2249, w_044_2251, w_044_2252, w_044_2253, w_044_2254, w_044_2255, w_044_2256, w_044_2257, w_044_2258, w_044_2259, w_044_2260, w_044_2261, w_044_2262, w_044_2263, w_044_2264, w_044_2268, w_044_2269, w_044_2271, w_044_2272, w_044_2273, w_044_2274, w_044_2275, w_044_2278, w_044_2279, w_044_2282, w_044_2284, w_044_2286, w_044_2287, w_044_2288, w_044_2289, w_044_2290, w_044_2291, w_044_2292, w_044_2293, w_044_2294, w_044_2295, w_044_2296, w_044_2297, w_044_2298, w_044_2301, w_044_2302, w_044_2304, w_044_2305, w_044_2309, w_044_2310, w_044_2314, w_044_2316, w_044_2317, w_044_2320, w_044_2321, w_044_2322, w_044_2323, w_044_2324, w_044_2325, w_044_2326, w_044_2327, w_044_2328, w_044_2329, w_044_2330, w_044_2331, w_044_2333, w_044_2334, w_044_2335, w_044_2337, w_044_2339, w_044_2341, w_044_2342, w_044_2343, w_044_2346, w_044_2347, w_044_2348, w_044_2349, w_044_2350, w_044_2351, w_044_2352, w_044_2354, w_044_2355, w_044_2356, w_044_2359, w_044_2360, w_044_2364, w_044_2365, w_044_2366, w_044_2367, w_044_2369, w_044_2370, w_044_2371, w_044_2373, w_044_2374, w_044_2375, w_044_2376, w_044_2378, w_044_2379, w_044_2380, w_044_2381, w_044_2382, w_044_2383, w_044_2385, w_044_2386, w_044_2387, w_044_2389, w_044_2394, w_044_2395, w_044_2397, w_044_2398, w_044_2399, w_044_2401, w_044_2402, w_044_2403, w_044_2410, w_044_2411, w_044_2412, w_044_2413, w_044_2414, w_044_2418, w_044_2419, w_044_2420, w_044_2422, w_044_2423, w_044_2424, w_044_2426, w_044_2427, w_044_2428, w_044_2429, w_044_2430, w_044_2431, w_044_2432, w_044_2433, w_044_2434, w_044_2435, w_044_2436, w_044_2438, w_044_2439, w_044_2440, w_044_2441, w_044_2442, w_044_2444, w_044_2445, w_044_2446, w_044_2448, w_044_2449, w_044_2450, w_044_2451, w_044_2452, w_044_2453, w_044_2454, w_044_2455, w_044_2458, w_044_2459, w_044_2461, w_044_2463, w_044_2464, w_044_2466, w_044_2467, w_044_2468, w_044_2472, w_044_2473, w_044_2474, w_044_2475, w_044_2476, w_044_2477, w_044_2479, w_044_2480, w_044_2481, w_044_2482, w_044_2483, w_044_2484, w_044_2485, w_044_2487, w_044_2488, w_044_2489, w_044_2491, w_044_2492, w_044_2493, w_044_2494, w_044_2495, w_044_2496, w_044_2497, w_044_2498, w_044_2499, w_044_2500, w_044_2501, w_044_2502, w_044_2504, w_044_2506, w_044_2508, w_044_2509, w_044_2511, w_044_2513, w_044_2515, w_044_2518, w_044_2520, w_044_2521, w_044_2523, w_044_2527, w_044_2528, w_044_2529, w_044_2531, w_044_2532, w_044_2534, w_044_2536, w_044_2537, w_044_2538, w_044_2541, w_044_2544, w_044_2545, w_044_2548, w_044_2553, w_044_2555, w_044_2557, w_044_2558, w_044_2559, w_044_2562, w_044_2563, w_044_2564, w_044_2565, w_044_2566, w_044_2568, w_044_2570, w_044_2571, w_044_2574, w_044_2575, w_044_2577, w_044_2578, w_044_2579, w_044_2581, w_044_2582, w_044_2583, w_044_2584, w_044_2586, w_044_2587, w_044_2589, w_044_2590, w_044_2591, w_044_2592, w_044_2595, w_044_2597, w_044_2603, w_044_2604, w_044_2605, w_044_2606, w_044_2607, w_044_2610, w_044_2611, w_044_2612, w_044_2613, w_044_2615, w_044_2616, w_044_2618, w_044_2619, w_044_2620, w_044_2621, w_044_2622, w_044_2623, w_044_2624, w_044_2626, w_044_2627, w_044_2630, w_044_2631, w_044_2632, w_044_2633, w_044_2634, w_044_2635, w_044_2636, w_044_2637, w_044_2638, w_044_2639, w_044_2641, w_044_2642, w_044_2645, w_044_2647, w_044_2648, w_044_2650, w_044_2651, w_044_2652, w_044_2656, w_044_2658, w_044_2659, w_044_2660, w_044_2661, w_044_2662, w_044_2663, w_044_2664, w_044_2665, w_044_2666, w_044_2667, w_044_2668, w_044_2669, w_044_2670, w_044_2671, w_044_2672, w_044_2673, w_044_2674, w_044_2675, w_044_2676, w_044_2677, w_044_2679, w_044_2681, w_044_2684, w_044_2685, w_044_2686, w_044_2687, w_044_2688, w_044_2689, w_044_2690, w_044_2691, w_044_2692, w_044_2694, w_044_2695, w_044_2697, w_044_2698, w_044_2700, w_044_2701, w_044_2703, w_044_2705, w_044_2706, w_044_2707, w_044_2708, w_044_2709, w_044_2710, w_044_2711, w_044_2717, w_044_2718, w_044_2719, w_044_2720, w_044_2721, w_044_2723, w_044_2724, w_044_2725, w_044_2726, w_044_2728, w_044_2729, w_044_2730, w_044_2731, w_044_2734, w_044_2735, w_044_2736, w_044_2737, w_044_2739, w_044_2740, w_044_2741, w_044_2742, w_044_2743, w_044_2744, w_044_2745, w_044_2746, w_044_2747, w_044_2748, w_044_2750, w_044_2751, w_044_2753, w_044_2754, w_044_2756, w_044_2758, w_044_2759, w_044_2760, w_044_2763, w_044_2764, w_044_2765, w_044_2766, w_044_2767, w_044_2768, w_044_2769, w_044_2772, w_044_2773, w_044_2774, w_044_2775, w_044_2776, w_044_2777, w_044_2780, w_044_2781, w_044_2782, w_044_2783, w_044_2785, w_044_2786, w_044_2787, w_044_2789, w_044_2790, w_044_2791, w_044_2792, w_044_2793, w_044_2795, w_044_2796, w_044_2797, w_044_2798, w_044_2799, w_044_2800, w_044_2801, w_044_2803, w_044_2804, w_044_2805, w_044_2806, w_044_2809, w_044_2810, w_044_2815, w_044_2816, w_044_2817, w_044_2818, w_044_2819, w_044_2823, w_044_2824, w_044_2826, w_044_2830, w_044_2831, w_044_2832, w_044_2833, w_044_2834, w_044_2835, w_044_2836, w_044_2837, w_044_2838, w_044_2839, w_044_2840, w_044_2841, w_044_2842, w_044_2843, w_044_2844, w_044_2845, w_044_2847, w_044_2848, w_044_2850, w_044_2851, w_044_2852, w_044_2853, w_044_2854, w_044_2855, w_044_2856, w_044_2857, w_044_2858, w_044_2859, w_044_2860, w_044_2861, w_044_2862, w_044_2863, w_044_2864, w_044_2867, w_044_2868, w_044_2869, w_044_2871, w_044_2872, w_044_2873, w_044_2874, w_044_2875, w_044_2876, w_044_2877, w_044_2878, w_044_2879, w_044_2881, w_044_2883, w_044_2885, w_044_2886, w_044_2887, w_044_2891, w_044_2893, w_044_2894, w_044_2896, w_044_2897, w_044_2898, w_044_2899, w_044_2900, w_044_2902, w_044_2906, w_044_2907, w_044_2911, w_044_2913, w_044_2914, w_044_2915, w_044_2919, w_044_2920, w_044_2921, w_044_2923, w_044_2925, w_044_2927, w_044_2930, w_044_2931, w_044_2932, w_044_2933, w_044_2935, w_044_2936, w_044_2937, w_044_2938, w_044_2939, w_044_2941, w_044_2942, w_044_2943, w_044_2945, w_044_2948, w_044_2950, w_044_2951, w_044_2952, w_044_2953, w_044_2954, w_044_2955, w_044_2956, w_044_2957, w_044_2959, w_044_2961, w_044_2963, w_044_2965, w_044_2966, w_044_2967, w_044_2968, w_044_2969, w_044_2970, w_044_2973, w_044_2975, w_044_2978, w_044_2979, w_044_2980, w_044_2981, w_044_2982, w_044_2984, w_044_2985, w_044_2987, w_044_2988, w_044_2990, w_044_2992, w_044_2994, w_044_2998, w_044_2999, w_044_3000, w_044_3001, w_044_3002, w_044_3003, w_044_3004, w_044_3005, w_044_3006, w_044_3008, w_044_3009, w_044_3011, w_044_3012, w_044_3013, w_044_3014, w_044_3016, w_044_3017, w_044_3018, w_044_3020, w_044_3021, w_044_3024, w_044_3025, w_044_3026, w_044_3027, w_044_3028, w_044_3029, w_044_3030, w_044_3031, w_044_3033, w_044_3034, w_044_3035, w_044_3036, w_044_3037, w_044_3038, w_044_3040, w_044_3042, w_044_3043, w_044_3044, w_044_3045, w_044_3046, w_044_3047, w_044_3049, w_044_3052, w_044_3053, w_044_3057, w_044_3058, w_044_3059, w_044_3062, w_044_3063, w_044_3064, w_044_3065, w_044_3066, w_044_3067, w_044_3068, w_044_3069, w_044_3071, w_044_3072, w_044_3073, w_044_3074, w_044_3075, w_044_3077, w_044_3078, w_044_3079, w_044_3083, w_044_3085, w_044_3086, w_044_3089, w_044_3091, w_044_3092, w_044_3093, w_044_3095, w_044_3097, w_044_3099, w_044_3101, w_044_3102, w_044_3105, w_044_3106, w_044_3107, w_044_3108, w_044_3109, w_044_3110, w_044_3111, w_044_3112, w_044_3113, w_044_3114, w_044_3116, w_044_3117, w_044_3119, w_044_3120, w_044_3122, w_044_3124, w_044_3126, w_044_3127, w_044_3128, w_044_3130, w_044_3131, w_044_3132, w_044_3134, w_044_3135, w_044_3136, w_044_3138, w_044_3139, w_044_3140, w_044_3141, w_044_3142, w_044_3145, w_044_3146, w_044_3149, w_044_3150, w_044_3151, w_044_3152, w_044_3153, w_044_3155, w_044_3156, w_044_3158, w_044_3159, w_044_3160, w_044_3161, w_044_3162, w_044_3164, w_044_3165, w_044_3166, w_044_3169, w_044_3171, w_044_3172, w_044_3173, w_044_3174, w_044_3177, w_044_3178, w_044_3179, w_044_3180, w_044_3181, w_044_3183, w_044_3184, w_044_3187, w_044_3188, w_044_3191, w_044_3192, w_044_3193, w_044_3194, w_044_3196, w_044_3197, w_044_3199, w_044_3201, w_044_3202, w_044_3203, w_044_3205, w_044_3206, w_044_3207, w_044_3208, w_044_3210, w_044_3212, w_044_3213, w_044_3215, w_044_3216, w_044_3217, w_044_3219, w_044_3220, w_044_3222, w_044_3223, w_044_3225, w_044_3226, w_044_3229, w_044_3230, w_044_3231, w_044_3232, w_044_3233, w_044_3234, w_044_3235, w_044_3236, w_044_3238, w_044_3239, w_044_3240, w_044_3241, w_044_3245, w_044_3246, w_044_3247, w_044_3248, w_044_3249, w_044_3250, w_044_3251, w_044_3253, w_044_3256, w_044_3259, w_044_3260, w_044_3263, w_044_3264, w_044_3265, w_044_3266, w_044_3267, w_044_3270, w_044_3271, w_044_3272, w_044_3273, w_044_3274, w_044_3275, w_044_3277, w_044_3278, w_044_3279, w_044_3280, w_044_3282, w_044_3283, w_044_3284, w_044_3285, w_044_3286, w_044_3288, w_044_3289, w_044_3290, w_044_3291, w_044_3293, w_044_3295, w_044_3297, w_044_3299, w_044_3300, w_044_3302, w_044_3303, w_044_3305, w_044_3306, w_044_3308, w_044_3309, w_044_3310, w_044_3311, w_044_3315, w_044_3317, w_044_3321, w_044_3322, w_044_3324, w_044_3325, w_044_3326, w_044_3327, w_044_3329, w_044_3331, w_044_3332, w_044_3333, w_044_3334, w_044_3335, w_044_3336, w_044_3337, w_044_3338, w_044_3339, w_044_3343, w_044_3344, w_044_3346, w_044_3347, w_044_3348, w_044_3351, w_044_3352, w_044_3353, w_044_3354, w_044_3355, w_044_3356, w_044_3358, w_044_3359, w_044_3360, w_044_3361, w_044_3362, w_044_3363, w_044_3364, w_044_3369, w_044_3372, w_044_3374, w_044_3377, w_044_3378, w_044_3379, w_044_3380, w_044_3381, w_044_3382, w_044_3385, w_044_3386, w_044_3387, w_044_3388, w_044_3389, w_044_3390, w_044_3391, w_044_3392, w_044_3393, w_044_3397, w_044_3398, w_044_3400, w_044_3402, w_044_3404, w_044_3406, w_044_3407, w_044_3409, w_044_3412, w_044_3413, w_044_3415, w_044_3417, w_044_3418, w_044_3419, w_044_3420, w_044_3422, w_044_3424, w_044_3425, w_044_3426, w_044_3427, w_044_3428, w_044_3429, w_044_3430, w_044_3432, w_044_3433, w_044_3434, w_044_3436, w_044_3438, w_044_3441, w_044_3443, w_044_3445, w_044_3446, w_044_3447, w_044_3449, w_044_3452, w_044_3456, w_044_3457, w_044_3458, w_044_3459, w_044_3461, w_044_3463, w_044_3464, w_044_3466, w_044_3468, w_044_3469, w_044_3472, w_044_3473, w_044_3475, w_044_3476, w_044_3477, w_044_3479, w_044_3480, w_044_3481, w_044_3482, w_044_3483, w_044_3484, w_044_3487, w_044_3488, w_044_3489, w_044_3490, w_044_3491, w_044_3493, w_044_3494, w_044_3495, w_044_3496, w_044_3497, w_044_3500, w_044_3501, w_044_3502, w_044_3503, w_044_3506, w_044_3507, w_044_3509, w_044_3512, w_044_3513, w_044_3514, w_044_3515, w_044_3519, w_044_3520, w_044_3521, w_044_3522, w_044_3524, w_044_3527, w_044_3528, w_044_3529, w_044_3532, w_044_3534, w_044_3535, w_044_3536, w_044_3537, w_044_3538, w_044_3539, w_044_3540, w_044_3544, w_044_3545, w_044_3546, w_044_3547, w_044_3548, w_044_3550, w_044_3551, w_044_3552, w_044_3553, w_044_3554, w_044_3556, w_044_3557, w_044_3558, w_044_3562, w_044_3563, w_044_3564, w_044_3568, w_044_3569, w_044_3570, w_044_3571, w_044_3572, w_044_3574, w_044_3577, w_044_3578, w_044_3579, w_044_3581, w_044_3582, w_044_3583, w_044_3584, w_044_3585, w_044_3588, w_044_3589, w_044_3590, w_044_3591, w_044_3592, w_044_3596, w_044_3599, w_044_3600, w_044_3603, w_044_3604, w_044_3605, w_044_3607, w_044_3608, w_044_3609, w_044_3610, w_044_3611, w_044_3612, w_044_3613, w_044_3614, w_044_3615, w_044_3616, w_044_3617, w_044_3618, w_044_3619, w_044_3621, w_044_3623, w_044_3624, w_044_3627, w_044_3629, w_044_3630, w_044_3631, w_044_3632, w_044_3633, w_044_3634, w_044_3636, w_044_3637, w_044_3638, w_044_3639, w_044_3641, w_044_3642, w_044_3643, w_044_3644, w_044_3645, w_044_3646, w_044_3647, w_044_3648, w_044_3650, w_044_3651, w_044_3653, w_044_3655, w_044_3656, w_044_3657, w_044_3658, w_044_3659, w_044_3661, w_044_3662, w_044_3663, w_044_3664, w_044_3665, w_044_3666, w_044_3668, w_044_3669, w_044_3671, w_044_3672, w_044_3675, w_044_3676, w_044_3677, w_044_3679, w_044_3680, w_044_3681, w_044_3682, w_044_3683, w_044_3684, w_044_3685, w_044_3686, w_044_3687, w_044_3690, w_044_3691, w_044_3693, w_044_3695, w_044_3696, w_044_3697, w_044_3698, w_044_3699, w_044_3700, w_044_3702, w_044_3703, w_044_3704, w_044_3705, w_044_3706, w_044_3708, w_044_3711, w_044_3713, w_044_3714, w_044_3715, w_044_3716, w_044_3717, w_044_3718, w_044_3720, w_044_3721, w_044_3722, w_044_3723, w_044_3724, w_044_3725, w_044_3726, w_044_3727, w_044_3729, w_044_3730, w_044_3731, w_044_3732, w_044_3733, w_044_3734, w_044_3735, w_044_3736, w_044_3737, w_044_3739, w_044_3740, w_044_3741, w_044_3742, w_044_3743, w_044_3744, w_044_3745, w_044_3749, w_044_3750, w_044_3753, w_044_3755, w_044_3756, w_044_3757, w_044_3759, w_044_3760, w_044_3761, w_044_3762, w_044_3766, w_044_3768, w_044_3771, w_044_3773, w_044_3776, w_044_3777, w_044_3778, w_044_3779, w_044_3780, w_044_3784, w_044_3789, w_044_3790, w_044_3791, w_044_3792, w_044_3793, w_044_3796, w_044_3797, w_044_3798, w_044_3799, w_044_3800, w_044_3801, w_044_3802, w_044_3804, w_044_3806, w_044_3807, w_044_3810, w_044_3812, w_044_3815, w_044_3818, w_044_3819, w_044_3820, w_044_3821, w_044_3824, w_044_3825, w_044_3826, w_044_3831, w_044_3834, w_044_3835, w_044_3838, w_044_3839, w_044_3840, w_044_3844, w_044_3845, w_044_3851, w_044_3853, w_044_3855, w_044_3858, w_044_3859, w_044_3860, w_044_3866, w_044_3867, w_044_3868, w_044_3872, w_044_3873, w_044_3876, w_044_3877, w_044_3880, w_044_3881, w_044_3883, w_044_3888, w_044_3893, w_044_3894, w_044_3896, w_044_3897, w_044_3901, w_044_3902, w_044_3903, w_044_3905, w_044_3906, w_044_3909, w_044_3912, w_044_3913, w_044_3915, w_044_3922, w_044_3923, w_044_3928, w_044_3930, w_044_3932, w_044_3934, w_044_3935, w_044_3937, w_044_3938, w_044_3939, w_044_3942, w_044_3948, w_044_3949, w_044_3951, w_044_3953, w_044_3954, w_044_3956, w_044_3957, w_044_3958, w_044_3960, w_044_3964, w_044_3966, w_044_3971, w_044_3975, w_044_3976, w_044_3977, w_044_3982, w_044_3984, w_044_3992, w_044_3994, w_044_3997, w_044_3998, w_044_3999, w_044_4001, w_044_4003, w_044_4006, w_044_4011, w_044_4012, w_044_4014, w_044_4021, w_044_4025, w_044_4027, w_044_4028, w_044_4030, w_044_4035, w_044_4036, w_044_4037, w_044_4040, w_044_4041, w_044_4044, w_044_4047, w_044_4048, w_044_4051, w_044_4053, w_044_4054, w_044_4056, w_044_4057, w_044_4058, w_044_4059, w_044_4060, w_044_4061, w_044_4064, w_044_4068, w_044_4069, w_044_4073, w_044_4075, w_044_4078, w_044_4086, w_044_4087, w_044_4097, w_044_4100, w_044_4101, w_044_4103, w_044_4104, w_044_4106, w_044_4112, w_044_4113, w_044_4120, w_044_4122, w_044_4123, w_044_4124, w_044_4136, w_044_4138, w_044_4142, w_044_4144, w_044_4146, w_044_4148, w_044_4150, w_044_4151, w_044_4154, w_044_4155, w_044_4156, w_044_4157, w_044_4161, w_044_4166, w_044_4170, w_044_4173, w_044_4175, w_044_4178, w_044_4179, w_044_4181, w_044_4186, w_044_4187, w_044_4188, w_044_4189, w_044_4190, w_044_4193, w_044_4198, w_044_4201, w_044_4203, w_044_4205, w_044_4206, w_044_4207, w_044_4209, w_044_4212, w_044_4213, w_044_4214, w_044_4215, w_044_4217, w_044_4218, w_044_4219, w_044_4220, w_044_4222, w_044_4223, w_044_4224, w_044_4225, w_044_4226, w_044_4227, w_044_4229, w_044_4230, w_044_4233, w_044_4234, w_044_4236, w_044_4237, w_044_4239, w_044_4240, w_044_4241, w_044_4243, w_044_4245, w_044_4249, w_044_4250, w_044_4251, w_044_4255, w_044_4256, w_044_4261, w_044_4262, w_044_4263, w_044_4265, w_044_4267, w_044_4268, w_044_4269, w_044_4270, w_044_4271, w_044_4272, w_044_4281, w_044_4284, w_044_4288, w_044_4290, w_044_4293, w_044_4295, w_044_4297, w_044_4298, w_044_4300, w_044_4302, w_044_4303, w_044_4304, w_044_4306, w_044_4311, w_044_4312, w_044_4313, w_044_4324, w_044_4326, w_044_4328, w_044_4329, w_044_4335, w_044_4336, w_044_4337, w_044_4338, w_044_4339, w_044_4340, w_044_4341, w_044_4342, w_044_4343, w_044_4345, w_044_4348, w_044_4349, w_044_4351, w_044_4352, w_044_4353, w_044_4355, w_044_4356, w_044_4357, w_044_4358, w_044_4360, w_044_4362, w_044_4364, w_044_4367, w_044_4370, w_044_4371, w_044_4380, w_044_4381, w_044_4382, w_044_4383, w_044_4384, w_044_4386, w_044_4387, w_044_4389, w_044_4391, w_044_4396, w_044_4398, w_044_4399, w_044_4401, w_044_4402, w_044_4403, w_044_4407, w_044_4409, w_044_4412, w_044_4416, w_044_4420, w_044_4422, w_044_4425, w_044_4426, w_044_4428, w_044_4429, w_044_4431, w_044_4432, w_044_4433, w_044_4435, w_044_4439, w_044_4441, w_044_4443, w_044_4445, w_044_4446, w_044_4447, w_044_4448, w_044_4450, w_044_4451, w_044_4453, w_044_4454, w_044_4457, w_044_4458, w_044_4459, w_044_4461, w_044_4463, w_044_4464, w_044_4465, w_044_4467, w_044_4468, w_044_4471, w_044_4480, w_044_4485, w_044_4487, w_044_4492, w_044_4496, w_044_4500, w_044_4502, w_044_4503, w_044_4505, w_044_4506, w_044_4513, w_044_4514, w_044_4518, w_044_4522, w_044_4525, w_044_4526, w_044_4530, w_044_4533, w_044_4538, w_044_4539, w_044_4541, w_044_4542, w_044_4543, w_044_4544, w_044_4545, w_044_4547, w_044_4548, w_044_4550, w_044_4555, w_044_4558, w_044_4560, w_044_4564, w_044_4565, w_044_4572, w_044_4573, w_044_4575, w_044_4576, w_044_4577, w_044_4581, w_044_4582, w_044_4583, w_044_4586, w_044_4587, w_044_4588, w_044_4590, w_044_4592, w_044_4594, w_044_4599, w_044_4602, w_044_4603, w_044_4604, w_044_4606, w_044_4608, w_044_4611, w_044_4612, w_044_4613, w_044_4616, w_044_4618, w_044_4619, w_044_4621, w_044_4625, w_044_4627, w_044_4628, w_044_4631, w_044_4634, w_044_4635, w_044_4637, w_044_4638, w_044_4641, w_044_4648, w_044_4651, w_044_4653, w_044_4654, w_044_4656, w_044_4657, w_044_4660, w_044_4661, w_044_4662, w_044_4663, w_044_4666, w_044_4668, w_044_4669, w_044_4670, w_044_4671, w_044_4673, w_044_4676, w_044_4677, w_044_4684, w_044_4686, w_044_4687, w_044_4688, w_044_4689, w_044_4690, w_044_4693, w_044_4697, w_044_4700, w_044_4702, w_044_4703, w_044_4705, w_044_4706, w_044_4710, w_044_4711, w_044_4712, w_044_4713, w_044_4715, w_044_4717, w_044_4718, w_044_4719, w_044_4724, w_044_4729, w_044_4732, w_044_4734, w_044_4735, w_044_4736, w_044_4739, w_044_4742, w_044_4743, w_044_4744, w_044_4745, w_044_4746, w_044_4747, w_044_4749, w_044_4751, w_044_4753, w_044_4755, w_044_4757, w_044_4758, w_044_4764, w_044_4769, w_044_4770, w_044_4774, w_044_4783, w_044_4785, w_044_4790, w_044_4791, w_044_4792, w_044_4794, w_044_4797, w_044_4798, w_044_4800, w_044_4801, w_044_4802, w_044_4803, w_044_4804, w_044_4805, w_044_4806, w_044_4809, w_044_4815, w_044_4816, w_044_4819, w_044_4821, w_044_4822, w_044_4823, w_044_4828, w_044_4830, w_044_4834, w_044_4835, w_044_4836, w_044_4839, w_044_4843, w_044_4845, w_044_4846, w_044_4847, w_044_4848, w_044_4851, w_044_4854, w_044_4856, w_044_4857, w_044_4863, w_044_4865, w_044_4869, w_044_4875, w_044_4876, w_044_4878, w_044_4882, w_044_4883, w_044_4884, w_044_4887, w_044_4889, w_044_4890, w_044_4891, w_044_4892, w_044_4894, w_044_4895, w_044_4898, w_044_4899, w_044_4900, w_044_4902, w_044_4903, w_044_4905, w_044_4906, w_044_4908, w_044_4909, w_044_4914, w_044_4916, w_044_4918, w_044_4919, w_044_4921, w_044_4922, w_044_4924, w_044_4925, w_044_4930, w_044_4932, w_044_4935, w_044_4937, w_044_4938, w_044_4941, w_044_4943, w_044_4945, w_044_4946, w_044_4947, w_044_4948, w_044_4949, w_044_4955, w_044_4957, w_044_4959, w_044_4960, w_044_4962, w_044_4963, w_044_4968, w_044_4972, w_044_4976, w_044_4977, w_044_4979, w_044_4985, w_044_4986, w_044_4987, w_044_4988, w_044_4989, w_044_4991, w_044_4992, w_044_4993, w_044_4995, w_044_4996, w_044_4997, w_044_4998, w_044_5002, w_044_5004, w_044_5007, w_044_5008, w_044_5014, w_044_5019, w_044_5022, w_044_5023, w_044_5024, w_044_5026, w_044_5028, w_044_5029, w_044_5030, w_044_5032, w_044_5035, w_044_5038, w_044_5039, w_044_5040, w_044_5041, w_044_5042, w_044_5043, w_044_5044, w_044_5045, w_044_5046, w_044_5048, w_044_5049, w_044_5051, w_044_5056, w_044_5057, w_044_5062, w_044_5065, w_044_5066, w_044_5068, w_044_5069, w_044_5072, w_044_5074, w_044_5075, w_044_5076, w_044_5077, w_044_5078, w_044_5080, w_044_5081, w_044_5083, w_044_5084, w_044_5085, w_044_5087, w_044_5088, w_044_5089, w_044_5091, w_044_5092, w_044_5093, w_044_5094, w_044_5095, w_044_5096, w_044_5097, w_044_5099, w_044_5100, w_044_5101, w_044_5102, w_044_5103, w_044_5104, w_044_5106, w_044_5108, w_044_5109, w_044_5113, w_044_5117, w_044_5121, w_044_5123, w_044_5125, w_044_5126, w_044_5130, w_044_5132, w_044_5140, w_044_5148, w_044_5150, w_044_5151, w_044_5157, w_044_5161, w_044_5164, w_044_5166, w_044_5168, w_044_5170, w_044_5171, w_044_5172, w_044_5173, w_044_5174, w_044_5175, w_044_5177, w_044_5178, w_044_5179, w_044_5183, w_044_5185, w_044_5187, w_044_5190, w_044_5192, w_044_5193, w_044_5195, w_044_5196, w_044_5200, w_044_5201, w_044_5202, w_044_5204, w_044_5210, w_044_5212, w_044_5214, w_044_5221, w_044_5222, w_044_5223, w_044_5224, w_044_5227, w_044_5228, w_044_5232, w_044_5233, w_044_5234, w_044_5237, w_044_5242, w_044_5245, w_044_5247, w_044_5248, w_044_5249, w_044_5250, w_044_5251, w_044_5254, w_044_5257, w_044_5259, w_044_5261, w_044_5262, w_044_5266, w_044_5268, w_044_5270, w_044_5271, w_044_5272, w_044_5273, w_044_5277, w_044_5281, w_044_5285, w_044_5290, w_044_5296, w_044_5297, w_044_5299, w_044_5300, w_044_5301, w_044_5304, w_044_5306, w_044_5307, w_044_5308, w_044_5310, w_044_5311, w_044_5312, w_044_5314, w_044_5315, w_044_5316, w_044_5327, w_044_5329, w_044_5335, w_044_5337, w_044_5341, w_044_5346, w_044_5348, w_044_5349, w_044_5351, w_044_5352, w_044_5353, w_044_5360, w_044_5365, w_044_5368, w_044_5369, w_044_5372, w_044_5374, w_044_5375, w_044_5376, w_044_5377, w_044_5378, w_044_5382, w_044_5384, w_044_5389, w_044_5391, w_044_5393, w_044_5394, w_044_5395, w_044_5396, w_044_5397, w_044_5398, w_044_5399, w_044_5405, w_044_5408, w_044_5410, w_044_5412, w_044_5415, w_044_5416, w_044_5418, w_044_5421, w_044_5423, w_044_5424, w_044_5425, w_044_5426, w_044_5430, w_044_5434, w_044_5435, w_044_5436, w_044_5438, w_044_5439, w_044_5440, w_044_5442, w_044_5443, w_044_5444, w_044_5452, w_044_5453, w_044_5458, w_044_5459, w_044_5462, w_044_5463, w_044_5467, w_044_5471, w_044_5472, w_044_5474, w_044_5475, w_044_5479, w_044_5481, w_044_5486, w_044_5487, w_044_5490, w_044_5498, w_044_5499, w_044_5500, w_044_5504, w_044_5508, w_044_5511, w_044_5512, w_044_5513, w_044_5517, w_044_5518, w_044_5519, w_044_5520, w_044_5522, w_044_5525, w_044_5527, w_044_5529, w_044_5530, w_044_5531, w_044_5537, w_044_5542, w_044_5545, w_044_5549, w_044_5550, w_044_5552, w_044_5555, w_044_5557, w_044_5558, w_044_5559, w_044_5564, w_044_5566, w_044_5570, w_044_5575, w_044_5576, w_044_5577, w_044_5578, w_044_5581, w_044_5582, w_044_5583, w_044_5586, w_044_5588, w_044_5590, w_044_5594, w_044_5595, w_044_5596, w_044_5597, w_044_5600, w_044_5602, w_044_5603, w_044_5606, w_044_5608, w_044_5609, w_044_5610, w_044_5611, w_044_5613, w_044_5615, w_044_5619, w_044_5620, w_044_5621, w_044_5622, w_044_5624, w_044_5629, w_044_5631, w_044_5638, w_044_5641, w_044_5642, w_044_5651, w_044_5655, w_044_5656, w_044_5657, w_044_5660, w_044_5661, w_044_5662, w_044_5663, w_044_5665, w_044_5666, w_044_5669, w_044_5670, w_044_5671, w_044_5672, w_044_5678, w_044_5682, w_044_5683, w_044_5684, w_044_5689, w_044_5694, w_044_5696, w_044_5699, w_044_5701, w_044_5705, w_044_5707, w_044_5710, w_044_5711, w_044_5713, w_044_5717, w_044_5719, w_044_5723, w_044_5730, w_044_5731, w_044_5733, w_044_5736, w_044_5744, w_044_5746, w_044_5750, w_044_5752, w_044_5754, w_044_5758, w_044_5759, w_044_5760, w_044_5761, w_044_5762, w_044_5767, w_044_5768, w_044_5770, w_044_5771, w_044_5772, w_044_5773, w_044_5779, w_044_5780, w_044_5783, w_044_5786, w_044_5787, w_044_5788, w_044_5790, w_044_5792, w_044_5797, w_044_5798, w_044_5800, w_044_5801, w_044_5802, w_044_5804, w_044_5806, w_044_5810, w_044_5812, w_044_5814, w_044_5817, w_044_5819, w_044_5821, w_044_5822, w_044_5827, w_044_5830, w_044_5831, w_044_5832, w_044_5833, w_044_5835, w_044_5837, w_044_5838, w_044_5840, w_044_5841, w_044_5842, w_044_5843, w_044_5844, w_044_5845, w_044_5846, w_044_5848, w_044_5849, w_044_5850, w_044_5853, w_044_5854, w_044_5855, w_044_5865, w_044_5867, w_044_5869, w_044_5871, w_044_5876, w_044_5877, w_044_5878, w_044_5879, w_044_5880, w_044_5890, w_044_5891, w_044_5894, w_044_5895, w_044_5896, w_044_5899, w_044_5900, w_044_5906, w_044_5907, w_044_5908, w_044_5911, w_044_5918, w_044_5920, w_044_5922, w_044_5923, w_044_5924, w_044_5925, w_044_5926, w_044_5928, w_044_5931, w_044_5935, w_044_5937, w_044_5941, w_044_5945, w_044_5947, w_044_5952, w_044_5953, w_044_5957, w_044_5960, w_044_5962, w_044_5963, w_044_5971, w_044_5972, w_044_5976, w_044_5977, w_044_5980, w_044_5981, w_044_5982, w_044_5983, w_044_5988, w_044_5990, w_044_6001, w_044_6005, w_044_6007, w_044_6008, w_044_6010, w_044_6011, w_044_6013, w_044_6015, w_044_6019, w_044_6022, w_044_6023, w_044_6030, w_044_6031, w_044_6032, w_044_6034, w_044_6035, w_044_6038, w_044_6041, w_044_6044, w_044_6046, w_044_6049, w_044_6050, w_044_6052, w_044_6058, w_044_6061, w_044_6062, w_044_6064, w_044_6065, w_044_6066, w_044_6067, w_044_6068, w_044_6069, w_044_6071, w_044_6072, w_044_6074, w_044_6079, w_044_6080, w_044_6081, w_044_6083, w_044_6091, w_044_6092, w_044_6096, w_044_6097, w_044_6098, w_044_6099, w_044_6101, w_044_6108, w_044_6112, w_044_6113, w_044_6114, w_044_6119, w_044_6120, w_044_6121, w_044_6122, w_044_6127, w_044_6128, w_044_6129, w_044_6131, w_044_6132, w_044_6138, w_044_6139, w_044_6148, w_044_6149, w_044_6153, w_044_6156, w_044_6158, w_044_6160, w_044_6162, w_044_6163, w_044_6167, w_044_6169, w_044_6170, w_044_6171, w_044_6172, w_044_6174, w_044_6175, w_044_6177, w_044_6178, w_044_6179, w_044_6180, w_044_6182, w_044_6184, w_044_6185;
  wire w_045_001, w_045_002, w_045_003, w_045_004, w_045_005, w_045_006, w_045_007, w_045_008, w_045_010, w_045_011, w_045_012, w_045_013, w_045_014, w_045_016, w_045_017, w_045_018, w_045_020, w_045_021, w_045_022, w_045_023, w_045_025, w_045_026, w_045_030, w_045_031, w_045_035, w_045_037, w_045_039, w_045_040, w_045_042, w_045_044, w_045_047, w_045_048, w_045_049, w_045_051, w_045_052, w_045_053, w_045_054, w_045_055, w_045_056, w_045_057, w_045_058, w_045_059, w_045_060, w_045_061, w_045_062, w_045_063, w_045_064, w_045_065, w_045_066, w_045_067, w_045_068, w_045_069, w_045_070, w_045_071, w_045_072, w_045_075, w_045_076, w_045_077, w_045_078, w_045_079, w_045_080, w_045_082, w_045_083, w_045_085, w_045_088, w_045_090, w_045_091, w_045_092, w_045_093, w_045_094, w_045_095, w_045_096, w_045_097, w_045_101, w_045_102, w_045_103, w_045_107, w_045_108, w_045_109, w_045_111, w_045_114, w_045_116, w_045_118, w_045_119, w_045_122, w_045_123, w_045_125, w_045_126, w_045_127, w_045_128, w_045_129, w_045_132, w_045_134, w_045_135, w_045_136, w_045_137, w_045_140, w_045_142, w_045_143, w_045_144, w_045_145, w_045_146, w_045_147, w_045_150, w_045_152, w_045_154, w_045_157, w_045_158, w_045_159, w_045_160, w_045_161, w_045_162, w_045_163, w_045_166, w_045_168, w_045_169, w_045_170, w_045_171, w_045_172, w_045_173, w_045_174, w_045_175, w_045_177, w_045_179, w_045_182, w_045_183, w_045_185, w_045_186, w_045_188, w_045_189, w_045_190, w_045_191, w_045_193, w_045_194, w_045_195, w_045_197, w_045_199, w_045_201, w_045_202, w_045_203, w_045_207, w_045_209, w_045_210, w_045_211, w_045_213, w_045_214, w_045_215, w_045_216, w_045_217, w_045_219, w_045_220, w_045_221, w_045_222, w_045_223, w_045_224, w_045_225, w_045_227, w_045_228, w_045_229, w_045_230, w_045_231, w_045_232, w_045_233, w_045_234, w_045_235, w_045_236, w_045_238, w_045_239, w_045_240, w_045_242, w_045_243, w_045_244, w_045_246, w_045_247, w_045_248, w_045_250, w_045_251, w_045_252, w_045_253, w_045_254, w_045_255, w_045_260, w_045_261, w_045_263, w_045_264, w_045_265, w_045_268, w_045_269, w_045_271, w_045_272, w_045_274, w_045_275, w_045_276, w_045_278, w_045_279, w_045_282, w_045_283, w_045_284, w_045_285, w_045_286, w_045_287, w_045_288, w_045_289, w_045_290, w_045_291, w_045_292, w_045_294, w_045_295, w_045_296, w_045_298, w_045_299, w_045_300, w_045_302, w_045_303, w_045_304, w_045_306, w_045_307, w_045_309, w_045_310, w_045_314, w_045_316, w_045_317, w_045_318, w_045_319, w_045_320, w_045_322, w_045_323, w_045_324, w_045_326, w_045_330, w_045_331, w_045_332, w_045_334, w_045_335, w_045_337, w_045_338, w_045_339, w_045_340, w_045_342, w_045_343, w_045_346, w_045_347, w_045_348, w_045_349, w_045_350, w_045_351, w_045_353, w_045_354, w_045_357, w_045_358, w_045_359, w_045_361, w_045_364, w_045_366, w_045_367, w_045_368, w_045_369, w_045_370, w_045_371, w_045_373, w_045_376, w_045_378, w_045_379, w_045_381, w_045_382, w_045_384, w_045_386, w_045_387, w_045_388, w_045_390, w_045_392, w_045_394, w_045_397, w_045_398, w_045_401, w_045_403, w_045_404, w_045_406, w_045_410, w_045_413, w_045_414, w_045_417, w_045_419, w_045_421, w_045_422, w_045_424, w_045_425, w_045_426, w_045_427, w_045_431, w_045_434, w_045_437, w_045_438, w_045_439, w_045_440, w_045_441, w_045_442, w_045_444, w_045_445, w_045_446, w_045_447, w_045_448, w_045_449, w_045_450, w_045_451, w_045_452, w_045_453, w_045_454, w_045_456, w_045_457, w_045_460, w_045_462, w_045_463, w_045_466, w_045_467, w_045_468, w_045_469, w_045_470, w_045_471, w_045_474, w_045_477, w_045_480, w_045_485, w_045_486, w_045_487, w_045_489, w_045_490, w_045_491, w_045_492, w_045_493, w_045_494, w_045_495, w_045_497, w_045_499, w_045_500, w_045_502, w_045_503, w_045_504, w_045_505, w_045_508, w_045_509, w_045_511, w_045_512, w_045_514, w_045_515, w_045_517, w_045_518, w_045_519, w_045_520, w_045_521, w_045_522, w_045_523, w_045_524, w_045_525, w_045_526, w_045_528, w_045_529, w_045_531, w_045_532, w_045_533, w_045_534, w_045_537, w_045_538, w_045_540, w_045_541, w_045_543, w_045_546, w_045_548, w_045_549, w_045_550, w_045_551, w_045_553, w_045_554, w_045_555, w_045_556, w_045_558, w_045_559, w_045_560, w_045_561, w_045_562, w_045_563, w_045_564, w_045_565, w_045_566, w_045_567, w_045_569, w_045_570, w_045_571, w_045_572, w_045_573, w_045_575, w_045_576, w_045_577, w_045_578, w_045_579, w_045_580, w_045_581, w_045_582, w_045_583, w_045_585, w_045_586, w_045_587, w_045_588, w_045_589, w_045_590, w_045_592, w_045_593, w_045_594, w_045_595, w_045_596, w_045_597, w_045_598, w_045_599, w_045_602, w_045_603, w_045_604, w_045_605, w_045_606, w_045_607, w_045_610, w_045_611, w_045_612, w_045_615, w_045_616, w_045_617, w_045_618, w_045_619, w_045_620, w_045_621, w_045_623, w_045_624, w_045_625, w_045_627, w_045_628, w_045_629, w_045_631, w_045_634, w_045_635, w_045_636, w_045_637, w_045_639, w_045_640, w_045_641, w_045_643, w_045_646, w_045_647, w_045_649, w_045_650, w_045_651, w_045_653, w_045_655, w_045_656, w_045_657, w_045_658, w_045_659, w_045_660, w_045_662, w_045_664, w_045_667, w_045_668, w_045_669, w_045_670, w_045_671, w_045_673, w_045_674, w_045_675, w_045_676, w_045_681, w_045_682, w_045_685, w_045_686, w_045_687, w_045_688, w_045_689, w_045_693, w_045_694, w_045_695, w_045_696, w_045_697, w_045_698, w_045_699, w_045_700, w_045_701, w_045_704, w_045_705, w_045_706, w_045_707, w_045_708, w_045_709, w_045_711, w_045_712, w_045_713, w_045_714, w_045_716, w_045_717, w_045_718, w_045_720, w_045_725, w_045_726, w_045_727, w_045_728, w_045_729, w_045_730, w_045_731, w_045_732, w_045_734, w_045_735, w_045_736, w_045_738, w_045_739, w_045_740, w_045_741, w_045_742, w_045_743, w_045_744, w_045_745, w_045_746, w_045_747, w_045_748, w_045_749, w_045_751, w_045_752, w_045_753, w_045_754, w_045_756, w_045_758, w_045_759, w_045_760, w_045_763, w_045_764, w_045_765, w_045_766, w_045_767, w_045_768, w_045_769, w_045_771, w_045_772, w_045_774, w_045_775, w_045_776, w_045_778, w_045_781, w_045_782, w_045_786, w_045_788, w_045_790, w_045_792, w_045_793, w_045_794, w_045_796, w_045_798, w_045_800, w_045_801, w_045_803, w_045_804, w_045_805, w_045_806, w_045_807, w_045_808, w_045_809, w_045_811, w_045_814, w_045_815, w_045_816, w_045_820, w_045_821, w_045_823, w_045_825, w_045_826, w_045_827, w_045_828, w_045_830, w_045_831, w_045_833, w_045_834, w_045_835, w_045_836, w_045_838, w_045_839, w_045_840, w_045_841, w_045_842, w_045_843, w_045_844, w_045_846, w_045_848, w_045_850, w_045_852, w_045_854, w_045_858, w_045_859, w_045_863, w_045_864, w_045_866, w_045_867, w_045_868, w_045_870, w_045_871, w_045_872, w_045_873, w_045_874, w_045_875, w_045_876, w_045_877, w_045_878, w_045_879, w_045_880, w_045_881, w_045_883, w_045_884, w_045_885, w_045_886, w_045_887, w_045_888, w_045_890, w_045_891, w_045_892, w_045_894, w_045_895, w_045_896, w_045_897, w_045_898, w_045_900, w_045_902, w_045_904, w_045_905, w_045_906, w_045_908, w_045_909, w_045_910, w_045_911, w_045_912, w_045_913, w_045_914, w_045_916, w_045_920, w_045_921, w_045_922, w_045_923, w_045_924, w_045_925, w_045_926, w_045_928, w_045_929, w_045_930, w_045_931, w_045_933, w_045_934, w_045_938, w_045_939, w_045_940, w_045_941, w_045_942, w_045_943, w_045_945, w_045_947, w_045_948, w_045_951, w_045_952, w_045_953, w_045_955, w_045_956, w_045_957, w_045_958, w_045_959, w_045_960, w_045_961, w_045_962, w_045_963, w_045_964, w_045_965, w_045_966, w_045_967, w_045_969, w_045_970, w_045_971, w_045_972, w_045_974, w_045_975, w_045_976, w_045_979, w_045_980, w_045_981, w_045_982, w_045_983, w_045_986, w_045_987, w_045_988, w_045_989, w_045_990, w_045_991, w_045_992, w_045_995, w_045_997, w_045_998, w_045_999, w_045_1000, w_045_1001, w_045_1003, w_045_1004, w_045_1005, w_045_1006, w_045_1007, w_045_1010, w_045_1011, w_045_1012, w_045_1013, w_045_1014, w_045_1015, w_045_1016, w_045_1017, w_045_1018, w_045_1019, w_045_1020, w_045_1021, w_045_1022, w_045_1023, w_045_1025, w_045_1026, w_045_1028, w_045_1029, w_045_1031, w_045_1035, w_045_1036, w_045_1037, w_045_1045, w_045_1046, w_045_1048, w_045_1049, w_045_1051, w_045_1052, w_045_1055, w_045_1056, w_045_1057, w_045_1058, w_045_1059, w_045_1060, w_045_1061, w_045_1062, w_045_1063, w_045_1064, w_045_1065, w_045_1067, w_045_1069, w_045_1070, w_045_1072, w_045_1073, w_045_1074, w_045_1076, w_045_1077, w_045_1078, w_045_1079, w_045_1082, w_045_1083, w_045_1085, w_045_1086, w_045_1087, w_045_1088, w_045_1089, w_045_1091, w_045_1092, w_045_1093, w_045_1094, w_045_1095, w_045_1096, w_045_1097, w_045_1098, w_045_1100, w_045_1101, w_045_1102, w_045_1103, w_045_1105, w_045_1107, w_045_1110, w_045_1112, w_045_1113, w_045_1114, w_045_1115, w_045_1116, w_045_1117, w_045_1118, w_045_1119, w_045_1121, w_045_1124, w_045_1127, w_045_1128, w_045_1129, w_045_1130, w_045_1131, w_045_1132, w_045_1134, w_045_1135, w_045_1139, w_045_1140, w_045_1141, w_045_1142, w_045_1144, w_045_1145, w_045_1147, w_045_1149, w_045_1150, w_045_1152, w_045_1154, w_045_1155, w_045_1158, w_045_1160, w_045_1161, w_045_1162, w_045_1164, w_045_1166, w_045_1167, w_045_1169, w_045_1170, w_045_1171, w_045_1172, w_045_1173, w_045_1175, w_045_1176, w_045_1178, w_045_1179, w_045_1180, w_045_1181, w_045_1184, w_045_1185, w_045_1187, w_045_1188, w_045_1189, w_045_1191, w_045_1193, w_045_1195, w_045_1196, w_045_1197, w_045_1198, w_045_1199, w_045_1200, w_045_1202, w_045_1203, w_045_1204, w_045_1207, w_045_1208, w_045_1209, w_045_1216, w_045_1217, w_045_1218, w_045_1220, w_045_1221, w_045_1222, w_045_1223, w_045_1225, w_045_1227, w_045_1228, w_045_1229, w_045_1231, w_045_1232, w_045_1233, w_045_1234, w_045_1236, w_045_1238, w_045_1239, w_045_1240, w_045_1243, w_045_1244, w_045_1245, w_045_1246, w_045_1249, w_045_1250, w_045_1251, w_045_1253, w_045_1254, w_045_1255, w_045_1257, w_045_1258, w_045_1260, w_045_1261, w_045_1262, w_045_1263, w_045_1264, w_045_1265, w_045_1266, w_045_1268, w_045_1271, w_045_1272, w_045_1273, w_045_1275, w_045_1276, w_045_1279, w_045_1281, w_045_1283, w_045_1284, w_045_1286, w_045_1287, w_045_1288, w_045_1290, w_045_1292, w_045_1293, w_045_1294, w_045_1295, w_045_1297, w_045_1298, w_045_1299, w_045_1301, w_045_1302, w_045_1303, w_045_1305, w_045_1308, w_045_1309, w_045_1310, w_045_1313, w_045_1316, w_045_1317, w_045_1318, w_045_1320, w_045_1324, w_045_1326, w_045_1327, w_045_1328, w_045_1332, w_045_1334, w_045_1338, w_045_1339, w_045_1341, w_045_1342, w_045_1343, w_045_1345, w_045_1346, w_045_1347, w_045_1350, w_045_1352, w_045_1354, w_045_1355, w_045_1356, w_045_1358, w_045_1359, w_045_1360, w_045_1361, w_045_1362, w_045_1365, w_045_1367, w_045_1368, w_045_1370, w_045_1371, w_045_1372, w_045_1373, w_045_1374, w_045_1378, w_045_1379, w_045_1380, w_045_1381, w_045_1382, w_045_1384, w_045_1387, w_045_1388, w_045_1389, w_045_1390, w_045_1391, w_045_1392, w_045_1394, w_045_1395, w_045_1396, w_045_1397, w_045_1398, w_045_1399, w_045_1400, w_045_1401, w_045_1403, w_045_1404, w_045_1407, w_045_1408, w_045_1409, w_045_1411, w_045_1414, w_045_1416, w_045_1417, w_045_1418, w_045_1421, w_045_1422, w_045_1423, w_045_1424, w_045_1425, w_045_1426, w_045_1428, w_045_1429, w_045_1431, w_045_1432, w_045_1433, w_045_1434, w_045_1435, w_045_1436, w_045_1437, w_045_1438, w_045_1439, w_045_1440, w_045_1441, w_045_1442, w_045_1444, w_045_1445, w_045_1446, w_045_1447, w_045_1448, w_045_1449, w_045_1450, w_045_1451, w_045_1453, w_045_1454, w_045_1456, w_045_1457, w_045_1459, w_045_1461, w_045_1462, w_045_1464, w_045_1466, w_045_1467, w_045_1469, w_045_1473, w_045_1474, w_045_1477, w_045_1478, w_045_1480, w_045_1481, w_045_1483, w_045_1484, w_045_1487, w_045_1488, w_045_1489, w_045_1492, w_045_1493, w_045_1495, w_045_1498, w_045_1499, w_045_1500, w_045_1501, w_045_1502, w_045_1504, w_045_1505, w_045_1508, w_045_1509, w_045_1510, w_045_1511, w_045_1513, w_045_1514, w_045_1515, w_045_1516, w_045_1518, w_045_1519, w_045_1520, w_045_1521, w_045_1522, w_045_1523, w_045_1524, w_045_1525, w_045_1526, w_045_1528, w_045_1529, w_045_1530, w_045_1531, w_045_1532, w_045_1534, w_045_1535, w_045_1536, w_045_1537, w_045_1538, w_045_1540, w_045_1541, w_045_1542, w_045_1543, w_045_1544, w_045_1545, w_045_1548, w_045_1549, w_045_1551, w_045_1553, w_045_1554, w_045_1555, w_045_1556, w_045_1557, w_045_1558, w_045_1559, w_045_1560, w_045_1562, w_045_1563, w_045_1564, w_045_1565, w_045_1566, w_045_1567, w_045_1570, w_045_1571, w_045_1574, w_045_1575, w_045_1576, w_045_1577, w_045_1582, w_045_1583, w_045_1584, w_045_1587, w_045_1588, w_045_1590, w_045_1593, w_045_1595, w_045_1596, w_045_1598, w_045_1601, w_045_1602, w_045_1604, w_045_1605, w_045_1606, w_045_1607, w_045_1608, w_045_1609, w_045_1610, w_045_1611, w_045_1612, w_045_1613, w_045_1614, w_045_1615, w_045_1616, w_045_1617, w_045_1618, w_045_1619, w_045_1620, w_045_1621, w_045_1623, w_045_1624, w_045_1625, w_045_1626, w_045_1627, w_045_1628, w_045_1629, w_045_1630, w_045_1632, w_045_1633, w_045_1635, w_045_1636, w_045_1637, w_045_1638, w_045_1639, w_045_1641, w_045_1642, w_045_1643, w_045_1644, w_045_1645, w_045_1646, w_045_1647, w_045_1648, w_045_1649, w_045_1650, w_045_1651, w_045_1652, w_045_1653, w_045_1655, w_045_1658, w_045_1659, w_045_1660, w_045_1661, w_045_1662, w_045_1665, w_045_1666, w_045_1667, w_045_1668, w_045_1669, w_045_1670, w_045_1671, w_045_1672, w_045_1673, w_045_1675, w_045_1676, w_045_1677, w_045_1678, w_045_1679, w_045_1680, w_045_1681, w_045_1682, w_045_1683, w_045_1688, w_045_1689, w_045_1690, w_045_1693, w_045_1694, w_045_1695, w_045_1696, w_045_1697, w_045_1698, w_045_1699, w_045_1701, w_045_1702, w_045_1704, w_045_1708, w_045_1709, w_045_1712, w_045_1713, w_045_1714, w_045_1715, w_045_1716, w_045_1718, w_045_1720, w_045_1721, w_045_1723, w_045_1724, w_045_1725, w_045_1726, w_045_1727, w_045_1730, w_045_1731, w_045_1732, w_045_1733, w_045_1737, w_045_1738, w_045_1740, w_045_1742, w_045_1743, w_045_1744, w_045_1745, w_045_1746, w_045_1747, w_045_1749, w_045_1750, w_045_1752, w_045_1753, w_045_1754, w_045_1755, w_045_1756, w_045_1758, w_045_1760, w_045_1761, w_045_1763, w_045_1764, w_045_1765, w_045_1766, w_045_1767, w_045_1768, w_045_1769, w_045_1770, w_045_1772, w_045_1773, w_045_1774, w_045_1776, w_045_1777, w_045_1778, w_045_1779, w_045_1782, w_045_1783, w_045_1784, w_045_1785, w_045_1787, w_045_1791, w_045_1792, w_045_1793, w_045_1794, w_045_1796, w_045_1800, w_045_1801, w_045_1802, w_045_1803, w_045_1804, w_045_1805, w_045_1807, w_045_1808, w_045_1812, w_045_1813, w_045_1814, w_045_1815, w_045_1817, w_045_1818, w_045_1820, w_045_1821, w_045_1822, w_045_1823, w_045_1824, w_045_1825, w_045_1827, w_045_1828, w_045_1829, w_045_1830, w_045_1831, w_045_1832, w_045_1834, w_045_1837, w_045_1840, w_045_1842, w_045_1845, w_045_1846, w_045_1847, w_045_1848, w_045_1849, w_045_1850, w_045_1851, w_045_1852, w_045_1853, w_045_1854, w_045_1855, w_045_1856, w_045_1859, w_045_1860, w_045_1861, w_045_1862, w_045_1863, w_045_1865, w_045_1866, w_045_1868, w_045_1870, w_045_1871, w_045_1872, w_045_1873, w_045_1874, w_045_1875, w_045_1877, w_045_1879, w_045_1880, w_045_1881, w_045_1884, w_045_1885, w_045_1886, w_045_1887, w_045_1888, w_045_1890, w_045_1891, w_045_1892, w_045_1893, w_045_1894, w_045_1898, w_045_1899, w_045_1900, w_045_1901, w_045_1902, w_045_1903, w_045_1904, w_045_1905, w_045_1906, w_045_1907, w_045_1908, w_045_1909, w_045_1910, w_045_1911, w_045_1912, w_045_1913, w_045_1915, w_045_1916, w_045_1917, w_045_1919, w_045_1920, w_045_1922, w_045_1923, w_045_1924, w_045_1925, w_045_1926, w_045_1928, w_045_1929, w_045_1930, w_045_1931, w_045_1932, w_045_1933, w_045_1936, w_045_1937, w_045_1939, w_045_1940, w_045_1941, w_045_1942, w_045_1943, w_045_1944, w_045_1946, w_045_1947, w_045_1948, w_045_1949, w_045_1950, w_045_1954, w_045_1955, w_045_1957, w_045_1961, w_045_1962, w_045_1963, w_045_1966, w_045_1967, w_045_1968, w_045_1970, w_045_1972, w_045_1975, w_045_1976, w_045_1977, w_045_1978, w_045_1979, w_045_1980, w_045_1981, w_045_1984, w_045_1985, w_045_1986, w_045_1987, w_045_1989, w_045_1990, w_045_1991, w_045_1993, w_045_1994, w_045_1995, w_045_1996, w_045_1997, w_045_2001, w_045_2003, w_045_2004, w_045_2005, w_045_2006, w_045_2007, w_045_2008, w_045_2009, w_045_2011, w_045_2013, w_045_2015, w_045_2016, w_045_2018, w_045_2019, w_045_2020, w_045_2021, w_045_2022, w_045_2023, w_045_2024, w_045_2025, w_045_2028, w_045_2029, w_045_2030, w_045_2031, w_045_2032, w_045_2033, w_045_2035, w_045_2037, w_045_2039, w_045_2040, w_045_2041, w_045_2042, w_045_2043, w_045_2044, w_045_2045, w_045_2046, w_045_2048, w_045_2050, w_045_2053, w_045_2054, w_045_2056, w_045_2057, w_045_2060, w_045_2061, w_045_2062, w_045_2063, w_045_2064, w_045_2065, w_045_2066, w_045_2067, w_045_2069, w_045_2070, w_045_2071, w_045_2072, w_045_2074, w_045_2076, w_045_2077, w_045_2078, w_045_2079, w_045_2086, w_045_2087, w_045_2089, w_045_2092, w_045_2094, w_045_2097, w_045_2099, w_045_2100, w_045_2101, w_045_2102, w_045_2103, w_045_2104, w_045_2106, w_045_2107, w_045_2108, w_045_2110, w_045_2111, w_045_2112, w_045_2113, w_045_2114, w_045_2118, w_045_2119, w_045_2120, w_045_2121, w_045_2122, w_045_2123, w_045_2124, w_045_2125, w_045_2129, w_045_2133, w_045_2134, w_045_2135, w_045_2136, w_045_2137, w_045_2138, w_045_2139, w_045_2140, w_045_2142, w_045_2145, w_045_2146, w_045_2147, w_045_2149, w_045_2150, w_045_2151, w_045_2152, w_045_2153, w_045_2154, w_045_2156, w_045_2157, w_045_2158, w_045_2159, w_045_2161, w_045_2162, w_045_2163, w_045_2164, w_045_2166, w_045_2167, w_045_2170, w_045_2171, w_045_2172, w_045_2173, w_045_2174, w_045_2175, w_045_2176, w_045_2177, w_045_2178, w_045_2179, w_045_2180, w_045_2181, w_045_2182, w_045_2183, w_045_2184, w_045_2185, w_045_2186, w_045_2187, w_045_2189, w_045_2190, w_045_2194, w_045_2195, w_045_2196, w_045_2198, w_045_2199, w_045_2200, w_045_2201, w_045_2202, w_045_2203, w_045_2205, w_045_2206, w_045_2207, w_045_2208, w_045_2209, w_045_2210, w_045_2211, w_045_2212, w_045_2213, w_045_2215, w_045_2216, w_045_2217, w_045_2218, w_045_2219, w_045_2221, w_045_2222, w_045_2225, w_045_2226, w_045_2227, w_045_2228, w_045_2229, w_045_2232, w_045_2234, w_045_2235, w_045_2236, w_045_2238, w_045_2239, w_045_2240, w_045_2242, w_045_2243, w_045_2244, w_045_2247, w_045_2248, w_045_2251, w_045_2252, w_045_2253, w_045_2255, w_045_2257, w_045_2258, w_045_2259, w_045_2262, w_045_2266, w_045_2268, w_045_2270, w_045_2271, w_045_2274, w_045_2275, w_045_2277, w_045_2279, w_045_2283, w_045_2284, w_045_2285, w_045_2288, w_045_2291, w_045_2294, w_045_2296, w_045_2299, w_045_2304, w_045_2309, w_045_2312, w_045_2316, w_045_2320, w_045_2325, w_045_2326, w_045_2327, w_045_2330, w_045_2331, w_045_2332, w_045_2333, w_045_2338, w_045_2339, w_045_2341, w_045_2348, w_045_2349, w_045_2351, w_045_2353, w_045_2355, w_045_2357, w_045_2361, w_045_2364, w_045_2367, w_045_2370, w_045_2372, w_045_2374, w_045_2380, w_045_2382, w_045_2383, w_045_2385, w_045_2386, w_045_2389, w_045_2390, w_045_2391, w_045_2393, w_045_2396, w_045_2398, w_045_2402, w_045_2405, w_045_2406, w_045_2408, w_045_2409, w_045_2412, w_045_2414, w_045_2420, w_045_2425, w_045_2427, w_045_2429, w_045_2430, w_045_2431, w_045_2432, w_045_2433, w_045_2435, w_045_2438, w_045_2444, w_045_2445, w_045_2446, w_045_2447, w_045_2454, w_045_2459, w_045_2460, w_045_2467, w_045_2468, w_045_2473, w_045_2474, w_045_2476, w_045_2477, w_045_2478, w_045_2479, w_045_2481, w_045_2484, w_045_2488, w_045_2490, w_045_2492, w_045_2493, w_045_2494, w_045_2498, w_045_2501, w_045_2503, w_045_2506, w_045_2508, w_045_2509, w_045_2510, w_045_2512, w_045_2516, w_045_2518, w_045_2519, w_045_2520, w_045_2522, w_045_2523, w_045_2525, w_045_2526, w_045_2527, w_045_2530, w_045_2533, w_045_2545, w_045_2547, w_045_2549, w_045_2550, w_045_2554, w_045_2555, w_045_2557, w_045_2558, w_045_2560, w_045_2563, w_045_2569, w_045_2572, w_045_2575, w_045_2576, w_045_2577, w_045_2578, w_045_2580, w_045_2582, w_045_2583, w_045_2589, w_045_2590, w_045_2592, w_045_2596, w_045_2597, w_045_2598, w_045_2602, w_045_2605, w_045_2607, w_045_2610, w_045_2612, w_045_2615, w_045_2616, w_045_2626, w_045_2627, w_045_2629, w_045_2630, w_045_2631, w_045_2637, w_045_2639, w_045_2643, w_045_2646, w_045_2649, w_045_2650, w_045_2653, w_045_2655, w_045_2660, w_045_2664, w_045_2668, w_045_2670, w_045_2672, w_045_2676, w_045_2677, w_045_2683, w_045_2684, w_045_2686, w_045_2687, w_045_2689, w_045_2693, w_045_2694, w_045_2695, w_045_2696, w_045_2699, w_045_2701, w_045_2704, w_045_2707, w_045_2711, w_045_2713, w_045_2716, w_045_2717, w_045_2720, w_045_2721, w_045_2722, w_045_2726, w_045_2729, w_045_2735, w_045_2739, w_045_2745, w_045_2747, w_045_2749, w_045_2750, w_045_2751, w_045_2752, w_045_2756, w_045_2757, w_045_2760, w_045_2761, w_045_2765, w_045_2766, w_045_2767, w_045_2769, w_045_2772, w_045_2775, w_045_2776, w_045_2778, w_045_2782, w_045_2788, w_045_2789, w_045_2790, w_045_2791, w_045_2792, w_045_2793, w_045_2794, w_045_2795, w_045_2797, w_045_2798, w_045_2802, w_045_2805, w_045_2806, w_045_2808, w_045_2813, w_045_2814, w_045_2815, w_045_2818, w_045_2824, w_045_2825, w_045_2828, w_045_2830, w_045_2832, w_045_2833, w_045_2834, w_045_2836, w_045_2837, w_045_2839, w_045_2840, w_045_2841, w_045_2844, w_045_2845, w_045_2846, w_045_2850, w_045_2853, w_045_2856, w_045_2857, w_045_2858, w_045_2859, w_045_2862, w_045_2864, w_045_2865, w_045_2867, w_045_2871, w_045_2873, w_045_2877, w_045_2882, w_045_2885, w_045_2886, w_045_2887, w_045_2889, w_045_2894, w_045_2895, w_045_2896, w_045_2899, w_045_2901, w_045_2904, w_045_2905, w_045_2906, w_045_2907, w_045_2908, w_045_2912, w_045_2914, w_045_2917, w_045_2918, w_045_2920, w_045_2921, w_045_2922, w_045_2925, w_045_2927, w_045_2928, w_045_2929, w_045_2931, w_045_2932, w_045_2935, w_045_2937, w_045_2938, w_045_2939, w_045_2942, w_045_2943, w_045_2944, w_045_2945, w_045_2949, w_045_2950, w_045_2955, w_045_2957, w_045_2959, w_045_2960, w_045_2967, w_045_2968, w_045_2969, w_045_2970, w_045_2972, w_045_2973, w_045_2974, w_045_2975, w_045_2978, w_045_2982, w_045_2983, w_045_2986, w_045_2988, w_045_2991, w_045_2992, w_045_2994, w_045_2997, w_045_3000, w_045_3004, w_045_3006, w_045_3008, w_045_3010, w_045_3011, w_045_3013, w_045_3014, w_045_3019, w_045_3020, w_045_3025, w_045_3026, w_045_3027, w_045_3028, w_045_3030, w_045_3034, w_045_3036, w_045_3039, w_045_3041, w_045_3042, w_045_3043, w_045_3044, w_045_3046, w_045_3047, w_045_3050, w_045_3052, w_045_3056, w_045_3064, w_045_3065, w_045_3066, w_045_3067, w_045_3069, w_045_3071, w_045_3075, w_045_3077, w_045_3078, w_045_3083, w_045_3085, w_045_3086, w_045_3087, w_045_3089, w_045_3092, w_045_3095, w_045_3099, w_045_3101, w_045_3102, w_045_3103, w_045_3107, w_045_3110, w_045_3118, w_045_3119, w_045_3126, w_045_3127, w_045_3128, w_045_3131, w_045_3132, w_045_3133, w_045_3134, w_045_3140, w_045_3141, w_045_3142, w_045_3143, w_045_3144, w_045_3147, w_045_3149, w_045_3150, w_045_3153, w_045_3154, w_045_3155, w_045_3158, w_045_3159, w_045_3161, w_045_3163, w_045_3164, w_045_3165, w_045_3166, w_045_3167, w_045_3172, w_045_3173, w_045_3179, w_045_3181, w_045_3182, w_045_3185, w_045_3186, w_045_3193, w_045_3203, w_045_3204, w_045_3206, w_045_3208, w_045_3209, w_045_3212, w_045_3213, w_045_3214, w_045_3217, w_045_3220, w_045_3222, w_045_3230, w_045_3234, w_045_3235, w_045_3236, w_045_3239, w_045_3241, w_045_3245, w_045_3249, w_045_3250, w_045_3252, w_045_3253, w_045_3254, w_045_3263, w_045_3266, w_045_3270, w_045_3276, w_045_3278, w_045_3281, w_045_3282, w_045_3284, w_045_3287, w_045_3289, w_045_3290, w_045_3291, w_045_3293, w_045_3294, w_045_3295, w_045_3299, w_045_3300, w_045_3304, w_045_3305, w_045_3306, w_045_3308, w_045_3309, w_045_3312, w_045_3318, w_045_3323, w_045_3324, w_045_3327, w_045_3328, w_045_3332, w_045_3335, w_045_3344, w_045_3346, w_045_3355, w_045_3359, w_045_3360, w_045_3362, w_045_3364, w_045_3365, w_045_3367, w_045_3371, w_045_3378, w_045_3379, w_045_3380, w_045_3383, w_045_3385, w_045_3386, w_045_3387, w_045_3388, w_045_3390, w_045_3393, w_045_3394, w_045_3395, w_045_3396, w_045_3397, w_045_3398, w_045_3400, w_045_3402, w_045_3405, w_045_3407, w_045_3410, w_045_3414, w_045_3418, w_045_3419, w_045_3425, w_045_3429, w_045_3431, w_045_3435, w_045_3436, w_045_3440, w_045_3443, w_045_3447, w_045_3448, w_045_3449, w_045_3450, w_045_3451, w_045_3452, w_045_3454, w_045_3455, w_045_3456, w_045_3461, w_045_3462, w_045_3463, w_045_3464, w_045_3465, w_045_3466, w_045_3467, w_045_3470, w_045_3471, w_045_3472, w_045_3474, w_045_3475, w_045_3476, w_045_3477, w_045_3478, w_045_3480, w_045_3484, w_045_3485, w_045_3487, w_045_3489, w_045_3490, w_045_3491, w_045_3493, w_045_3494, w_045_3499, w_045_3500, w_045_3505, w_045_3506, w_045_3507, w_045_3508, w_045_3511, w_045_3513, w_045_3514, w_045_3515, w_045_3516, w_045_3517, w_045_3519, w_045_3523, w_045_3524, w_045_3525, w_045_3526, w_045_3529, w_045_3534, w_045_3538, w_045_3539, w_045_3541, w_045_3542, w_045_3543, w_045_3544, w_045_3545, w_045_3546, w_045_3554, w_045_3555, w_045_3556, w_045_3558, w_045_3559, w_045_3562, w_045_3564, w_045_3569, w_045_3571, w_045_3574, w_045_3575, w_045_3580, w_045_3581, w_045_3582, w_045_3584, w_045_3585, w_045_3588, w_045_3589, w_045_3591, w_045_3592, w_045_3593, w_045_3594, w_045_3596, w_045_3600, w_045_3603, w_045_3606, w_045_3608, w_045_3610, w_045_3611, w_045_3614, w_045_3615, w_045_3617, w_045_3618, w_045_3624, w_045_3626, w_045_3627, w_045_3632, w_045_3634, w_045_3635, w_045_3636, w_045_3637, w_045_3640, w_045_3643, w_045_3645, w_045_3652, w_045_3655, w_045_3656, w_045_3657, w_045_3658, w_045_3659, w_045_3660, w_045_3662, w_045_3666, w_045_3669, w_045_3670, w_045_3672, w_045_3675, w_045_3676, w_045_3677, w_045_3678, w_045_3679, w_045_3680, w_045_3685, w_045_3686, w_045_3690, w_045_3691, w_045_3692, w_045_3693, w_045_3695, w_045_3697, w_045_3698, w_045_3699, w_045_3701, w_045_3704, w_045_3705, w_045_3706, w_045_3711, w_045_3715, w_045_3716, w_045_3720, w_045_3721, w_045_3722, w_045_3725, w_045_3728, w_045_3730, w_045_3731, w_045_3735, w_045_3736, w_045_3737, w_045_3740, w_045_3742, w_045_3747, w_045_3750, w_045_3751, w_045_3754, w_045_3757, w_045_3758, w_045_3759, w_045_3762, w_045_3764, w_045_3765, w_045_3771, w_045_3781, w_045_3782, w_045_3784, w_045_3786, w_045_3787, w_045_3790, w_045_3791, w_045_3792, w_045_3793, w_045_3794, w_045_3797, w_045_3798, w_045_3799, w_045_3802, w_045_3804, w_045_3805, w_045_3809, w_045_3820, w_045_3826, w_045_3827, w_045_3828, w_045_3830, w_045_3831, w_045_3835, w_045_3836, w_045_3837, w_045_3839, w_045_3843, w_045_3844, w_045_3845, w_045_3846, w_045_3851, w_045_3853, w_045_3856, w_045_3858, w_045_3859, w_045_3862, w_045_3866, w_045_3867, w_045_3869, w_045_3873, w_045_3876, w_045_3879, w_045_3881, w_045_3882, w_045_3884, w_045_3885, w_045_3886, w_045_3887, w_045_3888, w_045_3890, w_045_3891, w_045_3892, w_045_3896, w_045_3897, w_045_3898, w_045_3899, w_045_3902, w_045_3905, w_045_3907, w_045_3912, w_045_3914, w_045_3920, w_045_3921, w_045_3925, w_045_3928, w_045_3930, w_045_3932, w_045_3935, w_045_3937, w_045_3938, w_045_3939, w_045_3941, w_045_3943, w_045_3944, w_045_3948, w_045_3950, w_045_3951, w_045_3953, w_045_3955, w_045_3958, w_045_3960, w_045_3962, w_045_3963, w_045_3965, w_045_3966, w_045_3969, w_045_3974, w_045_3985, w_045_3986, w_045_3988, w_045_3990, w_045_3992, w_045_3994, w_045_4000, w_045_4006, w_045_4014, w_045_4023, w_045_4025, w_045_4027, w_045_4029, w_045_4030, w_045_4034, w_045_4035, w_045_4037, w_045_4040, w_045_4041, w_045_4044, w_045_4046, w_045_4048, w_045_4049, w_045_4050, w_045_4055, w_045_4056, w_045_4058, w_045_4059, w_045_4062, w_045_4064, w_045_4066, w_045_4069, w_045_4072, w_045_4075, w_045_4077, w_045_4079, w_045_4083, w_045_4085, w_045_4094, w_045_4096, w_045_4098, w_045_4101, w_045_4103, w_045_4104, w_045_4106, w_045_4107, w_045_4108, w_045_4109, w_045_4110, w_045_4116, w_045_4119, w_045_4120, w_045_4121, w_045_4122, w_045_4124, w_045_4127, w_045_4128, w_045_4130, w_045_4131, w_045_4134, w_045_4136, w_045_4137, w_045_4138, w_045_4141, w_045_4142, w_045_4143, w_045_4145, w_045_4148, w_045_4150, w_045_4155, w_045_4158, w_045_4159, w_045_4162, w_045_4163, w_045_4164, w_045_4169, w_045_4173, w_045_4174, w_045_4181, w_045_4182, w_045_4189, w_045_4190, w_045_4194, w_045_4197, w_045_4200, w_045_4201, w_045_4202, w_045_4203, w_045_4207, w_045_4210, w_045_4213, w_045_4215, w_045_4216, w_045_4218, w_045_4220, w_045_4226, w_045_4227, w_045_4233, w_045_4235, w_045_4237, w_045_4238, w_045_4240, w_045_4241, w_045_4242, w_045_4243, w_045_4244, w_045_4246, w_045_4248, w_045_4250, w_045_4251, w_045_4254, w_045_4256, w_045_4258, w_045_4265, w_045_4267, w_045_4268, w_045_4279, w_045_4280, w_045_4282, w_045_4283, w_045_4288, w_045_4290, w_045_4291, w_045_4292, w_045_4296, w_045_4297, w_045_4301, w_045_4303, w_045_4304, w_045_4316, w_045_4317, w_045_4320, w_045_4322, w_045_4323, w_045_4324, w_045_4327, w_045_4330, w_045_4334, w_045_4337, w_045_4340, w_045_4343, w_045_4346, w_045_4347, w_045_4348, w_045_4349, w_045_4351, w_045_4354, w_045_4355, w_045_4356, w_045_4359, w_045_4360, w_045_4361, w_045_4363, w_045_4365, w_045_4372, w_045_4375, w_045_4377, w_045_4378, w_045_4380, w_045_4382, w_045_4389, w_045_4394, w_045_4397, w_045_4401, w_045_4406, w_045_4409, w_045_4410, w_045_4414, w_045_4415, w_045_4416, w_045_4418, w_045_4419, w_045_4424, w_045_4425, w_045_4426, w_045_4429, w_045_4430, w_045_4431, w_045_4432, w_045_4437, w_045_4438, w_045_4439, w_045_4443, w_045_4444, w_045_4445, w_045_4447, w_045_4450, w_045_4452, w_045_4453, w_045_4454, w_045_4459, w_045_4462, w_045_4471, w_045_4473, w_045_4474, w_045_4475, w_045_4476, w_045_4480, w_045_4486, w_045_4488, w_045_4491, w_045_4494, w_045_4498, w_045_4500, w_045_4502, w_045_4503, w_045_4504, w_045_4506, w_045_4507, w_045_4508, w_045_4512, w_045_4514, w_045_4520, w_045_4521, w_045_4525, w_045_4527, w_045_4529, w_045_4531, w_045_4532, w_045_4533, w_045_4534, w_045_4536, w_045_4538, w_045_4542, w_045_4543, w_045_4546, w_045_4548, w_045_4549, w_045_4552, w_045_4556, w_045_4557, w_045_4558, w_045_4559, w_045_4561, w_045_4562, w_045_4564, w_045_4566, w_045_4568, w_045_4569, w_045_4571, w_045_4574, w_045_4575, w_045_4577, w_045_4578, w_045_4583, w_045_4584, w_045_4585, w_045_4587, w_045_4588, w_045_4589, w_045_4591, w_045_4594, w_045_4601, w_045_4604, w_045_4607, w_045_4608, w_045_4610, w_045_4615, w_045_4618, w_045_4621, w_045_4623, w_045_4628, w_045_4629, w_045_4632, w_045_4633, w_045_4635, w_045_4636, w_045_4637, w_045_4640, w_045_4641, w_045_4642, w_045_4643, w_045_4644, w_045_4650, w_045_4655, w_045_4662, w_045_4667, w_045_4669, w_045_4670, w_045_4672, w_045_4676, w_045_4677, w_045_4679, w_045_4682, w_045_4685, w_045_4686, w_045_4688, w_045_4692, w_045_4694, w_045_4695, w_045_4697, w_045_4698, w_045_4699, w_045_4701, w_045_4703, w_045_4704, w_045_4705, w_045_4707, w_045_4708, w_045_4709, w_045_4715, w_045_4716, w_045_4717, w_045_4718, w_045_4719, w_045_4721, w_045_4725, w_045_4728, w_045_4733, w_045_4738, w_045_4740, w_045_4744, w_045_4745, w_045_4747, w_045_4749, w_045_4752, w_045_4754, w_045_4759, w_045_4760, w_045_4761, w_045_4765, w_045_4767, w_045_4769, w_045_4774, w_045_4776, w_045_4779, w_045_4780, w_045_4782, w_045_4788, w_045_4790, w_045_4791, w_045_4792, w_045_4793, w_045_4794, w_045_4798, w_045_4802, w_045_4803, w_045_4807, w_045_4808, w_045_4812, w_045_4814, w_045_4816, w_045_4819, w_045_4820, w_045_4827, w_045_4831, w_045_4834, w_045_4835, w_045_4836, w_045_4839, w_045_4841, w_045_4842, w_045_4843, w_045_4851, w_045_4853, w_045_4856, w_045_4873, w_045_4874, w_045_4875, w_045_4882, w_045_4883, w_045_4884, w_045_4890, w_045_4891, w_045_4897, w_045_4899, w_045_4900, w_045_4901, w_045_4903, w_045_4905, w_045_4908, w_045_4910, w_045_4911, w_045_4913, w_045_4915, w_045_4918, w_045_4921, w_045_4924, w_045_4926, w_045_4929, w_045_4933, w_045_4934, w_045_4935, w_045_4936, w_045_4937, w_045_4938, w_045_4939, w_045_4941, w_045_4942, w_045_4943, w_045_4944, w_045_4945, w_045_4946, w_045_4949, w_045_4953, w_045_4955, w_045_4958, w_045_4959, w_045_4961, w_045_4967, w_045_4969, w_045_4971, w_045_4972, w_045_4973, w_045_4974, w_045_4975, w_045_4983, w_045_4984, w_045_4985, w_045_4986, w_045_4987, w_045_4991, w_045_4992, w_045_4994, w_045_4999, w_045_5000, w_045_5003, w_045_5004, w_045_5005, w_045_5011, w_045_5014, w_045_5015, w_045_5017, w_045_5018, w_045_5021, w_045_5022, w_045_5026, w_045_5030, w_045_5036, w_045_5037, w_045_5039, w_045_5041, w_045_5048, w_045_5049, w_045_5051, w_045_5052, w_045_5057, w_045_5058, w_045_5059, w_045_5062, w_045_5064, w_045_5069, w_045_5073, w_045_5074, w_045_5075, w_045_5076, w_045_5077, w_045_5079, w_045_5081, w_045_5083, w_045_5084, w_045_5087, w_045_5088, w_045_5091, w_045_5094, w_045_5096, w_045_5097, w_045_5100, w_045_5104, w_045_5106, w_045_5109, w_045_5111, w_045_5113, w_045_5114, w_045_5116, w_045_5117, w_045_5118, w_045_5121, w_045_5123, w_045_5127, w_045_5129, w_045_5130, w_045_5131, w_045_5132, w_045_5135, w_045_5138, w_045_5139, w_045_5141, w_045_5143, w_045_5144, w_045_5153, w_045_5157, w_045_5158, w_045_5159, w_045_5165, w_045_5166, w_045_5167, w_045_5168, w_045_5169, w_045_5173, w_045_5178, w_045_5182, w_045_5185, w_045_5186, w_045_5187, w_045_5188, w_045_5189, w_045_5191, w_045_5193, w_045_5194, w_045_5195, w_045_5198, w_045_5203, w_045_5205, w_045_5207, w_045_5210, w_045_5213, w_045_5217, w_045_5220, w_045_5221, w_045_5222, w_045_5227, w_045_5230, w_045_5232, w_045_5236, w_045_5240, w_045_5244, w_045_5246, w_045_5247, w_045_5251, w_045_5252, w_045_5255, w_045_5256, w_045_5258, w_045_5264, w_045_5271, w_045_5275, w_045_5277, w_045_5279, w_045_5280, w_045_5281, w_045_5283, w_045_5286, w_045_5295, w_045_5299, w_045_5301, w_045_5303, w_045_5305, w_045_5309, w_045_5310, w_045_5311, w_045_5313, w_045_5320, w_045_5322, w_045_5323, w_045_5327, w_045_5328, w_045_5330, w_045_5335, w_045_5336, w_045_5338, w_045_5342, w_045_5343, w_045_5344, w_045_5348, w_045_5350, w_045_5352, w_045_5354, w_045_5358, w_045_5361, w_045_5366, w_045_5370, w_045_5372, w_045_5375, w_045_5376, w_045_5381, w_045_5382, w_045_5384, w_045_5385, w_045_5387, w_045_5389, w_045_5392, w_045_5394, w_045_5395, w_045_5399, w_045_5401, w_045_5402, w_045_5405, w_045_5408, w_045_5411, w_045_5412, w_045_5414, w_045_5415, w_045_5416, w_045_5423, w_045_5425, w_045_5428, w_045_5430, w_045_5431, w_045_5435, w_045_5436, w_045_5438, w_045_5441, w_045_5442, w_045_5446, w_045_5449, w_045_5451, w_045_5455, w_045_5457, w_045_5458, w_045_5459, w_045_5461, w_045_5462, w_045_5465, w_045_5468, w_045_5469, w_045_5473, w_045_5477, w_045_5478, w_045_5481, w_045_5485, w_045_5486, w_045_5489, w_045_5490, w_045_5492, w_045_5493, w_045_5496, w_045_5501, w_045_5502, w_045_5503, w_045_5506, w_045_5507, w_045_5508, w_045_5509, w_045_5511, w_045_5512, w_045_5515, w_045_5517, w_045_5518, w_045_5520, w_045_5522, w_045_5524, w_045_5527, w_045_5529, w_045_5530, w_045_5531, w_045_5532, w_045_5535, w_045_5536, w_045_5538, w_045_5539, w_045_5540, w_045_5542, w_045_5544, w_045_5550, w_045_5551, w_045_5552, w_045_5553, w_045_5557, w_045_5558, w_045_5560, w_045_5563, w_045_5566, w_045_5567, w_045_5571, w_045_5572, w_045_5574, w_045_5577, w_045_5578, w_045_5581, w_045_5582, w_045_5584, w_045_5585, w_045_5586, w_045_5587, w_045_5589, w_045_5594, w_045_5595, w_045_5596, w_045_5597, w_045_5598, w_045_5602, w_045_5603, w_045_5605, w_045_5606, w_045_5607, w_045_5608, w_045_5612, w_045_5614, w_045_5615, w_045_5619, w_045_5620, w_045_5622, w_045_5623, w_045_5624, w_045_5630, w_045_5633, w_045_5636, w_045_5637, w_045_5638, w_045_5646, w_045_5647, w_045_5649, w_045_5653, w_045_5654, w_045_5655, w_045_5656, w_045_5658, w_045_5659, w_045_5660, w_045_5661, w_045_5663, w_045_5664, w_045_5666, w_045_5667, w_045_5669, w_045_5672, w_045_5673, w_045_5677, w_045_5678, w_045_5680, w_045_5682, w_045_5686, w_045_5687, w_045_5691, w_045_5692, w_045_5695, w_045_5703, w_045_5704, w_045_5707, w_045_5711, w_045_5713, w_045_5715, w_045_5716, w_045_5717, w_045_5718, w_045_5722, w_045_5723, w_045_5725, w_045_5726, w_045_5729, w_045_5730, w_045_5731, w_045_5732, w_045_5733, w_045_5736, w_045_5737, w_045_5739, w_045_5740, w_045_5741, w_045_5744, w_045_5745, w_045_5747, w_045_5749, w_045_5752, w_045_5754, w_045_5757, w_045_5758, w_045_5759, w_045_5761, w_045_5765, w_045_5766, w_045_5770, w_045_5772, w_045_5773, w_045_5779, w_045_5781, w_045_5783, w_045_5784, w_045_5787, w_045_5788, w_045_5789, w_045_5790, w_045_5791, w_045_5792, w_045_5794, w_045_5795, w_045_5797, w_045_5799, w_045_5800, w_045_5801, w_045_5804, w_045_5805, w_045_5806, w_045_5811, w_045_5815, w_045_5816, w_045_5818, w_045_5819, w_045_5820, w_045_5822, w_045_5823, w_045_5826, w_045_5829, w_045_5830, w_045_5831, w_045_5833, w_045_5834, w_045_5835, w_045_5836, w_045_5842, w_045_5850, w_045_5851, w_045_5852, w_045_5854, w_045_5857, w_045_5859, w_045_5863, w_045_5864, w_045_5865, w_045_5866, w_045_5867, w_045_5869, w_045_5870, w_045_5871, w_045_5874, w_045_5875, w_045_5877, w_045_5878, w_045_5879, w_045_5880, w_045_5881, w_045_5887, w_045_5888, w_045_5890, w_045_5895, w_045_5896, w_045_5899, w_045_5904, w_045_5910, w_045_5914, w_045_5915, w_045_5916, w_045_5917, w_045_5918, w_045_5919, w_045_5921, w_045_5922, w_045_5926, w_045_5928, w_045_5929, w_045_5930, w_045_5931, w_045_5939, w_045_5943, w_045_5945, w_045_5946, w_045_5947, w_045_5948, w_045_5954, w_045_5957, w_045_5958, w_045_5959, w_045_5960, w_045_5961, w_045_5964, w_045_5967, w_045_5968, w_045_5970, w_045_5972, w_045_5973, w_045_5978, w_045_5984, w_045_5985, w_045_5987, w_045_5988, w_045_5991, w_045_5993, w_045_5995, w_045_5997, w_045_5999, w_045_6004, w_045_6005, w_045_6006, w_045_6008, w_045_6010, w_045_6012, w_045_6020, w_045_6022, w_045_6023, w_045_6027, w_045_6028, w_045_6029, w_045_6031, w_045_6035, w_045_6040, w_045_6041, w_045_6043, w_045_6044, w_045_6045, w_045_6046, w_045_6047, w_045_6048, w_045_6049, w_045_6051, w_045_6056, w_045_6059, w_045_6064, w_045_6065, w_045_6066, w_045_6069, w_045_6072, w_045_6073, w_045_6077, w_045_6080, w_045_6082, w_045_6085, w_045_6087, w_045_6088, w_045_6089, w_045_6090, w_045_6091, w_045_6093, w_045_6094, w_045_6095, w_045_6096, w_045_6097, w_045_6098, w_045_6099, w_045_6100, w_045_6102, w_045_6104, w_045_6109, w_045_6110, w_045_6111, w_045_6114, w_045_6120, w_045_6126, w_045_6127, w_045_6129, w_045_6130, w_045_6136, w_045_6138, w_045_6139, w_045_6140, w_045_6145, w_045_6150, w_045_6151, w_045_6163, w_045_6167, w_045_6168, w_045_6169, w_045_6170, w_045_6176, w_045_6177, w_045_6178, w_045_6179, w_045_6182, w_045_6183, w_045_6186, w_045_6188, w_045_6189, w_045_6191, w_045_6192, w_045_6193, w_045_6195, w_045_6196, w_045_6202, w_045_6204, w_045_6205, w_045_6209, w_045_6215, w_045_6216, w_045_6217, w_045_6218, w_045_6219, w_045_6224, w_045_6225, w_045_6226, w_045_6227, w_045_6229, w_045_6233, w_045_6234, w_045_6235, w_045_6236, w_045_6239, w_045_6240, w_045_6241, w_045_6246, w_045_6249, w_045_6251, w_045_6254, w_045_6255, w_045_6259, w_045_6260, w_045_6262, w_045_6263, w_045_6267, w_045_6268, w_045_6272, w_045_6273, w_045_6274, w_045_6275, w_045_6278, w_045_6279, w_045_6282, w_045_6284, w_045_6285, w_045_6286, w_045_6288, w_045_6292, w_045_6296, w_045_6297, w_045_6298, w_045_6299, w_045_6301, w_045_6302, w_045_6304, w_045_6306, w_045_6307, w_045_6309, w_045_6310, w_045_6313, w_045_6314, w_045_6318, w_045_6326, w_045_6327, w_045_6328, w_045_6329, w_045_6330, w_045_6331, w_045_6334, w_045_6335, w_045_6336, w_045_6337, w_045_6340, w_045_6343, w_045_6346, w_045_6347, w_045_6349, w_045_6351, w_045_6354, w_045_6355, w_045_6358, w_045_6359, w_045_6362, w_045_6363, w_045_6364, w_045_6367, w_045_6368, w_045_6370, w_045_6372, w_045_6373, w_045_6374, w_045_6378, w_045_6379, w_045_6380, w_045_6382, w_045_6383, w_045_6384, w_045_6386, w_045_6387, w_045_6388, w_045_6389, w_045_6392, w_045_6393, w_045_6397, w_045_6399, w_045_6401, w_045_6403, w_045_6409, w_045_6410, w_045_6411, w_045_6414, w_045_6415, w_045_6419, w_045_6420, w_045_6421, w_045_6422, w_045_6425, w_045_6428, w_045_6429, w_045_6432, w_045_6436, w_045_6438, w_045_6440, w_045_6441, w_045_6442, w_045_6443, w_045_6445, w_045_6449, w_045_6450, w_045_6452, w_045_6453, w_045_6454, w_045_6455, w_045_6462, w_045_6465, w_045_6466, w_045_6469, w_045_6472, w_045_6473, w_045_6474, w_045_6482, w_045_6485, w_045_6489, w_045_6490, w_045_6499, w_045_6502, w_045_6503, w_045_6505, w_045_6506, w_045_6508, w_045_6509, w_045_6510, w_045_6511, w_045_6513, w_045_6514, w_045_6516, w_045_6517, w_045_6518, w_045_6523, w_045_6526, w_045_6531, w_045_6532, w_045_6534, w_045_6535, w_045_6539, w_045_6540, w_045_6541, w_045_6546, w_045_6547, w_045_6549, w_045_6550, w_045_6551, w_045_6557, w_045_6559, w_045_6567, w_045_6571, w_045_6574, w_045_6582, w_045_6585, w_045_6587, w_045_6589, w_045_6590, w_045_6591, w_045_6596, w_045_6601, w_045_6603, w_045_6607, w_045_6610, w_045_6614, w_045_6616, w_045_6619, w_045_6621, w_045_6622, w_045_6623, w_045_6624, w_045_6628, w_045_6630, w_045_6631, w_045_6634, w_045_6635, w_045_6638, w_045_6640, w_045_6641, w_045_6642, w_045_6644, w_045_6645, w_045_6648, w_045_6650, w_045_6651, w_045_6652, w_045_6653, w_045_6655, w_045_6656, w_045_6657, w_045_6660, w_045_6661, w_045_6663, w_045_6664, w_045_6667, w_045_6668, w_045_6669, w_045_6670, w_045_6671, w_045_6672, w_045_6674, w_045_6675, w_045_6676, w_045_6678, w_045_6679, w_045_6683, w_045_6684, w_045_6686, w_045_6687, w_045_6690, w_045_6691, w_045_6694, w_045_6696, w_045_6700, w_045_6701, w_045_6703, w_045_6705, w_045_6711, w_045_6715, w_045_6716, w_045_6722, w_045_6724, w_045_6726, w_045_6728, w_045_6729, w_045_6730, w_045_6733, w_045_6738, w_045_6739, w_045_6740, w_045_6742, w_045_6752, w_045_6753, w_045_6759, w_045_6760, w_045_6761, w_045_6762, w_045_6763, w_045_6766, w_045_6768, w_045_6769, w_045_6770, w_045_6772, w_045_6774, w_045_6776, w_045_6777, w_045_6788, w_045_6789, w_045_6791, w_045_6797, w_045_6798, w_045_6799, w_045_6800, w_045_6801, w_045_6802, w_045_6805, w_045_6806, w_045_6807, w_045_6810, w_045_6814, w_045_6817, w_045_6821, w_045_6823, w_045_6824, w_045_6826, w_045_6827, w_045_6829, w_045_6830, w_045_6834, w_045_6836, w_045_6837, w_045_6838, w_045_6842, w_045_6843, w_045_6850, w_045_6853, w_045_6856, w_045_6861, w_045_6864, w_045_6868, w_045_6876, w_045_6879, w_045_6881, w_045_6884, w_045_6885, w_045_6886, w_045_6889, w_045_6894, w_045_6897, w_045_6899, w_045_6900, w_045_6901, w_045_6902, w_045_6903, w_045_6904, w_045_6906, w_045_6909, w_045_6912, w_045_6913, w_045_6914, w_045_6916, w_045_6917, w_045_6920, w_045_6922, w_045_6924, w_045_6929, w_045_6932, w_045_6934, w_045_6938, w_045_6939, w_045_6940, w_045_6941, w_045_6942, w_045_6946, w_045_6950, w_045_6954, w_045_6955, w_045_6956, w_045_6957, w_045_6958, w_045_6959, w_045_6960, w_045_6962, w_045_6963, w_045_6964, w_045_6965, w_045_6966, w_045_6969, w_045_6974, w_045_6975, w_045_6976, w_045_6977, w_045_6980, w_045_6989, w_045_6994, w_045_6997, w_045_6998, w_045_7004, w_045_7008, w_045_7012, w_045_7013, w_045_7014, w_045_7016, w_045_7017, w_045_7019, w_045_7020, w_045_7022, w_045_7024, w_045_7026, w_045_7028, w_045_7030, w_045_7032, w_045_7035, w_045_7036, w_045_7037, w_045_7038, w_045_7039, w_045_7041, w_045_7045, w_045_7046, w_045_7047, w_045_7051, w_045_7053, w_045_7059, w_045_7062, w_045_7065, w_045_7066, w_045_7069, w_045_7072, w_045_7073, w_045_7075, w_045_7077, w_045_7078, w_045_7081, w_045_7092, w_045_7093, w_045_7094, w_045_7096, w_045_7100, w_045_7101, w_045_7103, w_045_7105, w_045_7106, w_045_7107, w_045_7109, w_045_7111, w_045_7115, w_045_7116, w_045_7121, w_045_7123, w_045_7124, w_045_7126, w_045_7127, w_045_7128, w_045_7130, w_045_7131, w_045_7133, w_045_7137, w_045_7140, w_045_7141, w_045_7142, w_045_7149, w_045_7150, w_045_7152, w_045_7160, w_045_7161, w_045_7162, w_045_7165, w_045_7167, w_045_7169, w_045_7171, w_045_7172, w_045_7173, w_045_7174, w_045_7176, w_045_7180, w_045_7183, w_045_7184, w_045_7186, w_045_7188, w_045_7192, w_045_7196, w_045_7207, w_045_7210, w_045_7212, w_045_7215, w_045_7216, w_045_7218, w_045_7221, w_045_7222, w_045_7225, w_045_7227, w_045_7228, w_045_7230, w_045_7232, w_045_7233, w_045_7236, w_045_7237, w_045_7239, w_045_7241, w_045_7244, w_045_7246, w_045_7248, w_045_7251, w_045_7253, w_045_7255, w_045_7256, w_045_7260, w_045_7261, w_045_7264, w_045_7266, w_045_7267, w_045_7269, w_045_7271, w_045_7272, w_045_7274, w_045_7276, w_045_7277, w_045_7279, w_045_7280, w_045_7285, w_045_7286, w_045_7287, w_045_7289, w_045_7294, w_045_7300, w_045_7302, w_045_7304, w_045_7310, w_045_7313, w_045_7314, w_045_7316, w_045_7317, w_045_7318, w_045_7319, w_045_7320, w_045_7323, w_045_7324, w_045_7325, w_045_7329, w_045_7332, w_045_7333, w_045_7334, w_045_7337, w_045_7338, w_045_7340, w_045_7341, w_045_7342, w_045_7346, w_045_7347, w_045_7348, w_045_7352, w_045_7353, w_045_7355, w_045_7357, w_045_7359, w_045_7364, w_045_7365, w_045_7367, w_045_7368, w_045_7373, w_045_7374, w_045_7376, w_045_7377, w_045_7378, w_045_7382, w_045_7383, w_045_7384, w_045_7385, w_045_7386, w_045_7387, w_045_7391, w_045_7392, w_045_7395, w_045_7398, w_045_7400, w_045_7404, w_045_7406, w_045_7407, w_045_7408, w_045_7414, w_045_7418, w_045_7419, w_045_7420, w_045_7421, w_045_7422, w_045_7425, w_045_7426, w_045_7428, w_045_7430, w_045_7431, w_045_7432, w_045_7435, w_045_7436, w_045_7438, w_045_7439, w_045_7440, w_045_7442, w_045_7443, w_045_7445, w_045_7449, w_045_7450, w_045_7452, w_045_7453, w_045_7455, w_045_7456, w_045_7457, w_045_7458, w_045_7459, w_045_7460, w_045_7462, w_045_7465, w_045_7467, w_045_7470, w_045_7471, w_045_7472, w_045_7483, w_045_7484, w_045_7486, w_045_7492, w_045_7493, w_045_7501, w_045_7502, w_045_7504, w_045_7507, w_045_7508, w_045_7510, w_045_7513, w_045_7518, w_045_7522, w_045_7525, w_045_7526, w_045_7527, w_045_7530, w_045_7531, w_045_7533, w_045_7534, w_045_7535, w_045_7536, w_045_7538, w_045_7539, w_045_7540, w_045_7543, w_045_7550, w_045_7553, w_045_7556, w_045_7558, w_045_7560, w_045_7561, w_045_7563, w_045_7569, w_045_7575, w_045_7581, w_045_7582, w_045_7583, w_045_7584, w_045_7588, w_045_7589, w_045_7590, w_045_7594, w_045_7596, w_045_7597, w_045_7599, w_045_7604, w_045_7606, w_045_7609, w_045_7610, w_045_7611, w_045_7613, w_045_7614, w_045_7616, w_045_7619, w_045_7620, w_045_7623, w_045_7626, w_045_7627, w_045_7628, w_045_7632, w_045_7633, w_045_7635, w_045_7636, w_045_7638, w_045_7641, w_045_7642, w_045_7644, w_045_7647, w_045_7649, w_045_7651, w_045_7654, w_045_7657, w_045_7658, w_045_7659, w_045_7660, w_045_7662, w_045_7665, w_045_7671, w_045_7673, w_045_7676, w_045_7680, w_045_7681, w_045_7682, w_045_7684, w_045_7686, w_045_7690, w_045_7692, w_045_7693, w_045_7696, w_045_7697, w_045_7701, w_045_7703, w_045_7705, w_045_7711, w_045_7714, w_045_7715, w_045_7717, w_045_7719, w_045_7721, w_045_7722, w_045_7723, w_045_7725, w_045_7727, w_045_7728, w_045_7730, w_045_7732, w_045_7735, w_045_7738, w_045_7739, w_045_7741, w_045_7744, w_045_7745, w_045_7747, w_045_7748, w_045_7749, w_045_7750, w_045_7751, w_045_7752, w_045_7755, w_045_7756, w_045_7759, w_045_7760;
  wire w_046_001, w_046_002, w_046_003, w_046_004, w_046_005, w_046_006, w_046_007, w_046_008, w_046_009, w_046_010, w_046_011, w_046_012, w_046_013, w_046_015, w_046_016, w_046_017, w_046_018, w_046_020, w_046_024, w_046_025, w_046_027, w_046_028, w_046_029, w_046_032, w_046_033, w_046_035, w_046_036, w_046_037, w_046_038, w_046_039, w_046_040, w_046_041, w_046_042, w_046_043, w_046_044, w_046_045, w_046_046, w_046_047, w_046_050, w_046_051, w_046_052, w_046_053, w_046_054, w_046_055, w_046_056, w_046_057, w_046_058, w_046_060, w_046_062, w_046_063, w_046_064, w_046_065, w_046_066, w_046_068, w_046_070, w_046_071, w_046_073, w_046_076, w_046_077, w_046_079, w_046_080, w_046_081, w_046_082, w_046_083, w_046_084, w_046_085, w_046_087, w_046_088, w_046_089, w_046_090, w_046_091, w_046_092, w_046_093, w_046_094, w_046_096, w_046_098, w_046_099, w_046_100, w_046_101, w_046_102, w_046_103, w_046_104, w_046_106, w_046_107, w_046_108, w_046_109, w_046_110, w_046_111, w_046_112, w_046_113, w_046_115, w_046_116, w_046_117, w_046_118, w_046_119, w_046_120, w_046_121, w_046_122, w_046_123, w_046_125, w_046_126, w_046_127, w_046_129, w_046_130, w_046_131, w_046_132, w_046_135, w_046_136, w_046_137, w_046_138, w_046_139, w_046_140, w_046_141, w_046_143, w_046_144, w_046_145, w_046_146, w_046_147, w_046_148, w_046_149, w_046_150, w_046_151, w_046_152, w_046_154, w_046_156, w_046_157, w_046_158, w_046_159, w_046_160, w_046_161, w_046_162, w_046_163, w_046_164, w_046_165, w_046_166, w_046_168, w_046_169, w_046_170, w_046_171, w_046_172, w_046_173, w_046_174, w_046_175, w_046_176, w_046_178, w_046_179, w_046_180, w_046_181, w_046_182, w_046_184, w_046_185, w_046_186, w_046_187, w_046_188, w_046_189, w_046_191, w_046_192, w_046_194, w_046_195, w_046_196, w_046_197, w_046_198, w_046_199, w_046_200, w_046_201, w_046_202, w_046_203, w_046_204, w_046_205, w_046_206, w_046_207, w_046_208, w_046_209, w_046_210, w_046_211, w_046_212, w_046_214, w_046_215, w_046_217, w_046_219, w_046_222, w_046_223, w_046_224, w_046_225, w_046_226, w_046_227, w_046_229, w_046_230, w_046_231, w_046_232, w_046_234, w_046_237, w_046_238, w_046_239, w_046_240, w_046_241, w_046_243, w_046_244, w_046_245, w_046_246, w_046_247, w_046_248, w_046_250, w_046_251, w_046_252, w_046_253, w_046_254, w_046_255, w_046_256, w_046_258, w_046_259, w_046_260, w_046_261, w_046_262, w_046_264, w_046_266, w_046_267, w_046_268, w_046_269, w_046_272, w_046_275, w_046_276, w_046_278, w_046_279, w_046_280, w_046_281, w_046_282, w_046_283, w_046_284, w_046_285, w_046_286, w_046_288, w_046_289, w_046_290, w_046_291, w_046_292, w_046_293, w_046_295, w_046_296, w_046_298, w_046_299, w_046_301, w_046_302, w_046_303, w_046_304, w_046_305, w_046_306, w_046_307, w_046_308, w_046_309, w_046_310, w_046_311, w_046_312, w_046_314, w_046_315, w_046_317, w_046_318, w_046_319, w_046_320, w_046_321, w_046_322, w_046_323, w_046_324, w_046_325, w_046_326, w_046_327, w_046_329, w_046_330, w_046_331, w_046_332, w_046_333, w_046_334, w_046_336, w_046_337, w_046_338, w_046_339, w_046_340, w_046_341, w_046_342, w_046_343, w_046_344, w_046_345, w_046_346, w_046_347, w_046_348, w_046_349, w_046_350, w_046_351, w_046_352, w_046_353, w_046_355, w_046_356, w_046_358, w_046_359, w_046_362, w_046_363, w_046_364, w_046_365, w_046_366, w_046_367, w_046_369, w_046_372, w_046_373, w_046_374, w_046_375, w_046_376, w_046_377, w_046_378, w_046_380, w_046_383, w_046_384, w_046_385, w_046_386, w_046_387, w_046_388, w_046_389, w_046_390, w_046_391, w_046_392, w_046_394, w_046_395, w_046_396, w_046_397, w_046_398, w_046_399, w_046_402, w_046_403, w_046_404, w_046_405, w_046_407, w_046_408, w_046_410, w_046_413, w_046_414, w_046_415, w_046_416, w_046_417, w_046_418, w_046_419, w_046_420, w_046_421, w_046_422, w_046_423, w_046_424, w_046_426, w_046_427, w_046_429, w_046_430, w_046_432, w_046_433, w_046_434, w_046_435, w_046_436, w_046_437, w_046_438, w_046_440, w_046_441, w_046_442, w_046_443, w_046_444, w_046_445, w_046_446, w_046_447, w_046_448, w_046_449, w_046_450, w_046_451, w_046_452, w_046_453, w_046_454, w_046_455, w_046_456, w_046_457, w_046_458, w_046_459, w_046_461, w_046_462, w_046_463, w_046_464, w_046_465, w_046_466, w_046_467, w_046_468, w_046_470, w_046_471, w_046_472, w_046_473, w_046_474, w_046_475, w_046_477, w_046_478, w_046_479, w_046_480, w_046_481, w_046_482, w_046_483, w_046_486, w_046_487, w_046_488, w_046_490, w_046_491, w_046_493, w_046_494, w_046_495, w_046_496, w_046_497, w_046_498, w_046_499, w_046_500, w_046_501, w_046_502, w_046_503, w_046_504, w_046_505, w_046_506, w_046_507, w_046_508, w_046_509, w_046_510, w_046_512, w_046_514, w_046_515, w_046_516, w_046_517, w_046_518, w_046_520, w_046_521, w_046_522, w_046_523, w_046_525, w_046_527, w_046_528, w_046_529, w_046_530, w_046_531, w_046_532, w_046_534, w_046_537, w_046_538, w_046_539, w_046_540, w_046_541, w_046_542, w_046_543, w_046_544, w_046_545, w_046_546, w_046_548, w_046_549, w_046_550, w_046_551, w_046_552, w_046_553, w_046_554, w_046_556, w_046_559, w_046_560, w_046_562, w_046_563, w_046_564, w_046_566, w_046_567, w_046_568, w_046_569, w_046_571, w_046_572, w_046_576, w_046_577, w_046_578, w_046_579, w_046_580, w_046_581, w_046_582, w_046_583, w_046_584, w_046_585, w_046_587, w_046_588, w_046_589, w_046_590, w_046_591, w_046_593, w_046_594, w_046_595, w_046_596, w_046_599, w_046_602, w_046_604, w_046_605, w_046_606, w_046_607, w_046_608, w_046_609, w_046_610, w_046_611, w_046_612, w_046_613, w_046_614, w_046_615, w_046_616, w_046_618, w_046_619, w_046_621, w_046_622, w_046_623, w_046_624, w_046_625, w_046_626, w_046_628, w_046_630, w_046_631, w_046_632, w_046_633, w_046_635, w_046_636, w_046_638, w_046_639, w_046_641, w_046_642, w_046_643, w_046_644, w_046_646, w_046_647, w_046_648, w_046_649, w_046_652, w_046_653, w_046_654, w_046_655, w_046_656, w_046_657, w_046_658, w_046_659, w_046_660, w_046_662, w_046_663, w_046_664, w_046_665, w_046_666, w_046_667, w_046_669, w_046_672, w_046_673, w_046_674, w_046_675, w_046_676, w_046_677, w_046_679, w_046_680, w_046_682, w_046_684, w_046_685, w_046_686, w_046_687, w_046_688, w_046_689, w_046_690, w_046_693, w_046_697, w_046_700, w_046_701, w_046_702, w_046_703, w_046_704, w_046_706, w_046_708, w_046_709, w_046_710, w_046_712, w_046_713, w_046_714, w_046_715, w_046_716, w_046_718, w_046_719, w_046_722, w_046_723, w_046_724, w_046_727, w_046_729, w_046_730, w_046_733, w_046_735, w_046_736, w_046_737, w_046_739, w_046_740, w_046_741, w_046_742, w_046_743, w_046_744, w_046_745, w_046_746, w_046_747, w_046_749, w_046_751, w_046_752, w_046_753, w_046_754, w_046_755, w_046_758, w_046_759, w_046_760, w_046_762, w_046_763, w_046_765, w_046_766, w_046_767, w_046_768, w_046_771, w_046_772, w_046_773, w_046_774, w_046_775, w_046_776, w_046_777, w_046_780, w_046_781, w_046_782, w_046_784, w_046_786, w_046_787, w_046_788, w_046_789, w_046_791, w_046_792, w_046_796, w_046_797, w_046_800, w_046_801, w_046_804, w_046_805, w_046_806, w_046_807, w_046_809, w_046_810, w_046_812, w_046_813, w_046_814, w_046_816, w_046_817, w_046_818, w_046_819, w_046_820, w_046_822, w_046_823, w_046_826, w_046_828, w_046_830, w_046_831, w_046_832, w_046_833, w_046_834, w_046_835, w_046_836, w_046_837, w_046_838, w_046_842, w_046_845, w_046_846, w_046_847, w_046_849, w_046_850, w_046_851, w_046_852, w_046_853, w_046_854, w_046_855, w_046_856, w_046_858, w_046_859, w_046_860, w_046_862, w_046_864, w_046_869, w_046_870, w_046_871, w_046_872, w_046_874, w_046_875, w_046_876, w_046_879, w_046_880, w_046_881, w_046_882, w_046_883, w_046_884, w_046_886, w_046_887, w_046_888, w_046_889, w_046_890, w_046_891, w_046_894, w_046_895, w_046_896, w_046_900, w_046_902, w_046_904, w_046_905, w_046_907, w_046_908, w_046_909, w_046_911, w_046_912, w_046_913, w_046_915, w_046_916, w_046_917, w_046_918, w_046_919, w_046_921, w_046_922, w_046_924, w_046_929, w_046_930, w_046_931, w_046_932, w_046_933, w_046_934, w_046_935, w_046_938, w_046_939, w_046_944, w_046_945, w_046_947, w_046_949, w_046_950, w_046_951, w_046_953, w_046_955, w_046_956, w_046_957, w_046_958, w_046_961, w_046_962, w_046_964, w_046_965, w_046_967, w_046_968, w_046_969, w_046_970, w_046_972, w_046_973, w_046_974, w_046_975, w_046_977, w_046_979, w_046_981, w_046_983, w_046_985, w_046_986, w_046_991, w_046_993, w_046_994, w_046_996, w_046_997, w_046_999, w_046_1001, w_046_1002, w_046_1003, w_046_1004, w_046_1007, w_046_1008, w_046_1009, w_046_1011, w_046_1012, w_046_1014, w_046_1015, w_046_1017, w_046_1018, w_046_1020, w_046_1021, w_046_1022, w_046_1025, w_046_1026, w_046_1027, w_046_1028, w_046_1030, w_046_1031, w_046_1032, w_046_1033, w_046_1034, w_046_1038, w_046_1044, w_046_1045, w_046_1048, w_046_1050, w_046_1055, w_046_1056, w_046_1059, w_046_1060, w_046_1062, w_046_1063, w_046_1064, w_046_1065, w_046_1067, w_046_1068, w_046_1069, w_046_1070, w_046_1071, w_046_1072, w_046_1074, w_046_1075, w_046_1077, w_046_1078, w_046_1079, w_046_1080, w_046_1083, w_046_1085, w_046_1088, w_046_1089, w_046_1090, w_046_1091, w_046_1092, w_046_1094, w_046_1096, w_046_1097, w_046_1099, w_046_1100, w_046_1101, w_046_1102, w_046_1103, w_046_1104, w_046_1106, w_046_1108, w_046_1109, w_046_1111, w_046_1112, w_046_1113, w_046_1114, w_046_1115, w_046_1116, w_046_1118, w_046_1120, w_046_1123, w_046_1124, w_046_1125, w_046_1127, w_046_1132, w_046_1134, w_046_1136, w_046_1137, w_046_1138, w_046_1139, w_046_1141, w_046_1142, w_046_1144, w_046_1145, w_046_1146, w_046_1147, w_046_1148, w_046_1150, w_046_1151, w_046_1152, w_046_1153, w_046_1154, w_046_1155, w_046_1156, w_046_1158, w_046_1163, w_046_1164, w_046_1167, w_046_1172, w_046_1175, w_046_1176, w_046_1177, w_046_1179, w_046_1180, w_046_1181, w_046_1186, w_046_1187, w_046_1188, w_046_1189, w_046_1190, w_046_1191, w_046_1192, w_046_1193, w_046_1194, w_046_1196, w_046_1197, w_046_1198, w_046_1200, w_046_1202, w_046_1203, w_046_1204, w_046_1205, w_046_1207, w_046_1208, w_046_1210, w_046_1211, w_046_1212, w_046_1213, w_046_1217, w_046_1218, w_046_1220, w_046_1222, w_046_1223, w_046_1224, w_046_1225, w_046_1226, w_046_1227, w_046_1229, w_046_1230, w_046_1231, w_046_1232, w_046_1233, w_046_1234, w_046_1235, w_046_1236, w_046_1237, w_046_1239, w_046_1240, w_046_1242, w_046_1245, w_046_1246, w_046_1247, w_046_1250, w_046_1251, w_046_1252, w_046_1253, w_046_1254, w_046_1255, w_046_1258, w_046_1259, w_046_1260, w_046_1262, w_046_1264, w_046_1265, w_046_1266, w_046_1267, w_046_1268, w_046_1269, w_046_1271, w_046_1272, w_046_1273, w_046_1276, w_046_1279, w_046_1280, w_046_1282, w_046_1283, w_046_1285, w_046_1286, w_046_1291, w_046_1292, w_046_1294, w_046_1296, w_046_1297, w_046_1298, w_046_1299, w_046_1301, w_046_1303, w_046_1304, w_046_1305, w_046_1306, w_046_1309, w_046_1310, w_046_1311, w_046_1312, w_046_1313, w_046_1314, w_046_1317, w_046_1318, w_046_1319, w_046_1320, w_046_1321, w_046_1322, w_046_1323, w_046_1324, w_046_1325, w_046_1326, w_046_1327, w_046_1329, w_046_1331, w_046_1334, w_046_1335, w_046_1336, w_046_1338, w_046_1339, w_046_1341, w_046_1342, w_046_1343, w_046_1345, w_046_1346, w_046_1347, w_046_1349, w_046_1350, w_046_1351, w_046_1352, w_046_1353, w_046_1354, w_046_1356, w_046_1357, w_046_1359, w_046_1360, w_046_1362, w_046_1365, w_046_1366, w_046_1367, w_046_1368, w_046_1370, w_046_1371, w_046_1372, w_046_1373, w_046_1374, w_046_1375, w_046_1376, w_046_1377, w_046_1378, w_046_1383, w_046_1384, w_046_1385, w_046_1387, w_046_1389, w_046_1390, w_046_1391, w_046_1392, w_046_1393, w_046_1394, w_046_1395, w_046_1396, w_046_1397, w_046_1401, w_046_1402, w_046_1404, w_046_1406, w_046_1407, w_046_1408, w_046_1409, w_046_1410, w_046_1411, w_046_1412, w_046_1413, w_046_1414, w_046_1415, w_046_1416, w_046_1417, w_046_1420, w_046_1423, w_046_1425, w_046_1426, w_046_1428, w_046_1429, w_046_1432, w_046_1433, w_046_1434, w_046_1435, w_046_1436, w_046_1437, w_046_1438, w_046_1440, w_046_1441, w_046_1443, w_046_1447, w_046_1448, w_046_1449, w_046_1450, w_046_1451, w_046_1453, w_046_1455, w_046_1456, w_046_1457, w_046_1458, w_046_1459, w_046_1462, w_046_1463, w_046_1464, w_046_1465, w_046_1466, w_046_1468, w_046_1469, w_046_1470, w_046_1471, w_046_1473, w_046_1475, w_046_1476, w_046_1478, w_046_1479, w_046_1480, w_046_1481, w_046_1482, w_046_1483, w_046_1484, w_046_1485, w_046_1486, w_046_1487, w_046_1488, w_046_1489, w_046_1490, w_046_1491, w_046_1492, w_046_1493, w_046_1494, w_046_1495, w_046_1496, w_046_1497, w_046_1498, w_046_1499, w_046_1500, w_046_1502, w_046_1503, w_046_1505, w_046_1506, w_046_1507, w_046_1508, w_046_1509, w_046_1510, w_046_1512, w_046_1513, w_046_1514, w_046_1515, w_046_1516, w_046_1517, w_046_1520, w_046_1522, w_046_1523, w_046_1524, w_046_1525, w_046_1526, w_046_1527, w_046_1530, w_046_1531, w_046_1532, w_046_1534, w_046_1535, w_046_1536, w_046_1537, w_046_1541, w_046_1542, w_046_1544, w_046_1545, w_046_1546, w_046_1548, w_046_1550, w_046_1551, w_046_1553, w_046_1555, w_046_1556, w_046_1557, w_046_1558, w_046_1559, w_046_1560, w_046_1561, w_046_1565, w_046_1568, w_046_1569, w_046_1570, w_046_1571, w_046_1572, w_046_1574, w_046_1575, w_046_1577, w_046_1579, w_046_1581, w_046_1582, w_046_1585, w_046_1586, w_046_1587, w_046_1588, w_046_1589, w_046_1590, w_046_1593, w_046_1594, w_046_1596, w_046_1597, w_046_1602, w_046_1604, w_046_1605, w_046_1606, w_046_1607, w_046_1608, w_046_1609, w_046_1611, w_046_1612, w_046_1613, w_046_1614, w_046_1616, w_046_1618, w_046_1620, w_046_1621, w_046_1622, w_046_1624, w_046_1625, w_046_1626, w_046_1627, w_046_1628, w_046_1630, w_046_1631, w_046_1633, w_046_1634, w_046_1635, w_046_1636, w_046_1637, w_046_1638, w_046_1639, w_046_1642, w_046_1644, w_046_1645, w_046_1646, w_046_1648, w_046_1649, w_046_1650, w_046_1651, w_046_1652, w_046_1653, w_046_1656, w_046_1659, w_046_1661, w_046_1662, w_046_1663, w_046_1665, w_046_1666, w_046_1667, w_046_1672, w_046_1674, w_046_1675, w_046_1677, w_046_1678, w_046_1679, w_046_1680, w_046_1683, w_046_1685, w_046_1686, w_046_1687, w_046_1688, w_046_1689, w_046_1690, w_046_1691, w_046_1693, w_046_1694, w_046_1695, w_046_1696, w_046_1697, w_046_1699, w_046_1700, w_046_1701, w_046_1702, w_046_1704, w_046_1705, w_046_1710, w_046_1712, w_046_1713, w_046_1714, w_046_1715, w_046_1717, w_046_1718, w_046_1719, w_046_1720, w_046_1723, w_046_1724, w_046_1725, w_046_1726, w_046_1727, w_046_1728, w_046_1729, w_046_1730, w_046_1731, w_046_1732, w_046_1734, w_046_1735, w_046_1736, w_046_1738, w_046_1739, w_046_1740, w_046_1741, w_046_1743, w_046_1746, w_046_1749, w_046_1751, w_046_1752, w_046_1754, w_046_1755, w_046_1756, w_046_1758, w_046_1760, w_046_1761, w_046_1762, w_046_1764, w_046_1765, w_046_1766, w_046_1767, w_046_1770, w_046_1771, w_046_1772, w_046_1773, w_046_1775, w_046_1780, w_046_1781, w_046_1782, w_046_1783, w_046_1784, w_046_1786, w_046_1787, w_046_1788, w_046_1789, w_046_1792, w_046_1793, w_046_1794, w_046_1796, w_046_1797, w_046_1798, w_046_1799, w_046_1801, w_046_1802, w_046_1804, w_046_1806, w_046_1808, w_046_1809, w_046_1811, w_046_1812, w_046_1817, w_046_1818, w_046_1819, w_046_1821, w_046_1822, w_046_1823, w_046_1824, w_046_1825, w_046_1826, w_046_1827, w_046_1829, w_046_1830, w_046_1831, w_046_1832, w_046_1834, w_046_1835, w_046_1836, w_046_1837, w_046_1838, w_046_1839, w_046_1840, w_046_1844, w_046_1845, w_046_1846, w_046_1847, w_046_1848, w_046_1849, w_046_1850, w_046_1851, w_046_1852, w_046_1853, w_046_1854, w_046_1856, w_046_1857, w_046_1858, w_046_1862, w_046_1863, w_046_1865, w_046_1866, w_046_1869, w_046_1870, w_046_1871, w_046_1873, w_046_1874, w_046_1875, w_046_1876, w_046_1877, w_046_1878, w_046_1879, w_046_1880, w_046_1881, w_046_1882, w_046_1883, w_046_1884, w_046_1885, w_046_1888, w_046_1889, w_046_1890, w_046_1891, w_046_1892, w_046_1893, w_046_1895, w_046_1898, w_046_1899, w_046_1900, w_046_1902, w_046_1903, w_046_1904, w_046_1905, w_046_1906, w_046_1907, w_046_1908, w_046_1910, w_046_1911, w_046_1913, w_046_1914, w_046_1916, w_046_1917, w_046_1919, w_046_1920, w_046_1921, w_046_1922, w_046_1923, w_046_1925, w_046_1926, w_046_1927, w_046_1928, w_046_1929, w_046_1931, w_046_1937, w_046_1940, w_046_1941, w_046_1942, w_046_1943, w_046_1944, w_046_1946, w_046_1947, w_046_1948, w_046_1949, w_046_1951, w_046_1953, w_046_1954, w_046_1955, w_046_1957, w_046_1958, w_046_1960, w_046_1961, w_046_1962, w_046_1963, w_046_1964, w_046_1965, w_046_1967, w_046_1968, w_046_1969, w_046_1970, w_046_1971, w_046_1972, w_046_1973, w_046_1974, w_046_1977, w_046_1978, w_046_1979, w_046_1980, w_046_1981, w_046_1982, w_046_1984, w_046_1985, w_046_1988, w_046_1989, w_046_1991, w_046_1993, w_046_1995, w_046_1996, w_046_1997, w_046_1999, w_046_2000, w_046_2001, w_046_2002, w_046_2003, w_046_2004, w_046_2005, w_046_2006, w_046_2007, w_046_2008, w_046_2009, w_046_2010, w_046_2013, w_046_2014, w_046_2015, w_046_2016, w_046_2017, w_046_2018, w_046_2019, w_046_2021, w_046_2023, w_046_2025, w_046_2027, w_046_2028, w_046_2029, w_046_2030, w_046_2032, w_046_2033, w_046_2034, w_046_2035, w_046_2036, w_046_2038, w_046_2039, w_046_2042, w_046_2043, w_046_2044, w_046_2045, w_046_2048, w_046_2049, w_046_2050, w_046_2052, w_046_2054, w_046_2055, w_046_2056, w_046_2057, w_046_2058, w_046_2060, w_046_2062, w_046_2063, w_046_2064, w_046_2065, w_046_2066, w_046_2067, w_046_2069, w_046_2070, w_046_2071, w_046_2073, w_046_2075, w_046_2076, w_046_2077, w_046_2078, w_046_2079, w_046_2080, w_046_2081, w_046_2085, w_046_2086, w_046_2087, w_046_2088, w_046_2090, w_046_2091, w_046_2092, w_046_2093, w_046_2094, w_046_2097, w_046_2098, w_046_2099, w_046_2101, w_046_2103, w_046_2104, w_046_2105, w_046_2106, w_046_2107, w_046_2108, w_046_2112, w_046_2114, w_046_2115, w_046_2116, w_046_2117, w_046_2118, w_046_2119, w_046_2120, w_046_2123, w_046_2124, w_046_2126, w_046_2127, w_046_2128, w_046_2129, w_046_2130, w_046_2131, w_046_2133, w_046_2135, w_046_2136, w_046_2137, w_046_2138, w_046_2139, w_046_2144, w_046_2146, w_046_2147, w_046_2150, w_046_2151, w_046_2153, w_046_2154, w_046_2157, w_046_2158, w_046_2160, w_046_2161, w_046_2162, w_046_2165, w_046_2166, w_046_2169, w_046_2170, w_046_2171, w_046_2172, w_046_2173, w_046_2174, w_046_2175, w_046_2176, w_046_2178, w_046_2179, w_046_2180, w_046_2181, w_046_2182, w_046_2183, w_046_2184, w_046_2185, w_046_2186, w_046_2187, w_046_2188, w_046_2189, w_046_2191, w_046_2194, w_046_2197, w_046_2198, w_046_2202, w_046_2203, w_046_2204, w_046_2205, w_046_2206, w_046_2209, w_046_2210, w_046_2212, w_046_2213, w_046_2215, w_046_2216, w_046_2217, w_046_2218, w_046_2219, w_046_2220, w_046_2221, w_046_2222, w_046_2224, w_046_2225, w_046_2226, w_046_2229, w_046_2230, w_046_2233, w_046_2235, w_046_2237, w_046_2238, w_046_2239, w_046_2240, w_046_2241, w_046_2242, w_046_2243, w_046_2244, w_046_2246, w_046_2247, w_046_2248, w_046_2250, w_046_2252, w_046_2253, w_046_2254, w_046_2256, w_046_2257, w_046_2258, w_046_2260, w_046_2262, w_046_2263, w_046_2264, w_046_2265, w_046_2268, w_046_2269, w_046_2270, w_046_2271, w_046_2272, w_046_2273, w_046_2274, w_046_2275, w_046_2276, w_046_2278, w_046_2280, w_046_2281, w_046_2282, w_046_2284, w_046_2286, w_046_2288, w_046_2289, w_046_2290, w_046_2291, w_046_2292, w_046_2293, w_046_2294, w_046_2295, w_046_2296, w_046_2299, w_046_2300, w_046_2301, w_046_2302, w_046_2304, w_046_2305, w_046_2306, w_046_2310, w_046_2311, w_046_2312, w_046_2313, w_046_2314, w_046_2315, w_046_2316, w_046_2317, w_046_2318, w_046_2320, w_046_2321, w_046_2322, w_046_2323, w_046_2324, w_046_2326, w_046_2328, w_046_2329, w_046_2330, w_046_2331, w_046_2332, w_046_2337, w_046_2340, w_046_2341, w_046_2342, w_046_2343, w_046_2344, w_046_2345, w_046_2348, w_046_2349, w_046_2350, w_046_2351, w_046_2352, w_046_2354, w_046_2357, w_046_2358, w_046_2359, w_046_2360, w_046_2361, w_046_2362, w_046_2363, w_046_2365, w_046_2369, w_046_2370, w_046_2371, w_046_2372, w_046_2373, w_046_2375, w_046_2376, w_046_2378, w_046_2379, w_046_2380, w_046_2381, w_046_2383, w_046_2384, w_046_2386, w_046_2387, w_046_2389, w_046_2390, w_046_2391, w_046_2394, w_046_2395, w_046_2396, w_046_2398, w_046_2399, w_046_2405, w_046_2406, w_046_2407, w_046_2410, w_046_2411, w_046_2412, w_046_2413, w_046_2415, w_046_2417, w_046_2419, w_046_2420, w_046_2421, w_046_2423, w_046_2424, w_046_2425, w_046_2426, w_046_2428, w_046_2429, w_046_2430, w_046_2431, w_046_2432, w_046_2433, w_046_2435, w_046_2437, w_046_2438, w_046_2439, w_046_2440, w_046_2441, w_046_2442, w_046_2443, w_046_2445, w_046_2446, w_046_2447, w_046_2448, w_046_2449, w_046_2451, w_046_2452, w_046_2453, w_046_2455, w_046_2456, w_046_2457, w_046_2458, w_046_2459, w_046_2460, w_046_2463, w_046_2464, w_046_2465, w_046_2466, w_046_2468, w_046_2469, w_046_2471, w_046_2472, w_046_2474, w_046_2475, w_046_2477, w_046_2478, w_046_2481, w_046_2484, w_046_2485, w_046_2486, w_046_2487, w_046_2489, w_046_2491, w_046_2492, w_046_2493, w_046_2494, w_046_2495, w_046_2496, w_046_2498, w_046_2500, w_046_2502, w_046_2503, w_046_2504, w_046_2506, w_046_2507, w_046_2508, w_046_2509, w_046_2511, w_046_2513, w_046_2516, w_046_2519, w_046_2520, w_046_2521, w_046_2522, w_046_2524, w_046_2525, w_046_2526, w_046_2528, w_046_2532, w_046_2533, w_046_2535, w_046_2537, w_046_2539, w_046_2540, w_046_2541, w_046_2542, w_046_2545, w_046_2549, w_046_2550, w_046_2551, w_046_2553, w_046_2554, w_046_2555, w_046_2556, w_046_2558, w_046_2560, w_046_2562, w_046_2563, w_046_2565, w_046_2566, w_046_2569, w_046_2572, w_046_2574, w_046_2575, w_046_2576, w_046_2578, w_046_2579, w_046_2580, w_046_2582, w_046_2583, w_046_2585, w_046_2587, w_046_2588, w_046_2589, w_046_2590, w_046_2591, w_046_2594, w_046_2596, w_046_2597, w_046_2598, w_046_2601, w_046_2602, w_046_2606, w_046_2607, w_046_2609, w_046_2610, w_046_2613, w_046_2614, w_046_2615, w_046_2617, w_046_2618, w_046_2620, w_046_2621, w_046_2622, w_046_2626, w_046_2627, w_046_2630, w_046_2632, w_046_2633, w_046_2634, w_046_2635, w_046_2638, w_046_2640, w_046_2642, w_046_2643, w_046_2644, w_046_2645, w_046_2646, w_046_2647, w_046_2648, w_046_2652, w_046_2653, w_046_2655, w_046_2656, w_046_2657, w_046_2659, w_046_2660, w_046_2662, w_046_2665, w_046_2668, w_046_2669, w_046_2670, w_046_2671, w_046_2672, w_046_2674, w_046_2675, w_046_2676, w_046_2677, w_046_2680, w_046_2681, w_046_2685, w_046_2688, w_046_2689, w_046_2692, w_046_2693, w_046_2694, w_046_2696, w_046_2698, w_046_2699, w_046_2700, w_046_2701, w_046_2702, w_046_2704, w_046_2708, w_046_2712, w_046_2714, w_046_2715, w_046_2716, w_046_2717, w_046_2718, w_046_2719, w_046_2720, w_046_2721, w_046_2722, w_046_2726, w_046_2729, w_046_2731, w_046_2732, w_046_2733, w_046_2734, w_046_2735, w_046_2736, w_046_2737, w_046_2738, w_046_2739, w_046_2740, w_046_2742, w_046_2745, w_046_2746, w_046_2747, w_046_2749, w_046_2750, w_046_2751, w_046_2755, w_046_2756, w_046_2758, w_046_2760, w_046_2761, w_046_2763, w_046_2764, w_046_2765, w_046_2766, w_046_2767, w_046_2768, w_046_2769, w_046_2770, w_046_2772, w_046_2773, w_046_2780, w_046_2781, w_046_2782, w_046_2784, w_046_2785, w_046_2786, w_046_2787, w_046_2789, w_046_2790, w_046_2791, w_046_2792, w_046_2795, w_046_2796, w_046_2797, w_046_2799, w_046_2800, w_046_2802, w_046_2804, w_046_2806, w_046_2807, w_046_2808, w_046_2810, w_046_2813, w_046_2814, w_046_2815, w_046_2816, w_046_2817, w_046_2819, w_046_2821, w_046_2822, w_046_2823, w_046_2825, w_046_2828, w_046_2829, w_046_2831, w_046_2833, w_046_2835, w_046_2836, w_046_2837, w_046_2839, w_046_2840, w_046_2841, w_046_2842, w_046_2844, w_046_2845, w_046_2846, w_046_2848, w_046_2849, w_046_2850, w_046_2851, w_046_2855, w_046_2857, w_046_2860, w_046_2864, w_046_2865, w_046_2866, w_046_2867, w_046_2868, w_046_2870, w_046_2873, w_046_2874, w_046_2875, w_046_2878, w_046_2879, w_046_2880, w_046_2883, w_046_2884, w_046_2885, w_046_2886, w_046_2887, w_046_2888, w_046_2889, w_046_2890, w_046_2891, w_046_2892, w_046_2893, w_046_2894, w_046_2895, w_046_2897, w_046_2898, w_046_2900, w_046_2901, w_046_2902, w_046_2905, w_046_2907, w_046_2908, w_046_2910, w_046_2911, w_046_2912, w_046_2913, w_046_2915, w_046_2917, w_046_2918, w_046_2919, w_046_2920, w_046_2922, w_046_2923, w_046_2924, w_046_2926, w_046_2927, w_046_2928, w_046_2929, w_046_2930, w_046_2931, w_046_2932, w_046_2933, w_046_2934, w_046_2935, w_046_2936, w_046_2939, w_046_2944, w_046_2945, w_046_2946, w_046_2947, w_046_2948, w_046_2949, w_046_2950, w_046_2951, w_046_2953, w_046_2955, w_046_2956, w_046_2957, w_046_2958, w_046_2959, w_046_2960, w_046_2962, w_046_2966, w_046_2967, w_046_2969, w_046_2970, w_046_2971, w_046_2972, w_046_2973, w_046_2974, w_046_2975, w_046_2976, w_046_2977, w_046_2978, w_046_2979, w_046_2981, w_046_2982, w_046_2986, w_046_2987, w_046_2990, w_046_2992, w_046_2993, w_046_2994, w_046_2995, w_046_2997, w_046_2998, w_046_2999, w_046_3001, w_046_3002, w_046_3003, w_046_3004, w_046_3005, w_046_3006, w_046_3007, w_046_3009, w_046_3010, w_046_3011, w_046_3012, w_046_3013, w_046_3014, w_046_3016, w_046_3017, w_046_3018, w_046_3019, w_046_3020, w_046_3021, w_046_3022, w_046_3024, w_046_3025, w_046_3026, w_046_3027, w_046_3029, w_046_3030, w_046_3031, w_046_3032, w_046_3033, w_046_3036, w_046_3037, w_046_3038, w_046_3039, w_046_3041, w_046_3042, w_046_3043, w_046_3044, w_046_3045, w_046_3047, w_046_3049, w_046_3050, w_046_3051, w_046_3052, w_046_3053, w_046_3055, w_046_3057, w_046_3061, w_046_3063, w_046_3065, w_046_3066, w_046_3067, w_046_3068, w_046_3069, w_046_3070, w_046_3071, w_046_3072, w_046_3073, w_046_3074, w_046_3075, w_046_3077, w_046_3078, w_046_3079, w_046_3081, w_046_3082, w_046_3085, w_046_3086, w_046_3087, w_046_3088, w_046_3089, w_046_3092, w_046_3093, w_046_3097, w_046_3098, w_046_3099, w_046_3100, w_046_3103, w_046_3104, w_046_3105, w_046_3106, w_046_3108, w_046_3111, w_046_3112, w_046_3113, w_046_3114, w_046_3116, w_046_3117, w_046_3120, w_046_3121, w_046_3122, w_046_3123, w_046_3125, w_046_3128, w_046_3129, w_046_3130, w_046_3132, w_046_3133, w_046_3134, w_046_3136, w_046_3139, w_046_3140, w_046_3141, w_046_3142, w_046_3144, w_046_3146, w_046_3147, w_046_3149, w_046_3151, w_046_3156, w_046_3158, w_046_3159, w_046_3160, w_046_3161, w_046_3162, w_046_3163, w_046_3165, w_046_3166, w_046_3168, w_046_3169, w_046_3170, w_046_3172, w_046_3173, w_046_3174, w_046_3176, w_046_3178, w_046_3179, w_046_3180, w_046_3181, w_046_3182, w_046_3183, w_046_3184, w_046_3185, w_046_3186, w_046_3187, w_046_3189, w_046_3190, w_046_3191, w_046_3192, w_046_3193, w_046_3195, w_046_3196, w_046_3198, w_046_3199, w_046_3200, w_046_3201, w_046_3203, w_046_3204, w_046_3205, w_046_3208, w_046_3209, w_046_3212, w_046_3213, w_046_3214, w_046_3215, w_046_3216, w_046_3219, w_046_3220, w_046_3222, w_046_3223, w_046_3224, w_046_3225, w_046_3226, w_046_3228, w_046_3230, w_046_3233, w_046_3236, w_046_3238, w_046_3239, w_046_3241, w_046_3242, w_046_3243, w_046_3246, w_046_3247, w_046_3249, w_046_3250, w_046_3254, w_046_3255, w_046_3256, w_046_3257, w_046_3258, w_046_3259, w_046_3261, w_046_3262, w_046_3263, w_046_3267, w_046_3271, w_046_3272, w_046_3274, w_046_3275, w_046_3276, w_046_3277, w_046_3280, w_046_3281, w_046_3282, w_046_3283, w_046_3284, w_046_3285, w_046_3286, w_046_3287, w_046_3289, w_046_3290, w_046_3291, w_046_3293, w_046_3294, w_046_3295, w_046_3296, w_046_3297, w_046_3298, w_046_3300, w_046_3303, w_046_3304, w_046_3305, w_046_3306, w_046_3307, w_046_3308, w_046_3309, w_046_3310, w_046_3311, w_046_3312, w_046_3313, w_046_3314, w_046_3315, w_046_3316, w_046_3319, w_046_3321, w_046_3322, w_046_3324, w_046_3325, w_046_3326, w_046_3327, w_046_3329, w_046_3330, w_046_3331, w_046_3332, w_046_3333, w_046_3335, w_046_3336, w_046_3337, w_046_3338, w_046_3339, w_046_3342, w_046_3343, w_046_3344, w_046_3345, w_046_3347, w_046_3348, w_046_3349, w_046_3352, w_046_3353, w_046_3354, w_046_3357, w_046_3360, w_046_3362, w_046_3364, w_046_3365, w_046_3366, w_046_3368, w_046_3371, w_046_3372, w_046_3373, w_046_3374, w_046_3376, w_046_3377, w_046_3379, w_046_3380, w_046_3381, w_046_3382, w_046_3383, w_046_3384, w_046_3388, w_046_3389, w_046_3390, w_046_3391, w_046_3392, w_046_3394, w_046_3395, w_046_3396, w_046_3398, w_046_3400, w_046_3401, w_046_3402, w_046_3403, w_046_3404, w_046_3406, w_046_3408, w_046_3409, w_046_3410, w_046_3411, w_046_3412, w_046_3413, w_046_3414, w_046_3415, w_046_3416, w_046_3417, w_046_3418, w_046_3419, w_046_3420, w_046_3421, w_046_3423, w_046_3424, w_046_3425, w_046_3426, w_046_3427, w_046_3428, w_046_3430, w_046_3431, w_046_3432, w_046_3434, w_046_3437, w_046_3438, w_046_3439, w_046_3440, w_046_3441, w_046_3443, w_046_3444, w_046_3445, w_046_3446, w_046_3447, w_046_3448, w_046_3449, w_046_3450, w_046_3451, w_046_3452, w_046_3453, w_046_3454, w_046_3457, w_046_3459, w_046_3460, w_046_3461, w_046_3462, w_046_3463, w_046_3465, w_046_3466, w_046_3467, w_046_3468, w_046_3469, w_046_3470, w_046_3472, w_046_3474, w_046_3475, w_046_3476, w_046_3477, w_046_3478, w_046_3481, w_046_3482, w_046_3484, w_046_3485, w_046_3488, w_046_3490, w_046_3491, w_046_3493, w_046_3494, w_046_3495, w_046_3496, w_046_3498, w_046_3499, w_046_3500, w_046_3501, w_046_3502, w_046_3503, w_046_3504, w_046_3505, w_046_3506, w_046_3507, w_046_3509, w_046_3510, w_046_3511, w_046_3512, w_046_3513, w_046_3514, w_046_3519, w_046_3520, w_046_3521, w_046_3522, w_046_3525, w_046_3526, w_046_3528, w_046_3529, w_046_3531, w_046_3534, w_046_3535, w_046_3536, w_046_3538, w_046_3540, w_046_3543, w_046_3546, w_046_3547, w_046_3548, w_046_3551, w_046_3552, w_046_3553, w_046_3555, w_046_3556, w_046_3557, w_046_3558, w_046_3559, w_046_3560, w_046_3561, w_046_3562, w_046_3563, w_046_3564, w_046_3565, w_046_3567, w_046_3569, w_046_3571, w_046_3572, w_046_3573, w_046_3574, w_046_3575, w_046_3577, w_046_3580, w_046_3582, w_046_3584, w_046_3585, w_046_3586, w_046_3587, w_046_3588, w_046_3589, w_046_3590, w_046_3592, w_046_3594, w_046_3595, w_046_3596, w_046_3598, w_046_3599, w_046_3601, w_046_3602, w_046_3604, w_046_3605, w_046_3606, w_046_3607, w_046_3608, w_046_3609, w_046_3612, w_046_3613, w_046_3614, w_046_3615, w_046_3617, w_046_3620, w_046_3621, w_046_3622, w_046_3623, w_046_3625, w_046_3626, w_046_3628, w_046_3630, w_046_3631, w_046_3632, w_046_3634, w_046_3636, w_046_3637, w_046_3639, w_046_3640, w_046_3643, w_046_3645, w_046_3646, w_046_3648, w_046_3650, w_046_3651, w_046_3652, w_046_3653, w_046_3655, w_046_3657, w_046_3659, w_046_3660, w_046_3661, w_046_3663, w_046_3664, w_046_3665, w_046_3666, w_046_3667, w_046_3671, w_046_3673, w_046_3674, w_046_3675, w_046_3677, w_046_3678, w_046_3679, w_046_3681, w_046_3682, w_046_3683, w_046_3684, w_046_3685, w_046_3686, w_046_3687, w_046_3688, w_046_3689, w_046_3690, w_046_3691, w_046_3693, w_046_3694, w_046_3697, w_046_3698, w_046_3699, w_046_3700, w_046_3701, w_046_3702, w_046_3703, w_046_3704, w_046_3705, w_046_3706, w_046_3708, w_046_3710, w_046_3711, w_046_3712, w_046_3713, w_046_3715, w_046_3716, w_046_3717, w_046_3720, w_046_3723, w_046_3724, w_046_3726, w_046_3727, w_046_3728, w_046_3729, w_046_3731, w_046_3734, w_046_3737, w_046_3738, w_046_3739, w_046_3741, w_046_3742, w_046_3744, w_046_3745, w_046_3747, w_046_3748, w_046_3750, w_046_3754, w_046_3755, w_046_3756, w_046_3757, w_046_3758, w_046_3759, w_046_3760, w_046_3761, w_046_3763, w_046_3764, w_046_3765, w_046_3766, w_046_3767, w_046_3768, w_046_3769, w_046_3770, w_046_3772, w_046_3773, w_046_3774, w_046_3775, w_046_3779, w_046_3780, w_046_3781, w_046_3782, w_046_3783, w_046_3784, w_046_3785, w_046_3786, w_046_3788, w_046_3789, w_046_3790, w_046_3791, w_046_3792, w_046_3793, w_046_3795, w_046_3796, w_046_3797, w_046_3798, w_046_3801, w_046_3802, w_046_3808, w_046_3809, w_046_3811, w_046_3813, w_046_3814, w_046_3816, w_046_3817, w_046_3818, w_046_3819, w_046_3820, w_046_3822, w_046_3823, w_046_3824, w_046_3826, w_046_3827, w_046_3828, w_046_3829, w_046_3830, w_046_3832, w_046_3833, w_046_3835, w_046_3838, w_046_3839, w_046_3840, w_046_3841, w_046_3842, w_046_3843, w_046_3844, w_046_3846, w_046_3849, w_046_3851, w_046_3852, w_046_3854, w_046_3855, w_046_3857, w_046_3858, w_046_3860, w_046_3861, w_046_3864, w_046_3865, w_046_3866, w_046_3867, w_046_3868, w_046_3869, w_046_3870, w_046_3871, w_046_3872, w_046_3874, w_046_3878, w_046_3879, w_046_3880, w_046_3881, w_046_3882, w_046_3883, w_046_3884, w_046_3885, w_046_3887, w_046_3888, w_046_3889, w_046_3890, w_046_3891, w_046_3892, w_046_3893, w_046_3894, w_046_3895, w_046_3896, w_046_3897, w_046_3898, w_046_3899, w_046_3901, w_046_3902, w_046_3903, w_046_3904, w_046_3905, w_046_3906, w_046_3908, w_046_3909, w_046_3911, w_046_3913, w_046_3915, w_046_3916, w_046_3918, w_046_3919, w_046_3920, w_046_3924, w_046_3927, w_046_3928, w_046_3929, w_046_3930, w_046_3931, w_046_3932, w_046_3933, w_046_3934, w_046_3935, w_046_3938, w_046_3939, w_046_3940, w_046_3941, w_046_3943, w_046_3946, w_046_3947, w_046_3948, w_046_3950, w_046_3951, w_046_3953, w_046_3955, w_046_3956, w_046_3958, w_046_3960, w_046_3961, w_046_3962, w_046_3965, w_046_3966, w_046_3968, w_046_3972, w_046_3973, w_046_3974, w_046_3976, w_046_3982, w_046_3983, w_046_3984, w_046_3985, w_046_3986, w_046_3987, w_046_3988, w_046_3990, w_046_3991, w_046_3992, w_046_3994, w_046_3995, w_046_3996, w_046_3997, w_046_3999, w_046_4000, w_046_4002, w_046_4004, w_046_4005, w_046_4006, w_046_4007, w_046_4008, w_046_4009, w_046_4010, w_046_4011, w_046_4012, w_046_4013, w_046_4014, w_046_4015, w_046_4017, w_046_4019, w_046_4020, w_046_4021, w_046_4024, w_046_4025, w_046_4027, w_046_4030, w_046_4031, w_046_4032, w_046_4034, w_046_4035, w_046_4036, w_046_4037, w_046_4038, w_046_4040, w_046_4042, w_046_4044, w_046_4045, w_046_4047, w_046_4049, w_046_4050, w_046_4053, w_046_4054, w_046_4056, w_046_4059, w_046_4060, w_046_4061, w_046_4063, w_046_4065, w_046_4066, w_046_4068, w_046_4069, w_046_4072, w_046_4074, w_046_4075, w_046_4077, w_046_4079, w_046_4080, w_046_4081, w_046_4082, w_046_4084, w_046_4086, w_046_4088, w_046_4090, w_046_4091, w_046_4092, w_046_4093, w_046_4094, w_046_4095, w_046_4096, w_046_4099, w_046_4100, w_046_4101, w_046_4104, w_046_4105, w_046_4106, w_046_4108, w_046_4109, w_046_4110, w_046_4111, w_046_4112, w_046_4113, w_046_4114, w_046_4115, w_046_4120, w_046_4121, w_046_4122, w_046_4123, w_046_4124, w_046_4125, w_046_4128, w_046_4132, w_046_4133, w_046_4134, w_046_4137, w_046_4140, w_046_4142, w_046_4143, w_046_4144, w_046_4145, w_046_4147, w_046_4148, w_046_4149, w_046_4151, w_046_4154, w_046_4155, w_046_4156, w_046_4157, w_046_4161, w_046_4162, w_046_4163, w_046_4166, w_046_4168, w_046_4169, w_046_4170, w_046_4171, w_046_4172, w_046_4174, w_046_4175, w_046_4176, w_046_4177, w_046_4178, w_046_4179, w_046_4180, w_046_4183, w_046_4184, w_046_4185, w_046_4186, w_046_4187, w_046_4188, w_046_4189, w_046_4190, w_046_4191, w_046_4193, w_046_4196, w_046_4198, w_046_4199, w_046_4200, w_046_4201, w_046_4202, w_046_4203, w_046_4204, w_046_4206, w_046_4207, w_046_4208, w_046_4209, w_046_4210, w_046_4211, w_046_4212, w_046_4213, w_046_4217, w_046_4220, w_046_4221, w_046_4224, w_046_4225, w_046_4226, w_046_4227, w_046_4228, w_046_4229, w_046_4230, w_046_4234, w_046_4237, w_046_4240, w_046_4242, w_046_4243, w_046_4245, w_046_4246, w_046_4247, w_046_4248, w_046_4250, w_046_4251, w_046_4252, w_046_4254, w_046_4255, w_046_4257, w_046_4260, w_046_4261, w_046_4262, w_046_4263, w_046_4264, w_046_4265, w_046_4267, w_046_4268, w_046_4271, w_046_4272, w_046_4273, w_046_4274, w_046_4276, w_046_4277, w_046_4279, w_046_4280, w_046_4283, w_046_4285, w_046_4286, w_046_4288, w_046_4289, w_046_4290, w_046_4291, w_046_4292, w_046_4293, w_046_4295, w_046_4297, w_046_4300, w_046_4301, w_046_4302, w_046_4303, w_046_4307, w_046_4308, w_046_4309, w_046_4310, w_046_4311, w_046_4313, w_046_4315, w_046_4316, w_046_4317, w_046_4319, w_046_4321, w_046_4323, w_046_4324, w_046_4326, w_046_4327, w_046_4329, w_046_4330, w_046_4331, w_046_4333, w_046_4334, w_046_4335, w_046_4336, w_046_4337, w_046_4338, w_046_4340, w_046_4341, w_046_4343, w_046_4344, w_046_4345, w_046_4346, w_046_4347, w_046_4348, w_046_4349, w_046_4350, w_046_4351, w_046_4353, w_046_4354, w_046_4356, w_046_4357, w_046_4358, w_046_4360, w_046_4361, w_046_4362, w_046_4368, w_046_4369, w_046_4370, w_046_4371, w_046_4374, w_046_4375, w_046_4377, w_046_4378, w_046_4379, w_046_4380, w_046_4381, w_046_4385, w_046_4386, w_046_4387, w_046_4390, w_046_4391, w_046_4392, w_046_4393, w_046_4395, w_046_4396, w_046_4397, w_046_4399, w_046_4401, w_046_4402, w_046_4403, w_046_4404, w_046_4406, w_046_4407, w_046_4408, w_046_4410, w_046_4411, w_046_4413, w_046_4414, w_046_4416, w_046_4417, w_046_4418, w_046_4419, w_046_4420, w_046_4422, w_046_4423, w_046_4425, w_046_4427, w_046_4428, w_046_4429, w_046_4433, w_046_4434, w_046_4439, w_046_4440, w_046_4442, w_046_4443, w_046_4444, w_046_4445, w_046_4446, w_046_4447, w_046_4448, w_046_4449, w_046_4450, w_046_4452, w_046_4453, w_046_4454, w_046_4455, w_046_4456, w_046_4457, w_046_4462, w_046_4465, w_046_4466, w_046_4467, w_046_4469, w_046_4470, w_046_4471, w_046_4473, w_046_4474, w_046_4475, w_046_4476, w_046_4477, w_046_4478, w_046_4479, w_046_4481, w_046_4482, w_046_4483, w_046_4486, w_046_4487, w_046_4488, w_046_4489, w_046_4490, w_046_4491, w_046_4492, w_046_4494, w_046_4495, w_046_4499, w_046_4500, w_046_4501, w_046_4502, w_046_4503, w_046_4504, w_046_4505, w_046_4506, w_046_4510, w_046_4511, w_046_4512, w_046_4513, w_046_4514, w_046_4515, w_046_4516, w_046_4518, w_046_4520, w_046_4521, w_046_4523, w_046_4524, w_046_4525, w_046_4526, w_046_4527, w_046_4528, w_046_4532, w_046_4534, w_046_4535, w_046_4536, w_046_4537, w_046_4538, w_046_4539, w_046_4540, w_046_4541, w_046_4542, w_046_4543, w_046_4547, w_046_4548, w_046_4550, w_046_4551, w_046_4552, w_046_4554, w_046_4555, w_046_4556, w_046_4557, w_046_4558, w_046_4560, w_046_4561, w_046_4562, w_046_4563, w_046_4564, w_046_4566, w_046_4568, w_046_4571, w_046_4573, w_046_4575, w_046_4576, w_046_4578, w_046_4579, w_046_4581, w_046_4583, w_046_4584, w_046_4586, w_046_4588, w_046_4589, w_046_4590, w_046_4591, w_046_4592, w_046_4594, w_046_4595, w_046_4598, w_046_4599, w_046_4602, w_046_4604, w_046_4605, w_046_4606, w_046_4609, w_046_4610, w_046_4611, w_046_4612, w_046_4614, w_046_4615, w_046_4617, w_046_4618, w_046_4620, w_046_4623, w_046_4624, w_046_4625, w_046_4626, w_046_4628, w_046_4629, w_046_4630, w_046_4631, w_046_4632, w_046_4635, w_046_4636, w_046_4639, w_046_4640, w_046_4642, w_046_4643, w_046_4645, w_046_4647, w_046_4651, w_046_4652, w_046_4653, w_046_4654, w_046_4655, w_046_4657, w_046_4658, w_046_4660, w_046_4661, w_046_4663, w_046_4665, w_046_4666, w_046_4667, w_046_4668, w_046_4669, w_046_4670, w_046_4674, w_046_4675, w_046_4678, w_046_4679, w_046_4680, w_046_4681, w_046_4684, w_046_4685;
  wire w_047_000, w_047_001, w_047_002, w_047_003, w_047_004, w_047_005, w_047_006, w_047_009, w_047_010, w_047_013, w_047_014, w_047_015, w_047_016, w_047_017, w_047_019, w_047_020, w_047_022, w_047_023, w_047_024, w_047_025, w_047_026, w_047_027, w_047_028, w_047_029, w_047_030, w_047_031, w_047_032, w_047_034, w_047_035, w_047_036, w_047_037, w_047_038, w_047_039, w_047_040, w_047_041, w_047_042, w_047_043, w_047_044, w_047_045, w_047_046, w_047_047, w_047_048, w_047_049, w_047_050, w_047_051, w_047_053, w_047_054, w_047_056, w_047_057, w_047_058, w_047_059, w_047_060, w_047_061, w_047_062, w_047_063, w_047_064, w_047_065, w_047_066, w_047_068, w_047_069, w_047_070, w_047_072, w_047_074, w_047_075, w_047_076, w_047_077, w_047_078, w_047_079, w_047_080, w_047_081, w_047_082, w_047_083, w_047_084, w_047_085, w_047_086, w_047_087, w_047_088, w_047_089, w_047_090, w_047_091, w_047_092, w_047_093, w_047_094, w_047_096, w_047_097, w_047_098, w_047_100, w_047_101, w_047_102, w_047_103, w_047_104, w_047_105, w_047_106, w_047_107, w_047_108, w_047_109, w_047_111, w_047_112, w_047_115, w_047_116, w_047_117, w_047_118, w_047_119, w_047_120, w_047_121, w_047_122, w_047_123, w_047_124, w_047_125, w_047_126, w_047_127, w_047_129, w_047_132, w_047_133, w_047_134, w_047_135, w_047_136, w_047_137, w_047_138, w_047_140, w_047_141, w_047_142, w_047_143, w_047_144, w_047_145, w_047_146, w_047_147, w_047_148, w_047_149, w_047_150, w_047_151, w_047_152, w_047_154, w_047_155, w_047_156, w_047_157, w_047_158, w_047_159, w_047_160, w_047_162, w_047_163, w_047_165, w_047_166, w_047_167, w_047_168, w_047_169, w_047_170, w_047_171, w_047_172, w_047_173, w_047_174, w_047_175, w_047_176, w_047_177, w_047_178, w_047_179, w_047_180, w_047_181, w_047_182, w_047_183, w_047_184, w_047_185, w_047_186, w_047_187, w_047_188, w_047_189, w_047_192, w_047_194, w_047_195, w_047_196, w_047_197, w_047_198, w_047_199, w_047_200, w_047_202, w_047_203, w_047_204, w_047_206, w_047_207, w_047_208, w_047_209, w_047_210, w_047_211, w_047_212, w_047_213, w_047_214, w_047_215, w_047_216, w_047_217, w_047_218, w_047_219, w_047_220, w_047_222, w_047_224, w_047_225, w_047_226, w_047_227, w_047_228, w_047_229, w_047_230, w_047_231, w_047_232, w_047_233, w_047_235, w_047_236, w_047_237, w_047_238, w_047_239, w_047_240, w_047_241, w_047_242, w_047_243, w_047_244, w_047_245, w_047_247, w_047_248, w_047_249, w_047_250, w_047_251, w_047_253, w_047_254, w_047_255, w_047_256, w_047_257, w_047_258, w_047_259, w_047_260, w_047_262, w_047_263, w_047_265, w_047_266, w_047_267, w_047_268, w_047_269, w_047_271, w_047_272, w_047_273, w_047_274, w_047_275, w_047_277, w_047_278, w_047_279, w_047_280, w_047_281, w_047_282, w_047_283, w_047_284, w_047_285, w_047_286, w_047_287, w_047_288, w_047_289, w_047_290, w_047_291, w_047_292, w_047_293, w_047_294, w_047_295, w_047_296, w_047_298, w_047_299, w_047_300, w_047_301, w_047_302, w_047_303, w_047_304, w_047_306, w_047_307, w_047_308, w_047_309, w_047_310, w_047_312, w_047_313, w_047_314, w_047_315, w_047_316, w_047_317, w_047_318, w_047_319, w_047_320, w_047_321, w_047_322, w_047_323, w_047_324, w_047_325, w_047_326, w_047_327, w_047_328, w_047_330, w_047_331, w_047_333, w_047_335, w_047_337, w_047_338, w_047_339, w_047_340, w_047_341, w_047_342, w_047_343, w_047_344, w_047_345, w_047_346, w_047_348, w_047_350, w_047_351, w_047_352, w_047_353, w_047_354, w_047_355, w_047_356, w_047_357, w_047_358, w_047_359, w_047_360, w_047_361, w_047_362, w_047_363, w_047_364, w_047_365, w_047_366, w_047_367, w_047_368, w_047_371, w_047_372, w_047_374, w_047_375, w_047_377, w_047_378, w_047_379, w_047_380, w_047_381, w_047_382, w_047_383, w_047_384, w_047_385, w_047_386, w_047_388, w_047_389, w_047_390, w_047_393, w_047_394, w_047_395, w_047_397, w_047_398, w_047_401, w_047_402, w_047_403, w_047_404, w_047_405, w_047_408, w_047_409, w_047_410, w_047_411, w_047_414, w_047_415, w_047_416, w_047_417, w_047_418, w_047_419, w_047_421, w_047_422, w_047_423, w_047_424, w_047_425, w_047_427, w_047_429, w_047_430, w_047_431, w_047_432, w_047_433, w_047_434, w_047_435, w_047_436, w_047_437, w_047_438, w_047_439, w_047_441, w_047_442, w_047_443, w_047_444, w_047_445, w_047_446, w_047_447, w_047_448, w_047_450, w_047_451, w_047_453, w_047_454, w_047_456, w_047_457, w_047_458, w_047_459, w_047_461, w_047_462, w_047_464, w_047_465, w_047_466, w_047_467, w_047_468, w_047_469, w_047_470, w_047_471, w_047_472, w_047_473, w_047_474, w_047_475, w_047_477, w_047_478, w_047_480, w_047_482, w_047_483, w_047_484, w_047_485, w_047_486, w_047_487, w_047_489, w_047_490, w_047_492, w_047_493, w_047_495, w_047_496, w_047_497, w_047_498, w_047_499, w_047_500, w_047_501, w_047_502, w_047_503, w_047_504, w_047_505, w_047_507, w_047_508, w_047_509, w_047_510, w_047_511, w_047_512, w_047_513, w_047_514, w_047_515, w_047_516, w_047_518, w_047_519, w_047_520, w_047_521, w_047_522, w_047_523, w_047_524, w_047_525, w_047_526, w_047_527, w_047_528, w_047_529, w_047_530, w_047_531, w_047_532, w_047_536, w_047_537, w_047_539, w_047_540, w_047_541, w_047_542, w_047_545, w_047_546, w_047_547, w_047_548, w_047_549, w_047_550, w_047_551, w_047_552, w_047_553, w_047_554, w_047_555, w_047_556, w_047_557, w_047_559, w_047_560, w_047_561, w_047_562, w_047_563, w_047_565, w_047_566, w_047_567, w_047_568, w_047_569, w_047_571, w_047_573, w_047_574, w_047_575, w_047_577, w_047_578, w_047_579, w_047_580, w_047_581, w_047_582, w_047_584, w_047_585, w_047_586, w_047_587, w_047_588, w_047_590, w_047_591, w_047_592, w_047_593, w_047_594, w_047_595, w_047_597, w_047_598, w_047_599, w_047_601, w_047_603, w_047_604, w_047_605, w_047_607, w_047_608, w_047_609, w_047_611, w_047_612, w_047_613, w_047_614, w_047_615, w_047_617, w_047_619, w_047_621, w_047_622, w_047_623, w_047_624, w_047_625, w_047_626, w_047_627, w_047_628, w_047_629, w_047_630, w_047_631, w_047_632, w_047_633, w_047_634, w_047_635, w_047_636, w_047_637, w_047_640, w_047_641, w_047_642, w_047_643, w_047_644, w_047_645, w_047_646, w_047_647, w_047_649, w_047_650, w_047_652, w_047_653, w_047_654, w_047_655, w_047_656, w_047_657, w_047_658, w_047_659, w_047_660, w_047_661, w_047_662, w_047_663, w_047_664, w_047_668, w_047_669, w_047_670, w_047_671, w_047_672, w_047_675, w_047_676, w_047_677, w_047_678, w_047_679, w_047_680, w_047_681, w_047_682, w_047_684, w_047_685, w_047_687, w_047_688, w_047_689, w_047_690, w_047_693, w_047_694, w_047_695, w_047_696, w_047_697, w_047_699, w_047_700, w_047_702, w_047_703, w_047_705, w_047_706, w_047_707, w_047_708, w_047_709, w_047_710, w_047_712, w_047_713, w_047_714, w_047_715, w_047_717, w_047_718, w_047_719, w_047_720, w_047_721, w_047_725, w_047_726, w_047_727, w_047_728, w_047_729, w_047_730, w_047_731, w_047_732, w_047_733, w_047_734, w_047_735, w_047_736, w_047_737, w_047_738, w_047_739, w_047_740, w_047_741, w_047_742, w_047_743, w_047_744, w_047_745, w_047_746, w_047_747, w_047_748, w_047_749, w_047_750, w_047_751, w_047_752, w_047_753, w_047_754, w_047_755, w_047_756, w_047_757, w_047_758, w_047_759, w_047_760, w_047_762, w_047_763, w_047_764, w_047_765, w_047_767, w_047_769, w_047_771, w_047_772, w_047_773, w_047_774, w_047_775, w_047_776, w_047_777, w_047_778, w_047_779, w_047_780, w_047_781, w_047_782, w_047_783, w_047_784, w_047_785, w_047_786, w_047_787, w_047_790, w_047_791, w_047_792, w_047_793, w_047_794, w_047_795, w_047_796, w_047_797, w_047_798, w_047_800, w_047_801, w_047_803, w_047_804, w_047_805, w_047_807, w_047_808, w_047_809, w_047_810, w_047_811, w_047_812, w_047_815, w_047_816, w_047_817, w_047_818, w_047_819, w_047_820, w_047_821, w_047_822, w_047_823, w_047_824, w_047_825, w_047_826, w_047_827, w_047_828, w_047_829, w_047_830, w_047_831, w_047_832, w_047_834, w_047_835, w_047_836, w_047_837, w_047_838, w_047_839, w_047_840, w_047_841, w_047_843, w_047_844, w_047_845, w_047_846, w_047_847, w_047_849, w_047_852, w_047_853, w_047_854, w_047_855, w_047_856, w_047_857, w_047_859, w_047_860, w_047_861, w_047_862, w_047_864, w_047_865, w_047_866, w_047_867, w_047_868, w_047_869, w_047_870, w_047_871, w_047_872, w_047_874, w_047_875, w_047_876, w_047_877, w_047_878, w_047_879, w_047_881, w_047_882, w_047_883, w_047_884, w_047_885, w_047_886, w_047_887, w_047_888, w_047_889, w_047_890, w_047_892, w_047_893, w_047_894, w_047_895, w_047_896, w_047_899, w_047_900, w_047_901, w_047_903, w_047_905, w_047_907, w_047_908, w_047_909, w_047_910, w_047_911, w_047_912, w_047_913, w_047_914, w_047_915, w_047_916, w_047_918, w_047_919, w_047_923, w_047_924, w_047_926, w_047_927, w_047_928, w_047_930, w_047_931, w_047_932, w_047_933, w_047_934, w_047_935, w_047_936, w_047_937, w_047_938, w_047_940, w_047_941, w_047_942, w_047_943, w_047_944, w_047_946, w_047_948, w_047_949, w_047_950, w_047_951, w_047_952, w_047_954, w_047_955, w_047_956, w_047_958, w_047_960, w_047_961, w_047_962, w_047_963, w_047_964, w_047_965, w_047_967, w_047_968, w_047_969, w_047_970, w_047_971, w_047_972, w_047_973, w_047_974, w_047_975, w_047_976, w_047_980, w_047_981, w_047_982, w_047_984, w_047_985, w_047_986, w_047_988, w_047_989, w_047_990, w_047_991, w_047_993, w_047_995, w_047_996, w_047_997, w_047_998, w_047_999, w_047_1000, w_047_1001, w_047_1003, w_047_1004, w_047_1006, w_047_1007, w_047_1008, w_047_1009, w_047_1010, w_047_1012, w_047_1014, w_047_1015, w_047_1016, w_047_1017, w_047_1018, w_047_1020, w_047_1022, w_047_1023, w_047_1024, w_047_1027, w_047_1028, w_047_1029, w_047_1030, w_047_1032, w_047_1034, w_047_1035, w_047_1037, w_047_1038, w_047_1039, w_047_1040, w_047_1041, w_047_1042, w_047_1043, w_047_1044, w_047_1045, w_047_1046, w_047_1048, w_047_1049, w_047_1050, w_047_1051, w_047_1052, w_047_1053, w_047_1054, w_047_1055, w_047_1056, w_047_1057, w_047_1058, w_047_1059, w_047_1060, w_047_1061, w_047_1062, w_047_1063, w_047_1065, w_047_1066, w_047_1067, w_047_1068, w_047_1069, w_047_1070, w_047_1071, w_047_1072, w_047_1073, w_047_1074, w_047_1075, w_047_1076, w_047_1077, w_047_1078, w_047_1079, w_047_1080, w_047_1081, w_047_1082, w_047_1083, w_047_1085, w_047_1086, w_047_1087, w_047_1089, w_047_1090, w_047_1091, w_047_1092, w_047_1093, w_047_1094, w_047_1095, w_047_1096, w_047_1097, w_047_1098, w_047_1099, w_047_1101, w_047_1103, w_047_1104, w_047_1105, w_047_1106, w_047_1108, w_047_1109, w_047_1110, w_047_1111, w_047_1112, w_047_1113, w_047_1114, w_047_1115, w_047_1116, w_047_1117, w_047_1118, w_047_1119, w_047_1120, w_047_1122, w_047_1123, w_047_1124, w_047_1125, w_047_1127, w_047_1128, w_047_1130, w_047_1131, w_047_1132, w_047_1133, w_047_1134, w_047_1135, w_047_1136, w_047_1138, w_047_1140, w_047_1141, w_047_1143, w_047_1144, w_047_1145, w_047_1146, w_047_1150, w_047_1151, w_047_1152, w_047_1153, w_047_1154, w_047_1155, w_047_1156, w_047_1158, w_047_1159, w_047_1160, w_047_1161, w_047_1162, w_047_1163, w_047_1165, w_047_1166, w_047_1167, w_047_1169, w_047_1170, w_047_1171, w_047_1172, w_047_1173, w_047_1175, w_047_1176, w_047_1179, w_047_1181, w_047_1182, w_047_1183, w_047_1184, w_047_1185, w_047_1186, w_047_1188, w_047_1190, w_047_1191, w_047_1193, w_047_1194, w_047_1195, w_047_1197, w_047_1198, w_047_1199, w_047_1201, w_047_1202, w_047_1203, w_047_1204, w_047_1205, w_047_1206, w_047_1208, w_047_1209, w_047_1210, w_047_1211, w_047_1212, w_047_1213, w_047_1214, w_047_1215, w_047_1216, w_047_1217, w_047_1220, w_047_1221, w_047_1222, w_047_1225, w_047_1226, w_047_1227, w_047_1229, w_047_1230, w_047_1231, w_047_1232, w_047_1233, w_047_1234, w_047_1235, w_047_1237, w_047_1238, w_047_1239, w_047_1241, w_047_1242, w_047_1243, w_047_1244, w_047_1245, w_047_1246, w_047_1248, w_047_1249, w_047_1250, w_047_1251, w_047_1252, w_047_1253, w_047_1257, w_047_1259, w_047_1260, w_047_1261, w_047_1262, w_047_1263, w_047_1265, w_047_1266, w_047_1267, w_047_1268, w_047_1269, w_047_1270, w_047_1271, w_047_1272, w_047_1273, w_047_1276, w_047_1277, w_047_1278, w_047_1279, w_047_1281, w_047_1282, w_047_1283, w_047_1284, w_047_1285, w_047_1286, w_047_1287, w_047_1288, w_047_1289, w_047_1290, w_047_1291, w_047_1293, w_047_1294, w_047_1295, w_047_1296, w_047_1298, w_047_1299, w_047_1301, w_047_1302, w_047_1304, w_047_1305, w_047_1306, w_047_1307, w_047_1309, w_047_1310, w_047_1311, w_047_1312, w_047_1313, w_047_1314, w_047_1315, w_047_1316, w_047_1318, w_047_1320, w_047_1321, w_047_1323, w_047_1324, w_047_1326, w_047_1327, w_047_1328, w_047_1330, w_047_1331, w_047_1333, w_047_1334, w_047_1335, w_047_1336, w_047_1337, w_047_1338, w_047_1339, w_047_1340, w_047_1342, w_047_1343, w_047_1344, w_047_1346, w_047_1347, w_047_1349, w_047_1350, w_047_1352, w_047_1354, w_047_1355, w_047_1356, w_047_1357, w_047_1358, w_047_1359, w_047_1360, w_047_1363, w_047_1364, w_047_1365, w_047_1366, w_047_1367, w_047_1368, w_047_1369, w_047_1370, w_047_1371, w_047_1372, w_047_1373, w_047_1375, w_047_1376, w_047_1378, w_047_1379, w_047_1380, w_047_1381, w_047_1382, w_047_1383, w_047_1384, w_047_1385, w_047_1386, w_047_1387, w_047_1389, w_047_1390, w_047_1393, w_047_1394, w_047_1396, w_047_1397, w_047_1398, w_047_1400, w_047_1401, w_047_1402, w_047_1404, w_047_1405, w_047_1406, w_047_1407, w_047_1408, w_047_1409, w_047_1410, w_047_1411, w_047_1412, w_047_1413, w_047_1414, w_047_1415, w_047_1417, w_047_1418, w_047_1420, w_047_1422, w_047_1423, w_047_1424, w_047_1425, w_047_1426, w_047_1427, w_047_1429, w_047_1430, w_047_1431, w_047_1432, w_047_1433, w_047_1435, w_047_1437, w_047_1438, w_047_1439, w_047_1440, w_047_1441, w_047_1443, w_047_1445, w_047_1446, w_047_1447, w_047_1449, w_047_1450, w_047_1451, w_047_1452, w_047_1453, w_047_1454, w_047_1456, w_047_1458, w_047_1459, w_047_1460, w_047_1461, w_047_1462, w_047_1463, w_047_1464, w_047_1465, w_047_1466, w_047_1467, w_047_1468, w_047_1469, w_047_1470, w_047_1471, w_047_1472, w_047_1473, w_047_1475, w_047_1477, w_047_1478, w_047_1479, w_047_1481, w_047_1482, w_047_1484, w_047_1485, w_047_1486, w_047_1487, w_047_1489, w_047_1490, w_047_1491, w_047_1492, w_047_1493, w_047_1494, w_047_1496, w_047_1497, w_047_1498, w_047_1499, w_047_1500, w_047_1501, w_047_1502, w_047_1503, w_047_1504, w_047_1506, w_047_1507, w_047_1509, w_047_1510, w_047_1511, w_047_1512, w_047_1513, w_047_1514, w_047_1515, w_047_1516, w_047_1517, w_047_1519, w_047_1520, w_047_1521, w_047_1522, w_047_1523, w_047_1524, w_047_1525, w_047_1526, w_047_1527, w_047_1528, w_047_1530, w_047_1532, w_047_1534, w_047_1535, w_047_1536, w_047_1537, w_047_1539, w_047_1540, w_047_1541, w_047_1542, w_047_1543, w_047_1544, w_047_1549, w_047_1551, w_047_1552, w_047_1553, w_047_1554, w_047_1555, w_047_1556, w_047_1557, w_047_1558, w_047_1559, w_047_1560, w_047_1561, w_047_1562, w_047_1563, w_047_1564, w_047_1565, w_047_1566, w_047_1567, w_047_1568, w_047_1569, w_047_1571, w_047_1572, w_047_1573, w_047_1574, w_047_1575, w_047_1576, w_047_1577, w_047_1579, w_047_1580, w_047_1581, w_047_1582, w_047_1583, w_047_1584, w_047_1585, w_047_1586, w_047_1587, w_047_1590, w_047_1591, w_047_1592, w_047_1594, w_047_1595, w_047_1596, w_047_1597, w_047_1598, w_047_1599, w_047_1601, w_047_1602, w_047_1603, w_047_1604, w_047_1608, w_047_1609, w_047_1611, w_047_1612, w_047_1613, w_047_1614, w_047_1615, w_047_1616, w_047_1617, w_047_1618, w_047_1619, w_047_1620, w_047_1622, w_047_1623, w_047_1624, w_047_1625, w_047_1626, w_047_1627, w_047_1628, w_047_1629, w_047_1630, w_047_1631, w_047_1632, w_047_1633, w_047_1634, w_047_1635, w_047_1636, w_047_1637, w_047_1638, w_047_1640, w_047_1641, w_047_1642, w_047_1643, w_047_1645, w_047_1646, w_047_1647, w_047_1648, w_047_1650, w_047_1651, w_047_1652, w_047_1654, w_047_1655, w_047_1656, w_047_1658, w_047_1659, w_047_1660, w_047_1662, w_047_1663, w_047_1664, w_047_1665, w_047_1666, w_047_1667, w_047_1668, w_047_1671, w_047_1672, w_047_1673, w_047_1674, w_047_1675, w_047_1677, w_047_1678, w_047_1681, w_047_1682, w_047_1683, w_047_1684, w_047_1685, w_047_1686, w_047_1687, w_047_1688, w_047_1689, w_047_1690, w_047_1691, w_047_1692, w_047_1693, w_047_1694, w_047_1695, w_047_1696, w_047_1697, w_047_1698, w_047_1699, w_047_1700, w_047_1701, w_047_1702, w_047_1703, w_047_1704, w_047_1706, w_047_1707, w_047_1708, w_047_1709, w_047_1710, w_047_1711, w_047_1712, w_047_1714, w_047_1715, w_047_1716, w_047_1717, w_047_1718, w_047_1719, w_047_1720, w_047_1721, w_047_1723, w_047_1724, w_047_1725, w_047_1726, w_047_1727, w_047_1728, w_047_1729, w_047_1730, w_047_1731, w_047_1732, w_047_1733, w_047_1735, w_047_1736, w_047_1737, w_047_1738, w_047_1739, w_047_1740, w_047_1742, w_047_1743, w_047_1744, w_047_1745, w_047_1746, w_047_1747, w_047_1748, w_047_1749, w_047_1751, w_047_1754, w_047_1755, w_047_1756, w_047_1757, w_047_1758, w_047_1761, w_047_1762, w_047_1763, w_047_1764, w_047_1765, w_047_1766, w_047_1767, w_047_1768, w_047_1769, w_047_1770, w_047_1772, w_047_1773, w_047_1774, w_047_1775, w_047_1777, w_047_1778, w_047_1779, w_047_1780, w_047_1781, w_047_1784, w_047_1785, w_047_1786, w_047_1787, w_047_1788, w_047_1789, w_047_1790, w_047_1791, w_047_1793, w_047_1794, w_047_1795, w_047_1796, w_047_1798, w_047_1799, w_047_1801, w_047_1802, w_047_1804, w_047_1805, w_047_1806, w_047_1807, w_047_1808, w_047_1809, w_047_1810, w_047_1811, w_047_1814, w_047_1815, w_047_1816, w_047_1817, w_047_1818, w_047_1819, w_047_1820, w_047_1821, w_047_1822, w_047_1823, w_047_1824, w_047_1825, w_047_1827, w_047_1829, w_047_1830, w_047_1831, w_047_1832, w_047_1833, w_047_1835, w_047_1836, w_047_1837, w_047_1839, w_047_1840, w_047_1841, w_047_1842, w_047_1843, w_047_1844, w_047_1845, w_047_1846, w_047_1847, w_047_1848, w_047_1849, w_047_1850, w_047_1851, w_047_1853, w_047_1854, w_047_1855, w_047_1856, w_047_1857, w_047_1858, w_047_1859, w_047_1860, w_047_1862, w_047_1864, w_047_1865, w_047_1866, w_047_1867, w_047_1869, w_047_1870, w_047_1871, w_047_1872, w_047_1873, w_047_1875, w_047_1876, w_047_1877, w_047_1879, w_047_1880, w_047_1882, w_047_1883, w_047_1884, w_047_1886, w_047_1888, w_047_1889, w_047_1890, w_047_1891, w_047_1893, w_047_1895, w_047_1896, w_047_1897, w_047_1898, w_047_1900, w_047_1901, w_047_1902, w_047_1904, w_047_1905, w_047_1906, w_047_1908, w_047_1909, w_047_1910, w_047_1912, w_047_1913, w_047_1914, w_047_1915, w_047_1917, w_047_1918, w_047_1919, w_047_1920, w_047_1921, w_047_1922, w_047_1923, w_047_1925, w_047_1926, w_047_1928, w_047_1929, w_047_1930, w_047_1931, w_047_1932, w_047_1933, w_047_1934, w_047_1935, w_047_1936, w_047_1937, w_047_1938, w_047_1939, w_047_1940, w_047_1941, w_047_1942, w_047_1943, w_047_1944, w_047_1945, w_047_1946, w_047_1947, w_047_1948, w_047_1949, w_047_1950, w_047_1951, w_047_1952, w_047_1953, w_047_1954, w_047_1955, w_047_1956, w_047_1957, w_047_1958, w_047_1959, w_047_1960, w_047_1961, w_047_1962, w_047_1963, w_047_1964, w_047_1965, w_047_1966, w_047_1967, w_047_1969, w_047_1970, w_047_1974, w_047_1975, w_047_1976, w_047_1977, w_047_1978, w_047_1980, w_047_1981, w_047_1982, w_047_1983, w_047_1984, w_047_1986, w_047_1988, w_047_1990, w_047_1991, w_047_1993, w_047_1994, w_047_1995, w_047_1997, w_047_1998, w_047_1999, w_047_2000, w_047_2001, w_047_2002, w_047_2003, w_047_2004, w_047_2006, w_047_2007, w_047_2008, w_047_2009, w_047_2011, w_047_2012, w_047_2014, w_047_2015, w_047_2017, w_047_2018, w_047_2019, w_047_2020, w_047_2021, w_047_2023, w_047_2024, w_047_2025, w_047_2027, w_047_2028, w_047_2029, w_047_2031, w_047_2032, w_047_2035, w_047_2036, w_047_2037, w_047_2038, w_047_2039, w_047_2040, w_047_2041, w_047_2042, w_047_2043, w_047_2044, w_047_2045, w_047_2046, w_047_2047, w_047_2048, w_047_2049, w_047_2050, w_047_2051, w_047_2052, w_047_2053, w_047_2054, w_047_2055, w_047_2057, w_047_2058, w_047_2059, w_047_2061, w_047_2064, w_047_2065, w_047_2066, w_047_2067, w_047_2068, w_047_2069, w_047_2070, w_047_2072, w_047_2073, w_047_2074, w_047_2075, w_047_2076, w_047_2077, w_047_2078, w_047_2079, w_047_2080, w_047_2081, w_047_2084, w_047_2085, w_047_2086, w_047_2087, w_047_2088, w_047_2089, w_047_2091, w_047_2092, w_047_2094, w_047_2095, w_047_2096, w_047_2097, w_047_2098, w_047_2099, w_047_2100, w_047_2101, w_047_2102, w_047_2103, w_047_2104, w_047_2105, w_047_2106, w_047_2107, w_047_2108, w_047_2109, w_047_2110, w_047_2111, w_047_2112, w_047_2113, w_047_2114, w_047_2116, w_047_2117, w_047_2119, w_047_2120, w_047_2121, w_047_2123, w_047_2124, w_047_2126, w_047_2128, w_047_2130, w_047_2132, w_047_2133, w_047_2135, w_047_2136, w_047_2137, w_047_2139, w_047_2141, w_047_2142, w_047_2144, w_047_2145, w_047_2147, w_047_2148, w_047_2149, w_047_2150, w_047_2151, w_047_2152, w_047_2153, w_047_2154, w_047_2155, w_047_2156, w_047_2157, w_047_2158, w_047_2159, w_047_2160, w_047_2161, w_047_2162, w_047_2163, w_047_2164, w_047_2165, w_047_2166, w_047_2167, w_047_2168, w_047_2169, w_047_2170, w_047_2171, w_047_2172, w_047_2173, w_047_2176, w_047_2177, w_047_2178, w_047_2179, w_047_2180, w_047_2182, w_047_2183, w_047_2184, w_047_2185, w_047_2186, w_047_2187, w_047_2188, w_047_2189, w_047_2190, w_047_2191, w_047_2192, w_047_2194, w_047_2196, w_047_2197, w_047_2199, w_047_2200, w_047_2202, w_047_2203, w_047_2204, w_047_2205, w_047_2207, w_047_2209, w_047_2210, w_047_2211, w_047_2213, w_047_2214, w_047_2215, w_047_2216, w_047_2217, w_047_2219, w_047_2220, w_047_2221, w_047_2223, w_047_2224, w_047_2225, w_047_2226, w_047_2227, w_047_2228, w_047_2229, w_047_2230, w_047_2231, w_047_2233, w_047_2234, w_047_2236, w_047_2237, w_047_2238, w_047_2241, w_047_2243, w_047_2244, w_047_2245, w_047_2246, w_047_2247, w_047_2249, w_047_2250, w_047_2251, w_047_2252, w_047_2253, w_047_2254, w_047_2255, w_047_2256, w_047_2257, w_047_2260, w_047_2261, w_047_2264, w_047_2265, w_047_2267, w_047_2268, w_047_2269, w_047_2271, w_047_2272, w_047_2273, w_047_2274, w_047_2276, w_047_2278, w_047_2279, w_047_2280, w_047_2281, w_047_2282, w_047_2283, w_047_2284, w_047_2285, w_047_2287, w_047_2288, w_047_2289, w_047_2291, w_047_2292, w_047_2296, w_047_2297, w_047_2298, w_047_2299, w_047_2300, w_047_2301, w_047_2303, w_047_2304, w_047_2305, w_047_2306, w_047_2309, w_047_2310, w_047_2311, w_047_2312, w_047_2314, w_047_2315, w_047_2316, w_047_2317, w_047_2318, w_047_2319, w_047_2320, w_047_2321, w_047_2323, w_047_2324, w_047_2325, w_047_2326, w_047_2327, w_047_2329, w_047_2330, w_047_2331, w_047_2332, w_047_2333, w_047_2334, w_047_2336, w_047_2337, w_047_2338, w_047_2339, w_047_2340, w_047_2341, w_047_2342, w_047_2343, w_047_2344, w_047_2345, w_047_2346, w_047_2347, w_047_2348, w_047_2349, w_047_2350, w_047_2351, w_047_2352, w_047_2353, w_047_2354, w_047_2355, w_047_2356, w_047_2357, w_047_2359, w_047_2362, w_047_2363, w_047_2364, w_047_2365, w_047_2366, w_047_2367, w_047_2368, w_047_2369, w_047_2370, w_047_2371, w_047_2372, w_047_2375, w_047_2376, w_047_2378, w_047_2379, w_047_2380, w_047_2381, w_047_2382, w_047_2383, w_047_2385, w_047_2387, w_047_2388, w_047_2389, w_047_2390, w_047_2391, w_047_2392, w_047_2393, w_047_2394, w_047_2395, w_047_2396, w_047_2397, w_047_2398, w_047_2399, w_047_2400, w_047_2401, w_047_2402, w_047_2404, w_047_2406, w_047_2407, w_047_2409, w_047_2411, w_047_2412, w_047_2415, w_047_2417, w_047_2419, w_047_2420, w_047_2421, w_047_2422, w_047_2423, w_047_2424, w_047_2426, w_047_2427, w_047_2428, w_047_2429, w_047_2431, w_047_2432, w_047_2435, w_047_2436, w_047_2437, w_047_2438, w_047_2440, w_047_2441, w_047_2443, w_047_2444, w_047_2445, w_047_2446, w_047_2447, w_047_2448, w_047_2449, w_047_2450, w_047_2451, w_047_2452, w_047_2453, w_047_2454, w_047_2455, w_047_2457, w_047_2458, w_047_2461, w_047_2462, w_047_2463, w_047_2464, w_047_2466, w_047_2467, w_047_2468, w_047_2469, w_047_2470, w_047_2472, w_047_2473, w_047_2475, w_047_2476, w_047_2477, w_047_2478, w_047_2480, w_047_2482, w_047_2483, w_047_2484, w_047_2485, w_047_2486, w_047_2487, w_047_2488, w_047_2489, w_047_2490, w_047_2492, w_047_2493, w_047_2494, w_047_2496, w_047_2497, w_047_2498, w_047_2499, w_047_2500, w_047_2501, w_047_2502, w_047_2503, w_047_2504, w_047_2505, w_047_2506, w_047_2507, w_047_2508, w_047_2509, w_047_2510, w_047_2511, w_047_2512, w_047_2514, w_047_2516, w_047_2519, w_047_2520, w_047_2522, w_047_2523, w_047_2526, w_047_2528, w_047_2529, w_047_2530, w_047_2531, w_047_2532, w_047_2533, w_047_2534, w_047_2535, w_047_2536, w_047_2537, w_047_2538, w_047_2539, w_047_2540, w_047_2541, w_047_2542, w_047_2543, w_047_2544, w_047_2545, w_047_2546, w_047_2547, w_047_2548, w_047_2549, w_047_2550, w_047_2551, w_047_2552, w_047_2554, w_047_2555, w_047_2556, w_047_2557, w_047_2558, w_047_2560, w_047_2561, w_047_2562, w_047_2563, w_047_2564, w_047_2565, w_047_2566, w_047_2567, w_047_2571, w_047_2572, w_047_2574, w_047_2575, w_047_2576, w_047_2577, w_047_2578, w_047_2579, w_047_2580, w_047_2581, w_047_2582, w_047_2583, w_047_2584, w_047_2586, w_047_2587, w_047_2590, w_047_2591, w_047_2592, w_047_2593, w_047_2594, w_047_2595, w_047_2596, w_047_2597, w_047_2598, w_047_2599, w_047_2600, w_047_2602, w_047_2603, w_047_2604, w_047_2606, w_047_2607, w_047_2608, w_047_2609, w_047_2610, w_047_2611, w_047_2612, w_047_2613, w_047_2614, w_047_2615, w_047_2616, w_047_2618, w_047_2620, w_047_2622, w_047_2623, w_047_2625, w_047_2626, w_047_2628, w_047_2629, w_047_2630, w_047_2631, w_047_2632, w_047_2633, w_047_2634, w_047_2635, w_047_2636, w_047_2637, w_047_2638, w_047_2639, w_047_2640, w_047_2642, w_047_2643, w_047_2644, w_047_2646, w_047_2647, w_047_2648, w_047_2649, w_047_2650, w_047_2651, w_047_2652, w_047_2653, w_047_2654, w_047_2655, w_047_2657, w_047_2658, w_047_2659, w_047_2660, w_047_2661, w_047_2662, w_047_2664, w_047_2665, w_047_2666, w_047_2667, w_047_2668, w_047_2669, w_047_2671, w_047_2672, w_047_2674, w_047_2675, w_047_2676, w_047_2677, w_047_2678, w_047_2679, w_047_2680, w_047_2682, w_047_2683, w_047_2684, w_047_2685, w_047_2686, w_047_2687, w_047_2689, w_047_2690, w_047_2691, w_047_2693, w_047_2694, w_047_2695, w_047_2696, w_047_2697, w_047_2698, w_047_2699, w_047_2700, w_047_2701, w_047_2702, w_047_2703, w_047_2704, w_047_2705, w_047_2706, w_047_2709, w_047_2710, w_047_2712, w_047_2713, w_047_2715, w_047_2716, w_047_2717, w_047_2718, w_047_2719, w_047_2720, w_047_2721, w_047_2722, w_047_2723, w_047_2724, w_047_2725, w_047_2726, w_047_2727, w_047_2728, w_047_2731, w_047_2732, w_047_2734, w_047_2735, w_047_2736, w_047_2737, w_047_2738, w_047_2739, w_047_2741, w_047_2742, w_047_2743, w_047_2744, w_047_2745, w_047_2746, w_047_2747, w_047_2748, w_047_2749, w_047_2750, w_047_2751, w_047_2752, w_047_2753, w_047_2754, w_047_2755, w_047_2756, w_047_2757, w_047_2758, w_047_2759, w_047_2762, w_047_2763, w_047_2764, w_047_2765, w_047_2767, w_047_2768, w_047_2771, w_047_2772, w_047_2773, w_047_2774, w_047_2775, w_047_2776, w_047_2777, w_047_2778, w_047_2779, w_047_2780, w_047_2782, w_047_2783, w_047_2784, w_047_2785, w_047_2786, w_047_2787, w_047_2788, w_047_2789, w_047_2791, w_047_2792, w_047_2793, w_047_2794, w_047_2795, w_047_2796, w_047_2797, w_047_2802, w_047_2803, w_047_2804, w_047_2805, w_047_2806, w_047_2807, w_047_2808, w_047_2809, w_047_2810, w_047_2811, w_047_2812, w_047_2813, w_047_2814, w_047_2815, w_047_2816, w_047_2817, w_047_2819, w_047_2820, w_047_2821, w_047_2822, w_047_2823, w_047_2824, w_047_2825, w_047_2826, w_047_2827, w_047_2828, w_047_2831, w_047_2832, w_047_2833, w_047_2835, w_047_2836, w_047_2837, w_047_2839, w_047_2840, w_047_2841, w_047_2842, w_047_2843, w_047_2844, w_047_2845, w_047_2846, w_047_2848, w_047_2849, w_047_2850, w_047_2851, w_047_2855, w_047_2856, w_047_2857, w_047_2858, w_047_2859, w_047_2860, w_047_2862, w_047_2864, w_047_2865, w_047_2866, w_047_2867, w_047_2868, w_047_2870, w_047_2871, w_047_2872, w_047_2873, w_047_2874, w_047_2875, w_047_2876, w_047_2877, w_047_2879, w_047_2881, w_047_2883, w_047_2885, w_047_2886, w_047_2887, w_047_2888, w_047_2889, w_047_2890, w_047_2891, w_047_2892, w_047_2893, w_047_2894, w_047_2895, w_047_2896, w_047_2899, w_047_2900, w_047_2901, w_047_2902, w_047_2903, w_047_2904, w_047_2906, w_047_2907, w_047_2909, w_047_2911, w_047_2912, w_047_2913, w_047_2914, w_047_2915, w_047_2916, w_047_2917, w_047_2919, w_047_2920, w_047_2921, w_047_2922, w_047_2923, w_047_2924, w_047_2925, w_047_2926, w_047_2927, w_047_2928, w_047_2930, w_047_2931, w_047_2932, w_047_2933, w_047_2935, w_047_2936, w_047_2937, w_047_2938, w_047_2939, w_047_2941, w_047_2942, w_047_2943, w_047_2944, w_047_2945, w_047_2947, w_047_2948, w_047_2949, w_047_2950, w_047_2951, w_047_2952, w_047_2953, w_047_2954, w_047_2955, w_047_2956, w_047_2957, w_047_2958, w_047_2961, w_047_2962, w_047_2963, w_047_2964, w_047_2965, w_047_2966, w_047_2967, w_047_2968, w_047_2969, w_047_2970, w_047_2971, w_047_2972, w_047_2973, w_047_2974, w_047_2975, w_047_2976, w_047_2977, w_047_2978, w_047_2979, w_047_2980, w_047_2981, w_047_2982, w_047_2984, w_047_2985, w_047_2986, w_047_2987, w_047_2988, w_047_2989, w_047_2990, w_047_2991, w_047_2992, w_047_2993, w_047_2994, w_047_2995, w_047_2997, w_047_2998, w_047_2999, w_047_3000, w_047_3001, w_047_3002, w_047_3003, w_047_3004, w_047_3005, w_047_3008, w_047_3010, w_047_3012, w_047_3013, w_047_3014, w_047_3015, w_047_3017, w_047_3018, w_047_3020, w_047_3021, w_047_3023, w_047_3025, w_047_3027, w_047_3028, w_047_3031, w_047_3033, w_047_3034, w_047_3035, w_047_3036, w_047_3038, w_047_3039, w_047_3041, w_047_3042, w_047_3043, w_047_3044, w_047_3045, w_047_3046, w_047_3047, w_047_3048, w_047_3049, w_047_3050, w_047_3052, w_047_3055, w_047_3056, w_047_3057, w_047_3060, w_047_3061, w_047_3062, w_047_3063, w_047_3065, w_047_3066, w_047_3068, w_047_3069, w_047_3070, w_047_3071, w_047_3072, w_047_3073, w_047_3074, w_047_3075, w_047_3076, w_047_3078, w_047_3080, w_047_3081, w_047_3083, w_047_3084, w_047_3085, w_047_3086, w_047_3087, w_047_3088, w_047_3089, w_047_3090, w_047_3092, w_047_3093, w_047_3094, w_047_3095, w_047_3096, w_047_3097, w_047_3098, w_047_3099, w_047_3100, w_047_3101, w_047_3102, w_047_3103, w_047_3104, w_047_3105, w_047_3106, w_047_3107, w_047_3108, w_047_3109, w_047_3110, w_047_3111, w_047_3112, w_047_3113, w_047_3114, w_047_3115, w_047_3116, w_047_3117, w_047_3118, w_047_3119, w_047_3120, w_047_3121, w_047_3122, w_047_3125, w_047_3126, w_047_3127, w_047_3128, w_047_3129, w_047_3130, w_047_3131, w_047_3132, w_047_3134, w_047_3136, w_047_3137, w_047_3138, w_047_3140, w_047_3141, w_047_3142, w_047_3143, w_047_3144, w_047_3145, w_047_3146, w_047_3147, w_047_3148, w_047_3150, w_047_3151, w_047_3153, w_047_3154, w_047_3156, w_047_3158, w_047_3159, w_047_3161, w_047_3162, w_047_3163, w_047_3164, w_047_3165, w_047_3166, w_047_3167, w_047_3168, w_047_3169, w_047_3170, w_047_3171, w_047_3172, w_047_3173, w_047_3174, w_047_3175, w_047_3176, w_047_3177, w_047_3178, w_047_3181, w_047_3182, w_047_3183, w_047_3184, w_047_3185, w_047_3186, w_047_3187, w_047_3188, w_047_3189, w_047_3190, w_047_3191, w_047_3192, w_047_3193, w_047_3194, w_047_3195, w_047_3196, w_047_3197, w_047_3198, w_047_3199, w_047_3200, w_047_3201, w_047_3202, w_047_3203, w_047_3204, w_047_3206, w_047_3207, w_047_3208, w_047_3209, w_047_3211, w_047_3212, w_047_3214;
  wire w_048_000, w_048_001, w_048_002, w_048_004, w_048_006, w_048_007, w_048_008, w_048_009, w_048_010, w_048_011, w_048_012, w_048_013, w_048_014, w_048_015, w_048_016, w_048_020, w_048_021, w_048_022, w_048_023, w_048_024, w_048_025, w_048_026, w_048_027, w_048_028, w_048_030, w_048_031, w_048_032, w_048_036, w_048_037, w_048_039, w_048_041, w_048_042, w_048_043, w_048_044, w_048_045, w_048_046, w_048_047, w_048_049, w_048_050, w_048_052, w_048_053, w_048_055, w_048_056, w_048_057, w_048_058, w_048_059, w_048_060, w_048_061, w_048_062, w_048_063, w_048_065, w_048_067, w_048_068, w_048_070, w_048_071, w_048_072, w_048_073, w_048_075, w_048_076, w_048_077, w_048_080, w_048_081, w_048_083, w_048_084, w_048_086, w_048_088, w_048_089, w_048_091, w_048_096, w_048_097, w_048_098, w_048_102, w_048_104, w_048_105, w_048_111, w_048_113, w_048_115, w_048_119, w_048_127, w_048_132, w_048_133, w_048_136, w_048_139, w_048_140, w_048_141, w_048_144, w_048_145, w_048_148, w_048_149, w_048_154, w_048_155, w_048_156, w_048_158, w_048_159, w_048_161, w_048_167, w_048_170, w_048_173, w_048_175, w_048_176, w_048_178, w_048_182, w_048_190, w_048_192, w_048_194, w_048_197, w_048_199, w_048_201, w_048_202, w_048_208, w_048_209, w_048_213, w_048_214, w_048_218, w_048_219, w_048_226, w_048_227, w_048_228, w_048_231, w_048_233, w_048_236, w_048_237, w_048_238, w_048_242, w_048_243, w_048_245, w_048_246, w_048_249, w_048_251, w_048_252, w_048_253, w_048_257, w_048_260, w_048_263, w_048_266, w_048_267, w_048_268, w_048_269, w_048_271, w_048_272, w_048_274, w_048_276, w_048_278, w_048_280, w_048_282, w_048_284, w_048_285, w_048_287, w_048_289, w_048_293, w_048_296, w_048_298, w_048_302, w_048_305, w_048_307, w_048_309, w_048_311, w_048_316, w_048_317, w_048_319, w_048_320, w_048_323, w_048_326, w_048_327, w_048_329, w_048_330, w_048_333, w_048_337, w_048_338, w_048_339, w_048_342, w_048_344, w_048_345, w_048_348, w_048_350, w_048_355, w_048_356, w_048_359, w_048_361, w_048_363, w_048_376, w_048_378, w_048_384, w_048_385, w_048_387, w_048_390, w_048_392, w_048_393, w_048_395, w_048_396, w_048_401, w_048_406, w_048_408, w_048_409, w_048_410, w_048_412, w_048_413, w_048_419, w_048_422, w_048_428, w_048_429, w_048_430, w_048_431, w_048_435, w_048_436, w_048_437, w_048_438, w_048_439, w_048_440, w_048_444, w_048_451, w_048_452, w_048_453, w_048_454, w_048_456, w_048_458, w_048_462, w_048_465, w_048_466, w_048_469, w_048_472, w_048_473, w_048_474, w_048_475, w_048_477, w_048_480, w_048_481, w_048_482, w_048_483, w_048_485, w_048_488, w_048_489, w_048_490, w_048_493, w_048_495, w_048_496, w_048_497, w_048_498, w_048_502, w_048_503, w_048_505, w_048_508, w_048_509, w_048_511, w_048_512, w_048_514, w_048_516, w_048_519, w_048_520, w_048_521, w_048_522, w_048_523, w_048_524, w_048_525, w_048_530, w_048_532, w_048_533, w_048_534, w_048_535, w_048_536, w_048_538, w_048_539, w_048_540, w_048_541, w_048_542, w_048_545, w_048_549, w_048_550, w_048_551, w_048_557, w_048_560, w_048_561, w_048_564, w_048_567, w_048_568, w_048_569, w_048_570, w_048_572, w_048_576, w_048_578, w_048_579, w_048_587, w_048_591, w_048_592, w_048_593, w_048_596, w_048_599, w_048_600, w_048_605, w_048_607, w_048_613, w_048_614, w_048_615, w_048_616, w_048_617, w_048_621, w_048_623, w_048_624, w_048_625, w_048_626, w_048_632, w_048_634, w_048_640, w_048_642, w_048_645, w_048_646, w_048_647, w_048_650, w_048_651, w_048_654, w_048_655, w_048_659, w_048_662, w_048_664, w_048_665, w_048_667, w_048_671, w_048_672, w_048_676, w_048_678, w_048_679, w_048_680, w_048_681, w_048_683, w_048_684, w_048_686, w_048_691, w_048_692, w_048_693, w_048_695, w_048_697, w_048_706, w_048_709, w_048_710, w_048_711, w_048_712, w_048_713, w_048_717, w_048_720, w_048_722, w_048_727, w_048_731, w_048_733, w_048_734, w_048_735, w_048_736, w_048_737, w_048_742, w_048_744, w_048_746, w_048_750, w_048_753, w_048_754, w_048_757, w_048_759, w_048_761, w_048_763, w_048_764, w_048_766, w_048_767, w_048_769, w_048_771, w_048_774, w_048_777, w_048_781, w_048_782, w_048_784, w_048_787, w_048_789, w_048_794, w_048_795, w_048_798, w_048_799, w_048_800, w_048_802, w_048_806, w_048_807, w_048_809, w_048_810, w_048_813, w_048_815, w_048_817, w_048_822, w_048_823, w_048_827, w_048_829, w_048_831, w_048_835, w_048_837, w_048_838, w_048_839, w_048_841, w_048_842, w_048_843, w_048_844, w_048_846, w_048_847, w_048_849, w_048_850, w_048_856, w_048_857, w_048_859, w_048_862, w_048_866, w_048_867, w_048_869, w_048_872, w_048_875, w_048_876, w_048_878, w_048_883, w_048_884, w_048_885, w_048_889, w_048_892, w_048_893, w_048_896, w_048_897, w_048_901, w_048_902, w_048_904, w_048_906, w_048_907, w_048_911, w_048_913, w_048_918, w_048_919, w_048_920, w_048_921, w_048_926, w_048_927, w_048_928, w_048_931, w_048_932, w_048_933, w_048_940, w_048_942, w_048_943, w_048_953, w_048_954, w_048_955, w_048_960, w_048_963, w_048_965, w_048_967, w_048_972, w_048_973, w_048_977, w_048_978, w_048_980, w_048_985, w_048_987, w_048_990, w_048_992, w_048_995, w_048_996, w_048_997, w_048_998, w_048_1000, w_048_1005, w_048_1008, w_048_1009, w_048_1010, w_048_1013, w_048_1015, w_048_1021, w_048_1029, w_048_1031, w_048_1032, w_048_1036, w_048_1037, w_048_1038, w_048_1039, w_048_1040, w_048_1041, w_048_1042, w_048_1045, w_048_1047, w_048_1048, w_048_1052, w_048_1059, w_048_1060, w_048_1062, w_048_1063, w_048_1065, w_048_1066, w_048_1069, w_048_1071, w_048_1073, w_048_1075, w_048_1076, w_048_1077, w_048_1078, w_048_1079, w_048_1083, w_048_1085, w_048_1089, w_048_1093, w_048_1095, w_048_1096, w_048_1098, w_048_1101, w_048_1102, w_048_1103, w_048_1105, w_048_1109, w_048_1111, w_048_1114, w_048_1115, w_048_1118, w_048_1119, w_048_1123, w_048_1124, w_048_1125, w_048_1127, w_048_1130, w_048_1132, w_048_1134, w_048_1136, w_048_1138, w_048_1139, w_048_1142, w_048_1145, w_048_1146, w_048_1147, w_048_1148, w_048_1149, w_048_1151, w_048_1152, w_048_1154, w_048_1157, w_048_1163, w_048_1165, w_048_1167, w_048_1168, w_048_1169, w_048_1171, w_048_1172, w_048_1174, w_048_1175, w_048_1177, w_048_1178, w_048_1179, w_048_1181, w_048_1182, w_048_1184, w_048_1185, w_048_1187, w_048_1188, w_048_1190, w_048_1195, w_048_1197, w_048_1199, w_048_1201, w_048_1203, w_048_1207, w_048_1208, w_048_1209, w_048_1212, w_048_1213, w_048_1216, w_048_1217, w_048_1220, w_048_1222, w_048_1223, w_048_1226, w_048_1228, w_048_1230, w_048_1233, w_048_1236, w_048_1240, w_048_1244, w_048_1246, w_048_1249, w_048_1250, w_048_1254, w_048_1256, w_048_1257, w_048_1258, w_048_1262, w_048_1263, w_048_1265, w_048_1268, w_048_1269, w_048_1271, w_048_1272, w_048_1273, w_048_1275, w_048_1282, w_048_1285, w_048_1292, w_048_1293, w_048_1296, w_048_1297, w_048_1298, w_048_1303, w_048_1304, w_048_1306, w_048_1307, w_048_1308, w_048_1310, w_048_1315, w_048_1319, w_048_1323, w_048_1327, w_048_1331, w_048_1332, w_048_1333, w_048_1335, w_048_1338, w_048_1343, w_048_1345, w_048_1346, w_048_1355, w_048_1359, w_048_1360, w_048_1369, w_048_1371, w_048_1372, w_048_1373, w_048_1374, w_048_1375, w_048_1377, w_048_1380, w_048_1383, w_048_1385, w_048_1388, w_048_1393, w_048_1397, w_048_1399, w_048_1401, w_048_1403, w_048_1405, w_048_1406, w_048_1409, w_048_1416, w_048_1417, w_048_1420, w_048_1422, w_048_1425, w_048_1426, w_048_1427, w_048_1428, w_048_1429, w_048_1431, w_048_1432, w_048_1435, w_048_1436, w_048_1438, w_048_1441, w_048_1446, w_048_1447, w_048_1450, w_048_1454, w_048_1456, w_048_1459, w_048_1461, w_048_1462, w_048_1463, w_048_1464, w_048_1468, w_048_1478, w_048_1479, w_048_1480, w_048_1486, w_048_1491, w_048_1494, w_048_1496, w_048_1497, w_048_1499, w_048_1501, w_048_1502, w_048_1503, w_048_1506, w_048_1508, w_048_1509, w_048_1511, w_048_1512, w_048_1513, w_048_1515, w_048_1516, w_048_1517, w_048_1518, w_048_1520, w_048_1523, w_048_1524, w_048_1527, w_048_1531, w_048_1533, w_048_1534, w_048_1537, w_048_1538, w_048_1539, w_048_1542, w_048_1551, w_048_1553, w_048_1554, w_048_1557, w_048_1560, w_048_1561, w_048_1565, w_048_1569, w_048_1570, w_048_1574, w_048_1576, w_048_1577, w_048_1587, w_048_1588, w_048_1590, w_048_1591, w_048_1592, w_048_1594, w_048_1595, w_048_1601, w_048_1602, w_048_1603, w_048_1605, w_048_1607, w_048_1615, w_048_1617, w_048_1619, w_048_1622, w_048_1628, w_048_1629, w_048_1630, w_048_1633, w_048_1637, w_048_1639, w_048_1641, w_048_1643, w_048_1644, w_048_1645, w_048_1647, w_048_1649, w_048_1652, w_048_1655, w_048_1656, w_048_1658, w_048_1659, w_048_1661, w_048_1668, w_048_1671, w_048_1672, w_048_1674, w_048_1675, w_048_1679, w_048_1681, w_048_1685, w_048_1686, w_048_1688, w_048_1689, w_048_1694, w_048_1696, w_048_1698, w_048_1699, w_048_1701, w_048_1702, w_048_1705, w_048_1709, w_048_1712, w_048_1713, w_048_1714, w_048_1715, w_048_1716, w_048_1719, w_048_1721, w_048_1724, w_048_1727, w_048_1728, w_048_1729, w_048_1731, w_048_1732, w_048_1733, w_048_1734, w_048_1738, w_048_1739, w_048_1744, w_048_1745, w_048_1748, w_048_1751, w_048_1752, w_048_1754, w_048_1756, w_048_1757, w_048_1758, w_048_1760, w_048_1762, w_048_1764, w_048_1765, w_048_1767, w_048_1768, w_048_1769, w_048_1772, w_048_1776, w_048_1777, w_048_1778, w_048_1782, w_048_1784, w_048_1792, w_048_1793, w_048_1795, w_048_1797, w_048_1807, w_048_1810, w_048_1815, w_048_1817, w_048_1820, w_048_1823, w_048_1826, w_048_1827, w_048_1829, w_048_1830, w_048_1833, w_048_1835, w_048_1836, w_048_1840, w_048_1847, w_048_1853, w_048_1857, w_048_1863, w_048_1865, w_048_1866, w_048_1867, w_048_1871, w_048_1872, w_048_1874, w_048_1875, w_048_1881, w_048_1884, w_048_1885, w_048_1887, w_048_1892, w_048_1893, w_048_1896, w_048_1897, w_048_1899, w_048_1900, w_048_1901, w_048_1902, w_048_1905, w_048_1907, w_048_1910, w_048_1912, w_048_1913, w_048_1915, w_048_1917, w_048_1918, w_048_1919, w_048_1920, w_048_1921, w_048_1922, w_048_1923, w_048_1925, w_048_1926, w_048_1931, w_048_1934, w_048_1935, w_048_1936, w_048_1938, w_048_1942, w_048_1943, w_048_1945, w_048_1948, w_048_1949, w_048_1950, w_048_1951, w_048_1953, w_048_1955, w_048_1956, w_048_1957, w_048_1961, w_048_1962, w_048_1964, w_048_1966, w_048_1968, w_048_1977, w_048_1979, w_048_1980, w_048_1992, w_048_1996, w_048_1998, w_048_1999, w_048_2000, w_048_2001, w_048_2006, w_048_2007, w_048_2008, w_048_2010, w_048_2014, w_048_2015, w_048_2017, w_048_2018, w_048_2019, w_048_2022, w_048_2026, w_048_2028, w_048_2033, w_048_2036, w_048_2037, w_048_2039, w_048_2046, w_048_2047, w_048_2050, w_048_2057, w_048_2058, w_048_2059, w_048_2063, w_048_2070, w_048_2072, w_048_2075, w_048_2077, w_048_2079, w_048_2080, w_048_2081, w_048_2082, w_048_2083, w_048_2084, w_048_2087, w_048_2088, w_048_2090, w_048_2096, w_048_2097, w_048_2099, w_048_2101, w_048_2113, w_048_2114, w_048_2118, w_048_2120, w_048_2124, w_048_2125, w_048_2130, w_048_2132, w_048_2133, w_048_2135, w_048_2136, w_048_2137, w_048_2138, w_048_2139, w_048_2141, w_048_2142, w_048_2143, w_048_2144, w_048_2148, w_048_2151, w_048_2153, w_048_2155, w_048_2168, w_048_2170, w_048_2171, w_048_2172, w_048_2173, w_048_2174, w_048_2175, w_048_2181, w_048_2182, w_048_2187, w_048_2188, w_048_2190, w_048_2192, w_048_2193, w_048_2196, w_048_2201, w_048_2204, w_048_2206, w_048_2208, w_048_2210, w_048_2214, w_048_2215, w_048_2217, w_048_2222, w_048_2224, w_048_2226, w_048_2227, w_048_2229, w_048_2230, w_048_2231, w_048_2234, w_048_2237, w_048_2238, w_048_2241, w_048_2245, w_048_2246, w_048_2247, w_048_2248, w_048_2249, w_048_2253, w_048_2255, w_048_2257, w_048_2258, w_048_2261, w_048_2262, w_048_2263, w_048_2267, w_048_2268, w_048_2276, w_048_2277, w_048_2280, w_048_2283, w_048_2285, w_048_2288, w_048_2289, w_048_2293, w_048_2294, w_048_2295, w_048_2296, w_048_2298, w_048_2302, w_048_2304, w_048_2309, w_048_2312, w_048_2321, w_048_2322, w_048_2325, w_048_2333, w_048_2335, w_048_2340, w_048_2341, w_048_2343, w_048_2349, w_048_2351, w_048_2352, w_048_2354, w_048_2355, w_048_2357, w_048_2358, w_048_2359, w_048_2362, w_048_2363, w_048_2367, w_048_2370, w_048_2371, w_048_2372, w_048_2373, w_048_2376, w_048_2378, w_048_2380, w_048_2381, w_048_2384, w_048_2385, w_048_2388, w_048_2389, w_048_2391, w_048_2393, w_048_2394, w_048_2395, w_048_2398, w_048_2401, w_048_2403, w_048_2407, w_048_2409, w_048_2411, w_048_2414, w_048_2416, w_048_2417, w_048_2418, w_048_2419, w_048_2421, w_048_2424, w_048_2428, w_048_2434, w_048_2435, w_048_2436, w_048_2438, w_048_2441, w_048_2445, w_048_2446, w_048_2448, w_048_2449, w_048_2454, w_048_2457, w_048_2458, w_048_2459, w_048_2461, w_048_2462, w_048_2463, w_048_2466, w_048_2467, w_048_2468, w_048_2469, w_048_2470, w_048_2471, w_048_2473, w_048_2475, w_048_2477, w_048_2479, w_048_2480, w_048_2482, w_048_2486, w_048_2488, w_048_2489, w_048_2492, w_048_2494, w_048_2495, w_048_2496, w_048_2498, w_048_2500, w_048_2507, w_048_2511, w_048_2513, w_048_2514, w_048_2515, w_048_2520, w_048_2521, w_048_2522, w_048_2524, w_048_2526, w_048_2528, w_048_2531, w_048_2539, w_048_2541, w_048_2542, w_048_2546, w_048_2550, w_048_2552, w_048_2554, w_048_2556, w_048_2558, w_048_2561, w_048_2563, w_048_2566, w_048_2569, w_048_2575, w_048_2579, w_048_2581, w_048_2586, w_048_2592, w_048_2595, w_048_2597, w_048_2599, w_048_2602, w_048_2603, w_048_2609, w_048_2610, w_048_2612, w_048_2618, w_048_2621, w_048_2625, w_048_2627, w_048_2629, w_048_2630, w_048_2631, w_048_2636, w_048_2638, w_048_2640, w_048_2646, w_048_2647, w_048_2648, w_048_2650, w_048_2652, w_048_2653, w_048_2654, w_048_2656, w_048_2658, w_048_2659, w_048_2661, w_048_2664, w_048_2665, w_048_2666, w_048_2668, w_048_2670, w_048_2675, w_048_2676, w_048_2677, w_048_2678, w_048_2679, w_048_2684, w_048_2686, w_048_2687, w_048_2688, w_048_2690, w_048_2692, w_048_2693, w_048_2699, w_048_2700, w_048_2701, w_048_2703, w_048_2706, w_048_2707, w_048_2711, w_048_2713, w_048_2716, w_048_2720, w_048_2721, w_048_2724, w_048_2727, w_048_2731, w_048_2743, w_048_2748, w_048_2750, w_048_2752, w_048_2754, w_048_2756, w_048_2759, w_048_2764, w_048_2766, w_048_2776, w_048_2784, w_048_2786, w_048_2791, w_048_2792, w_048_2793, w_048_2795, w_048_2797, w_048_2803, w_048_2806, w_048_2808, w_048_2812, w_048_2814, w_048_2815, w_048_2820, w_048_2821, w_048_2823, w_048_2824, w_048_2827, w_048_2830, w_048_2831, w_048_2836, w_048_2838, w_048_2840, w_048_2841, w_048_2843, w_048_2844, w_048_2846, w_048_2851, w_048_2853, w_048_2856, w_048_2857, w_048_2858, w_048_2860, w_048_2861, w_048_2862, w_048_2863, w_048_2864, w_048_2865, w_048_2867, w_048_2868, w_048_2869, w_048_2870, w_048_2871, w_048_2872, w_048_2873, w_048_2874, w_048_2883, w_048_2885, w_048_2887, w_048_2888, w_048_2894, w_048_2895, w_048_2901, w_048_2908, w_048_2913, w_048_2915, w_048_2916, w_048_2917, w_048_2918, w_048_2920, w_048_2921, w_048_2924, w_048_2925, w_048_2926, w_048_2927, w_048_2929, w_048_2935, w_048_2939, w_048_2940, w_048_2946, w_048_2949, w_048_2953, w_048_2955, w_048_2956, w_048_2958, w_048_2964, w_048_2965, w_048_2966, w_048_2971, w_048_2972, w_048_2973, w_048_2975, w_048_2977, w_048_2978, w_048_2980, w_048_2982, w_048_2983, w_048_2984, w_048_2987, w_048_2988, w_048_2989, w_048_2990, w_048_2994, w_048_2995, w_048_2998, w_048_3000, w_048_3003, w_048_3006, w_048_3009, w_048_3010, w_048_3011, w_048_3013, w_048_3015, w_048_3016, w_048_3018, w_048_3024, w_048_3026, w_048_3027, w_048_3028, w_048_3037, w_048_3040, w_048_3042, w_048_3047, w_048_3050, w_048_3051, w_048_3054, w_048_3056, w_048_3057, w_048_3059, w_048_3060, w_048_3063, w_048_3069, w_048_3070, w_048_3074, w_048_3076, w_048_3078, w_048_3079, w_048_3085, w_048_3097, w_048_3098, w_048_3100, w_048_3102, w_048_3103, w_048_3108, w_048_3110, w_048_3113, w_048_3117, w_048_3119, w_048_3121, w_048_3123, w_048_3124, w_048_3126, w_048_3127, w_048_3128, w_048_3130, w_048_3134, w_048_3137, w_048_3139, w_048_3142, w_048_3146, w_048_3148, w_048_3149, w_048_3150, w_048_3153, w_048_3164, w_048_3166, w_048_3167, w_048_3170, w_048_3171, w_048_3174, w_048_3175, w_048_3177, w_048_3178, w_048_3180, w_048_3181, w_048_3183, w_048_3184, w_048_3186, w_048_3190, w_048_3195, w_048_3196, w_048_3199, w_048_3204, w_048_3205, w_048_3207, w_048_3210, w_048_3213, w_048_3220, w_048_3222, w_048_3223, w_048_3225, w_048_3229, w_048_3230, w_048_3233, w_048_3234, w_048_3236, w_048_3237, w_048_3238, w_048_3239, w_048_3241, w_048_3243, w_048_3246, w_048_3249, w_048_3253, w_048_3254, w_048_3255, w_048_3258, w_048_3261, w_048_3262, w_048_3263, w_048_3265, w_048_3269, w_048_3271, w_048_3275, w_048_3277, w_048_3278, w_048_3281, w_048_3282, w_048_3285, w_048_3288, w_048_3289, w_048_3292, w_048_3293, w_048_3296, w_048_3297, w_048_3298, w_048_3299, w_048_3300, w_048_3305, w_048_3308, w_048_3309, w_048_3310, w_048_3311, w_048_3313, w_048_3317, w_048_3319, w_048_3320, w_048_3322, w_048_3323, w_048_3324, w_048_3326, w_048_3327, w_048_3328, w_048_3329, w_048_3330, w_048_3331, w_048_3335, w_048_3341, w_048_3342, w_048_3347, w_048_3348, w_048_3350, w_048_3351, w_048_3352, w_048_3353, w_048_3358, w_048_3359, w_048_3360, w_048_3361, w_048_3362, w_048_3364, w_048_3367, w_048_3370, w_048_3373, w_048_3375, w_048_3377, w_048_3383, w_048_3390, w_048_3391, w_048_3393, w_048_3396, w_048_3397, w_048_3398, w_048_3400, w_048_3402, w_048_3407, w_048_3409, w_048_3410, w_048_3411, w_048_3412, w_048_3417, w_048_3422, w_048_3424, w_048_3429, w_048_3430, w_048_3431, w_048_3433, w_048_3434, w_048_3435, w_048_3436, w_048_3437, w_048_3445, w_048_3451, w_048_3452, w_048_3453, w_048_3454, w_048_3458, w_048_3461, w_048_3462, w_048_3463, w_048_3466, w_048_3470, w_048_3472, w_048_3475, w_048_3476, w_048_3481, w_048_3483, w_048_3484, w_048_3485, w_048_3486, w_048_3492, w_048_3497, w_048_3498, w_048_3505, w_048_3508, w_048_3514, w_048_3517, w_048_3520, w_048_3523, w_048_3526, w_048_3532, w_048_3535, w_048_3545, w_048_3547, w_048_3548, w_048_3550, w_048_3552, w_048_3553, w_048_3556, w_048_3560, w_048_3561, w_048_3563, w_048_3565, w_048_3566, w_048_3570, w_048_3571, w_048_3574, w_048_3576, w_048_3579, w_048_3583, w_048_3586, w_048_3587, w_048_3591, w_048_3592, w_048_3596, w_048_3601, w_048_3604, w_048_3605, w_048_3609, w_048_3611, w_048_3612, w_048_3613, w_048_3614, w_048_3618, w_048_3620, w_048_3621, w_048_3623, w_048_3624, w_048_3630, w_048_3632, w_048_3633, w_048_3634, w_048_3638, w_048_3642, w_048_3643, w_048_3647, w_048_3650, w_048_3652, w_048_3653, w_048_3655, w_048_3657, w_048_3658, w_048_3661, w_048_3662, w_048_3665, w_048_3668, w_048_3670, w_048_3671, w_048_3678, w_048_3679, w_048_3682, w_048_3683, w_048_3688, w_048_3697, w_048_3699, w_048_3700, w_048_3701, w_048_3706, w_048_3707, w_048_3708, w_048_3711, w_048_3715, w_048_3717, w_048_3720, w_048_3722, w_048_3723, w_048_3731, w_048_3732, w_048_3735, w_048_3737, w_048_3740, w_048_3741, w_048_3744, w_048_3745, w_048_3746, w_048_3747, w_048_3750, w_048_3752, w_048_3755, w_048_3757, w_048_3759, w_048_3762, w_048_3765, w_048_3770, w_048_3771, w_048_3774, w_048_3780, w_048_3781, w_048_3783, w_048_3786, w_048_3789, w_048_3790, w_048_3793, w_048_3796, w_048_3799, w_048_3800, w_048_3803, w_048_3805, w_048_3806, w_048_3808, w_048_3809, w_048_3813, w_048_3814, w_048_3815, w_048_3820, w_048_3821, w_048_3824, w_048_3826, w_048_3829, w_048_3830, w_048_3831, w_048_3833, w_048_3834, w_048_3836, w_048_3837, w_048_3839, w_048_3842, w_048_3843, w_048_3845, w_048_3850, w_048_3851, w_048_3853, w_048_3854, w_048_3855, w_048_3856, w_048_3857, w_048_3858, w_048_3862, w_048_3864, w_048_3865, w_048_3866, w_048_3867, w_048_3868, w_048_3870, w_048_3873, w_048_3879, w_048_3881, w_048_3882, w_048_3883, w_048_3885, w_048_3886, w_048_3887, w_048_3889, w_048_3896, w_048_3899, w_048_3902, w_048_3904, w_048_3905, w_048_3906, w_048_3909, w_048_3910, w_048_3911, w_048_3916, w_048_3918, w_048_3919, w_048_3920, w_048_3927, w_048_3928, w_048_3929, w_048_3931, w_048_3934, w_048_3935, w_048_3936, w_048_3937, w_048_3939, w_048_3940, w_048_3943, w_048_3946, w_048_3947, w_048_3948, w_048_3949, w_048_3952, w_048_3954, w_048_3960, w_048_3962, w_048_3968, w_048_3972, w_048_3974, w_048_3975, w_048_3978, w_048_3979, w_048_3982, w_048_3983, w_048_3986, w_048_3987, w_048_3989, w_048_3990, w_048_3995, w_048_4000, w_048_4001, w_048_4009, w_048_4010, w_048_4011, w_048_4012, w_048_4016, w_048_4017, w_048_4018, w_048_4019, w_048_4020, w_048_4021, w_048_4022, w_048_4024, w_048_4028, w_048_4032, w_048_4034, w_048_4038, w_048_4041, w_048_4045, w_048_4049, w_048_4051, w_048_4052, w_048_4053, w_048_4054, w_048_4055, w_048_4064, w_048_4065, w_048_4068, w_048_4070, w_048_4072, w_048_4075, w_048_4077, w_048_4080, w_048_4081, w_048_4082, w_048_4083, w_048_4084, w_048_4085, w_048_4086, w_048_4093, w_048_4096, w_048_4100, w_048_4102, w_048_4106, w_048_4109, w_048_4112, w_048_4113, w_048_4116, w_048_4118, w_048_4123, w_048_4125, w_048_4130, w_048_4132, w_048_4133, w_048_4137, w_048_4139, w_048_4144, w_048_4158, w_048_4159, w_048_4160, w_048_4162, w_048_4167, w_048_4172, w_048_4173, w_048_4174, w_048_4175, w_048_4176, w_048_4178, w_048_4179, w_048_4181, w_048_4182, w_048_4184, w_048_4186, w_048_4187, w_048_4188, w_048_4189, w_048_4190, w_048_4191, w_048_4194, w_048_4195, w_048_4197, w_048_4198, w_048_4199, w_048_4203, w_048_4204, w_048_4206, w_048_4208, w_048_4214, w_048_4220, w_048_4221, w_048_4222, w_048_4225, w_048_4229, w_048_4231, w_048_4232, w_048_4233, w_048_4238, w_048_4240, w_048_4241, w_048_4242, w_048_4252, w_048_4255, w_048_4257, w_048_4260, w_048_4263, w_048_4264, w_048_4273, w_048_4274, w_048_4275, w_048_4276, w_048_4278, w_048_4279, w_048_4280, w_048_4282, w_048_4283, w_048_4285, w_048_4288, w_048_4289, w_048_4290, w_048_4292, w_048_4294, w_048_4295, w_048_4296, w_048_4298, w_048_4299, w_048_4305, w_048_4307, w_048_4308, w_048_4310, w_048_4314, w_048_4317, w_048_4319, w_048_4332, w_048_4335, w_048_4342, w_048_4343, w_048_4344, w_048_4348, w_048_4352, w_048_4354, w_048_4359, w_048_4360, w_048_4362, w_048_4363, w_048_4366, w_048_4370, w_048_4374, w_048_4376, w_048_4377, w_048_4378, w_048_4382, w_048_4384, w_048_4385, w_048_4387, w_048_4391, w_048_4392, w_048_4394, w_048_4397, w_048_4399, w_048_4401, w_048_4402, w_048_4409, w_048_4410, w_048_4411, w_048_4415, w_048_4416, w_048_4417, w_048_4421, w_048_4425, w_048_4426, w_048_4431, w_048_4432, w_048_4433, w_048_4434, w_048_4436, w_048_4437, w_048_4439, w_048_4442, w_048_4443, w_048_4447, w_048_4449, w_048_4450, w_048_4451, w_048_4452, w_048_4453, w_048_4454, w_048_4455, w_048_4456, w_048_4457, w_048_4458, w_048_4459, w_048_4461, w_048_4462, w_048_4472, w_048_4473, w_048_4475, w_048_4476, w_048_4478, w_048_4479, w_048_4482, w_048_4483, w_048_4484, w_048_4486, w_048_4490, w_048_4492, w_048_4497, w_048_4502, w_048_4508, w_048_4509, w_048_4513, w_048_4514, w_048_4520, w_048_4521, w_048_4523, w_048_4527, w_048_4528, w_048_4529, w_048_4531, w_048_4533, w_048_4536, w_048_4549, w_048_4550, w_048_4551, w_048_4553, w_048_4555, w_048_4556, w_048_4557, w_048_4566, w_048_4568, w_048_4569, w_048_4571, w_048_4573, w_048_4574, w_048_4577, w_048_4582, w_048_4583, w_048_4587, w_048_4589, w_048_4591, w_048_4593, w_048_4595, w_048_4600, w_048_4601, w_048_4602, w_048_4604, w_048_4607, w_048_4608, w_048_4611, w_048_4612, w_048_4616, w_048_4617, w_048_4621, w_048_4624, w_048_4627, w_048_4628, w_048_4629, w_048_4632, w_048_4634, w_048_4635, w_048_4636, w_048_4638, w_048_4640, w_048_4642, w_048_4643, w_048_4645, w_048_4646, w_048_4649, w_048_4650, w_048_4651, w_048_4652, w_048_4655, w_048_4658, w_048_4659, w_048_4660, w_048_4661, w_048_4662, w_048_4663, w_048_4666, w_048_4667, w_048_4669, w_048_4670, w_048_4671, w_048_4673, w_048_4675, w_048_4676, w_048_4678, w_048_4682, w_048_4684, w_048_4685, w_048_4687, w_048_4689, w_048_4690, w_048_4691, w_048_4692, w_048_4694, w_048_4695, w_048_4697, w_048_4698, w_048_4699, w_048_4700, w_048_4702, w_048_4704, w_048_4705, w_048_4708, w_048_4712, w_048_4716, w_048_4717, w_048_4722, w_048_4725, w_048_4739, w_048_4741, w_048_4742, w_048_4743, w_048_4747, w_048_4750, w_048_4751, w_048_4752, w_048_4753, w_048_4755, w_048_4756, w_048_4758, w_048_4761, w_048_4762, w_048_4764, w_048_4766, w_048_4767, w_048_4771, w_048_4774, w_048_4775, w_048_4778, w_048_4779, w_048_4783, w_048_4788, w_048_4791, w_048_4793, w_048_4794, w_048_4797, w_048_4800, w_048_4804, w_048_4805, w_048_4810, w_048_4813, w_048_4815, w_048_4816, w_048_4820, w_048_4826, w_048_4830, w_048_4832, w_048_4833, w_048_4834, w_048_4836, w_048_4838, w_048_4841, w_048_4843, w_048_4845, w_048_4847, w_048_4851, w_048_4852, w_048_4854, w_048_4858, w_048_4859, w_048_4860, w_048_4862, w_048_4863, w_048_4865, w_048_4866, w_048_4869, w_048_4870, w_048_4871, w_048_4873, w_048_4874, w_048_4876, w_048_4879, w_048_4882, w_048_4886, w_048_4887, w_048_4892, w_048_4894, w_048_4895, w_048_4896, w_048_4898, w_048_4899, w_048_4901, w_048_4903, w_048_4904, w_048_4910, w_048_4914, w_048_4918, w_048_4925, w_048_4926, w_048_4927, w_048_4931, w_048_4941, w_048_4942, w_048_4944, w_048_4947, w_048_4950, w_048_4952, w_048_4954, w_048_4956, w_048_4958, w_048_4959, w_048_4960, w_048_4961, w_048_4966, w_048_4968, w_048_4972, w_048_4975, w_048_4978, w_048_4979, w_048_4981, w_048_4983, w_048_4987, w_048_4989, w_048_4994, w_048_4999, w_048_5000, w_048_5002, w_048_5004, w_048_5005, w_048_5008, w_048_5009, w_048_5011, w_048_5014, w_048_5015, w_048_5016, w_048_5019, w_048_5020, w_048_5024, w_048_5026, w_048_5027, w_048_5031, w_048_5034, w_048_5035, w_048_5037, w_048_5039, w_048_5040, w_048_5042, w_048_5043, w_048_5044, w_048_5046, w_048_5051, w_048_5053, w_048_5054, w_048_5055, w_048_5057, w_048_5058, w_048_5060, w_048_5067, w_048_5068, w_048_5071, w_048_5072, w_048_5074, w_048_5081, w_048_5083, w_048_5085, w_048_5090, w_048_5095, w_048_5096, w_048_5097, w_048_5098, w_048_5099, w_048_5100, w_048_5104, w_048_5105, w_048_5109, w_048_5111, w_048_5114, w_048_5116, w_048_5119, w_048_5120, w_048_5121, w_048_5130, w_048_5131, w_048_5132, w_048_5133, w_048_5135, w_048_5138, w_048_5143, w_048_5144, w_048_5147, w_048_5149, w_048_5150, w_048_5152, w_048_5156, w_048_5158, w_048_5159, w_048_5167, w_048_5171, w_048_5174, w_048_5181, w_048_5182, w_048_5183, w_048_5185, w_048_5189, w_048_5192, w_048_5194, w_048_5197, w_048_5199, w_048_5201, w_048_5203, w_048_5204, w_048_5205, w_048_5206, w_048_5207, w_048_5209, w_048_5210, w_048_5211, w_048_5214, w_048_5216, w_048_5221, w_048_5222, w_048_5223, w_048_5224, w_048_5229, w_048_5233, w_048_5235, w_048_5236, w_048_5242, w_048_5249, w_048_5252, w_048_5255, w_048_5256, w_048_5259, w_048_5263, w_048_5264, w_048_5265, w_048_5266, w_048_5270, w_048_5274, w_048_5275, w_048_5276, w_048_5279, w_048_5283, w_048_5284, w_048_5285, w_048_5288, w_048_5290, w_048_5292, w_048_5294, w_048_5295, w_048_5299, w_048_5301, w_048_5306, w_048_5307, w_048_5308, w_048_5309, w_048_5310, w_048_5311, w_048_5312, w_048_5313, w_048_5315, w_048_5321, w_048_5323, w_048_5328, w_048_5330, w_048_5334, w_048_5337, w_048_5338, w_048_5341, w_048_5342, w_048_5343, w_048_5344, w_048_5345, w_048_5349, w_048_5352, w_048_5354, w_048_5356, w_048_5357, w_048_5359, w_048_5362, w_048_5363, w_048_5365, w_048_5366, w_048_5372, w_048_5374, w_048_5375, w_048_5383, w_048_5385, w_048_5387, w_048_5388, w_048_5389, w_048_5390, w_048_5391, w_048_5392, w_048_5395, w_048_5397, w_048_5398, w_048_5401, w_048_5403, w_048_5408, w_048_5410, w_048_5411, w_048_5412, w_048_5416, w_048_5418, w_048_5420, w_048_5422, w_048_5425, w_048_5426, w_048_5430, w_048_5433, w_048_5434, w_048_5435, w_048_5438, w_048_5439, w_048_5447, w_048_5449, w_048_5451, w_048_5453, w_048_5455, w_048_5460, w_048_5467, w_048_5468, w_048_5469, w_048_5473, w_048_5477, w_048_5481, w_048_5483, w_048_5485, w_048_5489, w_048_5491, w_048_5493, w_048_5494, w_048_5496, w_048_5498, w_048_5499, w_048_5505, w_048_5506, w_048_5507, w_048_5508, w_048_5514, w_048_5517, w_048_5518, w_048_5519, w_048_5524, w_048_5526, w_048_5527, w_048_5534, w_048_5535, w_048_5537, w_048_5540, w_048_5541, w_048_5552, w_048_5554, w_048_5556, w_048_5559, w_048_5561, w_048_5565, w_048_5569, w_048_5574, w_048_5575, w_048_5578, w_048_5579, w_048_5582, w_048_5583, w_048_5586, w_048_5594, w_048_5598, w_048_5599, w_048_5604, w_048_5606, w_048_5607, w_048_5609, w_048_5613, w_048_5614, w_048_5615, w_048_5620, w_048_5621, w_048_5624, w_048_5628, w_048_5631, w_048_5635, w_048_5641, w_048_5642, w_048_5644, w_048_5646, w_048_5648, w_048_5649, w_048_5650, w_048_5651, w_048_5653, w_048_5654, w_048_5655, w_048_5659, w_048_5661, w_048_5667, w_048_5668, w_048_5674, w_048_5679, w_048_5680, w_048_5681, w_048_5682, w_048_5683, w_048_5685, w_048_5686, w_048_5687, w_048_5688, w_048_5690, w_048_5694, w_048_5695, w_048_5696, w_048_5697, w_048_5700, w_048_5701, w_048_5703, w_048_5704, w_048_5706, w_048_5707, w_048_5714, w_048_5715, w_048_5722, w_048_5726, w_048_5728, w_048_5729, w_048_5733, w_048_5734, w_048_5737, w_048_5738, w_048_5741, w_048_5742, w_048_5743, w_048_5745, w_048_5754, w_048_5755, w_048_5758, w_048_5764, w_048_5771, w_048_5773, w_048_5779, w_048_5780, w_048_5782, w_048_5783, w_048_5785, w_048_5786, w_048_5791, w_048_5792, w_048_5793, w_048_5795, w_048_5796, w_048_5798, w_048_5800, w_048_5802, w_048_5808, w_048_5811, w_048_5814, w_048_5815, w_048_5817, w_048_5818, w_048_5819, w_048_5820, w_048_5823, w_048_5826, w_048_5827, w_048_5830, w_048_5831, w_048_5833, w_048_5834, w_048_5838, w_048_5842, w_048_5843, w_048_5845, w_048_5848, w_048_5849, w_048_5851, w_048_5853, w_048_5856, w_048_5857, w_048_5863, w_048_5867, w_048_5869, w_048_5870, w_048_5878, w_048_5881, w_048_5882, w_048_5883, w_048_5887, w_048_5888, w_048_5889, w_048_5890, w_048_5892, w_048_5893, w_048_5894, w_048_5895, w_048_5900, w_048_5902, w_048_5904, w_048_5907, w_048_5909, w_048_5910, w_048_5912, w_048_5913, w_048_5918, w_048_5928, w_048_5930, w_048_5932, w_048_5935, w_048_5937, w_048_5939, w_048_5945, w_048_5949, w_048_5951, w_048_5952, w_048_5957, w_048_5960, w_048_5962, w_048_5963, w_048_5965, w_048_5967, w_048_5968, w_048_5974, w_048_5976, w_048_5977, w_048_5978, w_048_5979, w_048_5980, w_048_5981, w_048_5983, w_048_5988, w_048_5994, w_048_5995, w_048_5996, w_048_5999, w_048_6001, w_048_6002, w_048_6004, w_048_6005, w_048_6015, w_048_6017, w_048_6018, w_048_6023, w_048_6024, w_048_6027, w_048_6028, w_048_6033, w_048_6036, w_048_6037, w_048_6040, w_048_6042, w_048_6043, w_048_6049, w_048_6054, w_048_6057, w_048_6059, w_048_6062, w_048_6065, w_048_6067, w_048_6070, w_048_6084, w_048_6089, w_048_6094, w_048_6097, w_048_6098, w_048_6102, w_048_6107, w_048_6108, w_048_6109, w_048_6112, w_048_6118, w_048_6119, w_048_6123, w_048_6126, w_048_6127, w_048_6129, w_048_6130, w_048_6135, w_048_6137, w_048_6140, w_048_6143, w_048_6145, w_048_6148, w_048_6150, w_048_6151, w_048_6152, w_048_6153, w_048_6155, w_048_6156, w_048_6158, w_048_6161, w_048_6162, w_048_6166, w_048_6171, w_048_6175, w_048_6186, w_048_6200, w_048_6205, w_048_6206, w_048_6209, w_048_6212, w_048_6214, w_048_6216, w_048_6223, w_048_6228, w_048_6234, w_048_6239, w_048_6240, w_048_6242, w_048_6244, w_048_6245, w_048_6248, w_048_6249, w_048_6251, w_048_6256, w_048_6257, w_048_6258, w_048_6259, w_048_6261, w_048_6264, w_048_6268, w_048_6271, w_048_6276, w_048_6281, w_048_6282, w_048_6287, w_048_6289, w_048_6293, w_048_6297, w_048_6298, w_048_6299, w_048_6301, w_048_6302, w_048_6306, w_048_6307, w_048_6309, w_048_6311, w_048_6312, w_048_6313, w_048_6316, w_048_6318, w_048_6321, w_048_6324, w_048_6325, w_048_6326, w_048_6327, w_048_6329, w_048_6333, w_048_6334, w_048_6337, w_048_6339, w_048_6340, w_048_6346, w_048_6347, w_048_6348, w_048_6349, w_048_6350, w_048_6354, w_048_6357, w_048_6360, w_048_6361, w_048_6362, w_048_6364, w_048_6365, w_048_6367, w_048_6370, w_048_6371, w_048_6375, w_048_6380, w_048_6382, w_048_6383, w_048_6390, w_048_6391, w_048_6394, w_048_6396, w_048_6402, w_048_6408, w_048_6412, w_048_6413, w_048_6416, w_048_6418, w_048_6421, w_048_6425, w_048_6426, w_048_6427, w_048_6430, w_048_6431, w_048_6433, w_048_6434, w_048_6436, w_048_6439, w_048_6442, w_048_6443, w_048_6446, w_048_6449, w_048_6453, w_048_6455, w_048_6456, w_048_6457, w_048_6463, w_048_6470, w_048_6471, w_048_6472, w_048_6473, w_048_6476, w_048_6477, w_048_6478, w_048_6480, w_048_6481, w_048_6482, w_048_6483, w_048_6486, w_048_6487, w_048_6490, w_048_6496, w_048_6499, w_048_6507, w_048_6514, w_048_6515, w_048_6516, w_048_6517, w_048_6518, w_048_6520, w_048_6523, w_048_6524, w_048_6525, w_048_6526, w_048_6527, w_048_6529, w_048_6530, w_048_6531, w_048_6536, w_048_6538, w_048_6539, w_048_6541, w_048_6543, w_048_6547, w_048_6549, w_048_6555, w_048_6557, w_048_6559, w_048_6561, w_048_6563, w_048_6564, w_048_6566, w_048_6567, w_048_6569, w_048_6570, w_048_6571, w_048_6573, w_048_6574, w_048_6579, w_048_6585, w_048_6587, w_048_6588, w_048_6592, w_048_6594, w_048_6597, w_048_6598, w_048_6599, w_048_6602, w_048_6604, w_048_6609, w_048_6610, w_048_6612, w_048_6615, w_048_6616, w_048_6618, w_048_6619, w_048_6620, w_048_6621, w_048_6622, w_048_6623, w_048_6626, w_048_6627, w_048_6628, w_048_6632, w_048_6633, w_048_6635, w_048_6636, w_048_6639, w_048_6641, w_048_6642, w_048_6646, w_048_6647, w_048_6649, w_048_6653, w_048_6657, w_048_6658, w_048_6661, w_048_6663, w_048_6664, w_048_6665, w_048_6667, w_048_6668, w_048_6672, w_048_6673, w_048_6674, w_048_6675, w_048_6676, w_048_6677, w_048_6680, w_048_6684, w_048_6685, w_048_6687, w_048_6691, w_048_6692, w_048_6695, w_048_6696, w_048_6698, w_048_6700, w_048_6702, w_048_6705, w_048_6706, w_048_6708, w_048_6709, w_048_6712, w_048_6713, w_048_6715, w_048_6716, w_048_6720, w_048_6721, w_048_6726, w_048_6727, w_048_6728, w_048_6729, w_048_6732, w_048_6737, w_048_6738, w_048_6739, w_048_6740, w_048_6741, w_048_6742, w_048_6744, w_048_6748, w_048_6750, w_048_6751, w_048_6754, w_048_6755, w_048_6758, w_048_6759, w_048_6761, w_048_6765, w_048_6766, w_048_6768, w_048_6770, w_048_6771, w_048_6775, w_048_6783, w_048_6789, w_048_6790, w_048_6791, w_048_6793, w_048_6796, w_048_6798, w_048_6802, w_048_6803, w_048_6804, w_048_6806, w_048_6807, w_048_6810, w_048_6814, w_048_6815, w_048_6817, w_048_6819, w_048_6822, w_048_6824, w_048_6830, w_048_6833, w_048_6835, w_048_6839, w_048_6842, w_048_6845, w_048_6848, w_048_6850, w_048_6851, w_048_6852, w_048_6857, w_048_6860, w_048_6862, w_048_6863, w_048_6864, w_048_6865, w_048_6869, w_048_6870, w_048_6873, w_048_6874, w_048_6877, w_048_6878, w_048_6879, w_048_6881, w_048_6885, w_048_6886, w_048_6895, w_048_6897, w_048_6900, w_048_6901, w_048_6902, w_048_6903, w_048_6904, w_048_6905, w_048_6906, w_048_6911, w_048_6916, w_048_6917, w_048_6919, w_048_6920, w_048_6922, w_048_6925, w_048_6929, w_048_6930, w_048_6932, w_048_6933, w_048_6939, w_048_6943, w_048_6944, w_048_6945, w_048_6946, w_048_6947, w_048_6948, w_048_6954, w_048_6957, w_048_6959, w_048_6962, w_048_6964, w_048_6966, w_048_6967, w_048_6968, w_048_6969, w_048_6970, w_048_6972, w_048_6974, w_048_6975, w_048_6977, w_048_6986, w_048_6992, w_048_6993, w_048_6996, w_048_6997, w_048_6998, w_048_6999, w_048_7001, w_048_7006, w_048_7020, w_048_7021, w_048_7022, w_048_7024, w_048_7025, w_048_7026, w_048_7028, w_048_7030, w_048_7031, w_048_7035, w_048_7036, w_048_7037, w_048_7041, w_048_7047, w_048_7049, w_048_7050, w_048_7052, w_048_7053, w_048_7055, w_048_7057, w_048_7058, w_048_7059, w_048_7061, w_048_7065, w_048_7066, w_048_7068, w_048_7071, w_048_7072, w_048_7076, w_048_7077, w_048_7078, w_048_7083, w_048_7088, w_048_7089, w_048_7090, w_048_7091, w_048_7092, w_048_7095, w_048_7097, w_048_7098, w_048_7099, w_048_7100, w_048_7101, w_048_7103, w_048_7104, w_048_7105, w_048_7107, w_048_7108, w_048_7109, w_048_7112, w_048_7118, w_048_7120, w_048_7138, w_048_7140, w_048_7141, w_048_7143, w_048_7145, w_048_7146, w_048_7148, w_048_7151, w_048_7152, w_048_7154, w_048_7155, w_048_7156, w_048_7162, w_048_7165, w_048_7166, w_048_7167, w_048_7175, w_048_7176, w_048_7178, w_048_7179, w_048_7183, w_048_7187, w_048_7190, w_048_7200, w_048_7201, w_048_7203, w_048_7205, w_048_7206, w_048_7209, w_048_7211, w_048_7212, w_048_7215, w_048_7216, w_048_7231, w_048_7232, w_048_7235, w_048_7236, w_048_7238, w_048_7239, w_048_7241, w_048_7242, w_048_7243, w_048_7247, w_048_7248, w_048_7250, w_048_7252, w_048_7253, w_048_7254, w_048_7256, w_048_7260, w_048_7261, w_048_7263, w_048_7266, w_048_7272, w_048_7273, w_048_7275, w_048_7276, w_048_7277, w_048_7279, w_048_7280, w_048_7283, w_048_7285, w_048_7287, w_048_7295, w_048_7296, w_048_7299, w_048_7300, w_048_7301, w_048_7302, w_048_7303, w_048_7306, w_048_7307, w_048_7310, w_048_7312, w_048_7315, w_048_7319, w_048_7320, w_048_7324, w_048_7327, w_048_7328, w_048_7330, w_048_7331, w_048_7334, w_048_7337, w_048_7338, w_048_7339, w_048_7346, w_048_7349, w_048_7354, w_048_7355, w_048_7360, w_048_7361, w_048_7363, w_048_7366, w_048_7372, w_048_7374, w_048_7375, w_048_7376, w_048_7378, w_048_7382, w_048_7388, w_048_7389, w_048_7391, w_048_7393, w_048_7397, w_048_7399, w_048_7401, w_048_7403, w_048_7408, w_048_7409, w_048_7411, w_048_7413, w_048_7414, w_048_7416, w_048_7418, w_048_7420, w_048_7421, w_048_7425, w_048_7427, w_048_7429, w_048_7433, w_048_7435, w_048_7436, w_048_7437, w_048_7438, w_048_7441, w_048_7442, w_048_7445, w_048_7446, w_048_7448, w_048_7449, w_048_7450, w_048_7451, w_048_7456, w_048_7458, w_048_7472, w_048_7473, w_048_7474, w_048_7476, w_048_7479, w_048_7481, w_048_7483, w_048_7486, w_048_7488, w_048_7490, w_048_7492, w_048_7495, w_048_7496, w_048_7501, w_048_7503, w_048_7508, w_048_7509, w_048_7510, w_048_7512, w_048_7518, w_048_7521, w_048_7522, w_048_7526, w_048_7529, w_048_7533, w_048_7538, w_048_7540, w_048_7543, w_048_7544, w_048_7548, w_048_7550, w_048_7556, w_048_7558, w_048_7559, w_048_7560, w_048_7561, w_048_7562, w_048_7563, w_048_7565, w_048_7571, w_048_7572, w_048_7573, w_048_7574, w_048_7576, w_048_7578, w_048_7579, w_048_7580, w_048_7583, w_048_7585, w_048_7586, w_048_7587, w_048_7591, w_048_7594, w_048_7596, w_048_7597, w_048_7598, w_048_7601, w_048_7605, w_048_7609, w_048_7610, w_048_7615, w_048_7617, w_048_7618, w_048_7620, w_048_7621, w_048_7622, w_048_7626, w_048_7629, w_048_7630, w_048_7633, w_048_7638, w_048_7648, w_048_7649, w_048_7653, w_048_7656, w_048_7658, w_048_7660, w_048_7661, w_048_7665, w_048_7666, w_048_7668, w_048_7677, w_048_7678, w_048_7679, w_048_7681, w_048_7682, w_048_7693, w_048_7696, w_048_7700, w_048_7701, w_048_7703, w_048_7704, w_048_7705, w_048_7708, w_048_7709, w_048_7712, w_048_7715, w_048_7716, w_048_7719, w_048_7723, w_048_7725, w_048_7727, w_048_7728, w_048_7729, w_048_7736, w_048_7739, w_048_7740, w_048_7741, w_048_7744, w_048_7746, w_048_7747, w_048_7749, w_048_7757, w_048_7758, w_048_7761, w_048_7762, w_048_7764, w_048_7765, w_048_7766, w_048_7771, w_048_7774, w_048_7778, w_048_7779, w_048_7780, w_048_7782, w_048_7785, w_048_7786, w_048_7787, w_048_7789, w_048_7790, w_048_7791, w_048_7803, w_048_7806, w_048_7807, w_048_7808, w_048_7809, w_048_7811, w_048_7812, w_048_7813, w_048_7814, w_048_7815, w_048_7816, w_048_7817, w_048_7823, w_048_7826, w_048_7828, w_048_7830, w_048_7832, w_048_7833, w_048_7835, w_048_7836, w_048_7840, w_048_7841, w_048_7844, w_048_7847, w_048_7853, w_048_7858, w_048_7862, w_048_7865, w_048_7868, w_048_7869, w_048_7870, w_048_7872, w_048_7875, w_048_7880, w_048_7883, w_048_7884, w_048_7890, w_048_7891, w_048_7893, w_048_7895, w_048_7897, w_048_7900, w_048_7901, w_048_7902, w_048_7903, w_048_7904, w_048_7906, w_048_7907, w_048_7909, w_048_7915, w_048_7928, w_048_7930, w_048_7931, w_048_7932, w_048_7935, w_048_7938, w_048_7942, w_048_7943, w_048_7946, w_048_7947, w_048_7954, w_048_7955, w_048_7957, w_048_7960, w_048_7964, w_048_7966, w_048_7971, w_048_7974, w_048_7978, w_048_7980, w_048_7981, w_048_7985, w_048_7988, w_048_7989, w_048_7991, w_048_7996, w_048_8002, w_048_8003, w_048_8004, w_048_8005, w_048_8006, w_048_8009, w_048_8016, w_048_8020, w_048_8022, w_048_8023, w_048_8024, w_048_8026, w_048_8028, w_048_8029, w_048_8032, w_048_8034, w_048_8037, w_048_8038, w_048_8042, w_048_8043, w_048_8044, w_048_8045, w_048_8047, w_048_8052, w_048_8054, w_048_8059, w_048_8060, w_048_8061, w_048_8062, w_048_8063, w_048_8065, w_048_8066, w_048_8067, w_048_8074, w_048_8079, w_048_8080, w_048_8081, w_048_8083, w_048_8084, w_048_8086, w_048_8089, w_048_8091, w_048_8095, w_048_8096, w_048_8097, w_048_8098, w_048_8100, w_048_8102, w_048_8103, w_048_8107, w_048_8108, w_048_8109, w_048_8110, w_048_8112, w_048_8114, w_048_8118, w_048_8126, w_048_8128, w_048_8130, w_048_8138, w_048_8139, w_048_8140, w_048_8141, w_048_8142, w_048_8144, w_048_8145, w_048_8146, w_048_8152, w_048_8156, w_048_8157, w_048_8161, w_048_8164, w_048_8166, w_048_8168, w_048_8170, w_048_8171, w_048_8174, w_048_8175, w_048_8177, w_048_8179, w_048_8181, w_048_8183, w_048_8186, w_048_8187, w_048_8189, w_048_8193, w_048_8197, w_048_8198, w_048_8200, w_048_8201, w_048_8202, w_048_8212, w_048_8214, w_048_8216, w_048_8217, w_048_8218, w_048_8221, w_048_8229, w_048_8231, w_048_8232, w_048_8234, w_048_8235, w_048_8240, w_048_8243, w_048_8247, w_048_8248, w_048_8249, w_048_8251, w_048_8252, w_048_8254, w_048_8255, w_048_8260, w_048_8262, w_048_8263, w_048_8264, w_048_8266, w_048_8269, w_048_8270, w_048_8274, w_048_8275, w_048_8277, w_048_8279, w_048_8280, w_048_8282, w_048_8287, w_048_8288, w_048_8289, w_048_8290, w_048_8293, w_048_8294, w_048_8295, w_048_8298, w_048_8300, w_048_8304, w_048_8305, w_048_8306, w_048_8310, w_048_8313, w_048_8314, w_048_8316, w_048_8319, w_048_8321, w_048_8328, w_048_8329, w_048_8336, w_048_8337, w_048_8339, w_048_8340, w_048_8344, w_048_8346, w_048_8347, w_048_8349, w_048_8353, w_048_8354, w_048_8355, w_048_8356, w_048_8357, w_048_8360, w_048_8361, w_048_8362, w_048_8363, w_048_8364, w_048_8365, w_048_8367, w_048_8370, w_048_8371, w_048_8374, w_048_8377, w_048_8378, w_048_8382, w_048_8383, w_048_8385, w_048_8388, w_048_8390, w_048_8394, w_048_8395, w_048_8397, w_048_8399, w_048_8401, w_048_8402, w_048_8403, w_048_8404, w_048_8407, w_048_8408, w_048_8413, w_048_8416, w_048_8418, w_048_8421, w_048_8422, w_048_8424, w_048_8425, w_048_8428, w_048_8429, w_048_8434, w_048_8436, w_048_8437, w_048_8438, w_048_8440, w_048_8441, w_048_8442, w_048_8443, w_048_8446, w_048_8450, w_048_8454, w_048_8460, w_048_8463, w_048_8468, w_048_8469, w_048_8470, w_048_8473, w_048_8478, w_048_8479, w_048_8481, w_048_8487, w_048_8490, w_048_8491, w_048_8493, w_048_8494, w_048_8497, w_048_8498, w_048_8499, w_048_8500, w_048_8505, w_048_8510, w_048_8511, w_048_8513, w_048_8515, w_048_8519, w_048_8520, w_048_8522, w_048_8527, w_048_8540, w_048_8543, w_048_8545, w_048_8547, w_048_8548, w_048_8552, w_048_8556, w_048_8557, w_048_8561, w_048_8562, w_048_8563, w_048_8564, w_048_8566, w_048_8569, w_048_8571, w_048_8572, w_048_8575, w_048_8576, w_048_8581, w_048_8583, w_048_8587, w_048_8589, w_048_8590, w_048_8594, w_048_8599, w_048_8600, w_048_8604, w_048_8605, w_048_8608, w_048_8610, w_048_8611, w_048_8614, w_048_8617, w_048_8618, w_048_8619, w_048_8621, w_048_8626, w_048_8628, w_048_8629, w_048_8630, w_048_8634, w_048_8635, w_048_8636, w_048_8638, w_048_8640, w_048_8641, w_048_8644, w_048_8646, w_048_8649, w_048_8650, w_048_8653, w_048_8654, w_048_8655, w_048_8656, w_048_8657, w_048_8658, w_048_8659, w_048_8669, w_048_8671, w_048_8672, w_048_8677, w_048_8681, w_048_8684, w_048_8685, w_048_8686, w_048_8687, w_048_8689, w_048_8691, w_048_8692, w_048_8694, w_048_8699, w_048_8702, w_048_8703, w_048_8705, w_048_8709, w_048_8711, w_048_8714, w_048_8715, w_048_8718, w_048_8720, w_048_8721, w_048_8722, w_048_8724, w_048_8730, w_048_8731, w_048_8733, w_048_8735, w_048_8736, w_048_8737, w_048_8743, w_048_8745, w_048_8747, w_048_8749, w_048_8750, w_048_8752, w_048_8754, w_048_8757, w_048_8759, w_048_8760, w_048_8762, w_048_8764, w_048_8765, w_048_8766, w_048_8775, w_048_8777, w_048_8778, w_048_8779, w_048_8782, w_048_8783, w_048_8784, w_048_8786, w_048_8787, w_048_8788, w_048_8792, w_048_8794, w_048_8795, w_048_8801, w_048_8803, w_048_8807, w_048_8809, w_048_8810, w_048_8812, w_048_8813, w_048_8816, w_048_8819, w_048_8823, w_048_8824, w_048_8825, w_048_8827, w_048_8828, w_048_8831, w_048_8832, w_048_8834, w_048_8837, w_048_8839, w_048_8843, w_048_8845, w_048_8847, w_048_8848, w_048_8850, w_048_8851, w_048_8855, w_048_8859, w_048_8861, w_048_8862, w_048_8863, w_048_8866, w_048_8867, w_048_8868, w_048_8875, w_048_8877, w_048_8886, w_048_8891, w_048_8892, w_048_8893, w_048_8897, w_048_8898, w_048_8900, w_048_8903, w_048_8904, w_048_8910, w_048_8915, w_048_8916, w_048_8918, w_048_8920, w_048_8923, w_048_8924, w_048_8928, w_048_8929, w_048_8936, w_048_8939, w_048_8942, w_048_8943, w_048_8944, w_048_8946, w_048_8949, w_048_8953, w_048_8956, w_048_8957, w_048_8963, w_048_8964, w_048_8966, w_048_8967, w_048_8969, w_048_8973, w_048_8977, w_048_8981, w_048_8983, w_048_8984, w_048_8989, w_048_8991, w_048_8992, w_048_8994, w_048_8998, w_048_8999, w_048_9006, w_048_9011, w_048_9012, w_048_9013, w_048_9018, w_048_9019, w_048_9021, w_048_9022, w_048_9025, w_048_9027, w_048_9028, w_048_9031, w_048_9032, w_048_9039, w_048_9040, w_048_9041, w_048_9043, w_048_9045, w_048_9046, w_048_9049, w_048_9050, w_048_9051, w_048_9052, w_048_9057, w_048_9060, w_048_9061, w_048_9062, w_048_9064, w_048_9065, w_048_9068, w_048_9070, w_048_9074, w_048_9075, w_048_9077, w_048_9081, w_048_9082, w_048_9083, w_048_9086, w_048_9089, w_048_9091, w_048_9092, w_048_9096, w_048_9099, w_048_9104, w_048_9105, w_048_9107, w_048_9108, w_048_9111, w_048_9112, w_048_9113, w_048_9116, w_048_9117, w_048_9118, w_048_9120, w_048_9124, w_048_9127, w_048_9131, w_048_9132, w_048_9133, w_048_9135, w_048_9136, w_048_9137, w_048_9138, w_048_9143, w_048_9145, w_048_9151, w_048_9154, w_048_9156, w_048_9157, w_048_9160, w_048_9161, w_048_9164, w_048_9165, w_048_9169, w_048_9173, w_048_9175, w_048_9179, w_048_9182, w_048_9187, w_048_9192, w_048_9193, w_048_9194, w_048_9197, w_048_9199, w_048_9202, w_048_9203, w_048_9204, w_048_9206, w_048_9210, w_048_9213, w_048_9215, w_048_9217, w_048_9224, w_048_9227, w_048_9228, w_048_9229, w_048_9231, w_048_9233, w_048_9235, w_048_9238, w_048_9242, w_048_9243, w_048_9245, w_048_9247, w_048_9248, w_048_9249, w_048_9253, w_048_9254, w_048_9255, w_048_9257, w_048_9259, w_048_9261, w_048_9267, w_048_9268, w_048_9274, w_048_9275, w_048_9282, w_048_9284, w_048_9288, w_048_9289, w_048_9290, w_048_9292, w_048_9293, w_048_9294, w_048_9296, w_048_9298, w_048_9299, w_048_9301, w_048_9303, w_048_9304, w_048_9305, w_048_9307, w_048_9308, w_048_9311, w_048_9315, w_048_9318, w_048_9319, w_048_9323, w_048_9326, w_048_9330, w_048_9331, w_048_9332, w_048_9333, w_048_9334, w_048_9335, w_048_9337, w_048_9339, w_048_9340, w_048_9342, w_048_9343, w_048_9347, w_048_9349, w_048_9352, w_048_9354, w_048_9355, w_048_9357, w_048_9361, w_048_9363, w_048_9364, w_048_9367, w_048_9370, w_048_9371, w_048_9378, w_048_9379, w_048_9380, w_048_9382, w_048_9384, w_048_9385, w_048_9388, w_048_9390, w_048_9392, w_048_9394, w_048_9397, w_048_9398, w_048_9399, w_048_9401, w_048_9403, w_048_9404, w_048_9408, w_048_9415, w_048_9422, w_048_9425, w_048_9433, w_048_9438, w_048_9441, w_048_9445, w_048_9448, w_048_9451, w_048_9454, w_048_9456, w_048_9458, w_048_9461, w_048_9463, w_048_9465, w_048_9466, w_048_9467, w_048_9472, w_048_9474, w_048_9475, w_048_9477, w_048_9478, w_048_9479, w_048_9481, w_048_9482, w_048_9485, w_048_9486, w_048_9487, w_048_9488, w_048_9490, w_048_9491, w_048_9494, w_048_9495, w_048_9498, w_048_9499, w_048_9502, w_048_9505, w_048_9508, w_048_9510, w_048_9515, w_048_9516, w_048_9518, w_048_9519, w_048_9522, w_048_9525, w_048_9527, w_048_9528, w_048_9533, w_048_9535, w_048_9536, w_048_9537, w_048_9538, w_048_9540, w_048_9542, w_048_9543, w_048_9544, w_048_9547, w_048_9548, w_048_9550, w_048_9553, w_048_9554, w_048_9555, w_048_9558, w_048_9560, w_048_9562, w_048_9569, w_048_9571, w_048_9574, w_048_9579, w_048_9581, w_048_9583, w_048_9584, w_048_9591, w_048_9593, w_048_9597, w_048_9598, w_048_9604, w_048_9605, w_048_9607, w_048_9611, w_048_9615, w_048_9618, w_048_9623, w_048_9625, w_048_9627, w_048_9629, w_048_9630, w_048_9631, w_048_9633, w_048_9639, w_048_9642, w_048_9644, w_048_9645, w_048_9646, w_048_9647, w_048_9648, w_048_9651, w_048_9652, w_048_9653, w_048_9659, w_048_9663, w_048_9665, w_048_9667, w_048_9669, w_048_9672, w_048_9673, w_048_9674, w_048_9676, w_048_9678, w_048_9679, w_048_9680, w_048_9685, w_048_9686, w_048_9690, w_048_9698, w_048_9701, w_048_9704, w_048_9705, w_048_9708, w_048_9710, w_048_9712, w_048_9714, w_048_9716, w_048_9719, w_048_9720, w_048_9722, w_048_9724, w_048_9726, w_048_9730, w_048_9734, w_048_9737, w_048_9741, w_048_9744, w_048_9745, w_048_9746, w_048_9747, w_048_9749, w_048_9754, w_048_9755, w_048_9757, w_048_9759, w_048_9760, w_048_9761, w_048_9762, w_048_9763, w_048_9767, w_048_9775, w_048_9776, w_048_9777, w_048_9779, w_048_9781, w_048_9784, w_048_9786, w_048_9787, w_048_9789, w_048_9791, w_048_9792, w_048_9793, w_048_9794, w_048_9796, w_048_9801, w_048_9802, w_048_9803, w_048_9806, w_048_9808, w_048_9811, w_048_9816, w_048_9822, w_048_9823, w_048_9825, w_048_9827, w_048_9828, w_048_9829, w_048_9831, w_048_9838, w_048_9841, w_048_9842, w_048_9845, w_048_9848, w_048_9851, w_048_9853, w_048_9854, w_048_9857, w_048_9859, w_048_9860, w_048_9863, w_048_9868, w_048_9871, w_048_9872, w_048_9874, w_048_9878, w_048_9881, w_048_9882, w_048_9886, w_048_9887, w_048_9888, w_048_9889, w_048_9895, w_048_9896, w_048_9900, w_048_9902, w_048_9904, w_048_9906, w_048_9913, w_048_9915;
  wire w_049_000, w_049_001, w_049_002, w_049_003, w_049_004, w_049_005, w_049_006, w_049_007, w_049_008, w_049_009, w_049_010, w_049_011, w_049_012, w_049_013, w_049_014, w_049_015, w_049_016, w_049_017, w_049_018, w_049_019, w_049_020, w_049_021, w_049_022, w_049_023, w_049_024, w_049_025, w_049_026, w_049_027, w_049_028, w_049_029, w_049_030, w_049_031, w_049_032, w_049_033, w_049_034, w_049_035, w_049_036, w_049_037, w_049_038, w_049_039, w_049_040, w_049_041, w_049_042, w_049_043, w_049_044, w_049_045, w_049_046, w_049_047, w_049_048, w_049_049, w_049_050, w_049_051, w_049_052, w_049_053, w_049_054, w_049_055, w_049_056, w_049_057, w_049_058, w_049_059, w_049_060, w_049_061, w_049_062, w_049_063, w_049_064, w_049_065, w_049_066, w_049_067, w_049_068, w_049_070, w_049_071, w_049_072, w_049_073, w_049_074, w_049_075, w_049_076, w_049_077, w_049_078, w_049_079, w_049_080, w_049_081, w_049_082, w_049_083, w_049_084, w_049_085, w_049_086, w_049_087, w_049_088, w_049_089, w_049_090, w_049_091, w_049_092, w_049_093, w_049_094, w_049_095, w_049_096, w_049_097, w_049_098, w_049_099, w_049_100, w_049_101, w_049_102, w_049_103, w_049_104, w_049_105, w_049_106, w_049_107, w_049_108, w_049_109, w_049_110, w_049_111, w_049_112, w_049_114, w_049_115, w_049_116, w_049_117, w_049_118, w_049_119, w_049_120, w_049_121, w_049_122, w_049_123, w_049_124, w_049_125, w_049_126, w_049_127, w_049_128, w_049_129, w_049_130, w_049_131, w_049_132, w_049_133, w_049_134, w_049_135, w_049_136, w_049_137, w_049_138, w_049_139, w_049_140, w_049_141, w_049_142, w_049_143, w_049_144, w_049_145, w_049_146, w_049_148, w_049_149, w_049_150, w_049_151, w_049_152, w_049_153, w_049_154, w_049_155, w_049_156, w_049_157, w_049_158, w_049_159, w_049_161, w_049_162, w_049_163, w_049_164, w_049_165, w_049_166, w_049_167, w_049_168, w_049_169, w_049_170, w_049_171, w_049_172, w_049_173, w_049_175, w_049_176, w_049_177, w_049_178, w_049_179, w_049_180, w_049_181, w_049_182, w_049_183, w_049_184, w_049_185, w_049_186, w_049_187, w_049_189, w_049_190, w_049_191, w_049_192, w_049_193, w_049_194, w_049_195, w_049_196, w_049_197, w_049_198, w_049_199, w_049_201, w_049_202, w_049_203, w_049_204, w_049_205, w_049_206, w_049_207, w_049_208, w_049_209, w_049_210, w_049_211, w_049_212, w_049_213, w_049_214, w_049_215, w_049_216, w_049_217, w_049_218, w_049_219, w_049_220, w_049_221, w_049_222, w_049_223, w_049_224, w_049_225, w_049_226, w_049_227, w_049_228, w_049_229, w_049_230, w_049_231, w_049_232, w_049_233, w_049_234, w_049_235, w_049_236, w_049_237, w_049_238, w_049_239, w_049_240, w_049_241, w_049_242, w_049_243, w_049_244, w_049_245, w_049_246, w_049_247, w_049_248, w_049_249, w_049_250, w_049_252, w_049_253, w_049_254, w_049_255, w_049_256, w_049_257, w_049_258, w_049_259, w_049_260, w_049_261, w_049_262, w_049_263, w_049_264, w_049_265, w_049_266, w_049_267, w_049_268, w_049_269, w_049_270, w_049_271, w_049_272, w_049_273, w_049_274, w_049_275, w_049_276, w_049_277, w_049_278, w_049_279, w_049_280, w_049_281, w_049_282, w_049_283, w_049_284, w_049_286, w_049_287, w_049_288, w_049_289, w_049_290, w_049_291, w_049_292, w_049_293, w_049_294, w_049_295, w_049_296, w_049_297, w_049_298, w_049_299, w_049_300, w_049_301, w_049_302, w_049_303, w_049_304, w_049_305, w_049_306, w_049_307, w_049_308, w_049_309, w_049_310, w_049_311, w_049_312, w_049_313, w_049_314, w_049_315, w_049_316, w_049_317, w_049_318, w_049_319, w_049_320, w_049_321, w_049_322, w_049_323, w_049_324, w_049_325, w_049_326, w_049_328, w_049_329, w_049_330, w_049_331, w_049_332, w_049_333, w_049_334, w_049_335, w_049_336, w_049_337, w_049_338, w_049_339, w_049_340, w_049_341, w_049_342, w_049_343, w_049_344, w_049_345, w_049_346, w_049_347, w_049_348, w_049_349, w_049_350, w_049_351, w_049_352, w_049_353, w_049_354, w_049_355, w_049_356, w_049_357, w_049_358, w_049_359, w_049_360, w_049_361, w_049_362, w_049_364, w_049_365, w_049_366, w_049_367, w_049_368, w_049_369, w_049_370, w_049_371, w_049_372, w_049_373, w_049_374, w_049_375, w_049_376, w_049_377, w_049_378, w_049_379, w_049_380, w_049_381, w_049_382, w_049_383, w_049_384, w_049_385, w_049_386, w_049_387, w_049_388, w_049_389, w_049_390, w_049_391, w_049_392, w_049_394, w_049_395, w_049_396, w_049_397, w_049_398, w_049_399, w_049_400, w_049_401, w_049_402, w_049_403, w_049_404, w_049_405, w_049_406, w_049_407, w_049_408, w_049_409, w_049_410, w_049_411, w_049_412, w_049_413, w_049_414, w_049_415, w_049_416, w_049_417, w_049_418, w_049_419, w_049_420, w_049_421, w_049_422, w_049_423, w_049_424, w_049_425, w_049_427, w_049_428, w_049_429, w_049_430, w_049_431, w_049_432, w_049_433, w_049_434, w_049_435, w_049_436, w_049_437, w_049_438, w_049_439, w_049_440, w_049_441, w_049_442, w_049_443, w_049_444, w_049_445, w_049_446, w_049_447, w_049_448, w_049_449, w_049_450, w_049_451, w_049_452, w_049_453, w_049_454, w_049_455, w_049_456, w_049_457, w_049_458, w_049_459, w_049_460, w_049_461, w_049_462, w_049_463, w_049_464, w_049_465, w_049_466, w_049_467, w_049_468, w_049_469, w_049_470, w_049_471, w_049_472, w_049_473, w_049_474, w_049_475, w_049_476, w_049_477, w_049_478, w_049_480, w_049_481, w_049_482, w_049_483, w_049_484, w_049_485, w_049_486, w_049_487, w_049_488, w_049_489, w_049_490, w_049_491, w_049_492, w_049_493, w_049_494, w_049_495, w_049_496, w_049_497, w_049_498, w_049_499, w_049_500, w_049_501, w_049_502, w_049_503, w_049_504, w_049_505, w_049_506, w_049_507, w_049_508, w_049_509, w_049_510, w_049_511, w_049_512, w_049_513, w_049_514, w_049_515, w_049_516, w_049_517, w_049_518, w_049_519, w_049_520, w_049_521, w_049_522, w_049_523, w_049_524, w_049_525, w_049_526, w_049_527, w_049_528, w_049_529, w_049_530, w_049_531, w_049_532, w_049_534, w_049_535, w_049_536, w_049_537, w_049_538, w_049_539, w_049_540, w_049_541, w_049_542, w_049_543, w_049_544, w_049_545, w_049_546, w_049_547, w_049_548, w_049_549, w_049_550, w_049_551, w_049_552, w_049_553, w_049_554, w_049_555, w_049_556, w_049_557, w_049_558, w_049_559, w_049_560, w_049_561, w_049_562, w_049_563, w_049_564, w_049_565, w_049_566, w_049_567, w_049_568, w_049_569, w_049_570, w_049_571, w_049_572, w_049_574, w_049_575, w_049_576, w_049_577, w_049_578, w_049_579, w_049_580, w_049_581, w_049_582, w_049_583, w_049_584, w_049_585, w_049_586, w_049_587, w_049_588, w_049_589, w_049_590, w_049_591, w_049_592, w_049_593, w_049_594, w_049_595, w_049_596, w_049_597, w_049_598, w_049_599, w_049_601, w_049_602, w_049_603, w_049_604, w_049_605, w_049_608, w_049_609, w_049_610, w_049_611, w_049_613, w_049_614, w_049_615, w_049_616, w_049_617, w_049_618, w_049_619, w_049_620, w_049_621, w_049_622, w_049_623, w_049_624, w_049_625, w_049_626, w_049_627, w_049_628, w_049_629, w_049_630, w_049_631, w_049_632, w_049_634, w_049_635, w_049_636, w_049_637, w_049_638, w_049_639, w_049_640, w_049_641, w_049_642, w_049_643, w_049_644, w_049_645, w_049_646, w_049_647, w_049_648, w_049_649, w_049_650, w_049_651, w_049_652, w_049_653, w_049_654, w_049_655, w_049_656, w_049_657, w_049_658, w_049_659, w_049_660, w_049_661, w_049_662, w_049_663, w_049_664, w_049_665, w_049_666, w_049_667, w_049_668, w_049_669, w_049_670, w_049_671, w_049_672, w_049_673, w_049_674, w_049_675, w_049_676, w_049_677, w_049_678, w_049_680, w_049_681, w_049_682, w_049_683, w_049_684, w_049_685, w_049_686, w_049_687, w_049_688, w_049_689, w_049_691, w_049_692, w_049_693, w_049_694, w_049_695, w_049_696, w_049_697, w_049_698, w_049_699, w_049_700, w_049_701, w_049_702, w_049_703, w_049_704, w_049_705, w_049_706, w_049_707, w_049_708, w_049_709, w_049_710, w_049_711, w_049_712, w_049_713, w_049_714, w_049_716, w_049_717, w_049_718, w_049_719, w_049_720, w_049_721, w_049_722, w_049_723, w_049_724, w_049_725, w_049_726, w_049_727, w_049_728, w_049_729, w_049_730, w_049_731, w_049_732, w_049_733, w_049_734, w_049_735, w_049_736, w_049_737, w_049_738, w_049_739, w_049_740, w_049_741, w_049_742, w_049_743, w_049_744, w_049_746, w_049_747, w_049_749, w_049_750, w_049_751, w_049_752, w_049_753, w_049_754, w_049_755, w_049_756, w_049_757, w_049_758, w_049_759, w_049_760, w_049_761, w_049_762, w_049_763, w_049_764, w_049_765, w_049_766, w_049_767, w_049_769, w_049_771, w_049_772, w_049_773, w_049_774, w_049_775, w_049_777, w_049_778, w_049_779, w_049_780, w_049_781, w_049_782, w_049_783, w_049_784, w_049_785, w_049_786, w_049_788, w_049_790, w_049_791, w_049_793, w_049_794, w_049_795, w_049_796, w_049_797, w_049_798, w_049_799, w_049_800, w_049_801, w_049_802, w_049_803, w_049_804, w_049_805, w_049_806, w_049_807, w_049_808, w_049_809, w_049_810, w_049_811, w_049_812, w_049_813, w_049_814, w_049_815, w_049_816, w_049_817, w_049_818, w_049_819, w_049_820, w_049_821, w_049_822, w_049_823, w_049_825, w_049_826, w_049_828, w_049_829, w_049_830, w_049_831, w_049_832, w_049_833, w_049_834, w_049_835, w_049_836, w_049_837, w_049_838, w_049_839, w_049_840, w_049_841, w_049_842, w_049_843, w_049_844, w_049_845, w_049_846, w_049_847, w_049_848, w_049_849, w_049_850, w_049_851, w_049_852, w_049_853, w_049_854, w_049_856, w_049_857, w_049_858, w_049_859, w_049_860, w_049_861, w_049_862, w_049_863, w_049_864, w_049_865, w_049_866, w_049_867, w_049_868, w_049_869, w_049_870, w_049_871, w_049_872, w_049_873, w_049_874, w_049_875, w_049_876, w_049_877, w_049_878, w_049_879, w_049_880, w_049_881, w_049_882, w_049_883, w_049_884, w_049_885, w_049_887, w_049_888, w_049_889, w_049_890, w_049_891, w_049_892, w_049_893, w_049_894, w_049_895, w_049_896, w_049_897, w_049_898, w_049_899, w_049_900, w_049_901, w_049_902, w_049_903, w_049_904, w_049_905, w_049_906, w_049_907, w_049_908, w_049_909, w_049_910, w_049_911, w_049_912, w_049_913, w_049_914, w_049_915, w_049_916, w_049_917, w_049_918, w_049_919, w_049_920, w_049_921, w_049_922, w_049_923, w_049_924, w_049_925, w_049_926, w_049_927, w_049_928, w_049_929, w_049_930, w_049_931, w_049_932, w_049_933, w_049_934, w_049_935, w_049_936, w_049_937, w_049_938, w_049_939, w_049_940, w_049_941, w_049_942, w_049_943, w_049_944, w_049_945, w_049_946, w_049_947, w_049_948, w_049_949, w_049_950, w_049_951, w_049_952, w_049_953, w_049_954, w_049_955, w_049_956, w_049_957, w_049_958, w_049_959, w_049_960, w_049_961, w_049_962, w_049_963, w_049_964, w_049_965, w_049_966, w_049_967, w_049_969, w_049_970, w_049_971, w_049_972, w_049_973, w_049_974, w_049_975, w_049_976, w_049_977, w_049_978, w_049_979, w_049_980, w_049_981, w_049_982, w_049_983, w_049_984, w_049_985, w_049_986, w_049_987, w_049_988, w_049_989, w_049_990, w_049_991, w_049_992, w_049_993, w_049_994, w_049_995, w_049_996, w_049_997, w_049_998, w_049_999, w_049_1000, w_049_1001, w_049_1002, w_049_1003, w_049_1004, w_049_1005, w_049_1006, w_049_1007, w_049_1008, w_049_1009, w_049_1010, w_049_1011, w_049_1012, w_049_1013, w_049_1014, w_049_1015, w_049_1016, w_049_1017, w_049_1018, w_049_1019, w_049_1020, w_049_1021, w_049_1022, w_049_1023, w_049_1024, w_049_1025, w_049_1026, w_049_1027, w_049_1028, w_049_1029, w_049_1030, w_049_1031, w_049_1032, w_049_1033, w_049_1034, w_049_1035, w_049_1036, w_049_1037, w_049_1038, w_049_1039, w_049_1040, w_049_1041, w_049_1042, w_049_1043, w_049_1044, w_049_1045, w_049_1046, w_049_1047, w_049_1048, w_049_1049, w_049_1050, w_049_1051, w_049_1052, w_049_1053, w_049_1054, w_049_1055, w_049_1056, w_049_1057, w_049_1058, w_049_1059, w_049_1060, w_049_1061, w_049_1062, w_049_1063, w_049_1064, w_049_1065, w_049_1066, w_049_1067, w_049_1068, w_049_1069, w_049_1070, w_049_1071, w_049_1072, w_049_1073, w_049_1074, w_049_1075, w_049_1076, w_049_1077, w_049_1078, w_049_1079, w_049_1080, w_049_1081, w_049_1082, w_049_1083, w_049_1084, w_049_1085, w_049_1087, w_049_1088, w_049_1089, w_049_1090, w_049_1091, w_049_1092, w_049_1093, w_049_1094, w_049_1095, w_049_1096, w_049_1097, w_049_1098, w_049_1099, w_049_1100, w_049_1102, w_049_1103, w_049_1104, w_049_1106, w_049_1107, w_049_1108, w_049_1109, w_049_1110, w_049_1111, w_049_1112, w_049_1113, w_049_1114, w_049_1115, w_049_1116, w_049_1117, w_049_1118, w_049_1119, w_049_1120, w_049_1121, w_049_1122, w_049_1123, w_049_1124, w_049_1125, w_049_1126, w_049_1127, w_049_1128, w_049_1129, w_049_1130, w_049_1131, w_049_1132, w_049_1133, w_049_1134, w_049_1135, w_049_1136, w_049_1137, w_049_1138, w_049_1139, w_049_1140, w_049_1141, w_049_1142, w_049_1143, w_049_1144, w_049_1145, w_049_1146, w_049_1147, w_049_1148, w_049_1150, w_049_1151, w_049_1152, w_049_1153, w_049_1154, w_049_1155, w_049_1156, w_049_1157, w_049_1158, w_049_1159, w_049_1160, w_049_1161, w_049_1162, w_049_1163, w_049_1164, w_049_1165, w_049_1166, w_049_1167, w_049_1168, w_049_1169, w_049_1170, w_049_1171, w_049_1172, w_049_1173, w_049_1174, w_049_1175, w_049_1176, w_049_1177, w_049_1178, w_049_1179, w_049_1180, w_049_1181, w_049_1182, w_049_1183, w_049_1184, w_049_1185, w_049_1186, w_049_1187, w_049_1188, w_049_1189, w_049_1190, w_049_1191, w_049_1192, w_049_1193, w_049_1194, w_049_1195, w_049_1196, w_049_1197, w_049_1198, w_049_1199, w_049_1200, w_049_1201, w_049_1202, w_049_1203, w_049_1204, w_049_1205, w_049_1206, w_049_1207, w_049_1208, w_049_1209, w_049_1210, w_049_1211, w_049_1212, w_049_1213, w_049_1214, w_049_1215, w_049_1217, w_049_1218, w_049_1219, w_049_1220, w_049_1221, w_049_1222, w_049_1223, w_049_1224, w_049_1225, w_049_1226, w_049_1227, w_049_1228, w_049_1229, w_049_1230, w_049_1231, w_049_1232, w_049_1233, w_049_1234, w_049_1235, w_049_1236, w_049_1237, w_049_1238, w_049_1239, w_049_1240, w_049_1241, w_049_1242, w_049_1243, w_049_1244, w_049_1245, w_049_1246, w_049_1247, w_049_1248, w_049_1249, w_049_1250, w_049_1251, w_049_1252, w_049_1253, w_049_1254, w_049_1255, w_049_1256, w_049_1257, w_049_1258, w_049_1259, w_049_1261, w_049_1262, w_049_1263, w_049_1264, w_049_1265, w_049_1266, w_049_1267, w_049_1268, w_049_1269, w_049_1270, w_049_1272, w_049_1273, w_049_1274, w_049_1275, w_049_1276, w_049_1277, w_049_1278, w_049_1279, w_049_1281, w_049_1282, w_049_1283, w_049_1284, w_049_1285, w_049_1286, w_049_1287, w_049_1288, w_049_1289, w_049_1290, w_049_1291, w_049_1292, w_049_1293, w_049_1294, w_049_1295, w_049_1296, w_049_1297, w_049_1298, w_049_1299, w_049_1300, w_049_1301, w_049_1302, w_049_1303, w_049_1304, w_049_1305, w_049_1306, w_049_1307, w_049_1308, w_049_1309, w_049_1310, w_049_1311, w_049_1312, w_049_1313, w_049_1314, w_049_1315, w_049_1316, w_049_1317, w_049_1318, w_049_1319, w_049_1320, w_049_1321, w_049_1322, w_049_1323, w_049_1324, w_049_1325, w_049_1326, w_049_1327, w_049_1328, w_049_1329, w_049_1330, w_049_1331, w_049_1332, w_049_1333, w_049_1334, w_049_1335, w_049_1336, w_049_1337, w_049_1338, w_049_1339, w_049_1340, w_049_1341, w_049_1342, w_049_1343, w_049_1344, w_049_1345, w_049_1346, w_049_1347, w_049_1348, w_049_1349, w_049_1350, w_049_1351, w_049_1352, w_049_1353, w_049_1354, w_049_1355, w_049_1356, w_049_1357, w_049_1358, w_049_1359, w_049_1360, w_049_1361, w_049_1362, w_049_1363, w_049_1364, w_049_1365, w_049_1366, w_049_1367, w_049_1368, w_049_1369, w_049_1370, w_049_1371, w_049_1372, w_049_1373, w_049_1374, w_049_1375, w_049_1376, w_049_1377, w_049_1378, w_049_1379, w_049_1380, w_049_1381, w_049_1382, w_049_1383, w_049_1384, w_049_1385, w_049_1386, w_049_1387, w_049_1388, w_049_1389, w_049_1390, w_049_1391, w_049_1392, w_049_1393, w_049_1394, w_049_1395, w_049_1396, w_049_1397, w_049_1398, w_049_1399, w_049_1400, w_049_1401, w_049_1402, w_049_1403, w_049_1404, w_049_1405, w_049_1406, w_049_1407, w_049_1408, w_049_1409, w_049_1410, w_049_1411, w_049_1412, w_049_1413, w_049_1414, w_049_1415, w_049_1416, w_049_1417, w_049_1418, w_049_1419, w_049_1420, w_049_1421, w_049_1422, w_049_1423, w_049_1424, w_049_1426, w_049_1427, w_049_1428, w_049_1429, w_049_1430, w_049_1431, w_049_1432, w_049_1433, w_049_1434, w_049_1435, w_049_1436, w_049_1437, w_049_1438, w_049_1440, w_049_1441, w_049_1442, w_049_1443, w_049_1444, w_049_1445, w_049_1446, w_049_1447, w_049_1448, w_049_1449, w_049_1450, w_049_1451, w_049_1452, w_049_1453, w_049_1454, w_049_1455, w_049_1456, w_049_1457, w_049_1458, w_049_1459, w_049_1460, w_049_1461, w_049_1462, w_049_1463, w_049_1464, w_049_1465, w_049_1466, w_049_1467, w_049_1468, w_049_1469, w_049_1470, w_049_1471, w_049_1472, w_049_1473, w_049_1474, w_049_1475, w_049_1476, w_049_1477, w_049_1478, w_049_1479, w_049_1480, w_049_1481, w_049_1482, w_049_1483, w_049_1484, w_049_1485, w_049_1486, w_049_1487, w_049_1488, w_049_1489, w_049_1490, w_049_1491, w_049_1492, w_049_1493, w_049_1494, w_049_1495, w_049_1496, w_049_1497, w_049_1498, w_049_1499, w_049_1500, w_049_1501, w_049_1502, w_049_1503, w_049_1504, w_049_1505, w_049_1506, w_049_1507, w_049_1508, w_049_1509, w_049_1510, w_049_1511, w_049_1512, w_049_1513, w_049_1514, w_049_1515, w_049_1516, w_049_1517, w_049_1518, w_049_1520, w_049_1521, w_049_1522, w_049_1523, w_049_1524, w_049_1525, w_049_1526, w_049_1527, w_049_1528, w_049_1529, w_049_1530, w_049_1531, w_049_1532, w_049_1533, w_049_1534, w_049_1535, w_049_1536, w_049_1537, w_049_1538, w_049_1539, w_049_1540, w_049_1541, w_049_1542, w_049_1543, w_049_1544, w_049_1545, w_049_1546, w_049_1547, w_049_1548, w_049_1549, w_049_1550, w_049_1551, w_049_1552, w_049_1553, w_049_1554, w_049_1555, w_049_1556, w_049_1557, w_049_1558, w_049_1559, w_049_1560, w_049_1561, w_049_1562, w_049_1563, w_049_1564, w_049_1565, w_049_1566, w_049_1567, w_049_1568, w_049_1569, w_049_1570, w_049_1571, w_049_1572, w_049_1573, w_049_1574, w_049_1575, w_049_1576, w_049_1577, w_049_1578, w_049_1579, w_049_1580, w_049_1581, w_049_1582, w_049_1583, w_049_1584, w_049_1585, w_049_1586, w_049_1587, w_049_1588, w_049_1589, w_049_1590, w_049_1591, w_049_1592, w_049_1593, w_049_1594, w_049_1595, w_049_1596, w_049_1597, w_049_1598, w_049_1599, w_049_1600, w_049_1601, w_049_1602, w_049_1603, w_049_1604, w_049_1605, w_049_1606, w_049_1607, w_049_1608, w_049_1609, w_049_1610, w_049_1611, w_049_1612, w_049_1613, w_049_1614, w_049_1615, w_049_1616, w_049_1617, w_049_1618, w_049_1619, w_049_1620, w_049_1621, w_049_1622, w_049_1623, w_049_1624, w_049_1625, w_049_1626, w_049_1627, w_049_1628, w_049_1629, w_049_1630, w_049_1631, w_049_1632, w_049_1634, w_049_1635, w_049_1636, w_049_1637, w_049_1638, w_049_1639, w_049_1641, w_049_1642, w_049_1643, w_049_1644, w_049_1645, w_049_1646, w_049_1647, w_049_1648, w_049_1649, w_049_1650, w_049_1651, w_049_1652, w_049_1653, w_049_1654, w_049_1655, w_049_1656, w_049_1657, w_049_1658, w_049_1659, w_049_1660, w_049_1661, w_049_1662, w_049_1663, w_049_1664, w_049_1665, w_049_1666, w_049_1667, w_049_1668, w_049_1669, w_049_1670, w_049_1671, w_049_1672, w_049_1673, w_049_1674, w_049_1675, w_049_1676, w_049_1677, w_049_1678, w_049_1679;
  wire w_050_000, w_050_001, w_050_002, w_050_004, w_050_005, w_050_006, w_050_008, w_050_009, w_050_010, w_050_011, w_050_014, w_050_015, w_050_016, w_050_020, w_050_024, w_050_026, w_050_027, w_050_028, w_050_029, w_050_031, w_050_035, w_050_036, w_050_038, w_050_040, w_050_041, w_050_042, w_050_046, w_050_048, w_050_049, w_050_050, w_050_051, w_050_053, w_050_054, w_050_056, w_050_057, w_050_058, w_050_060, w_050_065, w_050_066, w_050_067, w_050_068, w_050_075, w_050_076, w_050_077, w_050_078, w_050_079, w_050_080, w_050_083, w_050_085, w_050_086, w_050_087, w_050_088, w_050_090, w_050_091, w_050_093, w_050_095, w_050_096, w_050_098, w_050_099, w_050_100, w_050_102, w_050_103, w_050_104, w_050_105, w_050_108, w_050_109, w_050_110, w_050_111, w_050_113, w_050_114, w_050_115, w_050_116, w_050_118, w_050_119, w_050_120, w_050_122, w_050_125, w_050_126, w_050_128, w_050_129, w_050_132, w_050_133, w_050_134, w_050_135, w_050_136, w_050_137, w_050_138, w_050_141, w_050_143, w_050_144, w_050_145, w_050_146, w_050_148, w_050_150, w_050_151, w_050_152, w_050_153, w_050_155, w_050_160, w_050_161, w_050_162, w_050_163, w_050_164, w_050_165, w_050_166, w_050_167, w_050_170, w_050_171, w_050_172, w_050_173, w_050_174, w_050_176, w_050_177, w_050_179, w_050_182, w_050_183, w_050_184, w_050_189, w_050_190, w_050_191, w_050_192, w_050_193, w_050_195, w_050_197, w_050_199, w_050_201, w_050_202, w_050_203, w_050_204, w_050_207, w_050_208, w_050_209, w_050_210, w_050_211, w_050_212, w_050_213, w_050_215, w_050_216, w_050_217, w_050_218, w_050_219, w_050_221, w_050_222, w_050_224, w_050_226, w_050_227, w_050_228, w_050_230, w_050_231, w_050_232, w_050_234, w_050_235, w_050_236, w_050_237, w_050_239, w_050_240, w_050_241, w_050_244, w_050_245, w_050_246, w_050_247, w_050_249, w_050_252, w_050_253, w_050_254, w_050_255, w_050_256, w_050_257, w_050_258, w_050_260, w_050_261, w_050_263, w_050_264, w_050_265, w_050_266, w_050_267, w_050_269, w_050_270, w_050_272, w_050_273, w_050_275, w_050_276, w_050_278, w_050_279, w_050_280, w_050_281, w_050_283, w_050_284, w_050_285, w_050_289, w_050_291, w_050_294, w_050_295, w_050_296, w_050_297, w_050_299, w_050_300, w_050_301, w_050_302, w_050_304, w_050_305, w_050_306, w_050_307, w_050_308, w_050_311, w_050_312, w_050_316, w_050_317, w_050_318, w_050_320, w_050_321, w_050_323, w_050_324, w_050_325, w_050_328, w_050_330, w_050_331, w_050_333, w_050_334, w_050_336, w_050_337, w_050_339, w_050_343, w_050_344, w_050_346, w_050_348, w_050_349, w_050_352, w_050_356, w_050_357, w_050_359, w_050_362, w_050_363, w_050_364, w_050_365, w_050_367, w_050_369, w_050_370, w_050_372, w_050_374, w_050_375, w_050_376, w_050_386, w_050_388, w_050_389, w_050_391, w_050_393, w_050_394, w_050_395, w_050_396, w_050_397, w_050_398, w_050_399, w_050_401, w_050_403, w_050_404, w_050_405, w_050_406, w_050_407, w_050_408, w_050_410, w_050_411, w_050_412, w_050_414, w_050_416, w_050_417, w_050_419, w_050_420, w_050_421, w_050_423, w_050_424, w_050_427, w_050_428, w_050_429, w_050_430, w_050_431, w_050_435, w_050_436, w_050_440, w_050_441, w_050_442, w_050_443, w_050_444, w_050_447, w_050_448, w_050_449, w_050_450, w_050_451, w_050_453, w_050_454, w_050_455, w_050_456, w_050_457, w_050_458, w_050_459, w_050_460, w_050_462, w_050_463, w_050_464, w_050_465, w_050_466, w_050_468, w_050_469, w_050_471, w_050_472, w_050_473, w_050_474, w_050_475, w_050_478, w_050_481, w_050_482, w_050_484, w_050_485, w_050_486, w_050_488, w_050_490, w_050_491, w_050_495, w_050_497, w_050_498, w_050_500, w_050_502, w_050_504, w_050_505, w_050_506, w_050_507, w_050_508, w_050_509, w_050_510, w_050_512, w_050_513, w_050_516, w_050_518, w_050_519, w_050_520, w_050_522, w_050_523, w_050_524, w_050_527, w_050_528, w_050_529, w_050_531, w_050_532, w_050_533, w_050_534, w_050_536, w_050_538, w_050_539, w_050_540, w_050_541, w_050_543, w_050_544, w_050_546, w_050_547, w_050_548, w_050_549, w_050_550, w_050_554, w_050_557, w_050_560, w_050_561, w_050_562, w_050_563, w_050_564, w_050_566, w_050_569, w_050_571, w_050_572, w_050_575, w_050_577, w_050_579, w_050_580, w_050_581, w_050_582, w_050_584, w_050_586, w_050_587, w_050_589, w_050_590, w_050_591, w_050_592, w_050_595, w_050_596, w_050_597, w_050_599, w_050_600, w_050_602, w_050_603, w_050_605, w_050_607, w_050_608, w_050_609, w_050_611, w_050_614, w_050_615, w_050_616, w_050_617, w_050_618, w_050_619, w_050_620, w_050_621, w_050_623, w_050_628, w_050_630, w_050_631, w_050_634, w_050_635, w_050_636, w_050_637, w_050_638, w_050_639, w_050_640, w_050_641, w_050_642, w_050_643, w_050_644, w_050_645, w_050_646, w_050_647, w_050_648, w_050_649, w_050_651, w_050_652, w_050_653, w_050_654, w_050_655, w_050_656, w_050_658, w_050_660, w_050_662, w_050_664, w_050_668, w_050_670, w_050_671, w_050_672, w_050_673, w_050_674, w_050_675, w_050_676, w_050_678, w_050_682, w_050_683, w_050_684, w_050_687, w_050_689, w_050_691, w_050_693, w_050_694, w_050_695, w_050_696, w_050_698, w_050_700, w_050_704, w_050_705, w_050_706, w_050_707, w_050_711, w_050_712, w_050_713, w_050_715, w_050_718, w_050_719, w_050_720, w_050_722, w_050_723, w_050_724, w_050_725, w_050_726, w_050_727, w_050_729, w_050_730, w_050_731, w_050_732, w_050_733, w_050_734, w_050_735, w_050_736, w_050_737, w_050_739, w_050_741, w_050_742, w_050_743, w_050_747, w_050_748, w_050_749, w_050_750, w_050_751, w_050_752, w_050_753, w_050_754, w_050_756, w_050_757, w_050_758, w_050_759, w_050_761, w_050_762, w_050_764, w_050_766, w_050_767, w_050_770, w_050_771, w_050_772, w_050_773, w_050_777, w_050_778, w_050_779, w_050_780, w_050_782, w_050_783, w_050_785, w_050_787, w_050_788, w_050_791, w_050_793, w_050_794, w_050_795, w_050_796, w_050_799, w_050_800, w_050_802, w_050_806, w_050_807, w_050_808, w_050_811, w_050_812, w_050_814, w_050_816, w_050_818, w_050_819, w_050_820, w_050_821, w_050_823, w_050_826, w_050_828, w_050_829, w_050_830, w_050_831, w_050_832, w_050_835, w_050_838, w_050_839, w_050_842, w_050_843, w_050_844, w_050_845, w_050_848, w_050_851, w_050_855, w_050_856, w_050_857, w_050_860, w_050_862, w_050_863, w_050_864, w_050_865, w_050_867, w_050_868, w_050_871, w_050_872, w_050_873, w_050_875, w_050_877, w_050_878, w_050_879, w_050_880, w_050_882, w_050_884, w_050_885, w_050_886, w_050_887, w_050_891, w_050_894, w_050_895, w_050_896, w_050_899, w_050_900, w_050_901, w_050_902, w_050_903, w_050_907, w_050_908, w_050_909, w_050_911, w_050_912, w_050_914, w_050_915, w_050_916, w_050_917, w_050_918, w_050_920, w_050_921, w_050_923, w_050_925, w_050_926, w_050_927, w_050_928, w_050_929, w_050_931, w_050_934, w_050_936, w_050_937, w_050_938, w_050_940, w_050_942, w_050_943, w_050_944, w_050_946, w_050_947, w_050_950, w_050_951, w_050_952, w_050_953, w_050_955, w_050_956, w_050_957, w_050_958, w_050_961, w_050_962, w_050_963, w_050_964, w_050_966, w_050_968, w_050_969, w_050_970, w_050_971, w_050_972, w_050_973, w_050_974, w_050_975, w_050_976, w_050_977, w_050_979, w_050_980, w_050_981, w_050_982, w_050_983, w_050_985, w_050_987, w_050_988, w_050_989, w_050_990, w_050_992, w_050_993, w_050_995, w_050_996, w_050_998, w_050_1000, w_050_1001, w_050_1002, w_050_1003, w_050_1004, w_050_1005, w_050_1006, w_050_1007, w_050_1010, w_050_1011, w_050_1012, w_050_1013, w_050_1014, w_050_1015, w_050_1016, w_050_1020, w_050_1023, w_050_1024, w_050_1025, w_050_1026, w_050_1028, w_050_1029, w_050_1032, w_050_1033, w_050_1035, w_050_1036, w_050_1037, w_050_1041, w_050_1042, w_050_1043, w_050_1044, w_050_1045, w_050_1046, w_050_1047, w_050_1048, w_050_1050, w_050_1051, w_050_1054, w_050_1056, w_050_1057, w_050_1058, w_050_1062, w_050_1063, w_050_1067, w_050_1068, w_050_1069, w_050_1072, w_050_1074, w_050_1077, w_050_1078, w_050_1079, w_050_1080, w_050_1084, w_050_1086, w_050_1091, w_050_1094, w_050_1095, w_050_1097, w_050_1098, w_050_1102, w_050_1107, w_050_1108, w_050_1109, w_050_1114, w_050_1116, w_050_1119, w_050_1122, w_050_1123, w_050_1124, w_050_1126, w_050_1129, w_050_1131, w_050_1132, w_050_1133, w_050_1135, w_050_1136, w_050_1138, w_050_1139, w_050_1140, w_050_1141, w_050_1143, w_050_1145, w_050_1146, w_050_1147, w_050_1148, w_050_1149, w_050_1150, w_050_1151, w_050_1152, w_050_1153, w_050_1154, w_050_1158, w_050_1159, w_050_1160, w_050_1165, w_050_1167, w_050_1168, w_050_1169, w_050_1170, w_050_1172, w_050_1175, w_050_1176, w_050_1177, w_050_1178, w_050_1179, w_050_1180, w_050_1182, w_050_1183, w_050_1186, w_050_1188, w_050_1189, w_050_1190, w_050_1191, w_050_1192, w_050_1193, w_050_1194, w_050_1196, w_050_1198, w_050_1201, w_050_1202, w_050_1203, w_050_1204, w_050_1208, w_050_1209, w_050_1212, w_050_1213, w_050_1217, w_050_1218, w_050_1219, w_050_1220, w_050_1221, w_050_1224, w_050_1225, w_050_1229, w_050_1230, w_050_1232, w_050_1233, w_050_1235, w_050_1236, w_050_1238, w_050_1239, w_050_1240, w_050_1241, w_050_1243, w_050_1244, w_050_1247, w_050_1249, w_050_1252, w_050_1253, w_050_1255, w_050_1256, w_050_1260, w_050_1261, w_050_1262, w_050_1263, w_050_1265, w_050_1266, w_050_1269, w_050_1273, w_050_1274, w_050_1275, w_050_1276, w_050_1277, w_050_1279, w_050_1280, w_050_1281, w_050_1282, w_050_1284, w_050_1285, w_050_1287, w_050_1288, w_050_1289, w_050_1290, w_050_1291, w_050_1292, w_050_1293, w_050_1294, w_050_1295, w_050_1296, w_050_1297, w_050_1300, w_050_1304, w_050_1305, w_050_1306, w_050_1307, w_050_1308, w_050_1309, w_050_1311, w_050_1313, w_050_1314, w_050_1315, w_050_1316, w_050_1318, w_050_1319, w_050_1323, w_050_1324, w_050_1325, w_050_1329, w_050_1330, w_050_1332, w_050_1333, w_050_1335, w_050_1338, w_050_1339, w_050_1341, w_050_1342, w_050_1343, w_050_1346, w_050_1347, w_050_1351, w_050_1352, w_050_1353, w_050_1354, w_050_1355, w_050_1356, w_050_1357, w_050_1359, w_050_1360, w_050_1361, w_050_1363, w_050_1365, w_050_1366, w_050_1367, w_050_1368, w_050_1369, w_050_1372, w_050_1373, w_050_1374, w_050_1375, w_050_1376, w_050_1377, w_050_1378, w_050_1379, w_050_1382, w_050_1383, w_050_1384, w_050_1385, w_050_1387, w_050_1390, w_050_1391, w_050_1392, w_050_1395, w_050_1398, w_050_1399, w_050_1400, w_050_1402, w_050_1403, w_050_1404, w_050_1405, w_050_1407, w_050_1408, w_050_1410, w_050_1412, w_050_1413, w_050_1414, w_050_1417, w_050_1419, w_050_1421, w_050_1422, w_050_1423, w_050_1424, w_050_1425, w_050_1426, w_050_1427, w_050_1428, w_050_1429, w_050_1431, w_050_1432, w_050_1433, w_050_1434, w_050_1436, w_050_1439, w_050_1440, w_050_1441, w_050_1443, w_050_1444, w_050_1445, w_050_1447, w_050_1448, w_050_1450, w_050_1452, w_050_1453, w_050_1454, w_050_1455, w_050_1456, w_050_1457, w_050_1459, w_050_1462, w_050_1464, w_050_1465, w_050_1466, w_050_1468, w_050_1469, w_050_1470, w_050_1472, w_050_1473, w_050_1475, w_050_1477, w_050_1480, w_050_1481, w_050_1483, w_050_1484, w_050_1485, w_050_1486, w_050_1487, w_050_1488, w_050_1491, w_050_1493, w_050_1494, w_050_1495, w_050_1497, w_050_1499, w_050_1500, w_050_1501, w_050_1503, w_050_1507, w_050_1508, w_050_1509, w_050_1510, w_050_1511, w_050_1512, w_050_1513, w_050_1514, w_050_1515, w_050_1516, w_050_1517, w_050_1518, w_050_1520, w_050_1521, w_050_1522, w_050_1523, w_050_1524, w_050_1525, w_050_1526, w_050_1527, w_050_1529, w_050_1530, w_050_1531, w_050_1532, w_050_1534, w_050_1535, w_050_1536, w_050_1537, w_050_1538, w_050_1544, w_050_1546, w_050_1547, w_050_1549, w_050_1550, w_050_1551, w_050_1552, w_050_1554, w_050_1555, w_050_1556, w_050_1558, w_050_1559, w_050_1561, w_050_1562, w_050_1563, w_050_1564, w_050_1565, w_050_1566, w_050_1568, w_050_1569, w_050_1571, w_050_1572, w_050_1574, w_050_1575, w_050_1576, w_050_1578, w_050_1580, w_050_1582, w_050_1584, w_050_1586, w_050_1588, w_050_1590, w_050_1591, w_050_1592, w_050_1593, w_050_1594, w_050_1596, w_050_1600, w_050_1601, w_050_1602, w_050_1604, w_050_1605, w_050_1606, w_050_1608, w_050_1609, w_050_1610, w_050_1612, w_050_1613, w_050_1614, w_050_1615, w_050_1618, w_050_1620, w_050_1621, w_050_1623, w_050_1624, w_050_1625, w_050_1626, w_050_1627, w_050_1632, w_050_1633, w_050_1634, w_050_1636, w_050_1637, w_050_1638, w_050_1640, w_050_1646, w_050_1647, w_050_1648, w_050_1649, w_050_1652, w_050_1654, w_050_1655, w_050_1656, w_050_1658, w_050_1659, w_050_1660, w_050_1662, w_050_1664, w_050_1667, w_050_1668, w_050_1669, w_050_1672, w_050_1673, w_050_1674, w_050_1678, w_050_1679, w_050_1682, w_050_1683, w_050_1685, w_050_1686, w_050_1687, w_050_1689, w_050_1690, w_050_1692, w_050_1693, w_050_1694, w_050_1695, w_050_1697, w_050_1698, w_050_1700, w_050_1701, w_050_1703, w_050_1704, w_050_1705, w_050_1706, w_050_1707, w_050_1708, w_050_1709, w_050_1710, w_050_1711, w_050_1713, w_050_1714, w_050_1715, w_050_1719, w_050_1720, w_050_1722, w_050_1723, w_050_1724, w_050_1725, w_050_1726, w_050_1728, w_050_1729, w_050_1730, w_050_1731, w_050_1732, w_050_1733, w_050_1734, w_050_1735, w_050_1736, w_050_1737, w_050_1738, w_050_1739, w_050_1740, w_050_1742, w_050_1743, w_050_1744, w_050_1745, w_050_1746, w_050_1747, w_050_1750, w_050_1751, w_050_1754, w_050_1755, w_050_1756, w_050_1757, w_050_1759, w_050_1760, w_050_1761, w_050_1762, w_050_1763, w_050_1764, w_050_1766, w_050_1767, w_050_1768, w_050_1769, w_050_1772, w_050_1773, w_050_1774, w_050_1775, w_050_1776, w_050_1777, w_050_1778, w_050_1781, w_050_1782, w_050_1783, w_050_1785, w_050_1786, w_050_1788, w_050_1789, w_050_1790, w_050_1791, w_050_1792, w_050_1797, w_050_1799, w_050_1801, w_050_1802, w_050_1803, w_050_1804, w_050_1805, w_050_1808, w_050_1809, w_050_1811, w_050_1812, w_050_1814, w_050_1815, w_050_1816, w_050_1818, w_050_1819, w_050_1821, w_050_1822, w_050_1823, w_050_1826, w_050_1829, w_050_1830, w_050_1834, w_050_1839, w_050_1840, w_050_1841, w_050_1843, w_050_1845, w_050_1847, w_050_1848, w_050_1849, w_050_1850, w_050_1851, w_050_1852, w_050_1853, w_050_1854, w_050_1861, w_050_1862, w_050_1865, w_050_1868, w_050_1869, w_050_1870, w_050_1872, w_050_1873, w_050_1874, w_050_1880, w_050_1881, w_050_1882, w_050_1883, w_050_1884, w_050_1885, w_050_1887, w_050_1888, w_050_1890, w_050_1891, w_050_1892, w_050_1893, w_050_1894, w_050_1895, w_050_1896, w_050_1898, w_050_1899, w_050_1900, w_050_1902, w_050_1903, w_050_1905, w_050_1906, w_050_1910, w_050_1911, w_050_1912, w_050_1913, w_050_1914, w_050_1915, w_050_1916, w_050_1919, w_050_1920, w_050_1921, w_050_1922, w_050_1923, w_050_1927, w_050_1929, w_050_1930, w_050_1931, w_050_1932, w_050_1933, w_050_1934, w_050_1935, w_050_1936, w_050_1938, w_050_1939, w_050_1941, w_050_1943, w_050_1944, w_050_1945, w_050_1946, w_050_1947, w_050_1948, w_050_1949, w_050_1953, w_050_1957, w_050_1958, w_050_1959, w_050_1960, w_050_1962, w_050_1963, w_050_1965, w_050_1967, w_050_1968, w_050_1970, w_050_1972, w_050_1973, w_050_1975, w_050_1976, w_050_1977, w_050_1978, w_050_1979, w_050_1980, w_050_1982, w_050_1983, w_050_1984, w_050_1985, w_050_1987, w_050_1988, w_050_1989, w_050_1990, w_050_1991, w_050_1992, w_050_1993, w_050_1994, w_050_1995, w_050_1996, w_050_1997, w_050_2001, w_050_2002, w_050_2004, w_050_2005, w_050_2006, w_050_2009, w_050_2012, w_050_2013, w_050_2016, w_050_2018, w_050_2019, w_050_2021, w_050_2022, w_050_2023, w_050_2024, w_050_2025, w_050_2026, w_050_2027, w_050_2028, w_050_2030, w_050_2032, w_050_2033, w_050_2035, w_050_2036, w_050_2039, w_050_2042, w_050_2043, w_050_2045, w_050_2046, w_050_2047, w_050_2048, w_050_2049, w_050_2051, w_050_2053, w_050_2054, w_050_2056, w_050_2057, w_050_2058, w_050_2059, w_050_2064, w_050_2066, w_050_2068, w_050_2070, w_050_2072, w_050_2078, w_050_2080, w_050_2081, w_050_2082, w_050_2083, w_050_2084, w_050_2085, w_050_2088, w_050_2090, w_050_2091, w_050_2094, w_050_2095, w_050_2096, w_050_2097, w_050_2098, w_050_2101, w_050_2103, w_050_2104, w_050_2105, w_050_2106, w_050_2107, w_050_2109, w_050_2110, w_050_2111, w_050_2113, w_050_2114, w_050_2115, w_050_2116, w_050_2117, w_050_2118, w_050_2121, w_050_2122, w_050_2123, w_050_2125, w_050_2126, w_050_2127, w_050_2133, w_050_2134, w_050_2137, w_050_2139, w_050_2140, w_050_2141, w_050_2143, w_050_2144, w_050_2145, w_050_2146, w_050_2147, w_050_2148, w_050_2150, w_050_2151, w_050_2153, w_050_2154, w_050_2156, w_050_2157, w_050_2158, w_050_2160, w_050_2161, w_050_2162, w_050_2164, w_050_2165, w_050_2166, w_050_2167, w_050_2168, w_050_2173, w_050_2176, w_050_2182, w_050_2184, w_050_2185, w_050_2188, w_050_2190, w_050_2191, w_050_2192, w_050_2195, w_050_2197, w_050_2198, w_050_2201, w_050_2203, w_050_2204, w_050_2206, w_050_2207, w_050_2208, w_050_2209, w_050_2210, w_050_2214, w_050_2216, w_050_2217, w_050_2219, w_050_2221, w_050_2222, w_050_2224, w_050_2225, w_050_2226, w_050_2228, w_050_2229, w_050_2231, w_050_2232, w_050_2235, w_050_2236, w_050_2237, w_050_2238, w_050_2239, w_050_2243, w_050_2244, w_050_2246, w_050_2247, w_050_2252, w_050_2253, w_050_2254, w_050_2256, w_050_2257, w_050_2258, w_050_2260, w_050_2262, w_050_2263, w_050_2267, w_050_2268, w_050_2271, w_050_2272, w_050_2274, w_050_2275, w_050_2276, w_050_2278, w_050_2280, w_050_2281, w_050_2282, w_050_2285, w_050_2287, w_050_2288, w_050_2289, w_050_2290, w_050_2291, w_050_2292, w_050_2293, w_050_2295, w_050_2296, w_050_2297, w_050_2298, w_050_2300, w_050_2301, w_050_2302, w_050_2306, w_050_2307, w_050_2310, w_050_2311, w_050_2313, w_050_2316, w_050_2318, w_050_2319, w_050_2320, w_050_2321, w_050_2322, w_050_2323, w_050_2326, w_050_2329, w_050_2330, w_050_2332, w_050_2333, w_050_2334, w_050_2335, w_050_2337, w_050_2339, w_050_2341, w_050_2342, w_050_2343, w_050_2344, w_050_2345, w_050_2347, w_050_2348, w_050_2349, w_050_2351, w_050_2352, w_050_2353, w_050_2355, w_050_2356, w_050_2357, w_050_2358, w_050_2359, w_050_2360, w_050_2362, w_050_2364, w_050_2365, w_050_2368, w_050_2371, w_050_2373, w_050_2374, w_050_2375, w_050_2376, w_050_2379, w_050_2380, w_050_2381, w_050_2383, w_050_2384, w_050_2385, w_050_2386, w_050_2387, w_050_2388, w_050_2392, w_050_2393, w_050_2396, w_050_2398, w_050_2399, w_050_2402, w_050_2403, w_050_2404, w_050_2405, w_050_2406, w_050_2408, w_050_2409, w_050_2411, w_050_2412, w_050_2413, w_050_2414, w_050_2415, w_050_2417, w_050_2419, w_050_2421, w_050_2423, w_050_2424, w_050_2429, w_050_2430, w_050_2431, w_050_2432, w_050_2434, w_050_2438, w_050_2439, w_050_2442, w_050_2443, w_050_2444, w_050_2445, w_050_2446, w_050_2451, w_050_2453, w_050_2454, w_050_2457, w_050_2458, w_050_2461, w_050_2462, w_050_2463, w_050_2464, w_050_2465, w_050_2466, w_050_2468, w_050_2469, w_050_2471, w_050_2473, w_050_2474, w_050_2477, w_050_2478, w_050_2479, w_050_2480, w_050_2481, w_050_2482, w_050_2485, w_050_2486, w_050_2487, w_050_2488, w_050_2489, w_050_2491, w_050_2492, w_050_2493, w_050_2494, w_050_2498, w_050_2501, w_050_2502, w_050_2503, w_050_2504, w_050_2508, w_050_2511, w_050_2513, w_050_2515, w_050_2516, w_050_2517, w_050_2519, w_050_2520, w_050_2521, w_050_2522, w_050_2526, w_050_2527, w_050_2528, w_050_2530, w_050_2531, w_050_2533, w_050_2534, w_050_2536, w_050_2537, w_050_2539, w_050_2540, w_050_2541, w_050_2542, w_050_2543, w_050_2544, w_050_2545, w_050_2546, w_050_2547, w_050_2548, w_050_2550, w_050_2551, w_050_2553, w_050_2554, w_050_2556, w_050_2557, w_050_2558, w_050_2560, w_050_2561, w_050_2562, w_050_2565, w_050_2566, w_050_2567, w_050_2570, w_050_2571, w_050_2572, w_050_2574, w_050_2576, w_050_2577, w_050_2580, w_050_2581, w_050_2582, w_050_2584, w_050_2585, w_050_2586, w_050_2588, w_050_2589, w_050_2591, w_050_2592, w_050_2594, w_050_2595, w_050_2597, w_050_2598, w_050_2599, w_050_2600, w_050_2602, w_050_2603, w_050_2606, w_050_2609, w_050_2610, w_050_2612, w_050_2614, w_050_2615, w_050_2617, w_050_2618, w_050_2619, w_050_2622, w_050_2623, w_050_2627, w_050_2628, w_050_2629, w_050_2630, w_050_2631, w_050_2633, w_050_2634, w_050_2636, w_050_2639, w_050_2641, w_050_2646, w_050_2648, w_050_2649, w_050_2650, w_050_2651, w_050_2653, w_050_2654, w_050_2655, w_050_2658, w_050_2659, w_050_2660, w_050_2662, w_050_2663, w_050_2665, w_050_2668, w_050_2669, w_050_2670, w_050_2671, w_050_2672, w_050_2675, w_050_2676, w_050_2678, w_050_2679, w_050_2680, w_050_2681, w_050_2682, w_050_2684, w_050_2685, w_050_2686, w_050_2688, w_050_2692, w_050_2693, w_050_2695, w_050_2696, w_050_2697, w_050_2698, w_050_2700, w_050_2701, w_050_2702, w_050_2703, w_050_2704, w_050_2705, w_050_2706, w_050_2709, w_050_2711, w_050_2712, w_050_2714, w_050_2715, w_050_2723, w_050_2724, w_050_2725, w_050_2727, w_050_2728, w_050_2729, w_050_2732, w_050_2734, w_050_2735, w_050_2736, w_050_2737, w_050_2738, w_050_2739, w_050_2740, w_050_2741, w_050_2742, w_050_2743, w_050_2744, w_050_2755, w_050_2756, w_050_2757, w_050_2760, w_050_2761, w_050_2762, w_050_2764, w_050_2765, w_050_2767, w_050_2768, w_050_2769, w_050_2770, w_050_2771, w_050_2772, w_050_2773, w_050_2774, w_050_2776, w_050_2778, w_050_2779, w_050_2780, w_050_2781, w_050_2782, w_050_2783, w_050_2784, w_050_2787, w_050_2788, w_050_2789, w_050_2790, w_050_2791, w_050_2792, w_050_2794, w_050_2795, w_050_2796, w_050_2797, w_050_2799, w_050_2800, w_050_2801, w_050_2802, w_050_2803, w_050_2804, w_050_2809, w_050_2811, w_050_2812, w_050_2813, w_050_2814, w_050_2816, w_050_2817, w_050_2818, w_050_2822, w_050_2823, w_050_2824, w_050_2825, w_050_2826, w_050_2828, w_050_2829, w_050_2831, w_050_2832, w_050_2833, w_050_2835, w_050_2836, w_050_2837, w_050_2839, w_050_2840, w_050_2841, w_050_2842, w_050_2843, w_050_2844, w_050_2845, w_050_2847, w_050_2848, w_050_2851, w_050_2852, w_050_2855, w_050_2856, w_050_2857, w_050_2860, w_050_2862, w_050_2864, w_050_2870, w_050_2871, w_050_2872, w_050_2874, w_050_2875, w_050_2877, w_050_2878, w_050_2879, w_050_2883, w_050_2884, w_050_2885, w_050_2886, w_050_2887, w_050_2889, w_050_2891, w_050_2892, w_050_2893, w_050_2894, w_050_2900, w_050_2901, w_050_2903, w_050_2905, w_050_2906, w_050_2907, w_050_2908, w_050_2910, w_050_2911, w_050_2913, w_050_2917, w_050_2918, w_050_2920, w_050_2922, w_050_2923, w_050_2926, w_050_2927, w_050_2929, w_050_2930, w_050_2932, w_050_2933, w_050_2934, w_050_2935, w_050_2938, w_050_2939, w_050_2941, w_050_2942, w_050_2943, w_050_2944, w_050_2945, w_050_2947, w_050_2948, w_050_2950, w_050_2951, w_050_2952, w_050_2954, w_050_2955, w_050_2957, w_050_2958, w_050_2959, w_050_2961, w_050_2963, w_050_2964, w_050_2965, w_050_2966, w_050_2970, w_050_2972, w_050_2975, w_050_2976, w_050_2979, w_050_2980, w_050_2981, w_050_2982, w_050_2983, w_050_2984, w_050_2985, w_050_2986, w_050_2987, w_050_2988, w_050_2989, w_050_2990, w_050_2991, w_050_2992, w_050_2994, w_050_2996, w_050_2997, w_050_2999, w_050_3001, w_050_3002, w_050_3004, w_050_3006, w_050_3007, w_050_3008, w_050_3009, w_050_3011, w_050_3014, w_050_3016, w_050_3020, w_050_3021, w_050_3025, w_050_3026, w_050_3027, w_050_3028, w_050_3029, w_050_3031, w_050_3032, w_050_3033, w_050_3034, w_050_3037, w_050_3038, w_050_3040, w_050_3041, w_050_3043, w_050_3045, w_050_3047, w_050_3049, w_050_3051, w_050_3052, w_050_3053, w_050_3055, w_050_3056, w_050_3057, w_050_3059, w_050_3060, w_050_3061, w_050_3062, w_050_3063, w_050_3069, w_050_3070, w_050_3071, w_050_3072, w_050_3075, w_050_3076, w_050_3078, w_050_3079, w_050_3080, w_050_3083, w_050_3088, w_050_3089, w_050_3090, w_050_3091, w_050_3093, w_050_3094, w_050_3095, w_050_3096, w_050_3098, w_050_3099, w_050_3100, w_050_3101, w_050_3104, w_050_3105, w_050_3106, w_050_3107, w_050_3108, w_050_3111, w_050_3112, w_050_3113, w_050_3116, w_050_3118, w_050_3119, w_050_3120, w_050_3121, w_050_3122, w_050_3125, w_050_3126, w_050_3127, w_050_3128, w_050_3129, w_050_3130, w_050_3131, w_050_3133, w_050_3134, w_050_3138, w_050_3139, w_050_3142, w_050_3145, w_050_3146, w_050_3148, w_050_3149, w_050_3150, w_050_3151, w_050_3154, w_050_3156, w_050_3157, w_050_3159, w_050_3160, w_050_3161, w_050_3162, w_050_3163, w_050_3164, w_050_3168, w_050_3169, w_050_3170, w_050_3171, w_050_3172, w_050_3173, w_050_3175, w_050_3178, w_050_3179, w_050_3181, w_050_3187, w_050_3188, w_050_3191, w_050_3192, w_050_3194, w_050_3195, w_050_3196, w_050_3197, w_050_3198, w_050_3199, w_050_3200, w_050_3201, w_050_3203, w_050_3205, w_050_3206, w_050_3207, w_050_3209, w_050_3212, w_050_3213, w_050_3214, w_050_3215, w_050_3216, w_050_3218, w_050_3219, w_050_3221, w_050_3223, w_050_3224, w_050_3226, w_050_3227, w_050_3229, w_050_3230, w_050_3231, w_050_3234, w_050_3237, w_050_3238, w_050_3240, w_050_3241, w_050_3243, w_050_3244, w_050_3246, w_050_3247, w_050_3248, w_050_3249, w_050_3254, w_050_3255, w_050_3258, w_050_3262, w_050_3263, w_050_3265, w_050_3266, w_050_3268, w_050_3269, w_050_3270, w_050_3272, w_050_3273, w_050_3274, w_050_3275, w_050_3278, w_050_3279, w_050_3280, w_050_3281, w_050_3282, w_050_3283, w_050_3284, w_050_3285, w_050_3288, w_050_3293, w_050_3294, w_050_3295, w_050_3296, w_050_3298, w_050_3299, w_050_3300, w_050_3301, w_050_3303, w_050_3304, w_050_3306, w_050_3310, w_050_3311, w_050_3313, w_050_3314, w_050_3318, w_050_3319, w_050_3320, w_050_3322, w_050_3323, w_050_3325, w_050_3329, w_050_3331, w_050_3332, w_050_3333, w_050_3334, w_050_3335, w_050_3336, w_050_3340, w_050_3341, w_050_3342, w_050_3345, w_050_3346, w_050_3347, w_050_3348, w_050_3350, w_050_3352, w_050_3353, w_050_3354, w_050_3356, w_050_3357, w_050_3363, w_050_3364, w_050_3368, w_050_3369, w_050_3370, w_050_3371, w_050_3372, w_050_3373, w_050_3377, w_050_3378, w_050_3379, w_050_3381, w_050_3382, w_050_3385, w_050_3389, w_050_3391, w_050_3393, w_050_3394, w_050_3396, w_050_3397, w_050_3398, w_050_3399, w_050_3401, w_050_3403, w_050_3404, w_050_3405, w_050_3406, w_050_3407, w_050_3408, w_050_3409, w_050_3410, w_050_3411, w_050_3413, w_050_3414, w_050_3415, w_050_3417, w_050_3418, w_050_3420, w_050_3421, w_050_3423, w_050_3425, w_050_3429, w_050_3430, w_050_3431, w_050_3432, w_050_3434, w_050_3437, w_050_3439, w_050_3440, w_050_3441, w_050_3444, w_050_3445, w_050_3446, w_050_3447, w_050_3450, w_050_3452, w_050_3453, w_050_3454, w_050_3459, w_050_3462, w_050_3463, w_050_3464, w_050_3465, w_050_3466, w_050_3468, w_050_3470, w_050_3471, w_050_3473, w_050_3475, w_050_3476, w_050_3478, w_050_3479, w_050_3480, w_050_3481, w_050_3483, w_050_3487, w_050_3489, w_050_3493, w_050_3499, w_050_3500, w_050_3503, w_050_3505, w_050_3511, w_050_3513, w_050_3514, w_050_3517, w_050_3521, w_050_3526, w_050_3528, w_050_3529, w_050_3530, w_050_3533, w_050_3535, w_050_3538, w_050_3540, w_050_3544, w_050_3545, w_050_3546, w_050_3549, w_050_3554, w_050_3560, w_050_3563, w_050_3564, w_050_3565, w_050_3567, w_050_3569, w_050_3570, w_050_3574, w_050_3575, w_050_3577, w_050_3587, w_050_3589, w_050_3591, w_050_3598, w_050_3599, w_050_3600, w_050_3604, w_050_3608, w_050_3609, w_050_3612, w_050_3613, w_050_3615, w_050_3617, w_050_3618, w_050_3620, w_050_3622, w_050_3630, w_050_3631, w_050_3632, w_050_3638, w_050_3640, w_050_3641, w_050_3645, w_050_3646, w_050_3647, w_050_3649, w_050_3652, w_050_3653, w_050_3657, w_050_3659, w_050_3660, w_050_3661, w_050_3665, w_050_3666, w_050_3668, w_050_3671, w_050_3672, w_050_3673, w_050_3674, w_050_3681, w_050_3683, w_050_3686, w_050_3690, w_050_3691, w_050_3694, w_050_3695, w_050_3698, w_050_3701, w_050_3702, w_050_3703, w_050_3705, w_050_3706, w_050_3710, w_050_3714, w_050_3715, w_050_3717, w_050_3719, w_050_3721, w_050_3728, w_050_3732, w_050_3733, w_050_3735, w_050_3737, w_050_3740, w_050_3746, w_050_3748, w_050_3749, w_050_3752, w_050_3757, w_050_3759, w_050_3761, w_050_3766, w_050_3767, w_050_3770, w_050_3773, w_050_3774, w_050_3776, w_050_3777, w_050_3778, w_050_3781, w_050_3784, w_050_3786, w_050_3788, w_050_3789, w_050_3798, w_050_3799, w_050_3806, w_050_3810, w_050_3811, w_050_3813, w_050_3816, w_050_3819, w_050_3821, w_050_3824, w_050_3828, w_050_3829, w_050_3830, w_050_3831, w_050_3833, w_050_3834, w_050_3837, w_050_3839, w_050_3840, w_050_3841, w_050_3844, w_050_3845, w_050_3853, w_050_3857, w_050_3858, w_050_3859, w_050_3860, w_050_3866, w_050_3867, w_050_3869, w_050_3870, w_050_3883, w_050_3889, w_050_3890, w_050_3892, w_050_3895, w_050_3896, w_050_3898, w_050_3900, w_050_3903, w_050_3905, w_050_3912, w_050_3913, w_050_3919, w_050_3921, w_050_3923, w_050_3925, w_050_3930, w_050_3934, w_050_3936, w_050_3942, w_050_3945, w_050_3946, w_050_3947, w_050_3949, w_050_3950, w_050_3955, w_050_3957, w_050_3958, w_050_3959, w_050_3963, w_050_3966, w_050_3969, w_050_3973, w_050_3975, w_050_3976, w_050_3983, w_050_3984, w_050_3985, w_050_3988, w_050_3990, w_050_3992, w_050_3993, w_050_3994, w_050_3997, w_050_3999, w_050_4000, w_050_4001, w_050_4003, w_050_4004, w_050_4005, w_050_4006, w_050_4008, w_050_4009, w_050_4010, w_050_4011, w_050_4013, w_050_4026, w_050_4030, w_050_4033, w_050_4036, w_050_4038, w_050_4039, w_050_4040, w_050_4042, w_050_4043, w_050_4045, w_050_4049, w_050_4050, w_050_4052, w_050_4053, w_050_4056, w_050_4057, w_050_4058, w_050_4059, w_050_4062, w_050_4065, w_050_4067, w_050_4070, w_050_4071, w_050_4073, w_050_4074, w_050_4075, w_050_4081, w_050_4082, w_050_4083, w_050_4085, w_050_4087, w_050_4092, w_050_4096, w_050_4097, w_050_4100, w_050_4106, w_050_4108, w_050_4109, w_050_4113, w_050_4115, w_050_4116, w_050_4119, w_050_4123, w_050_4126, w_050_4127, w_050_4128, w_050_4129, w_050_4131, w_050_4133, w_050_4134, w_050_4139, w_050_4140, w_050_4141, w_050_4144, w_050_4145, w_050_4146, w_050_4149, w_050_4150, w_050_4152, w_050_4153, w_050_4154, w_050_4157, w_050_4160, w_050_4162, w_050_4164, w_050_4165, w_050_4170, w_050_4172, w_050_4173, w_050_4174, w_050_4179, w_050_4186, w_050_4191, w_050_4192, w_050_4193, w_050_4195, w_050_4196, w_050_4197, w_050_4201, w_050_4204, w_050_4206, w_050_4207, w_050_4210, w_050_4211, w_050_4215, w_050_4217, w_050_4218, w_050_4219, w_050_4220, w_050_4221, w_050_4222, w_050_4223, w_050_4224, w_050_4229, w_050_4233, w_050_4234, w_050_4235, w_050_4236, w_050_4238, w_050_4239, w_050_4244, w_050_4245, w_050_4246, w_050_4247, w_050_4249, w_050_4250, w_050_4251, w_050_4253, w_050_4255, w_050_4256, w_050_4259, w_050_4260, w_050_4263, w_050_4267, w_050_4271, w_050_4272, w_050_4283, w_050_4285, w_050_4287, w_050_4288, w_050_4292, w_050_4298, w_050_4301, w_050_4303, w_050_4306, w_050_4309, w_050_4310, w_050_4312, w_050_4315, w_050_4316, w_050_4321, w_050_4324, w_050_4329, w_050_4333, w_050_4339, w_050_4340, w_050_4341, w_050_4342, w_050_4343, w_050_4348, w_050_4350, w_050_4351, w_050_4354, w_050_4355, w_050_4358, w_050_4359, w_050_4361, w_050_4363, w_050_4366, w_050_4368, w_050_4371, w_050_4373, w_050_4374, w_050_4375, w_050_4379, w_050_4392, w_050_4395, w_050_4397, w_050_4406, w_050_4407, w_050_4409, w_050_4412, w_050_4414, w_050_4418, w_050_4422, w_050_4424, w_050_4427, w_050_4428, w_050_4431, w_050_4433, w_050_4435, w_050_4441, w_050_4445, w_050_4446, w_050_4448, w_050_4449, w_050_4450, w_050_4451, w_050_4454, w_050_4455, w_050_4458, w_050_4459, w_050_4460, w_050_4463, w_050_4467, w_050_4470, w_050_4472, w_050_4474, w_050_4476, w_050_4480, w_050_4485, w_050_4486, w_050_4487, w_050_4488, w_050_4491, w_050_4494, w_050_4495, w_050_4496, w_050_4498, w_050_4500, w_050_4502, w_050_4507, w_050_4515, w_050_4517, w_050_4520, w_050_4522, w_050_4524, w_050_4525, w_050_4526, w_050_4527, w_050_4528, w_050_4532, w_050_4533, w_050_4534, w_050_4539, w_050_4540, w_050_4541, w_050_4543, w_050_4544, w_050_4547, w_050_4548, w_050_4549, w_050_4550, w_050_4551, w_050_4552, w_050_4553, w_050_4554, w_050_4555, w_050_4556, w_050_4557, w_050_4562, w_050_4563, w_050_4566, w_050_4567, w_050_4568, w_050_4570, w_050_4571, w_050_4572, w_050_4574, w_050_4577, w_050_4581, w_050_4582, w_050_4583, w_050_4589, w_050_4590, w_050_4592, w_050_4597, w_050_4598, w_050_4602, w_050_4604, w_050_4609, w_050_4611, w_050_4612, w_050_4615, w_050_4617, w_050_4619, w_050_4620, w_050_4622, w_050_4631, w_050_4635, w_050_4636, w_050_4639, w_050_4641, w_050_4642, w_050_4644, w_050_4645, w_050_4647, w_050_4650, w_050_4651, w_050_4652, w_050_4653, w_050_4654, w_050_4655, w_050_4664, w_050_4666, w_050_4667, w_050_4671, w_050_4675, w_050_4676, w_050_4678, w_050_4685, w_050_4690, w_050_4691, w_050_4693, w_050_4694, w_050_4695, w_050_4696, w_050_4701, w_050_4707, w_050_4716, w_050_4723, w_050_4725, w_050_4726, w_050_4728, w_050_4729, w_050_4732, w_050_4735, w_050_4738, w_050_4739, w_050_4742, w_050_4746, w_050_4751, w_050_4754, w_050_4755, w_050_4757, w_050_4759, w_050_4761, w_050_4762, w_050_4763, w_050_4766, w_050_4773, w_050_4774, w_050_4775, w_050_4780, w_050_4782, w_050_4784, w_050_4785, w_050_4786, w_050_4789, w_050_4791, w_050_4796, w_050_4798, w_050_4801, w_050_4802, w_050_4811, w_050_4816, w_050_4818, w_050_4819, w_050_4822, w_050_4824, w_050_4825, w_050_4826, w_050_4827, w_050_4829, w_050_4830, w_050_4831, w_050_4836, w_050_4837, w_050_4838, w_050_4839, w_050_4843, w_050_4844, w_050_4846, w_050_4847, w_050_4851, w_050_4853, w_050_4854, w_050_4856, w_050_4862, w_050_4864, w_050_4865, w_050_4866, w_050_4868, w_050_4870, w_050_4872, w_050_4874, w_050_4875, w_050_4877, w_050_4878, w_050_4879, w_050_4880, w_050_4882, w_050_4886, w_050_4887, w_050_4888, w_050_4889, w_050_4890, w_050_4892, w_050_4893, w_050_4895, w_050_4896, w_050_4900, w_050_4901, w_050_4902, w_050_4903, w_050_4906, w_050_4907, w_050_4912, w_050_4918, w_050_4919, w_050_4921, w_050_4923, w_050_4924, w_050_4925, w_050_4927, w_050_4928, w_050_4930, w_050_4933, w_050_4937, w_050_4940, w_050_4941, w_050_4946, w_050_4951, w_050_4953, w_050_4954, w_050_4955, w_050_4959, w_050_4960, w_050_4961, w_050_4965, w_050_4970, w_050_4971, w_050_4974, w_050_4975, w_050_4976, w_050_4978, w_050_4979, w_050_4981, w_050_4983, w_050_4984, w_050_4992, w_050_4993, w_050_4998, w_050_5000, w_050_5002, w_050_5003, w_050_5005, w_050_5007, w_050_5009, w_050_5014, w_050_5018, w_050_5020, w_050_5021, w_050_5022, w_050_5027, w_050_5031, w_050_5032, w_050_5036, w_050_5038, w_050_5039, w_050_5040, w_050_5042, w_050_5044, w_050_5045, w_050_5048, w_050_5049, w_050_5051, w_050_5054, w_050_5057, w_050_5061, w_050_5067, w_050_5069, w_050_5072, w_050_5074, w_050_5078, w_050_5080, w_050_5081, w_050_5084, w_050_5086, w_050_5087, w_050_5088, w_050_5089, w_050_5091, w_050_5092, w_050_5093, w_050_5095, w_050_5096, w_050_5097, w_050_5100, w_050_5102, w_050_5105, w_050_5106, w_050_5109, w_050_5113, w_050_5114, w_050_5115, w_050_5118, w_050_5119, w_050_5120, w_050_5121, w_050_5123, w_050_5126, w_050_5138, w_050_5139, w_050_5143, w_050_5144, w_050_5145, w_050_5147, w_050_5149, w_050_5151, w_050_5152, w_050_5153, w_050_5154, w_050_5156, w_050_5157, w_050_5159, w_050_5161, w_050_5163, w_050_5167, w_050_5168, w_050_5181, w_050_5182, w_050_5187, w_050_5188, w_050_5189, w_050_5191, w_050_5192, w_050_5194, w_050_5196, w_050_5202, w_050_5204, w_050_5205, w_050_5207, w_050_5208, w_050_5209, w_050_5210, w_050_5213, w_050_5219, w_050_5221, w_050_5223, w_050_5225, w_050_5226, w_050_5231, w_050_5234, w_050_5235, w_050_5238, w_050_5239, w_050_5240, w_050_5245, w_050_5250, w_050_5253, w_050_5255, w_050_5260, w_050_5262, w_050_5268, w_050_5272, w_050_5276, w_050_5280, w_050_5281, w_050_5283, w_050_5286, w_050_5288, w_050_5290, w_050_5295, w_050_5297, w_050_5299, w_050_5300, w_050_5304, w_050_5307, w_050_5308, w_050_5309, w_050_5311, w_050_5313, w_050_5314, w_050_5315, w_050_5317, w_050_5319, w_050_5322, w_050_5333, w_050_5335, w_050_5336, w_050_5339, w_050_5340, w_050_5341, w_050_5342, w_050_5343, w_050_5347, w_050_5351, w_050_5352, w_050_5353, w_050_5356, w_050_5357, w_050_5364, w_050_5365, w_050_5366, w_050_5370, w_050_5374, w_050_5377, w_050_5380, w_050_5382, w_050_5384, w_050_5386, w_050_5387, w_050_5388, w_050_5389, w_050_5392, w_050_5393, w_050_5395, w_050_5396, w_050_5399, w_050_5400, w_050_5401, w_050_5402, w_050_5405, w_050_5407, w_050_5409, w_050_5412, w_050_5421, w_050_5422, w_050_5431, w_050_5436, w_050_5437, w_050_5438, w_050_5439, w_050_5440, w_050_5443, w_050_5446, w_050_5449, w_050_5450, w_050_5458, w_050_5459, w_050_5460, w_050_5470, w_050_5476, w_050_5485, w_050_5487, w_050_5488, w_050_5489, w_050_5490, w_050_5496, w_050_5497, w_050_5498, w_050_5503, w_050_5509, w_050_5512, w_050_5520, w_050_5521, w_050_5522, w_050_5524, w_050_5527, w_050_5528, w_050_5531, w_050_5534, w_050_5537, w_050_5538, w_050_5541, w_050_5542, w_050_5543, w_050_5544, w_050_5550, w_050_5551, w_050_5555, w_050_5557, w_050_5564, w_050_5565, w_050_5566, w_050_5567, w_050_5568, w_050_5572, w_050_5574, w_050_5575, w_050_5576, w_050_5577, w_050_5580, w_050_5582, w_050_5583, w_050_5584, w_050_5589, w_050_5591, w_050_5592, w_050_5594, w_050_5595, w_050_5599, w_050_5600, w_050_5602, w_050_5603, w_050_5608, w_050_5611, w_050_5612, w_050_5613, w_050_5617, w_050_5618, w_050_5621, w_050_5623, w_050_5627, w_050_5628, w_050_5629, w_050_5630, w_050_5631, w_050_5633, w_050_5637, w_050_5640, w_050_5643, w_050_5645, w_050_5647, w_050_5648, w_050_5649, w_050_5651, w_050_5652, w_050_5656, w_050_5657, w_050_5659, w_050_5662, w_050_5664, w_050_5665, w_050_5668, w_050_5669, w_050_5672, w_050_5673, w_050_5674, w_050_5675, w_050_5678, w_050_5680, w_050_5684, w_050_5685, w_050_5688, w_050_5690, w_050_5693, w_050_5694, w_050_5695, w_050_5697, w_050_5701, w_050_5703, w_050_5705, w_050_5706, w_050_5707, w_050_5709, w_050_5710, w_050_5711, w_050_5714, w_050_5715, w_050_5716, w_050_5717, w_050_5718, w_050_5720, w_050_5722, w_050_5725, w_050_5729, w_050_5732, w_050_5733, w_050_5734, w_050_5735, w_050_5738, w_050_5741, w_050_5742, w_050_5743, w_050_5745, w_050_5751, w_050_5757, w_050_5758, w_050_5761, w_050_5763, w_050_5766, w_050_5771, w_050_5773, w_050_5774, w_050_5775, w_050_5776, w_050_5778, w_050_5779, w_050_5780, w_050_5782, w_050_5783, w_050_5787, w_050_5791, w_050_5795, w_050_5796, w_050_5801, w_050_5803, w_050_5804, w_050_5805, w_050_5806, w_050_5807, w_050_5810, w_050_5812, w_050_5813, w_050_5814, w_050_5818, w_050_5821, w_050_5822, w_050_5824, w_050_5825, w_050_5828, w_050_5832, w_050_5833, w_050_5838, w_050_5839, w_050_5842, w_050_5844, w_050_5845, w_050_5847, w_050_5849, w_050_5857, w_050_5860, w_050_5862, w_050_5863, w_050_5864, w_050_5865, w_050_5867, w_050_5868, w_050_5869, w_050_5870, w_050_5874, w_050_5875, w_050_5877, w_050_5878, w_050_5880, w_050_5888, w_050_5889, w_050_5890, w_050_5891, w_050_5892, w_050_5894, w_050_5897, w_050_5899, w_050_5903, w_050_5904, w_050_5905, w_050_5907, w_050_5910, w_050_5911, w_050_5913, w_050_5918, w_050_5919, w_050_5921, w_050_5922, w_050_5924, w_050_5925, w_050_5930, w_050_5933, w_050_5934, w_050_5939, w_050_5940, w_050_5942, w_050_5943, w_050_5945, w_050_5946, w_050_5948, w_050_5953, w_050_5955, w_050_5957, w_050_5964, w_050_5965, w_050_5967, w_050_5968, w_050_5969, w_050_5970, w_050_5972, w_050_5977, w_050_5980, w_050_5981, w_050_5988, w_050_5991, w_050_5992, w_050_5993, w_050_5998, w_050_6000, w_050_6001, w_050_6004, w_050_6006, w_050_6009, w_050_6011, w_050_6012, w_050_6013, w_050_6015, w_050_6016, w_050_6017, w_050_6018, w_050_6020, w_050_6021, w_050_6022, w_050_6023, w_050_6026, w_050_6027, w_050_6028, w_050_6030, w_050_6033, w_050_6035, w_050_6037, w_050_6038, w_050_6039, w_050_6044, w_050_6046, w_050_6048, w_050_6051, w_050_6052, w_050_6055, w_050_6056, w_050_6057, w_050_6060, w_050_6061, w_050_6062, w_050_6063, w_050_6065, w_050_6066, w_050_6072, w_050_6082, w_050_6087, w_050_6090, w_050_6091, w_050_6096, w_050_6099, w_050_6100, w_050_6102, w_050_6106, w_050_6107, w_050_6113, w_050_6114, w_050_6117, w_050_6118, w_050_6119, w_050_6122, w_050_6126, w_050_6130, w_050_6133, w_050_6135, w_050_6138, w_050_6141, w_050_6142, w_050_6145, w_050_6146, w_050_6148, w_050_6151, w_050_6152, w_050_6153, w_050_6155, w_050_6156, w_050_6158, w_050_6159, w_050_6160, w_050_6161, w_050_6162, w_050_6163, w_050_6175, w_050_6181, w_050_6182, w_050_6183, w_050_6185, w_050_6186, w_050_6188, w_050_6190, w_050_6192, w_050_6193, w_050_6194, w_050_6197, w_050_6202, w_050_6203, w_050_6205, w_050_6206, w_050_6207, w_050_6208, w_050_6210, w_050_6212, w_050_6215, w_050_6216, w_050_6219, w_050_6223, w_050_6225, w_050_6226, w_050_6230, w_050_6231, w_050_6232, w_050_6235, w_050_6236, w_050_6237, w_050_6238, w_050_6239, w_050_6240, w_050_6244, w_050_6248, w_050_6250, w_050_6251, w_050_6255, w_050_6256, w_050_6259, w_050_6261, w_050_6264, w_050_6266, w_050_6269, w_050_6274, w_050_6277, w_050_6278, w_050_6282, w_050_6284, w_050_6285, w_050_6288, w_050_6289, w_050_6290, w_050_6292, w_050_6296, w_050_6298, w_050_6299, w_050_6302, w_050_6304, w_050_6305, w_050_6310, w_050_6312, w_050_6313, w_050_6316, w_050_6317, w_050_6318, w_050_6319, w_050_6322, w_050_6325, w_050_6329, w_050_6331, w_050_6333, w_050_6335, w_050_6337, w_050_6339, w_050_6343, w_050_6348, w_050_6349, w_050_6350, w_050_6351, w_050_6352, w_050_6353, w_050_6356, w_050_6364, w_050_6368, w_050_6372, w_050_6377, w_050_6378, w_050_6380, w_050_6381, w_050_6382, w_050_6383, w_050_6384, w_050_6391, w_050_6392, w_050_6401, w_050_6403, w_050_6408, w_050_6409, w_050_6410, w_050_6412, w_050_6413, w_050_6415, w_050_6418, w_050_6419, w_050_6424, w_050_6425, w_050_6426, w_050_6427, w_050_6428, w_050_6434, w_050_6435, w_050_6436, w_050_6437, w_050_6438, w_050_6439, w_050_6442, w_050_6443, w_050_6447, w_050_6451, w_050_6461, w_050_6462, w_050_6464, w_050_6467, w_050_6468, w_050_6469, w_050_6471, w_050_6472, w_050_6473, w_050_6478, w_050_6479, w_050_6495, w_050_6496, w_050_6498, w_050_6499, w_050_6502, w_050_6503, w_050_6505, w_050_6507, w_050_6512, w_050_6515;
  wire w_051_000, w_051_001, w_051_002, w_051_003, w_051_004, w_051_005, w_051_006, w_051_007, w_051_011, w_051_012, w_051_014, w_051_015, w_051_016, w_051_017, w_051_020, w_051_021, w_051_024, w_051_026, w_051_028, w_051_029, w_051_030, w_051_031, w_051_032, w_051_033, w_051_036, w_051_037, w_051_038, w_051_039, w_051_040, w_051_042, w_051_043, w_051_044, w_051_045, w_051_046, w_051_047, w_051_050, w_051_052, w_051_053, w_051_057, w_051_058, w_051_059, w_051_061, w_051_062, w_051_063, w_051_064, w_051_065, w_051_066, w_051_067, w_051_068, w_051_069, w_051_070, w_051_074, w_051_076, w_051_077, w_051_078, w_051_080, w_051_084, w_051_085, w_051_086, w_051_089, w_051_090, w_051_091, w_051_093, w_051_095, w_051_097, w_051_098, w_051_100, w_051_101, w_051_104, w_051_106, w_051_107, w_051_109, w_051_112, w_051_114, w_051_115, w_051_116, w_051_119, w_051_122, w_051_123, w_051_125, w_051_127, w_051_128, w_051_130, w_051_131, w_051_133, w_051_134, w_051_135, w_051_136, w_051_140, w_051_142, w_051_143, w_051_146, w_051_147, w_051_148, w_051_149, w_051_151, w_051_152, w_051_155, w_051_157, w_051_159, w_051_160, w_051_161, w_051_162, w_051_163, w_051_164, w_051_167, w_051_168, w_051_169, w_051_171, w_051_172, w_051_173, w_051_174, w_051_176, w_051_177, w_051_181, w_051_182, w_051_183, w_051_185, w_051_187, w_051_189, w_051_190, w_051_191, w_051_192, w_051_195, w_051_196, w_051_200, w_051_201, w_051_202, w_051_204, w_051_206, w_051_209, w_051_210, w_051_213, w_051_214, w_051_216, w_051_217, w_051_219, w_051_220, w_051_222, w_051_223, w_051_225, w_051_226, w_051_227, w_051_228, w_051_230, w_051_231, w_051_234, w_051_236, w_051_237, w_051_238, w_051_239, w_051_241, w_051_243, w_051_244, w_051_245, w_051_246, w_051_247, w_051_249, w_051_252, w_051_254, w_051_255, w_051_256, w_051_257, w_051_259, w_051_260, w_051_263, w_051_264, w_051_266, w_051_267, w_051_269, w_051_271, w_051_272, w_051_273, w_051_274, w_051_275, w_051_276, w_051_279, w_051_280, w_051_281, w_051_283, w_051_285, w_051_286, w_051_287, w_051_288, w_051_290, w_051_291, w_051_293, w_051_295, w_051_297, w_051_299, w_051_300, w_051_301, w_051_304, w_051_305, w_051_306, w_051_307, w_051_308, w_051_309, w_051_310, w_051_311, w_051_312, w_051_313, w_051_314, w_051_316, w_051_317, w_051_318, w_051_319, w_051_321, w_051_322, w_051_323, w_051_324, w_051_325, w_051_327, w_051_328, w_051_329, w_051_333, w_051_334, w_051_336, w_051_337, w_051_338, w_051_339, w_051_340, w_051_341, w_051_344, w_051_345, w_051_346, w_051_347, w_051_348, w_051_349, w_051_351, w_051_352, w_051_353, w_051_354, w_051_356, w_051_357, w_051_359, w_051_360, w_051_362, w_051_363, w_051_365, w_051_367, w_051_368, w_051_370, w_051_371, w_051_372, w_051_373, w_051_374, w_051_376, w_051_377, w_051_378, w_051_380, w_051_382, w_051_383, w_051_384, w_051_385, w_051_386, w_051_387, w_051_388, w_051_389, w_051_390, w_051_391, w_051_392, w_051_394, w_051_395, w_051_396, w_051_397, w_051_398, w_051_399, w_051_401, w_051_402, w_051_403, w_051_405, w_051_406, w_051_407, w_051_408, w_051_409, w_051_411, w_051_412, w_051_413, w_051_414, w_051_415, w_051_416, w_051_417, w_051_418, w_051_421, w_051_422, w_051_424, w_051_425, w_051_426, w_051_427, w_051_428, w_051_429, w_051_430, w_051_432, w_051_435, w_051_436, w_051_438, w_051_439, w_051_441, w_051_442, w_051_444, w_051_445, w_051_449, w_051_450, w_051_451, w_051_452, w_051_453, w_051_455, w_051_460, w_051_462, w_051_463, w_051_465, w_051_466, w_051_467, w_051_468, w_051_471, w_051_472, w_051_473, w_051_476, w_051_477, w_051_478, w_051_479, w_051_483, w_051_484, w_051_485, w_051_486, w_051_488, w_051_489, w_051_490, w_051_496, w_051_498, w_051_499, w_051_503, w_051_504, w_051_506, w_051_509, w_051_510, w_051_511, w_051_513, w_051_514, w_051_516, w_051_517, w_051_520, w_051_522, w_051_523, w_051_524, w_051_525, w_051_526, w_051_528, w_051_529, w_051_530, w_051_538, w_051_542, w_051_544, w_051_547, w_051_550, w_051_551, w_051_552, w_051_557, w_051_558, w_051_559, w_051_561, w_051_563, w_051_564, w_051_568, w_051_570, w_051_571, w_051_572, w_051_573, w_051_574, w_051_578, w_051_579, w_051_580, w_051_582, w_051_583, w_051_584, w_051_585, w_051_586, w_051_587, w_051_588, w_051_589, w_051_591, w_051_592, w_051_595, w_051_596, w_051_600, w_051_601, w_051_603, w_051_604, w_051_606, w_051_607, w_051_609, w_051_610, w_051_612, w_051_613, w_051_614, w_051_615, w_051_616, w_051_617, w_051_619, w_051_620, w_051_621, w_051_622, w_051_623, w_051_624, w_051_625, w_051_626, w_051_627, w_051_628, w_051_630, w_051_631, w_051_632, w_051_633, w_051_635, w_051_637, w_051_638, w_051_641, w_051_643, w_051_646, w_051_648, w_051_649, w_051_650, w_051_651, w_051_652, w_051_653, w_051_654, w_051_655, w_051_656, w_051_657, w_051_658, w_051_659, w_051_660, w_051_661, w_051_662, w_051_663, w_051_665, w_051_666, w_051_667, w_051_668, w_051_669, w_051_670, w_051_671, w_051_674, w_051_675, w_051_676, w_051_677, w_051_679, w_051_680, w_051_681, w_051_682, w_051_683, w_051_684, w_051_685, w_051_686, w_051_687, w_051_688, w_051_690, w_051_692, w_051_693, w_051_694, w_051_695, w_051_697, w_051_698, w_051_699, w_051_700, w_051_702, w_051_703, w_051_705, w_051_706, w_051_708, w_051_709, w_051_712, w_051_714, w_051_715, w_051_716, w_051_717, w_051_720, w_051_722, w_051_725, w_051_726, w_051_728, w_051_730, w_051_731, w_051_732, w_051_733, w_051_734, w_051_735, w_051_738, w_051_741, w_051_742, w_051_744, w_051_745, w_051_746, w_051_747, w_051_749, w_051_750, w_051_752, w_051_753, w_051_754, w_051_755, w_051_756, w_051_757, w_051_759, w_051_762, w_051_763, w_051_764, w_051_767, w_051_769, w_051_770, w_051_771, w_051_773, w_051_774, w_051_775, w_051_776, w_051_777, w_051_778, w_051_779, w_051_780, w_051_781, w_051_783, w_051_784, w_051_785, w_051_786, w_051_791, w_051_792, w_051_793, w_051_794, w_051_797, w_051_799, w_051_800, w_051_801, w_051_802, w_051_806, w_051_807, w_051_809, w_051_810, w_051_812, w_051_813, w_051_814, w_051_815, w_051_817, w_051_820, w_051_821, w_051_823, w_051_824, w_051_827, w_051_830, w_051_831, w_051_835, w_051_836, w_051_840, w_051_841, w_051_842, w_051_846, w_051_848, w_051_849, w_051_850, w_051_851, w_051_853, w_051_855, w_051_857, w_051_859, w_051_863, w_051_865, w_051_866, w_051_867, w_051_871, w_051_872, w_051_875, w_051_877, w_051_878, w_051_881, w_051_882, w_051_883, w_051_884, w_051_885, w_051_886, w_051_887, w_051_889, w_051_890, w_051_893, w_051_894, w_051_896, w_051_897, w_051_898, w_051_900, w_051_901, w_051_905, w_051_906, w_051_907, w_051_908, w_051_910, w_051_912, w_051_913, w_051_914, w_051_917, w_051_919, w_051_921, w_051_922, w_051_923, w_051_924, w_051_925, w_051_926, w_051_927, w_051_928, w_051_929, w_051_933, w_051_934, w_051_936, w_051_937, w_051_938, w_051_939, w_051_940, w_051_941, w_051_942, w_051_943, w_051_946, w_051_949, w_051_950, w_051_952, w_051_953, w_051_954, w_051_956, w_051_957, w_051_960, w_051_963, w_051_964, w_051_965, w_051_966, w_051_971, w_051_975, w_051_977, w_051_981, w_051_986, w_051_987, w_051_989, w_051_990, w_051_996, w_051_998, w_051_999, w_051_1001, w_051_1002, w_051_1004, w_051_1005, w_051_1006, w_051_1008, w_051_1009, w_051_1010, w_051_1011, w_051_1012, w_051_1013, w_051_1014, w_051_1015, w_051_1016, w_051_1017, w_051_1020, w_051_1021, w_051_1022, w_051_1023, w_051_1026, w_051_1028, w_051_1029, w_051_1031, w_051_1032, w_051_1035, w_051_1036, w_051_1037, w_051_1038, w_051_1039, w_051_1041, w_051_1042, w_051_1043, w_051_1044, w_051_1045, w_051_1047, w_051_1050, w_051_1051, w_051_1052, w_051_1053, w_051_1054, w_051_1061, w_051_1062, w_051_1064, w_051_1065, w_051_1066, w_051_1067, w_051_1069, w_051_1071, w_051_1072, w_051_1075, w_051_1076, w_051_1078, w_051_1082, w_051_1083, w_051_1084, w_051_1085, w_051_1086, w_051_1088, w_051_1089, w_051_1092, w_051_1093, w_051_1095, w_051_1096, w_051_1097, w_051_1098, w_051_1099, w_051_1100, w_051_1101, w_051_1102, w_051_1103, w_051_1108, w_051_1110, w_051_1111, w_051_1112, w_051_1115, w_051_1116, w_051_1117, w_051_1118, w_051_1119, w_051_1120, w_051_1122, w_051_1124, w_051_1125, w_051_1126, w_051_1127, w_051_1128, w_051_1129, w_051_1132, w_051_1133, w_051_1134, w_051_1136, w_051_1139, w_051_1140, w_051_1141, w_051_1144, w_051_1145, w_051_1146, w_051_1147, w_051_1148, w_051_1150, w_051_1151, w_051_1154, w_051_1156, w_051_1157, w_051_1158, w_051_1159, w_051_1161, w_051_1162, w_051_1165, w_051_1166, w_051_1167, w_051_1169, w_051_1170, w_051_1171, w_051_1173, w_051_1175, w_051_1176, w_051_1177, w_051_1178, w_051_1179, w_051_1180, w_051_1181, w_051_1182, w_051_1184, w_051_1187, w_051_1188, w_051_1189, w_051_1190, w_051_1192, w_051_1193, w_051_1194, w_051_1196, w_051_1200, w_051_1201, w_051_1202, w_051_1203, w_051_1204, w_051_1205, w_051_1206, w_051_1207, w_051_1215, w_051_1216, w_051_1217, w_051_1219, w_051_1220, w_051_1221, w_051_1222, w_051_1223, w_051_1224, w_051_1225, w_051_1227, w_051_1228, w_051_1229, w_051_1230, w_051_1231, w_051_1232, w_051_1234, w_051_1235, w_051_1236, w_051_1238, w_051_1240, w_051_1241, w_051_1242, w_051_1243, w_051_1245, w_051_1246, w_051_1247, w_051_1248, w_051_1249, w_051_1250, w_051_1251, w_051_1253, w_051_1254, w_051_1255, w_051_1256, w_051_1258, w_051_1259, w_051_1260, w_051_1261, w_051_1262, w_051_1264, w_051_1266, w_051_1267, w_051_1268, w_051_1269, w_051_1271, w_051_1272, w_051_1275, w_051_1276, w_051_1278, w_051_1279, w_051_1280, w_051_1281, w_051_1282, w_051_1283, w_051_1285, w_051_1286, w_051_1287, w_051_1288, w_051_1289, w_051_1290, w_051_1292, w_051_1295, w_051_1296, w_051_1297, w_051_1298, w_051_1299, w_051_1300, w_051_1301, w_051_1302, w_051_1303, w_051_1305, w_051_1306, w_051_1307, w_051_1310, w_051_1311, w_051_1315, w_051_1316, w_051_1317, w_051_1318, w_051_1319, w_051_1320, w_051_1321, w_051_1322, w_051_1324, w_051_1325, w_051_1326, w_051_1327, w_051_1328, w_051_1329, w_051_1330, w_051_1331, w_051_1332, w_051_1333, w_051_1334, w_051_1335, w_051_1338, w_051_1339, w_051_1340, w_051_1342, w_051_1346, w_051_1348, w_051_1349, w_051_1351, w_051_1352, w_051_1354, w_051_1356, w_051_1359, w_051_1360, w_051_1362, w_051_1366, w_051_1368, w_051_1369, w_051_1371, w_051_1373, w_051_1375, w_051_1377, w_051_1379, w_051_1380, w_051_1381, w_051_1382, w_051_1384, w_051_1387, w_051_1389, w_051_1390, w_051_1391, w_051_1393, w_051_1396, w_051_1398, w_051_1399, w_051_1400, w_051_1402, w_051_1403, w_051_1404, w_051_1405, w_051_1407, w_051_1408, w_051_1411, w_051_1412, w_051_1414, w_051_1416, w_051_1417, w_051_1419, w_051_1420, w_051_1421, w_051_1422, w_051_1423, w_051_1424, w_051_1425, w_051_1426, w_051_1427, w_051_1428, w_051_1429, w_051_1430, w_051_1432, w_051_1433, w_051_1434, w_051_1435, w_051_1436, w_051_1437, w_051_1440, w_051_1441, w_051_1443, w_051_1445, w_051_1447, w_051_1448, w_051_1449, w_051_1453, w_051_1455, w_051_1457, w_051_1459, w_051_1461, w_051_1463, w_051_1464, w_051_1465, w_051_1467, w_051_1468, w_051_1469, w_051_1470, w_051_1472, w_051_1473, w_051_1475, w_051_1476, w_051_1477, w_051_1478, w_051_1479, w_051_1480, w_051_1483, w_051_1484, w_051_1485, w_051_1489, w_051_1490, w_051_1491, w_051_1492, w_051_1493, w_051_1494, w_051_1496, w_051_1497, w_051_1500, w_051_1501, w_051_1502, w_051_1503, w_051_1504, w_051_1506, w_051_1510, w_051_1511, w_051_1512, w_051_1513, w_051_1514, w_051_1515, w_051_1516, w_051_1517, w_051_1519, w_051_1520, w_051_1521, w_051_1522, w_051_1524, w_051_1525, w_051_1526, w_051_1527, w_051_1529, w_051_1530, w_051_1531, w_051_1532, w_051_1535, w_051_1536, w_051_1537, w_051_1538, w_051_1539, w_051_1540, w_051_1541, w_051_1544, w_051_1546, w_051_1547, w_051_1549, w_051_1550, w_051_1551, w_051_1554, w_051_1555, w_051_1556, w_051_1558, w_051_1559, w_051_1561, w_051_1562, w_051_1565, w_051_1566, w_051_1567, w_051_1573, w_051_1574, w_051_1575, w_051_1576, w_051_1577, w_051_1578, w_051_1579, w_051_1580, w_051_1581, w_051_1582, w_051_1583, w_051_1584, w_051_1586, w_051_1587, w_051_1589, w_051_1590, w_051_1591, w_051_1593, w_051_1594, w_051_1598, w_051_1599, w_051_1601, w_051_1602, w_051_1604, w_051_1608, w_051_1609, w_051_1612, w_051_1615, w_051_1617, w_051_1618, w_051_1619, w_051_1621, w_051_1622, w_051_1624, w_051_1625, w_051_1626, w_051_1628, w_051_1629, w_051_1631, w_051_1632, w_051_1634, w_051_1636, w_051_1637, w_051_1639, w_051_1640, w_051_1643, w_051_1645, w_051_1646, w_051_1647, w_051_1648, w_051_1651, w_051_1653, w_051_1657, w_051_1659, w_051_1660, w_051_1661, w_051_1664, w_051_1665, w_051_1666, w_051_1667, w_051_1668, w_051_1670, w_051_1671, w_051_1674, w_051_1681, w_051_1682, w_051_1683, w_051_1684, w_051_1685, w_051_1687, w_051_1690, w_051_1691, w_051_1692, w_051_1693, w_051_1694, w_051_1695, w_051_1698, w_051_1699, w_051_1700, w_051_1702, w_051_1703, w_051_1704, w_051_1706, w_051_1707, w_051_1709, w_051_1711, w_051_1713, w_051_1715, w_051_1716, w_051_1717, w_051_1718, w_051_1720, w_051_1721, w_051_1723, w_051_1724, w_051_1728, w_051_1732, w_051_1735, w_051_1736, w_051_1737, w_051_1738, w_051_1739, w_051_1740, w_051_1742, w_051_1743, w_051_1745, w_051_1746, w_051_1747, w_051_1748, w_051_1750, w_051_1751, w_051_1752, w_051_1753, w_051_1756, w_051_1758, w_051_1759, w_051_1760, w_051_1762, w_051_1763, w_051_1764, w_051_1765, w_051_1767, w_051_1769, w_051_1772, w_051_1776, w_051_1777, w_051_1778, w_051_1779, w_051_1780, w_051_1781, w_051_1782, w_051_1783, w_051_1784, w_051_1786, w_051_1787, w_051_1788, w_051_1789, w_051_1792, w_051_1795, w_051_1796, w_051_1797, w_051_1799, w_051_1801, w_051_1804, w_051_1808, w_051_1809, w_051_1810, w_051_1812, w_051_1813, w_051_1814, w_051_1815, w_051_1816, w_051_1817, w_051_1819, w_051_1820, w_051_1823, w_051_1824, w_051_1826, w_051_1827, w_051_1828, w_051_1829, w_051_1833, w_051_1835, w_051_1836, w_051_1837, w_051_1838, w_051_1839, w_051_1840, w_051_1842, w_051_1844, w_051_1845, w_051_1847, w_051_1850, w_051_1851, w_051_1854, w_051_1856, w_051_1858, w_051_1859, w_051_1860, w_051_1864, w_051_1865, w_051_1868, w_051_1869, w_051_1870, w_051_1871, w_051_1872, w_051_1873, w_051_1874, w_051_1877, w_051_1879, w_051_1880, w_051_1881, w_051_1883, w_051_1886, w_051_1887, w_051_1888, w_051_1889, w_051_1891, w_051_1892, w_051_1893, w_051_1895, w_051_1896, w_051_1897, w_051_1898, w_051_1899, w_051_1902, w_051_1905, w_051_1908, w_051_1909, w_051_1910, w_051_1911, w_051_1914, w_051_1916, w_051_1918, w_051_1919, w_051_1920, w_051_1921, w_051_1925, w_051_1926, w_051_1928, w_051_1929, w_051_1930, w_051_1931, w_051_1932, w_051_1934, w_051_1936, w_051_1940, w_051_1942, w_051_1944, w_051_1946, w_051_1947, w_051_1949, w_051_1953, w_051_1957, w_051_1959, w_051_1960, w_051_1965, w_051_1966, w_051_1969, w_051_1970, w_051_1972, w_051_1974, w_051_1975, w_051_1976, w_051_1977, w_051_1979, w_051_1981, w_051_1984, w_051_1985, w_051_1988, w_051_1992, w_051_1996, w_051_1997, w_051_2001, w_051_2003, w_051_2006, w_051_2007, w_051_2011, w_051_2012, w_051_2013, w_051_2014, w_051_2015, w_051_2016, w_051_2019, w_051_2020, w_051_2021, w_051_2024, w_051_2026, w_051_2027, w_051_2028, w_051_2029, w_051_2031, w_051_2033, w_051_2036, w_051_2037, w_051_2038, w_051_2040, w_051_2041, w_051_2042, w_051_2043, w_051_2044, w_051_2045, w_051_2046, w_051_2047, w_051_2048, w_051_2049, w_051_2053, w_051_2054, w_051_2056, w_051_2057, w_051_2058, w_051_2059, w_051_2060, w_051_2062, w_051_2063, w_051_2064, w_051_2065, w_051_2066, w_051_2067, w_051_2070, w_051_2072, w_051_2073, w_051_2074, w_051_2078, w_051_2079, w_051_2080, w_051_2081, w_051_2082, w_051_2083, w_051_2084, w_051_2085, w_051_2086, w_051_2088, w_051_2089, w_051_2092, w_051_2094, w_051_2096, w_051_2097, w_051_2098, w_051_2101, w_051_2102, w_051_2103, w_051_2104, w_051_2105, w_051_2106, w_051_2107, w_051_2108, w_051_2109, w_051_2110, w_051_2111, w_051_2113, w_051_2114, w_051_2116, w_051_2119, w_051_2121, w_051_2122, w_051_2123, w_051_2124, w_051_2126, w_051_2129, w_051_2130, w_051_2133, w_051_2134, w_051_2135, w_051_2136, w_051_2138, w_051_2141, w_051_2142, w_051_2143, w_051_2144, w_051_2145, w_051_2146, w_051_2147, w_051_2148, w_051_2149, w_051_2150, w_051_2151, w_051_2152, w_051_2153, w_051_2154, w_051_2156, w_051_2157, w_051_2158, w_051_2159, w_051_2160, w_051_2164, w_051_2166, w_051_2167, w_051_2168, w_051_2170, w_051_2171, w_051_2172, w_051_2174, w_051_2175, w_051_2178, w_051_2180, w_051_2182, w_051_2184, w_051_2185, w_051_2188, w_051_2189, w_051_2191, w_051_2192, w_051_2193, w_051_2194, w_051_2195, w_051_2196, w_051_2197, w_051_2198, w_051_2202, w_051_2203, w_051_2205, w_051_2206, w_051_2207, w_051_2208, w_051_2210, w_051_2211, w_051_2213, w_051_2214, w_051_2215, w_051_2216, w_051_2219, w_051_2221, w_051_2222, w_051_2224, w_051_2225, w_051_2226, w_051_2227, w_051_2229, w_051_2230, w_051_2232, w_051_2233, w_051_2236, w_051_2237, w_051_2238, w_051_2239, w_051_2241, w_051_2243, w_051_2244, w_051_2246, w_051_2247, w_051_2249, w_051_2250, w_051_2251, w_051_2253, w_051_2254, w_051_2255, w_051_2256, w_051_2257, w_051_2258, w_051_2259, w_051_2260, w_051_2263, w_051_2264, w_051_2265, w_051_2266, w_051_2268, w_051_2269, w_051_2271, w_051_2272, w_051_2273, w_051_2274, w_051_2275, w_051_2276, w_051_2277, w_051_2278, w_051_2279, w_051_2280, w_051_2281, w_051_2282, w_051_2286, w_051_2287, w_051_2289, w_051_2290, w_051_2291, w_051_2292, w_051_2293, w_051_2294, w_051_2295, w_051_2296, w_051_2299, w_051_2300, w_051_2301, w_051_2302, w_051_2303, w_051_2305, w_051_2307, w_051_2308, w_051_2310, w_051_2311, w_051_2312, w_051_2313, w_051_2315, w_051_2316, w_051_2320, w_051_2322, w_051_2324, w_051_2326, w_051_2327, w_051_2328, w_051_2330, w_051_2331, w_051_2332, w_051_2335, w_051_2337, w_051_2338, w_051_2339, w_051_2340, w_051_2342, w_051_2344, w_051_2346, w_051_2351, w_051_2352, w_051_2353, w_051_2354, w_051_2355, w_051_2358, w_051_2360, w_051_2361, w_051_2364, w_051_2365, w_051_2366, w_051_2368, w_051_2372, w_051_2374, w_051_2376, w_051_2378, w_051_2379, w_051_2381, w_051_2383, w_051_2386, w_051_2387, w_051_2388, w_051_2389, w_051_2390, w_051_2391, w_051_2392, w_051_2396, w_051_2397, w_051_2398, w_051_2399, w_051_2400, w_051_2401, w_051_2402, w_051_2404, w_051_2405, w_051_2406, w_051_2407, w_051_2408, w_051_2409, w_051_2410, w_051_2412, w_051_2414, w_051_2415, w_051_2416, w_051_2418, w_051_2419, w_051_2420, w_051_2421, w_051_2422, w_051_2423, w_051_2424, w_051_2425, w_051_2426, w_051_2427, w_051_2428, w_051_2429, w_051_2432, w_051_2433, w_051_2434, w_051_2435, w_051_2436, w_051_2437, w_051_2438, w_051_2439, w_051_2442, w_051_2443, w_051_2446, w_051_2448, w_051_2449, w_051_2450, w_051_2451, w_051_2452, w_051_2454, w_051_2455, w_051_2457, w_051_2459, w_051_2460, w_051_2461, w_051_2462, w_051_2463, w_051_2465, w_051_2466, w_051_2467, w_051_2468, w_051_2472, w_051_2473, w_051_2474, w_051_2475, w_051_2476, w_051_2477, w_051_2478, w_051_2480, w_051_2482, w_051_2483, w_051_2484, w_051_2485, w_051_2486, w_051_2487, w_051_2490, w_051_2492, w_051_2494, w_051_2498, w_051_2501, w_051_2503, w_051_2504, w_051_2505, w_051_2506, w_051_2507, w_051_2508, w_051_2510, w_051_2511, w_051_2512, w_051_2513, w_051_2514, w_051_2515, w_051_2517, w_051_2519, w_051_2520, w_051_2522, w_051_2523, w_051_2524, w_051_2526, w_051_2528, w_051_2529, w_051_2531, w_051_2533, w_051_2534, w_051_2535, w_051_2536, w_051_2537, w_051_2542, w_051_2544, w_051_2545, w_051_2549, w_051_2551, w_051_2552, w_051_2553, w_051_2555, w_051_2558, w_051_2559, w_051_2561, w_051_2562, w_051_2564, w_051_2566, w_051_2567, w_051_2570, w_051_2571, w_051_2572, w_051_2576, w_051_2577, w_051_2578, w_051_2579, w_051_2580, w_051_2581, w_051_2582, w_051_2583, w_051_2585, w_051_2586, w_051_2587, w_051_2588, w_051_2591, w_051_2592, w_051_2593, w_051_2594, w_051_2595, w_051_2597, w_051_2598, w_051_2599, w_051_2600, w_051_2601, w_051_2602, w_051_2604, w_051_2605, w_051_2606, w_051_2607, w_051_2608, w_051_2609, w_051_2610, w_051_2611, w_051_2613, w_051_2615, w_051_2616, w_051_2617, w_051_2619, w_051_2620, w_051_2621, w_051_2624, w_051_2625, w_051_2626, w_051_2627, w_051_2628, w_051_2630, w_051_2631, w_051_2632, w_051_2633, w_051_2636, w_051_2639, w_051_2640, w_051_2641, w_051_2642, w_051_2644, w_051_2645, w_051_2646, w_051_2649, w_051_2650, w_051_2651, w_051_2652, w_051_2653, w_051_2654, w_051_2655, w_051_2657, w_051_2658, w_051_2659, w_051_2661, w_051_2662, w_051_2664, w_051_2665, w_051_2667, w_051_2668, w_051_2669, w_051_2670, w_051_2671, w_051_2674, w_051_2676, w_051_2677, w_051_2678, w_051_2679, w_051_2680, w_051_2681, w_051_2682, w_051_2683, w_051_2684, w_051_2687, w_051_2691, w_051_2692, w_051_2694, w_051_2695, w_051_2696, w_051_2698, w_051_2699, w_051_2700, w_051_2702, w_051_2706, w_051_2707, w_051_2708, w_051_2709, w_051_2710, w_051_2711, w_051_2712, w_051_2714, w_051_2715, w_051_2716, w_051_2718, w_051_2722, w_051_2723, w_051_2724, w_051_2725, w_051_2727, w_051_2729, w_051_2730, w_051_2731, w_051_2732, w_051_2733, w_051_2734, w_051_2735, w_051_2736, w_051_2737, w_051_2739, w_051_2742, w_051_2744, w_051_2746, w_051_2747, w_051_2757, w_051_2759, w_051_2761, w_051_2762, w_051_2764, w_051_2765, w_051_2768, w_051_2770, w_051_2774, w_051_2775, w_051_2776, w_051_2777, w_051_2780, w_051_2781, w_051_2783, w_051_2784, w_051_2785, w_051_2786, w_051_2788, w_051_2789, w_051_2791, w_051_2796, w_051_2798, w_051_2799, w_051_2801, w_051_2802, w_051_2803, w_051_2804, w_051_2805, w_051_2806, w_051_2808, w_051_2813, w_051_2814, w_051_2816, w_051_2817, w_051_2818, w_051_2821, w_051_2822, w_051_2824, w_051_2825, w_051_2826, w_051_2827, w_051_2829, w_051_2830, w_051_2832, w_051_2833, w_051_2834, w_051_2835, w_051_2837, w_051_2839, w_051_2841, w_051_2843, w_051_2845, w_051_2847, w_051_2850, w_051_2851, w_051_2852, w_051_2857, w_051_2858, w_051_2859, w_051_2860, w_051_2861, w_051_2862, w_051_2863, w_051_2864, w_051_2866, w_051_2868, w_051_2869, w_051_2870, w_051_2871, w_051_2872, w_051_2873, w_051_2874, w_051_2876, w_051_2878, w_051_2879, w_051_2886, w_051_2887, w_051_2888, w_051_2889, w_051_2891, w_051_2893, w_051_2894, w_051_2895, w_051_2897, w_051_2898, w_051_2899, w_051_2901, w_051_2902, w_051_2903, w_051_2904, w_051_2905, w_051_2906, w_051_2907, w_051_2908, w_051_2909, w_051_2910, w_051_2912, w_051_2916, w_051_2917, w_051_2918, w_051_2920, w_051_2921, w_051_2922, w_051_2923, w_051_2926, w_051_2927, w_051_2930, w_051_2931, w_051_2932, w_051_2934, w_051_2936, w_051_2939, w_051_2940, w_051_2941, w_051_2943, w_051_2945, w_051_2946, w_051_2948, w_051_2949, w_051_2950, w_051_2951, w_051_2952, w_051_2955, w_051_2956, w_051_2957, w_051_2959, w_051_2963, w_051_2964, w_051_2966, w_051_2967, w_051_2968, w_051_2971, w_051_2972, w_051_2974, w_051_2979, w_051_2980, w_051_2983, w_051_2985, w_051_2986, w_051_2988, w_051_2989, w_051_2992, w_051_2993, w_051_2995, w_051_2997, w_051_2998, w_051_2999, w_051_3000, w_051_3001, w_051_3002, w_051_3003, w_051_3004, w_051_3007, w_051_3008, w_051_3009, w_051_3011, w_051_3012, w_051_3013, w_051_3014, w_051_3016, w_051_3017, w_051_3018, w_051_3019, w_051_3020, w_051_3021, w_051_3022, w_051_3023, w_051_3024, w_051_3025, w_051_3026, w_051_3027, w_051_3031, w_051_3032, w_051_3033, w_051_3034, w_051_3036, w_051_3037, w_051_3040, w_051_3041, w_051_3042, w_051_3043, w_051_3046, w_051_3048, w_051_3051, w_051_3052, w_051_3053, w_051_3054, w_051_3055, w_051_3056, w_051_3057, w_051_3058, w_051_3061, w_051_3063, w_051_3064, w_051_3065, w_051_3066, w_051_3067, w_051_3068, w_051_3069, w_051_3071, w_051_3072, w_051_3073, w_051_3074, w_051_3075, w_051_3079, w_051_3080, w_051_3084, w_051_3086, w_051_3088, w_051_3089, w_051_3090, w_051_3092, w_051_3095, w_051_3096, w_051_3097, w_051_3101, w_051_3103, w_051_3104, w_051_3105, w_051_3107, w_051_3108, w_051_3109, w_051_3111, w_051_3112, w_051_3113, w_051_3114, w_051_3115, w_051_3116, w_051_3118, w_051_3119, w_051_3120, w_051_3121, w_051_3122, w_051_3123, w_051_3126, w_051_3128, w_051_3129, w_051_3130, w_051_3131, w_051_3132, w_051_3135, w_051_3138, w_051_3139, w_051_3140, w_051_3142, w_051_3143, w_051_3144, w_051_3145, w_051_3146, w_051_3147, w_051_3149, w_051_3150, w_051_3151, w_051_3152, w_051_3153, w_051_3155, w_051_3156, w_051_3158, w_051_3159, w_051_3160, w_051_3161, w_051_3162, w_051_3163, w_051_3164, w_051_3167, w_051_3168, w_051_3170, w_051_3171, w_051_3172, w_051_3173, w_051_3174, w_051_3176, w_051_3177, w_051_3178, w_051_3180, w_051_3183, w_051_3184, w_051_3185, w_051_3186, w_051_3187, w_051_3190, w_051_3191, w_051_3192, w_051_3193, w_051_3194, w_051_3196, w_051_3198, w_051_3200, w_051_3203, w_051_3204, w_051_3207, w_051_3208, w_051_3209, w_051_3213, w_051_3214, w_051_3215, w_051_3217, w_051_3218, w_051_3220, w_051_3223, w_051_3224, w_051_3230, w_051_3231, w_051_3234, w_051_3235, w_051_3237, w_051_3238, w_051_3239, w_051_3241, w_051_3243, w_051_3244, w_051_3246, w_051_3247, w_051_3248, w_051_3249, w_051_3250, w_051_3252, w_051_3257, w_051_3258, w_051_3260, w_051_3267, w_051_3268, w_051_3271, w_051_3273, w_051_3274, w_051_3276, w_051_3277, w_051_3278, w_051_3281, w_051_3282, w_051_3283, w_051_3285, w_051_3286, w_051_3287, w_051_3290, w_051_3291, w_051_3292, w_051_3293, w_051_3294, w_051_3296, w_051_3297, w_051_3298, w_051_3299, w_051_3301, w_051_3306, w_051_3307, w_051_3308, w_051_3312, w_051_3313, w_051_3314, w_051_3320, w_051_3321, w_051_3322, w_051_3323, w_051_3324, w_051_3325, w_051_3326, w_051_3327, w_051_3329, w_051_3330, w_051_3331, w_051_3332, w_051_3333, w_051_3334, w_051_3335, w_051_3336, w_051_3338, w_051_3340, w_051_3341, w_051_3343, w_051_3346, w_051_3348, w_051_3349, w_051_3350, w_051_3353, w_051_3354, w_051_3356, w_051_3357, w_051_3360, w_051_3361, w_051_3362, w_051_3363, w_051_3364, w_051_3365, w_051_3366, w_051_3367, w_051_3368, w_051_3369, w_051_3370, w_051_3373, w_051_3374, w_051_3375, w_051_3378, w_051_3379, w_051_3382, w_051_3383, w_051_3385, w_051_3387, w_051_3388, w_051_3389, w_051_3391, w_051_3392, w_051_3393, w_051_3394, w_051_3395, w_051_3396, w_051_3397, w_051_3398, w_051_3399, w_051_3403, w_051_3404, w_051_3405, w_051_3406, w_051_3407, w_051_3409, w_051_3411, w_051_3413, w_051_3414, w_051_3416, w_051_3417, w_051_3418, w_051_3419, w_051_3421, w_051_3422, w_051_3423, w_051_3424, w_051_3425, w_051_3426, w_051_3427, w_051_3428, w_051_3430, w_051_3431, w_051_3432, w_051_3433, w_051_3434, w_051_3435, w_051_3436, w_051_3437, w_051_3438, w_051_3439, w_051_3440, w_051_3442, w_051_3443, w_051_3445, w_051_3447, w_051_3448, w_051_3449, w_051_3452, w_051_3453, w_051_3454, w_051_3455, w_051_3456, w_051_3459, w_051_3460, w_051_3463, w_051_3465, w_051_3466, w_051_3467, w_051_3469, w_051_3470, w_051_3471, w_051_3473, w_051_3477, w_051_3478, w_051_3479, w_051_3480, w_051_3482, w_051_3483, w_051_3484, w_051_3485, w_051_3487, w_051_3489, w_051_3490, w_051_3491, w_051_3492, w_051_3493, w_051_3494, w_051_3495, w_051_3496, w_051_3497, w_051_3498, w_051_3500, w_051_3503, w_051_3507, w_051_3508, w_051_3512, w_051_3514, w_051_3515, w_051_3516, w_051_3518, w_051_3520, w_051_3521, w_051_3522, w_051_3523, w_051_3524, w_051_3525, w_051_3526, w_051_3527, w_051_3529, w_051_3530, w_051_3533, w_051_3534, w_051_3536, w_051_3537, w_051_3538, w_051_3540, w_051_3541, w_051_3543, w_051_3544, w_051_3545, w_051_3547, w_051_3549, w_051_3550, w_051_3551, w_051_3552, w_051_3553, w_051_3554, w_051_3555, w_051_3557, w_051_3558, w_051_3562, w_051_3563, w_051_3565, w_051_3566, w_051_3571, w_051_3572, w_051_3574, w_051_3575, w_051_3576, w_051_3577, w_051_3579, w_051_3581, w_051_3583, w_051_3584, w_051_3587, w_051_3588, w_051_3589, w_051_3592, w_051_3593, w_051_3594, w_051_3595, w_051_3597, w_051_3600, w_051_3602, w_051_3604, w_051_3605, w_051_3607, w_051_3608, w_051_3609, w_051_3610, w_051_3611, w_051_3613, w_051_3614, w_051_3615, w_051_3616, w_051_3617, w_051_3618, w_051_3621, w_051_3622, w_051_3623, w_051_3624, w_051_3628, w_051_3629, w_051_3630, w_051_3635, w_051_3636, w_051_3639, w_051_3640, w_051_3641, w_051_3642, w_051_3643, w_051_3648, w_051_3651, w_051_3653, w_051_3654, w_051_3656, w_051_3657, w_051_3659, w_051_3660, w_051_3661, w_051_3662, w_051_3665, w_051_3666, w_051_3668, w_051_3674, w_051_3676, w_051_3677, w_051_3678, w_051_3679, w_051_3680, w_051_3681, w_051_3682, w_051_3683, w_051_3686, w_051_3687, w_051_3688, w_051_3689, w_051_3690, w_051_3691, w_051_3693, w_051_3694, w_051_3696, w_051_3697, w_051_3698, w_051_3699, w_051_3701, w_051_3702, w_051_3703, w_051_3704, w_051_3705, w_051_3706, w_051_3708, w_051_3709, w_051_3710, w_051_3713, w_051_3714, w_051_3715, w_051_3717, w_051_3718, w_051_3719, w_051_3721, w_051_3724, w_051_3727, w_051_3728, w_051_3732, w_051_3733, w_051_3734, w_051_3735, w_051_3737, w_051_3738, w_051_3740, w_051_3741, w_051_3742, w_051_3743, w_051_3744, w_051_3746, w_051_3748, w_051_3749, w_051_3750, w_051_3752, w_051_3753, w_051_3755, w_051_3756, w_051_3757, w_051_3758, w_051_3760, w_051_3761, w_051_3762, w_051_3763, w_051_3764, w_051_3765, w_051_3767, w_051_3768, w_051_3769, w_051_3770, w_051_3771, w_051_3772, w_051_3776, w_051_3778, w_051_3780, w_051_3781, w_051_3782, w_051_3783, w_051_3787, w_051_3788, w_051_3789, w_051_3790, w_051_3792, w_051_3794, w_051_3795, w_051_3796, w_051_3797, w_051_3798, w_051_3799, w_051_3804, w_051_3805, w_051_3806, w_051_3807, w_051_3813, w_051_3814, w_051_3815, w_051_3821, w_051_3822, w_051_3823, w_051_3824, w_051_3826, w_051_3827, w_051_3830, w_051_3831, w_051_3833, w_051_3834, w_051_3836, w_051_3840, w_051_3841, w_051_3842, w_051_3846, w_051_3847, w_051_3848, w_051_3849, w_051_3851, w_051_3854, w_051_3856, w_051_3857, w_051_3858, w_051_3861, w_051_3863, w_051_3864, w_051_3867, w_051_3871, w_051_3872, w_051_3876, w_051_3877, w_051_3880, w_051_3881, w_051_3882, w_051_3885, w_051_3886, w_051_3888, w_051_3892, w_051_3895, w_051_3896, w_051_3897, w_051_3898, w_051_3899, w_051_3900, w_051_3905, w_051_3906, w_051_3907, w_051_3908, w_051_3910, w_051_3911, w_051_3913, w_051_3914, w_051_3918, w_051_3919, w_051_3920, w_051_3921, w_051_3923, w_051_3924, w_051_3926, w_051_3929, w_051_3930, w_051_3931, w_051_3933, w_051_3934, w_051_3937, w_051_3938, w_051_3941, w_051_3942, w_051_3944, w_051_3945, w_051_3946, w_051_3947, w_051_3951, w_051_3953, w_051_3954, w_051_3958, w_051_3959, w_051_3960, w_051_3961, w_051_3962, w_051_3963, w_051_3964, w_051_3966, w_051_3967, w_051_3970, w_051_3971, w_051_3973, w_051_3975, w_051_3976, w_051_3977, w_051_3978, w_051_3980, w_051_3982, w_051_3983, w_051_3985, w_051_3986, w_051_3987, w_051_3989, w_051_3991, w_051_3993, w_051_3994, w_051_3996, w_051_3997, w_051_3998, w_051_4001, w_051_4002, w_051_4003, w_051_4004, w_051_4005, w_051_4006, w_051_4007, w_051_4009, w_051_4011, w_051_4014, w_051_4015, w_051_4018, w_051_4020, w_051_4021, w_051_4022, w_051_4023, w_051_4024, w_051_4026, w_051_4027, w_051_4030, w_051_4031, w_051_4033, w_051_4034, w_051_4035, w_051_4036, w_051_4037, w_051_4038, w_051_4040, w_051_4041, w_051_4042, w_051_4047, w_051_4049, w_051_4050, w_051_4053, w_051_4054, w_051_4055, w_051_4056, w_051_4059, w_051_4060, w_051_4061, w_051_4062, w_051_4063, w_051_4064, w_051_4065, w_051_4066, w_051_4067, w_051_4068, w_051_4070, w_051_4071, w_051_4072, w_051_4073, w_051_4074, w_051_4075, w_051_4077, w_051_4078, w_051_4079, w_051_4080, w_051_4081, w_051_4082, w_051_4083, w_051_4084, w_051_4085, w_051_4087, w_051_4088, w_051_4089, w_051_4090, w_051_4091, w_051_4092, w_051_4093, w_051_4094, w_051_4096, w_051_4097, w_051_4098, w_051_4100, w_051_4101, w_051_4103, w_051_4104, w_051_4108, w_051_4111, w_051_4112, w_051_4113, w_051_4115, w_051_4117, w_051_4118, w_051_4119, w_051_4120, w_051_4121, w_051_4122, w_051_4124, w_051_4126, w_051_4127, w_051_4128, w_051_4129, w_051_4130, w_051_4131, w_051_4132, w_051_4133, w_051_4134, w_051_4135, w_051_4136, w_051_4137, w_051_4139, w_051_4140, w_051_4142, w_051_4143, w_051_4144, w_051_4145, w_051_4146, w_051_4147, w_051_4148, w_051_4152, w_051_4155, w_051_4156, w_051_4157, w_051_4159, w_051_4160, w_051_4161, w_051_4163, w_051_4165, w_051_4166, w_051_4169, w_051_4170, w_051_4171, w_051_4174, w_051_4175, w_051_4176, w_051_4177, w_051_4178, w_051_4179, w_051_4180, w_051_4182, w_051_4183, w_051_4185, w_051_4186, w_051_4189, w_051_4191, w_051_4194, w_051_4195, w_051_4196, w_051_4197, w_051_4199, w_051_4200, w_051_4201, w_051_4202, w_051_4203, w_051_4206, w_051_4207, w_051_4208, w_051_4209, w_051_4210, w_051_4211, w_051_4212, w_051_4213, w_051_4215, w_051_4217, w_051_4219, w_051_4221, w_051_4223, w_051_4226, w_051_4227, w_051_4228, w_051_4232, w_051_4233, w_051_4234, w_051_4238, w_051_4240, w_051_4241, w_051_4242, w_051_4244, w_051_4245, w_051_4247, w_051_4249, w_051_4250, w_051_4251, w_051_4253, w_051_4255, w_051_4256, w_051_4257, w_051_4259, w_051_4261, w_051_4262, w_051_4263, w_051_4264, w_051_4265, w_051_4266, w_051_4268, w_051_4271, w_051_4272, w_051_4273, w_051_4274, w_051_4276, w_051_4278, w_051_4279, w_051_4280, w_051_4282, w_051_4283, w_051_4284, w_051_4285, w_051_4286, w_051_4287, w_051_4289, w_051_4291, w_051_4292, w_051_4294, w_051_4295, w_051_4297, w_051_4299, w_051_4301, w_051_4302, w_051_4304, w_051_4307, w_051_4308, w_051_4309, w_051_4310, w_051_4311, w_051_4312, w_051_4314, w_051_4315, w_051_4316, w_051_4317, w_051_4318, w_051_4319, w_051_4320, w_051_4321, w_051_4325, w_051_4326, w_051_4328, w_051_4330, w_051_4331, w_051_4332, w_051_4333, w_051_4337, w_051_4339, w_051_4340, w_051_4341, w_051_4342, w_051_4344, w_051_4345, w_051_4346, w_051_4347, w_051_4348, w_051_4349, w_051_4350, w_051_4353, w_051_4354, w_051_4356, w_051_4357, w_051_4359, w_051_4360, w_051_4361, w_051_4362, w_051_4366, w_051_4368, w_051_4370, w_051_4372, w_051_4373, w_051_4374, w_051_4375, w_051_4376, w_051_4377, w_051_4378, w_051_4380, w_051_4381, w_051_4382, w_051_4383, w_051_4384, w_051_4385, w_051_4386, w_051_4387, w_051_4391, w_051_4393, w_051_4399, w_051_4401, w_051_4407, w_051_4410, w_051_4415, w_051_4419, w_051_4421, w_051_4423, w_051_4425, w_051_4426, w_051_4427, w_051_4428, w_051_4430, w_051_4442, w_051_4444, w_051_4445, w_051_4447, w_051_4452, w_051_4454, w_051_4456, w_051_4464, w_051_4468, w_051_4473, w_051_4483, w_051_4484, w_051_4488, w_051_4490, w_051_4491, w_051_4492, w_051_4493, w_051_4502, w_051_4503, w_051_4508, w_051_4511, w_051_4512, w_051_4515, w_051_4519, w_051_4520, w_051_4523, w_051_4525, w_051_4527, w_051_4529, w_051_4532, w_051_4534, w_051_4539, w_051_4544, w_051_4545, w_051_4549, w_051_4550, w_051_4551, w_051_4552, w_051_4555, w_051_4562, w_051_4567, w_051_4569, w_051_4570, w_051_4571, w_051_4577, w_051_4579, w_051_4583, w_051_4585, w_051_4589, w_051_4591, w_051_4592, w_051_4593, w_051_4600, w_051_4601, w_051_4603, w_051_4605, w_051_4606, w_051_4610, w_051_4613, w_051_4618, w_051_4619, w_051_4621, w_051_4623, w_051_4627, w_051_4628, w_051_4629, w_051_4637, w_051_4639, w_051_4645, w_051_4646, w_051_4647, w_051_4648, w_051_4650, w_051_4651, w_051_4653, w_051_4654, w_051_4656, w_051_4658, w_051_4659, w_051_4663, w_051_4667, w_051_4671, w_051_4674, w_051_4682, w_051_4685, w_051_4687, w_051_4692, w_051_4695, w_051_4701, w_051_4702, w_051_4707, w_051_4709, w_051_4711, w_051_4714, w_051_4715, w_051_4720, w_051_4723, w_051_4724, w_051_4725, w_051_4727, w_051_4730, w_051_4734, w_051_4735, w_051_4739, w_051_4740, w_051_4741, w_051_4742, w_051_4749, w_051_4755, w_051_4758, w_051_4763, w_051_4766, w_051_4771, w_051_4772, w_051_4773, w_051_4779, w_051_4780, w_051_4781, w_051_4785, w_051_4787, w_051_4789, w_051_4793, w_051_4797, w_051_4799, w_051_4800, w_051_4804, w_051_4805, w_051_4807, w_051_4808, w_051_4809, w_051_4810, w_051_4815, w_051_4818, w_051_4820, w_051_4822, w_051_4823, w_051_4824, w_051_4826, w_051_4827, w_051_4830, w_051_4831, w_051_4851, w_051_4854, w_051_4855, w_051_4856, w_051_4858, w_051_4860, w_051_4861, w_051_4865, w_051_4866, w_051_4867, w_051_4870, w_051_4872, w_051_4873, w_051_4876, w_051_4877, w_051_4878, w_051_4879, w_051_4881, w_051_4882, w_051_4884, w_051_4885, w_051_4886, w_051_4887, w_051_4889, w_051_4894, w_051_4896, w_051_4897, w_051_4898, w_051_4900, w_051_4902, w_051_4905, w_051_4910, w_051_4913, w_051_4916, w_051_4918, w_051_4920, w_051_4922, w_051_4924, w_051_4925, w_051_4931, w_051_4932, w_051_4934, w_051_4936, w_051_4945, w_051_4946, w_051_4948, w_051_4951, w_051_4957, w_051_4959, w_051_4960, w_051_4964, w_051_4967, w_051_4968, w_051_4970, w_051_4973, w_051_4974, w_051_4976, w_051_4978, w_051_4983, w_051_4987, w_051_4993, w_051_4994, w_051_4995, w_051_4999, w_051_5001, w_051_5006, w_051_5007, w_051_5012, w_051_5014, w_051_5023, w_051_5024, w_051_5026, w_051_5027, w_051_5028, w_051_5030, w_051_5037, w_051_5038, w_051_5041, w_051_5047, w_051_5051, w_051_5052, w_051_5054, w_051_5055, w_051_5056, w_051_5057, w_051_5062, w_051_5063, w_051_5064, w_051_5066, w_051_5073, w_051_5076, w_051_5077, w_051_5078, w_051_5079, w_051_5080, w_051_5083, w_051_5084, w_051_5087, w_051_5088, w_051_5089, w_051_5093, w_051_5095, w_051_5099, w_051_5100, w_051_5101, w_051_5102, w_051_5107, w_051_5108, w_051_5116, w_051_5117, w_051_5118, w_051_5121, w_051_5124, w_051_5125, w_051_5133, w_051_5136, w_051_5137, w_051_5138, w_051_5140, w_051_5143, w_051_5146, w_051_5147, w_051_5151, w_051_5153, w_051_5160, w_051_5161, w_051_5168, w_051_5169, w_051_5170, w_051_5173, w_051_5174, w_051_5180, w_051_5185, w_051_5186, w_051_5192, w_051_5195, w_051_5196, w_051_5198, w_051_5200, w_051_5201, w_051_5202, w_051_5204, w_051_5209, w_051_5213, w_051_5219, w_051_5224, w_051_5226, w_051_5227, w_051_5228, w_051_5231, w_051_5233, w_051_5234, w_051_5237, w_051_5238, w_051_5241, w_051_5242, w_051_5243, w_051_5244, w_051_5248, w_051_5250, w_051_5253, w_051_5255, w_051_5261, w_051_5262, w_051_5268, w_051_5269, w_051_5270, w_051_5272, w_051_5273, w_051_5274, w_051_5275, w_051_5277, w_051_5278, w_051_5289, w_051_5290, w_051_5291, w_051_5294, w_051_5296, w_051_5297, w_051_5300, w_051_5301, w_051_5304, w_051_5306, w_051_5310, w_051_5313, w_051_5316, w_051_5317, w_051_5318, w_051_5321, w_051_5322, w_051_5324, w_051_5326, w_051_5328, w_051_5329, w_051_5330, w_051_5335, w_051_5339, w_051_5345, w_051_5348, w_051_5349, w_051_5351, w_051_5352, w_051_5353, w_051_5354, w_051_5357, w_051_5358, w_051_5365, w_051_5366, w_051_5368, w_051_5369, w_051_5370, w_051_5372, w_051_5374, w_051_5383, w_051_5386, w_051_5387, w_051_5388, w_051_5391, w_051_5392, w_051_5399, w_051_5401, w_051_5408, w_051_5409, w_051_5412, w_051_5417, w_051_5418, w_051_5419, w_051_5422, w_051_5424, w_051_5425, w_051_5426, w_051_5428, w_051_5430, w_051_5432, w_051_5436, w_051_5437, w_051_5438, w_051_5439, w_051_5440, w_051_5441, w_051_5443, w_051_5444, w_051_5445, w_051_5451, w_051_5457, w_051_5459, w_051_5464, w_051_5466, w_051_5467, w_051_5469, w_051_5478, w_051_5479, w_051_5480, w_051_5488, w_051_5490, w_051_5491, w_051_5495, w_051_5503, w_051_5504, w_051_5507, w_051_5512, w_051_5514, w_051_5520, w_051_5526, w_051_5530, w_051_5531, w_051_5532, w_051_5534, w_051_5535, w_051_5536, w_051_5537, w_051_5539, w_051_5549, w_051_5551, w_051_5552, w_051_5555, w_051_5556, w_051_5561, w_051_5563, w_051_5564, w_051_5570, w_051_5578, w_051_5579, w_051_5581, w_051_5585, w_051_5586, w_051_5587, w_051_5591, w_051_5593, w_051_5594, w_051_5595, w_051_5596, w_051_5598, w_051_5599, w_051_5600, w_051_5604, w_051_5607, w_051_5609, w_051_5610;
  wire w_052_000, w_052_001, w_052_002, w_052_003, w_052_004, w_052_005, w_052_006, w_052_007, w_052_009, w_052_010, w_052_011, w_052_012, w_052_013, w_052_014, w_052_015, w_052_016, w_052_018, w_052_019, w_052_020, w_052_022, w_052_023, w_052_024, w_052_025, w_052_026, w_052_027, w_052_028, w_052_029, w_052_030, w_052_031, w_052_032, w_052_033, w_052_034, w_052_035, w_052_036, w_052_037, w_052_038, w_052_039, w_052_040, w_052_041, w_052_042, w_052_043, w_052_044, w_052_045, w_052_046, w_052_047, w_052_049, w_052_050, w_052_051, w_052_052, w_052_053, w_052_055, w_052_056, w_052_057, w_052_058, w_052_059, w_052_060, w_052_061, w_052_062, w_052_063, w_052_064, w_052_065, w_052_066, w_052_067, w_052_068, w_052_069, w_052_070, w_052_071, w_052_072, w_052_073, w_052_074, w_052_075, w_052_076, w_052_078, w_052_079, w_052_080, w_052_081, w_052_082, w_052_083, w_052_084, w_052_085, w_052_086, w_052_087, w_052_088, w_052_089, w_052_090, w_052_091, w_052_092, w_052_093, w_052_094, w_052_095, w_052_096, w_052_097, w_052_098, w_052_099, w_052_100, w_052_101, w_052_102, w_052_103, w_052_104, w_052_105, w_052_106, w_052_107, w_052_108, w_052_109, w_052_110, w_052_111, w_052_112, w_052_113, w_052_114, w_052_115, w_052_116, w_052_117, w_052_118, w_052_119, w_052_120, w_052_121, w_052_122, w_052_123, w_052_124, w_052_125, w_052_126, w_052_127, w_052_128, w_052_129, w_052_130, w_052_131, w_052_132, w_052_133, w_052_134, w_052_135, w_052_136, w_052_137, w_052_138, w_052_139, w_052_140, w_052_141, w_052_143, w_052_144, w_052_145, w_052_146, w_052_147, w_052_148, w_052_149, w_052_150, w_052_151, w_052_152, w_052_154, w_052_155, w_052_156, w_052_157, w_052_158, w_052_159, w_052_160, w_052_161, w_052_162, w_052_163, w_052_164, w_052_165, w_052_166, w_052_167, w_052_168, w_052_169, w_052_170, w_052_171, w_052_172, w_052_173, w_052_174, w_052_175, w_052_176, w_052_177, w_052_178, w_052_179, w_052_180, w_052_181, w_052_182, w_052_183, w_052_184, w_052_185, w_052_186, w_052_187, w_052_188, w_052_189, w_052_190, w_052_191, w_052_192, w_052_193, w_052_194, w_052_195, w_052_196, w_052_197, w_052_198, w_052_199, w_052_200, w_052_201, w_052_202, w_052_203, w_052_204, w_052_205, w_052_206, w_052_207, w_052_208, w_052_209, w_052_210, w_052_211, w_052_213, w_052_214, w_052_215, w_052_216, w_052_217, w_052_218, w_052_219, w_052_220, w_052_221, w_052_222, w_052_223, w_052_225, w_052_226, w_052_227, w_052_228, w_052_229, w_052_230, w_052_231, w_052_232, w_052_233, w_052_234, w_052_235, w_052_236, w_052_237, w_052_238, w_052_239, w_052_240, w_052_241, w_052_242, w_052_243, w_052_244, w_052_246, w_052_247, w_052_248, w_052_249, w_052_250, w_052_251, w_052_252, w_052_253, w_052_254, w_052_255, w_052_256, w_052_257, w_052_258, w_052_259, w_052_260, w_052_261, w_052_262, w_052_263, w_052_264, w_052_265, w_052_266, w_052_267, w_052_268, w_052_269, w_052_270, w_052_271, w_052_272, w_052_273, w_052_274, w_052_275, w_052_276, w_052_277, w_052_278, w_052_279, w_052_280, w_052_281, w_052_282, w_052_283, w_052_284, w_052_285, w_052_286, w_052_287, w_052_288, w_052_289, w_052_290, w_052_291, w_052_292, w_052_293, w_052_294, w_052_295, w_052_296, w_052_297, w_052_298, w_052_300, w_052_301, w_052_302, w_052_303, w_052_304, w_052_306, w_052_307, w_052_309, w_052_310, w_052_311, w_052_312, w_052_313, w_052_314, w_052_315, w_052_316, w_052_317, w_052_318, w_052_319, w_052_320, w_052_321, w_052_322, w_052_323, w_052_324, w_052_325, w_052_326, w_052_327, w_052_328, w_052_329, w_052_330, w_052_331, w_052_332, w_052_333, w_052_334, w_052_335, w_052_336, w_052_337, w_052_338, w_052_339, w_052_340, w_052_341, w_052_342, w_052_343, w_052_344, w_052_345, w_052_346, w_052_347, w_052_348, w_052_349, w_052_350, w_052_351, w_052_352, w_052_353, w_052_356, w_052_357, w_052_358, w_052_360, w_052_361, w_052_362, w_052_363, w_052_364, w_052_365, w_052_366, w_052_367, w_052_368, w_052_369, w_052_370, w_052_371, w_052_372, w_052_374, w_052_375, w_052_376, w_052_377, w_052_378, w_052_379, w_052_380, w_052_381, w_052_382, w_052_383, w_052_384, w_052_385, w_052_386, w_052_387, w_052_388, w_052_389, w_052_390, w_052_391, w_052_392, w_052_393, w_052_394, w_052_395, w_052_396, w_052_397, w_052_398, w_052_400, w_052_401, w_052_402, w_052_403, w_052_404, w_052_405, w_052_406, w_052_407, w_052_408, w_052_409, w_052_410, w_052_411, w_052_412, w_052_413, w_052_414, w_052_415, w_052_416, w_052_417, w_052_418, w_052_419, w_052_420, w_052_422, w_052_423, w_052_424, w_052_425, w_052_426, w_052_427, w_052_428, w_052_429, w_052_430, w_052_431, w_052_432, w_052_434, w_052_436, w_052_437, w_052_438, w_052_439, w_052_440, w_052_441, w_052_442, w_052_443, w_052_444, w_052_445, w_052_446, w_052_447, w_052_448, w_052_449, w_052_450, w_052_451, w_052_452, w_052_453, w_052_454, w_052_455, w_052_456, w_052_457, w_052_458, w_052_459, w_052_460, w_052_461, w_052_462, w_052_463, w_052_464, w_052_465, w_052_466, w_052_467, w_052_468, w_052_469, w_052_470, w_052_471, w_052_472, w_052_474, w_052_475, w_052_476, w_052_477, w_052_478, w_052_479, w_052_480, w_052_481, w_052_482, w_052_483, w_052_484, w_052_485, w_052_486, w_052_487, w_052_488, w_052_489, w_052_490, w_052_491, w_052_492, w_052_493, w_052_494, w_052_496, w_052_497, w_052_498, w_052_499, w_052_500, w_052_501, w_052_502, w_052_503, w_052_504, w_052_505, w_052_506, w_052_507, w_052_509, w_052_510, w_052_511, w_052_512, w_052_513, w_052_514, w_052_515, w_052_516, w_052_517, w_052_518, w_052_519, w_052_520, w_052_521, w_052_522, w_052_523, w_052_524, w_052_525, w_052_526, w_052_527, w_052_528, w_052_529, w_052_530, w_052_531, w_052_532, w_052_533, w_052_534, w_052_535, w_052_536, w_052_537, w_052_538, w_052_539, w_052_540, w_052_541, w_052_542, w_052_543, w_052_544, w_052_545, w_052_546, w_052_547, w_052_548, w_052_549, w_052_550, w_052_551, w_052_552, w_052_553, w_052_554, w_052_555, w_052_556, w_052_557, w_052_558, w_052_559, w_052_560, w_052_561, w_052_562, w_052_563, w_052_564, w_052_565, w_052_566, w_052_567, w_052_568, w_052_569, w_052_570, w_052_571, w_052_572, w_052_573, w_052_574, w_052_575, w_052_576, w_052_577, w_052_578, w_052_579, w_052_580, w_052_581, w_052_582, w_052_583, w_052_584, w_052_585, w_052_586, w_052_587, w_052_588, w_052_589, w_052_590, w_052_591, w_052_592, w_052_593, w_052_594, w_052_595, w_052_596, w_052_597, w_052_598, w_052_599, w_052_600, w_052_601, w_052_602, w_052_603, w_052_604, w_052_605, w_052_606, w_052_607, w_052_608, w_052_609, w_052_610, w_052_611, w_052_613, w_052_614, w_052_615, w_052_616, w_052_617, w_052_618, w_052_619, w_052_620, w_052_622, w_052_623, w_052_624, w_052_625, w_052_626, w_052_627, w_052_628, w_052_629, w_052_630, w_052_631, w_052_632, w_052_633, w_052_634, w_052_635, w_052_636, w_052_637, w_052_638, w_052_639, w_052_640, w_052_642, w_052_643, w_052_644, w_052_645, w_052_646, w_052_647, w_052_648, w_052_649, w_052_650, w_052_651, w_052_653, w_052_654, w_052_655, w_052_656, w_052_657, w_052_658, w_052_659, w_052_660, w_052_661, w_052_662, w_052_663, w_052_664, w_052_665, w_052_666, w_052_668, w_052_669, w_052_670, w_052_671, w_052_672, w_052_673, w_052_674, w_052_675, w_052_676, w_052_677, w_052_678, w_052_679, w_052_680, w_052_681, w_052_682, w_052_683, w_052_684, w_052_685, w_052_686, w_052_688, w_052_689, w_052_690, w_052_691, w_052_692, w_052_693, w_052_694, w_052_695, w_052_696, w_052_697, w_052_698, w_052_700, w_052_701, w_052_702, w_052_704, w_052_706, w_052_707, w_052_708, w_052_709, w_052_710, w_052_711, w_052_712, w_052_713, w_052_714, w_052_715, w_052_716, w_052_717, w_052_718, w_052_719, w_052_720, w_052_721, w_052_722, w_052_723, w_052_724, w_052_725, w_052_726, w_052_727, w_052_728, w_052_729, w_052_730, w_052_731, w_052_732, w_052_733, w_052_734, w_052_735, w_052_736, w_052_737, w_052_738, w_052_739, w_052_740, w_052_741, w_052_742, w_052_743, w_052_745, w_052_747, w_052_748, w_052_749, w_052_750, w_052_751, w_052_752, w_052_753, w_052_754, w_052_755, w_052_756, w_052_757, w_052_758, w_052_759, w_052_760, w_052_761, w_052_762, w_052_763, w_052_764, w_052_765, w_052_766, w_052_767, w_052_768, w_052_769, w_052_770, w_052_771, w_052_773, w_052_774, w_052_775, w_052_776, w_052_777, w_052_778, w_052_779, w_052_780, w_052_781, w_052_782, w_052_783, w_052_784, w_052_785, w_052_786, w_052_787, w_052_788, w_052_789, w_052_790, w_052_791, w_052_792, w_052_793, w_052_794, w_052_795, w_052_796, w_052_797, w_052_798, w_052_799, w_052_800, w_052_801, w_052_802, w_052_803, w_052_804, w_052_805, w_052_806, w_052_807, w_052_808, w_052_809, w_052_810, w_052_811, w_052_812, w_052_814, w_052_815, w_052_816, w_052_817, w_052_819, w_052_820, w_052_822, w_052_823, w_052_824, w_052_825, w_052_827, w_052_828, w_052_829, w_052_830, w_052_833, w_052_834, w_052_835, w_052_836, w_052_837, w_052_838, w_052_839, w_052_840, w_052_841, w_052_842, w_052_843, w_052_844, w_052_845, w_052_846, w_052_847, w_052_848, w_052_849, w_052_850, w_052_851, w_052_852, w_052_853, w_052_854, w_052_856, w_052_857, w_052_859, w_052_860, w_052_861, w_052_862, w_052_863, w_052_864, w_052_865, w_052_866, w_052_867, w_052_868, w_052_869, w_052_870, w_052_871, w_052_872, w_052_873, w_052_874, w_052_875, w_052_876, w_052_877, w_052_878, w_052_879, w_052_880, w_052_881, w_052_882, w_052_883, w_052_884, w_052_885, w_052_886, w_052_887, w_052_888, w_052_889, w_052_890, w_052_891, w_052_892, w_052_893, w_052_894, w_052_895, w_052_897, w_052_898, w_052_899, w_052_900, w_052_901, w_052_902, w_052_903, w_052_904, w_052_905, w_052_906, w_052_908, w_052_909, w_052_910, w_052_911, w_052_912, w_052_913, w_052_914, w_052_915, w_052_916, w_052_918, w_052_919, w_052_920, w_052_922, w_052_923, w_052_924, w_052_925, w_052_926, w_052_927, w_052_928, w_052_929, w_052_930, w_052_931, w_052_932, w_052_934, w_052_935, w_052_936, w_052_937, w_052_938, w_052_939, w_052_940, w_052_941, w_052_942, w_052_943, w_052_944, w_052_945, w_052_946, w_052_947, w_052_948, w_052_949, w_052_950, w_052_951, w_052_952, w_052_953, w_052_954, w_052_955, w_052_956, w_052_957, w_052_958, w_052_959, w_052_960, w_052_961, w_052_962, w_052_963, w_052_964, w_052_965, w_052_966, w_052_968, w_052_969, w_052_970, w_052_971, w_052_972, w_052_973, w_052_974, w_052_976, w_052_977, w_052_978, w_052_979, w_052_980, w_052_981, w_052_982, w_052_983, w_052_986, w_052_987, w_052_988, w_052_989, w_052_990, w_052_991, w_052_992, w_052_993, w_052_994, w_052_995, w_052_996, w_052_997, w_052_998, w_052_999, w_052_1001, w_052_1002, w_052_1003, w_052_1004, w_052_1005, w_052_1006, w_052_1007, w_052_1008, w_052_1009, w_052_1010, w_052_1011, w_052_1012, w_052_1013, w_052_1014, w_052_1016, w_052_1017, w_052_1018, w_052_1019, w_052_1020, w_052_1021, w_052_1022, w_052_1023, w_052_1024, w_052_1026, w_052_1027, w_052_1028, w_052_1029, w_052_1030, w_052_1031, w_052_1032, w_052_1033, w_052_1034, w_052_1035, w_052_1036, w_052_1037, w_052_1038, w_052_1039, w_052_1040, w_052_1041, w_052_1042, w_052_1043, w_052_1044, w_052_1045, w_052_1047, w_052_1048, w_052_1050, w_052_1051, w_052_1052, w_052_1053, w_052_1054, w_052_1056, w_052_1057, w_052_1058, w_052_1060, w_052_1062, w_052_1063, w_052_1066, w_052_1067, w_052_1068, w_052_1069, w_052_1070, w_052_1071, w_052_1072, w_052_1073, w_052_1074, w_052_1075, w_052_1076, w_052_1077, w_052_1078, w_052_1079, w_052_1080, w_052_1081, w_052_1082, w_052_1083, w_052_1084, w_052_1085, w_052_1087, w_052_1088, w_052_1089, w_052_1090, w_052_1092, w_052_1093, w_052_1094, w_052_1095, w_052_1096, w_052_1097, w_052_1098, w_052_1101, w_052_1102, w_052_1103, w_052_1104, w_052_1105, w_052_1106, w_052_1107, w_052_1108, w_052_1109, w_052_1110, w_052_1111, w_052_1112, w_052_1113, w_052_1114, w_052_1115, w_052_1116, w_052_1117, w_052_1118, w_052_1119, w_052_1120, w_052_1121, w_052_1122, w_052_1123, w_052_1124, w_052_1126, w_052_1127, w_052_1128, w_052_1129, w_052_1130, w_052_1131, w_052_1132, w_052_1133, w_052_1134, w_052_1135, w_052_1136, w_052_1137, w_052_1138, w_052_1139, w_052_1140, w_052_1141, w_052_1142, w_052_1143, w_052_1144, w_052_1145, w_052_1146, w_052_1147, w_052_1148, w_052_1149, w_052_1150, w_052_1151, w_052_1152, w_052_1153, w_052_1154, w_052_1155, w_052_1156, w_052_1157, w_052_1158, w_052_1159, w_052_1160, w_052_1161, w_052_1162, w_052_1163, w_052_1164, w_052_1165, w_052_1166, w_052_1167, w_052_1168, w_052_1169, w_052_1170, w_052_1171, w_052_1172, w_052_1173, w_052_1175, w_052_1176, w_052_1177, w_052_1178, w_052_1179, w_052_1180, w_052_1181, w_052_1182, w_052_1183, w_052_1184, w_052_1185, w_052_1186, w_052_1187, w_052_1188, w_052_1189, w_052_1191, w_052_1192, w_052_1193, w_052_1194, w_052_1195, w_052_1197, w_052_1198, w_052_1199, w_052_1200, w_052_1202, w_052_1203, w_052_1204, w_052_1205, w_052_1206, w_052_1207, w_052_1208, w_052_1209, w_052_1210, w_052_1211, w_052_1212, w_052_1213, w_052_1214, w_052_1215, w_052_1216, w_052_1217, w_052_1218, w_052_1221, w_052_1222, w_052_1223, w_052_1224, w_052_1225, w_052_1226, w_052_1227, w_052_1228, w_052_1229, w_052_1230, w_052_1232, w_052_1233, w_052_1234, w_052_1235, w_052_1237, w_052_1238, w_052_1239, w_052_1241, w_052_1242, w_052_1243, w_052_1244, w_052_1245, w_052_1246, w_052_1247, w_052_1248, w_052_1249, w_052_1250, w_052_1251, w_052_1252, w_052_1253, w_052_1255, w_052_1256, w_052_1257, w_052_1258, w_052_1259, w_052_1260, w_052_1261, w_052_1262, w_052_1263, w_052_1264, w_052_1265, w_052_1266, w_052_1267, w_052_1269, w_052_1270, w_052_1271, w_052_1272, w_052_1273, w_052_1274, w_052_1275, w_052_1276, w_052_1277, w_052_1278, w_052_1279, w_052_1280, w_052_1281, w_052_1282, w_052_1283, w_052_1284, w_052_1286, w_052_1287, w_052_1289, w_052_1291, w_052_1292, w_052_1293, w_052_1294, w_052_1295, w_052_1296, w_052_1297, w_052_1298, w_052_1299, w_052_1300, w_052_1301, w_052_1302, w_052_1303, w_052_1304, w_052_1305, w_052_1306, w_052_1307, w_052_1308, w_052_1309, w_052_1311, w_052_1312, w_052_1313, w_052_1314, w_052_1315, w_052_1316, w_052_1317, w_052_1318, w_052_1319, w_052_1320, w_052_1321, w_052_1322, w_052_1324, w_052_1325, w_052_1326, w_052_1327, w_052_1328, w_052_1329, w_052_1330, w_052_1331, w_052_1332, w_052_1333, w_052_1334, w_052_1336, w_052_1337, w_052_1338, w_052_1339, w_052_1340, w_052_1341, w_052_1342, w_052_1343, w_052_1345, w_052_1346, w_052_1347, w_052_1348, w_052_1349, w_052_1350, w_052_1351, w_052_1352, w_052_1353, w_052_1354, w_052_1355, w_052_1357, w_052_1358, w_052_1360, w_052_1361, w_052_1362, w_052_1363, w_052_1364, w_052_1365, w_052_1366, w_052_1367, w_052_1368, w_052_1369, w_052_1370, w_052_1372, w_052_1373, w_052_1374, w_052_1375, w_052_1376, w_052_1377, w_052_1378, w_052_1379, w_052_1380, w_052_1381, w_052_1382, w_052_1383, w_052_1384, w_052_1386, w_052_1387, w_052_1388, w_052_1389, w_052_1390, w_052_1391, w_052_1392, w_052_1393, w_052_1394, w_052_1395, w_052_1396, w_052_1397, w_052_1398, w_052_1399, w_052_1400, w_052_1401, w_052_1402, w_052_1403, w_052_1404, w_052_1405, w_052_1406, w_052_1407, w_052_1408, w_052_1409, w_052_1410, w_052_1411, w_052_1412, w_052_1413, w_052_1414, w_052_1415, w_052_1416, w_052_1417, w_052_1418, w_052_1419, w_052_1420, w_052_1421, w_052_1422, w_052_1423, w_052_1424, w_052_1425, w_052_1426, w_052_1427, w_052_1428, w_052_1429, w_052_1430, w_052_1431, w_052_1432, w_052_1434, w_052_1435, w_052_1436, w_052_1437, w_052_1438, w_052_1439, w_052_1440, w_052_1441, w_052_1442, w_052_1443, w_052_1444, w_052_1445, w_052_1446, w_052_1447, w_052_1448, w_052_1449, w_052_1450, w_052_1451, w_052_1452, w_052_1453, w_052_1454, w_052_1455, w_052_1456, w_052_1457, w_052_1458, w_052_1459, w_052_1460, w_052_1461, w_052_1462, w_052_1463, w_052_1464, w_052_1465, w_052_1466, w_052_1467, w_052_1468, w_052_1469, w_052_1470, w_052_1471, w_052_1472, w_052_1473, w_052_1475, w_052_1476, w_052_1477, w_052_1479, w_052_1480, w_052_1481, w_052_1482, w_052_1483, w_052_1485, w_052_1487, w_052_1488, w_052_1489, w_052_1490, w_052_1491, w_052_1492, w_052_1493, w_052_1494, w_052_1495, w_052_1496, w_052_1497, w_052_1498, w_052_1499, w_052_1500, w_052_1501, w_052_1502, w_052_1503, w_052_1504, w_052_1505, w_052_1506, w_052_1508, w_052_1509, w_052_1510, w_052_1511, w_052_1512, w_052_1513, w_052_1515, w_052_1516, w_052_1517, w_052_1518, w_052_1519, w_052_1520, w_052_1521, w_052_1522, w_052_1523, w_052_1524, w_052_1526, w_052_1527, w_052_1528, w_052_1529, w_052_1530, w_052_1531, w_052_1532, w_052_1533, w_052_1534, w_052_1536, w_052_1537, w_052_1538, w_052_1540, w_052_1541, w_052_1543, w_052_1544, w_052_1545, w_052_1546, w_052_1547, w_052_1548, w_052_1549, w_052_1550, w_052_1551, w_052_1552, w_052_1553, w_052_1554, w_052_1555, w_052_1556, w_052_1557, w_052_1558, w_052_1559, w_052_1560, w_052_1561, w_052_1562, w_052_1563, w_052_1564, w_052_1565, w_052_1566, w_052_1567, w_052_1568, w_052_1569, w_052_1570, w_052_1571, w_052_1572, w_052_1573, w_052_1574, w_052_1576, w_052_1577, w_052_1578, w_052_1579, w_052_1580, w_052_1582, w_052_1583, w_052_1584, w_052_1585, w_052_1586, w_052_1587, w_052_1588, w_052_1589, w_052_1590, w_052_1591, w_052_1592, w_052_1593, w_052_1594, w_052_1595, w_052_1596, w_052_1597, w_052_1598, w_052_1599, w_052_1600, w_052_1601, w_052_1602, w_052_1603, w_052_1604, w_052_1605, w_052_1606, w_052_1607, w_052_1608, w_052_1609, w_052_1610, w_052_1611, w_052_1612, w_052_1613, w_052_1614, w_052_1615, w_052_1616, w_052_1617, w_052_1618, w_052_1619, w_052_1620, w_052_1621, w_052_1622, w_052_1623, w_052_1624, w_052_1625, w_052_1626, w_052_1627, w_052_1628, w_052_1629, w_052_1630, w_052_1631, w_052_1632, w_052_1633, w_052_1634, w_052_1635, w_052_1636, w_052_1637, w_052_1638, w_052_1639, w_052_1640, w_052_1641, w_052_1642, w_052_1643, w_052_1644, w_052_1645, w_052_1646, w_052_1647, w_052_1648, w_052_1649, w_052_1650, w_052_1651, w_052_1652, w_052_1653, w_052_1654, w_052_1655, w_052_1656, w_052_1657, w_052_1658, w_052_1659, w_052_1660, w_052_1661, w_052_1662, w_052_1663, w_052_1664, w_052_1665, w_052_1666, w_052_1668, w_052_1669, w_052_1670, w_052_1671, w_052_1672, w_052_1673, w_052_1674, w_052_1675, w_052_1677, w_052_1678, w_052_1679, w_052_1680, w_052_1681, w_052_1682, w_052_1683, w_052_1684, w_052_1685, w_052_1686, w_052_1687, w_052_1688, w_052_1689, w_052_1690, w_052_1692, w_052_1693, w_052_1694, w_052_1695, w_052_1696, w_052_1697, w_052_1698, w_052_1699, w_052_1700, w_052_1701, w_052_1702, w_052_1703, w_052_1704, w_052_1705, w_052_1706, w_052_1707, w_052_1708, w_052_1709, w_052_1710, w_052_1711, w_052_1712, w_052_1713, w_052_1714, w_052_1716, w_052_1717, w_052_1719, w_052_1720, w_052_1721, w_052_1722, w_052_1723, w_052_1724, w_052_1725, w_052_1726, w_052_1727, w_052_1728, w_052_1729, w_052_1731, w_052_1732, w_052_1733, w_052_1734, w_052_1735, w_052_1737, w_052_1738, w_052_1739, w_052_1740, w_052_1741, w_052_1743, w_052_1744, w_052_1745, w_052_1746, w_052_1747, w_052_1748, w_052_1750, w_052_1752, w_052_1753, w_052_1754, w_052_1756, w_052_1757, w_052_1758, w_052_1759, w_052_1760, w_052_1761, w_052_1763, w_052_1764, w_052_1765, w_052_1766, w_052_1767, w_052_1768, w_052_1769, w_052_1770, w_052_1771, w_052_1772, w_052_1773, w_052_1774, w_052_1775, w_052_1776, w_052_1778, w_052_1779, w_052_1780, w_052_1781, w_052_1782, w_052_1783, w_052_1784, w_052_1785, w_052_1787, w_052_1788, w_052_1789, w_052_1790, w_052_1791, w_052_1793, w_052_1794, w_052_1795, w_052_1796, w_052_1797, w_052_1798, w_052_1799, w_052_1800, w_052_1801, w_052_1802, w_052_1803, w_052_1804, w_052_1805, w_052_1806, w_052_1807, w_052_1808, w_052_1809, w_052_1810, w_052_1811, w_052_1812, w_052_1813, w_052_1814, w_052_1815, w_052_1816, w_052_1817, w_052_1819, w_052_1821, w_052_1822, w_052_1823, w_052_1824, w_052_1825, w_052_1826, w_052_1827, w_052_1828, w_052_1830, w_052_1831, w_052_1832, w_052_1833, w_052_1834, w_052_1835, w_052_1836, w_052_1837, w_052_1838, w_052_1839, w_052_1840, w_052_1841, w_052_1842, w_052_1843, w_052_1844, w_052_1845, w_052_1846, w_052_1847, w_052_1848, w_052_1849, w_052_1850, w_052_1851, w_052_1852, w_052_1854, w_052_1855, w_052_1856, w_052_1857, w_052_1858, w_052_1859, w_052_1860, w_052_1861, w_052_1862, w_052_1863, w_052_1864, w_052_1865, w_052_1866, w_052_1867, w_052_1868, w_052_1869, w_052_1870, w_052_1871, w_052_1872, w_052_1873, w_052_1874, w_052_1875, w_052_1876, w_052_1877, w_052_1878, w_052_1879, w_052_1880, w_052_1881, w_052_1882, w_052_1883, w_052_1885, w_052_1886, w_052_1887, w_052_1888, w_052_1889, w_052_1890, w_052_1891, w_052_1892, w_052_1893, w_052_1894, w_052_1895, w_052_1896, w_052_1897, w_052_1898, w_052_1899, w_052_1900, w_052_1901, w_052_1902, w_052_1903, w_052_1904, w_052_1905, w_052_1908, w_052_1909, w_052_1910, w_052_1911, w_052_1912, w_052_1913, w_052_1914, w_052_1915, w_052_1916, w_052_1917, w_052_1918, w_052_1919, w_052_1920, w_052_1921, w_052_1922, w_052_1923, w_052_1924, w_052_1925, w_052_1926, w_052_1927, w_052_1928, w_052_1929, w_052_1930, w_052_1931, w_052_1932, w_052_1933;
  wire w_053_001, w_053_002, w_053_003, w_053_004, w_053_006, w_053_007, w_053_008, w_053_009, w_053_012, w_053_013, w_053_014, w_053_016, w_053_017, w_053_020, w_053_021, w_053_022, w_053_025, w_053_027, w_053_030, w_053_031, w_053_032, w_053_035, w_053_036, w_053_037, w_053_038, w_053_040, w_053_042, w_053_044, w_053_046, w_053_047, w_053_048, w_053_049, w_053_050, w_053_052, w_053_053, w_053_055, w_053_056, w_053_057, w_053_059, w_053_061, w_053_064, w_053_065, w_053_067, w_053_069, w_053_070, w_053_071, w_053_072, w_053_074, w_053_077, w_053_078, w_053_080, w_053_081, w_053_082, w_053_085, w_053_086, w_053_087, w_053_089, w_053_090, w_053_091, w_053_092, w_053_093, w_053_097, w_053_099, w_053_100, w_053_101, w_053_103, w_053_104, w_053_105, w_053_106, w_053_110, w_053_113, w_053_114, w_053_116, w_053_117, w_053_118, w_053_121, w_053_123, w_053_124, w_053_125, w_053_126, w_053_127, w_053_129, w_053_130, w_053_131, w_053_132, w_053_133, w_053_135, w_053_136, w_053_137, w_053_138, w_053_140, w_053_141, w_053_142, w_053_143, w_053_146, w_053_147, w_053_149, w_053_152, w_053_154, w_053_155, w_053_157, w_053_161, w_053_162, w_053_163, w_053_164, w_053_165, w_053_166, w_053_169, w_053_170, w_053_172, w_053_173, w_053_174, w_053_175, w_053_177, w_053_180, w_053_184, w_053_185, w_053_186, w_053_187, w_053_188, w_053_192, w_053_193, w_053_197, w_053_199, w_053_200, w_053_201, w_053_202, w_053_203, w_053_204, w_053_205, w_053_206, w_053_207, w_053_208, w_053_209, w_053_210, w_053_211, w_053_212, w_053_213, w_053_214, w_053_215, w_053_216, w_053_217, w_053_218, w_053_220, w_053_223, w_053_224, w_053_228, w_053_229, w_053_230, w_053_232, w_053_234, w_053_236, w_053_239, w_053_241, w_053_243, w_053_245, w_053_247, w_053_248, w_053_251, w_053_252, w_053_254, w_053_256, w_053_257, w_053_259, w_053_260, w_053_261, w_053_262, w_053_265, w_053_266, w_053_268, w_053_269, w_053_270, w_053_271, w_053_272, w_053_273, w_053_274, w_053_275, w_053_277, w_053_278, w_053_279, w_053_281, w_053_282, w_053_283, w_053_284, w_053_286, w_053_288, w_053_289, w_053_291, w_053_292, w_053_295, w_053_296, w_053_298, w_053_299, w_053_300, w_053_302, w_053_304, w_053_305, w_053_306, w_053_309, w_053_310, w_053_314, w_053_317, w_053_318, w_053_319, w_053_322, w_053_323, w_053_326, w_053_327, w_053_328, w_053_330, w_053_331, w_053_332, w_053_336, w_053_338, w_053_339, w_053_342, w_053_345, w_053_347, w_053_350, w_053_351, w_053_353, w_053_354, w_053_355, w_053_356, w_053_357, w_053_358, w_053_359, w_053_361, w_053_363, w_053_367, w_053_369, w_053_371, w_053_373, w_053_374, w_053_375, w_053_377, w_053_378, w_053_380, w_053_381, w_053_382, w_053_383, w_053_386, w_053_393, w_053_397, w_053_398, w_053_400, w_053_401, w_053_403, w_053_405, w_053_406, w_053_408, w_053_410, w_053_412, w_053_419, w_053_422, w_053_423, w_053_424, w_053_425, w_053_430, w_053_431, w_053_432, w_053_438, w_053_439, w_053_441, w_053_442, w_053_443, w_053_444, w_053_445, w_053_449, w_053_450, w_053_452, w_053_453, w_053_455, w_053_457, w_053_458, w_053_459, w_053_460, w_053_462, w_053_463, w_053_464, w_053_467, w_053_469, w_053_470, w_053_472, w_053_473, w_053_475, w_053_476, w_053_477, w_053_478, w_053_479, w_053_480, w_053_482, w_053_483, w_053_486, w_053_488, w_053_490, w_053_493, w_053_495, w_053_496, w_053_497, w_053_498, w_053_499, w_053_500, w_053_502, w_053_504, w_053_505, w_053_507, w_053_508, w_053_509, w_053_510, w_053_515, w_053_516, w_053_518, w_053_519, w_053_520, w_053_524, w_053_525, w_053_533, w_053_534, w_053_535, w_053_537, w_053_538, w_053_540, w_053_541, w_053_543, w_053_546, w_053_547, w_053_548, w_053_549, w_053_550, w_053_552, w_053_553, w_053_555, w_053_556, w_053_557, w_053_558, w_053_561, w_053_563, w_053_564, w_053_565, w_053_568, w_053_569, w_053_571, w_053_572, w_053_573, w_053_574, w_053_575, w_053_576, w_053_577, w_053_579, w_053_580, w_053_581, w_053_583, w_053_584, w_053_585, w_053_586, w_053_587, w_053_589, w_053_590, w_053_591, w_053_592, w_053_593, w_053_594, w_053_595, w_053_597, w_053_598, w_053_599, w_053_601, w_053_603, w_053_604, w_053_607, w_053_608, w_053_609, w_053_610, w_053_612, w_053_613, w_053_614, w_053_615, w_053_616, w_053_617, w_053_619, w_053_620, w_053_623, w_053_624, w_053_625, w_053_626, w_053_629, w_053_630, w_053_633, w_053_634, w_053_635, w_053_636, w_053_637, w_053_638, w_053_640, w_053_641, w_053_642, w_053_643, w_053_645, w_053_646, w_053_647, w_053_648, w_053_649, w_053_650, w_053_651, w_053_652, w_053_656, w_053_659, w_053_660, w_053_661, w_053_662, w_053_663, w_053_664, w_053_665, w_053_666, w_053_668, w_053_669, w_053_670, w_053_671, w_053_672, w_053_673, w_053_674, w_053_675, w_053_677, w_053_679, w_053_680, w_053_681, w_053_682, w_053_686, w_053_689, w_053_691, w_053_693, w_053_695, w_053_697, w_053_699, w_053_700, w_053_702, w_053_703, w_053_704, w_053_705, w_053_706, w_053_707, w_053_709, w_053_710, w_053_711, w_053_713, w_053_718, w_053_719, w_053_721, w_053_722, w_053_723, w_053_724, w_053_726, w_053_727, w_053_731, w_053_733, w_053_734, w_053_736, w_053_738, w_053_739, w_053_740, w_053_741, w_053_743, w_053_744, w_053_745, w_053_746, w_053_748, w_053_750, w_053_753, w_053_755, w_053_757, w_053_758, w_053_759, w_053_760, w_053_761, w_053_762, w_053_763, w_053_764, w_053_765, w_053_767, w_053_768, w_053_770, w_053_773, w_053_774, w_053_776, w_053_778, w_053_779, w_053_781, w_053_782, w_053_783, w_053_784, w_053_786, w_053_787, w_053_789, w_053_790, w_053_791, w_053_792, w_053_794, w_053_795, w_053_796, w_053_797, w_053_799, w_053_800, w_053_803, w_053_804, w_053_806, w_053_808, w_053_809, w_053_810, w_053_811, w_053_812, w_053_815, w_053_816, w_053_817, w_053_820, w_053_821, w_053_822, w_053_823, w_053_824, w_053_825, w_053_826, w_053_827, w_053_828, w_053_829, w_053_830, w_053_831, w_053_834, w_053_836, w_053_838, w_053_840, w_053_841, w_053_842, w_053_843, w_053_844, w_053_848, w_053_849, w_053_850, w_053_852, w_053_855, w_053_856, w_053_857, w_053_859, w_053_860, w_053_861, w_053_862, w_053_863, w_053_865, w_053_866, w_053_867, w_053_868, w_053_869, w_053_872, w_053_874, w_053_875, w_053_877, w_053_878, w_053_879, w_053_880, w_053_882, w_053_883, w_053_887, w_053_888, w_053_890, w_053_892, w_053_893, w_053_895, w_053_897, w_053_899, w_053_901, w_053_903, w_053_905, w_053_907, w_053_908, w_053_912, w_053_913, w_053_914, w_053_916, w_053_918, w_053_922, w_053_923, w_053_924, w_053_925, w_053_927, w_053_929, w_053_930, w_053_933, w_053_934, w_053_937, w_053_938, w_053_939, w_053_940, w_053_941, w_053_942, w_053_945, w_053_946, w_053_947, w_053_948, w_053_950, w_053_952, w_053_953, w_053_954, w_053_956, w_053_957, w_053_959, w_053_960, w_053_961, w_053_962, w_053_963, w_053_966, w_053_967, w_053_968, w_053_969, w_053_970, w_053_975, w_053_976, w_053_977, w_053_980, w_053_983, w_053_984, w_053_985, w_053_986, w_053_988, w_053_989, w_053_993, w_053_994, w_053_996, w_053_998, w_053_1000, w_053_1001, w_053_1002, w_053_1004, w_053_1005, w_053_1006, w_053_1007, w_053_1008, w_053_1009, w_053_1010, w_053_1011, w_053_1012, w_053_1016, w_053_1018, w_053_1019, w_053_1020, w_053_1022, w_053_1023, w_053_1026, w_053_1029, w_053_1031, w_053_1032, w_053_1033, w_053_1034, w_053_1037, w_053_1040, w_053_1041, w_053_1042, w_053_1044, w_053_1045, w_053_1047, w_053_1048, w_053_1049, w_053_1050, w_053_1052, w_053_1056, w_053_1057, w_053_1060, w_053_1061, w_053_1062, w_053_1063, w_053_1065, w_053_1066, w_053_1067, w_053_1068, w_053_1069, w_053_1070, w_053_1071, w_053_1072, w_053_1073, w_053_1075, w_053_1076, w_053_1077, w_053_1081, w_053_1082, w_053_1087, w_053_1089, w_053_1090, w_053_1091, w_053_1094, w_053_1098, w_053_1100, w_053_1102, w_053_1104, w_053_1105, w_053_1106, w_053_1110, w_053_1111, w_053_1114, w_053_1115, w_053_1119, w_053_1121, w_053_1122, w_053_1123, w_053_1124, w_053_1125, w_053_1126, w_053_1129, w_053_1131, w_053_1132, w_053_1138, w_053_1140, w_053_1143, w_053_1145, w_053_1146, w_053_1148, w_053_1150, w_053_1154, w_053_1156, w_053_1158, w_053_1159, w_053_1161, w_053_1162, w_053_1164, w_053_1165, w_053_1167, w_053_1169, w_053_1171, w_053_1172, w_053_1174, w_053_1175, w_053_1181, w_053_1182, w_053_1183, w_053_1184, w_053_1185, w_053_1186, w_053_1189, w_053_1190, w_053_1191, w_053_1192, w_053_1193, w_053_1194, w_053_1196, w_053_1199, w_053_1200, w_053_1201, w_053_1202, w_053_1205, w_053_1207, w_053_1209, w_053_1212, w_053_1220, w_053_1221, w_053_1222, w_053_1226, w_053_1227, w_053_1228, w_053_1231, w_053_1232, w_053_1233, w_053_1235, w_053_1238, w_053_1239, w_053_1241, w_053_1242, w_053_1244, w_053_1245, w_053_1249, w_053_1250, w_053_1251, w_053_1252, w_053_1253, w_053_1254, w_053_1255, w_053_1257, w_053_1258, w_053_1261, w_053_1262, w_053_1266, w_053_1268, w_053_1269, w_053_1270, w_053_1271, w_053_1272, w_053_1273, w_053_1274, w_053_1275, w_053_1276, w_053_1277, w_053_1279, w_053_1280, w_053_1283, w_053_1284, w_053_1287, w_053_1288, w_053_1289, w_053_1290, w_053_1291, w_053_1292, w_053_1295, w_053_1296, w_053_1297, w_053_1298, w_053_1300, w_053_1301, w_053_1302, w_053_1303, w_053_1304, w_053_1305, w_053_1306, w_053_1307, w_053_1308, w_053_1309, w_053_1310, w_053_1311, w_053_1313, w_053_1314, w_053_1316, w_053_1317, w_053_1318, w_053_1319, w_053_1320, w_053_1321, w_053_1322, w_053_1323, w_053_1324, w_053_1325, w_053_1327, w_053_1328, w_053_1329, w_053_1331, w_053_1333, w_053_1335, w_053_1336, w_053_1338, w_053_1340, w_053_1342, w_053_1343, w_053_1344, w_053_1347, w_053_1348, w_053_1349, w_053_1350, w_053_1351, w_053_1353, w_053_1354, w_053_1357, w_053_1361, w_053_1363, w_053_1365, w_053_1366, w_053_1367, w_053_1368, w_053_1374, w_053_1377, w_053_1379, w_053_1380, w_053_1381, w_053_1382, w_053_1387, w_053_1388, w_053_1389, w_053_1390, w_053_1393, w_053_1395, w_053_1399, w_053_1400, w_053_1401, w_053_1402, w_053_1403, w_053_1404, w_053_1405, w_053_1406, w_053_1407, w_053_1409, w_053_1410, w_053_1411, w_053_1413, w_053_1415, w_053_1418, w_053_1419, w_053_1422, w_053_1423, w_053_1424, w_053_1426, w_053_1427, w_053_1429, w_053_1431, w_053_1432, w_053_1433, w_053_1434, w_053_1435, w_053_1437, w_053_1442, w_053_1443, w_053_1444, w_053_1446, w_053_1447, w_053_1448, w_053_1449, w_053_1453, w_053_1454, w_053_1455, w_053_1457, w_053_1458, w_053_1459, w_053_1460, w_053_1461, w_053_1462, w_053_1463, w_053_1464, w_053_1467, w_053_1470, w_053_1471, w_053_1472, w_053_1473, w_053_1474, w_053_1477, w_053_1479, w_053_1484, w_053_1485, w_053_1489, w_053_1490, w_053_1491, w_053_1493, w_053_1494, w_053_1495, w_053_1496, w_053_1498, w_053_1499, w_053_1500, w_053_1501, w_053_1503, w_053_1504, w_053_1505, w_053_1507, w_053_1508, w_053_1509, w_053_1510, w_053_1514, w_053_1515, w_053_1516, w_053_1518, w_053_1519, w_053_1520, w_053_1521, w_053_1522, w_053_1524, w_053_1526, w_053_1530, w_053_1531, w_053_1532, w_053_1533, w_053_1535, w_053_1536, w_053_1540, w_053_1541, w_053_1543, w_053_1551, w_053_1552, w_053_1553, w_053_1554, w_053_1555, w_053_1557, w_053_1559, w_053_1561, w_053_1562, w_053_1563, w_053_1564, w_053_1566, w_053_1569, w_053_1573, w_053_1576, w_053_1577, w_053_1578, w_053_1579, w_053_1581, w_053_1582, w_053_1584, w_053_1585, w_053_1586, w_053_1587, w_053_1591, w_053_1594, w_053_1596, w_053_1600, w_053_1602, w_053_1603, w_053_1605, w_053_1607, w_053_1610, w_053_1613, w_053_1615, w_053_1616, w_053_1618, w_053_1619, w_053_1620, w_053_1625, w_053_1626, w_053_1628, w_053_1629, w_053_1630, w_053_1631, w_053_1633, w_053_1634, w_053_1635, w_053_1639, w_053_1640, w_053_1643, w_053_1644, w_053_1645, w_053_1646, w_053_1647, w_053_1648, w_053_1649, w_053_1652, w_053_1653, w_053_1654, w_053_1655, w_053_1656, w_053_1657, w_053_1658, w_053_1659, w_053_1661, w_053_1662, w_053_1663, w_053_1664, w_053_1665, w_053_1667, w_053_1668, w_053_1669, w_053_1670, w_053_1671, w_053_1673, w_053_1678, w_053_1679, w_053_1682, w_053_1683, w_053_1684, w_053_1685, w_053_1686, w_053_1688, w_053_1689, w_053_1693, w_053_1695, w_053_1697, w_053_1699, w_053_1700, w_053_1701, w_053_1702, w_053_1703, w_053_1704, w_053_1705, w_053_1708, w_053_1709, w_053_1710, w_053_1713, w_053_1714, w_053_1716, w_053_1717, w_053_1718, w_053_1719, w_053_1721, w_053_1722, w_053_1723, w_053_1724, w_053_1725, w_053_1726, w_053_1729, w_053_1731, w_053_1732, w_053_1734, w_053_1736, w_053_1739, w_053_1740, w_053_1744, w_053_1745, w_053_1746, w_053_1747, w_053_1748, w_053_1749, w_053_1750, w_053_1751, w_053_1752, w_053_1753, w_053_1756, w_053_1759, w_053_1762, w_053_1763, w_053_1765, w_053_1766, w_053_1767, w_053_1769, w_053_1770, w_053_1771, w_053_1773, w_053_1774, w_053_1775, w_053_1778, w_053_1779, w_053_1780, w_053_1781, w_053_1782, w_053_1785, w_053_1786, w_053_1788, w_053_1789, w_053_1790, w_053_1791, w_053_1792, w_053_1793, w_053_1794, w_053_1796, w_053_1797, w_053_1798, w_053_1799, w_053_1801, w_053_1802, w_053_1803, w_053_1805, w_053_1806, w_053_1807, w_053_1810, w_053_1811, w_053_1812, w_053_1813, w_053_1814, w_053_1818, w_053_1820, w_053_1821, w_053_1824, w_053_1825, w_053_1827, w_053_1832, w_053_1833, w_053_1834, w_053_1836, w_053_1839, w_053_1840, w_053_1841, w_053_1842, w_053_1845, w_053_1847, w_053_1848, w_053_1849, w_053_1850, w_053_1851, w_053_1853, w_053_1854, w_053_1857, w_053_1858, w_053_1859, w_053_1860, w_053_1861, w_053_1863, w_053_1864, w_053_1865, w_053_1866, w_053_1868, w_053_1870, w_053_1871, w_053_1872, w_053_1875, w_053_1876, w_053_1877, w_053_1878, w_053_1881, w_053_1883, w_053_1886, w_053_1887, w_053_1888, w_053_1892, w_053_1893, w_053_1894, w_053_1896, w_053_1897, w_053_1898, w_053_1900, w_053_1902, w_053_1903, w_053_1904, w_053_1905, w_053_1906, w_053_1907, w_053_1908, w_053_1909, w_053_1910, w_053_1911, w_053_1912, w_053_1913, w_053_1914, w_053_1915, w_053_1918, w_053_1919, w_053_1920, w_053_1921, w_053_1924, w_053_1925, w_053_1927, w_053_1928, w_053_1929, w_053_1931, w_053_1933, w_053_1935, w_053_1936, w_053_1939, w_053_1940, w_053_1942, w_053_1944, w_053_1948, w_053_1949, w_053_1950, w_053_1951, w_053_1954, w_053_1955, w_053_1956, w_053_1957, w_053_1959, w_053_1961, w_053_1962, w_053_1963, w_053_1965, w_053_1966, w_053_1969, w_053_1971, w_053_1972, w_053_1973, w_053_1974, w_053_1975, w_053_1976, w_053_1979, w_053_1981, w_053_1982, w_053_1987, w_053_1988, w_053_1989, w_053_1991, w_053_1992, w_053_1994, w_053_1997, w_053_1998, w_053_1999, w_053_2000, w_053_2002, w_053_2003, w_053_2004, w_053_2005, w_053_2009, w_053_2011, w_053_2014, w_053_2015, w_053_2016, w_053_2017, w_053_2018, w_053_2019, w_053_2021, w_053_2022, w_053_2023, w_053_2024, w_053_2025, w_053_2028, w_053_2029, w_053_2030, w_053_2031, w_053_2032, w_053_2033, w_053_2034, w_053_2035, w_053_2036, w_053_2037, w_053_2038, w_053_2041, w_053_2042, w_053_2044, w_053_2046, w_053_2047, w_053_2048, w_053_2050, w_053_2052, w_053_2053, w_053_2054, w_053_2055, w_053_2057, w_053_2058, w_053_2059, w_053_2061, w_053_2063, w_053_2064, w_053_2065, w_053_2067, w_053_2068, w_053_2071, w_053_2072, w_053_2073, w_053_2074, w_053_2076, w_053_2077, w_053_2078, w_053_2080, w_053_2081, w_053_2083, w_053_2084, w_053_2085, w_053_2086, w_053_2087, w_053_2088, w_053_2089, w_053_2090, w_053_2091, w_053_2092, w_053_2093, w_053_2094, w_053_2095, w_053_2096, w_053_2097, w_053_2099, w_053_2100, w_053_2101, w_053_2102, w_053_2103, w_053_2104, w_053_2105, w_053_2107, w_053_2109, w_053_2110, w_053_2111, w_053_2114, w_053_2119, w_053_2120, w_053_2123, w_053_2124, w_053_2129, w_053_2130, w_053_2131, w_053_2133, w_053_2139, w_053_2140, w_053_2141, w_053_2142, w_053_2143, w_053_2144, w_053_2145, w_053_2147, w_053_2148, w_053_2151, w_053_2152, w_053_2154, w_053_2155, w_053_2156, w_053_2157, w_053_2161, w_053_2162, w_053_2163, w_053_2167, w_053_2168, w_053_2170, w_053_2171, w_053_2173, w_053_2174, w_053_2175, w_053_2176, w_053_2177, w_053_2178, w_053_2179, w_053_2180, w_053_2182, w_053_2183, w_053_2184, w_053_2186, w_053_2190, w_053_2191, w_053_2192, w_053_2193, w_053_2194, w_053_2195, w_053_2196, w_053_2197, w_053_2198, w_053_2199, w_053_2200, w_053_2201, w_053_2202, w_053_2203, w_053_2208, w_053_2209, w_053_2210, w_053_2211, w_053_2213, w_053_2215, w_053_2216, w_053_2217, w_053_2218, w_053_2220, w_053_2222, w_053_2224, w_053_2227, w_053_2228, w_053_2229, w_053_2231, w_053_2234, w_053_2235, w_053_2236, w_053_2237, w_053_2238, w_053_2239, w_053_2243, w_053_2246, w_053_2248, w_053_2249, w_053_2251, w_053_2254, w_053_2255, w_053_2256, w_053_2257, w_053_2259, w_053_2260, w_053_2261, w_053_2264, w_053_2265, w_053_2266, w_053_2267, w_053_2271, w_053_2272, w_053_2274, w_053_2275, w_053_2276, w_053_2277, w_053_2278, w_053_2282, w_053_2283, w_053_2285, w_053_2290, w_053_2291, w_053_2292, w_053_2295, w_053_2297, w_053_2298, w_053_2299, w_053_2300, w_053_2302, w_053_2306, w_053_2308, w_053_2309, w_053_2310, w_053_2311, w_053_2313, w_053_2314, w_053_2316, w_053_2317, w_053_2320, w_053_2322, w_053_2323, w_053_2325, w_053_2326, w_053_2327, w_053_2329, w_053_2332, w_053_2333, w_053_2335, w_053_2336, w_053_2337, w_053_2338, w_053_2339, w_053_2340, w_053_2341, w_053_2342, w_053_2343, w_053_2344, w_053_2345, w_053_2346, w_053_2347, w_053_2349, w_053_2350, w_053_2351, w_053_2353, w_053_2354, w_053_2358, w_053_2361, w_053_2362, w_053_2363, w_053_2365, w_053_2366, w_053_2367, w_053_2368, w_053_2370, w_053_2371, w_053_2372, w_053_2373, w_053_2374, w_053_2376, w_053_2377, w_053_2380, w_053_2384, w_053_2386, w_053_2387, w_053_2390, w_053_2392, w_053_2393, w_053_2394, w_053_2395, w_053_2397, w_053_2398, w_053_2401, w_053_2403, w_053_2404, w_053_2406, w_053_2407, w_053_2408, w_053_2410, w_053_2411, w_053_2413, w_053_2414, w_053_2415, w_053_2416, w_053_2420, w_053_2421, w_053_2422, w_053_2423, w_053_2426, w_053_2428, w_053_2432, w_053_2435, w_053_2437, w_053_2440, w_053_2443, w_053_2444, w_053_2445, w_053_2446, w_053_2447, w_053_2453, w_053_2454, w_053_2455, w_053_2456, w_053_2461, w_053_2462, w_053_2463, w_053_2464, w_053_2466, w_053_2467, w_053_2468, w_053_2469, w_053_2470, w_053_2472, w_053_2473, w_053_2474, w_053_2476, w_053_2477, w_053_2478, w_053_2482, w_053_2486, w_053_2491, w_053_2492, w_053_2494, w_053_2495, w_053_2498, w_053_2499, w_053_2500, w_053_2501, w_053_2502, w_053_2503, w_053_2506, w_053_2507, w_053_2508, w_053_2509, w_053_2510, w_053_2511, w_053_2512, w_053_2515, w_053_2516, w_053_2517, w_053_2518, w_053_2519, w_053_2521, w_053_2523, w_053_2524, w_053_2525, w_053_2527, w_053_2528, w_053_2529, w_053_2531, w_053_2532, w_053_2534, w_053_2536, w_053_2537, w_053_2538, w_053_2539, w_053_2540, w_053_2542, w_053_2544, w_053_2546, w_053_2547, w_053_2551, w_053_2552, w_053_2553, w_053_2555, w_053_2556, w_053_2557, w_053_2559, w_053_2560, w_053_2562, w_053_2564, w_053_2565, w_053_2568, w_053_2569, w_053_2573, w_053_2575, w_053_2578, w_053_2580, w_053_2582, w_053_2583, w_053_2584, w_053_2586, w_053_2587, w_053_2588, w_053_2589, w_053_2590, w_053_2591, w_053_2595, w_053_2597, w_053_2598, w_053_2599, w_053_2600, w_053_2601, w_053_2604, w_053_2605, w_053_2607, w_053_2608, w_053_2610, w_053_2611, w_053_2612, w_053_2614, w_053_2616, w_053_2618, w_053_2619, w_053_2621, w_053_2622, w_053_2625, w_053_2627, w_053_2629, w_053_2632, w_053_2635, w_053_2636, w_053_2637, w_053_2638, w_053_2639, w_053_2640, w_053_2641, w_053_2642, w_053_2643, w_053_2645, w_053_2646, w_053_2648, w_053_2649, w_053_2650, w_053_2651, w_053_2652, w_053_2655, w_053_2657, w_053_2658, w_053_2660, w_053_2661, w_053_2662, w_053_2664, w_053_2665, w_053_2666, w_053_2667, w_053_2669, w_053_2673, w_053_2674, w_053_2675, w_053_2677, w_053_2678, w_053_2679, w_053_2680, w_053_2681, w_053_2683, w_053_2684, w_053_2685, w_053_2689, w_053_2690, w_053_2692, w_053_2693, w_053_2695, w_053_2698, w_053_2700, w_053_2705, w_053_2707, w_053_2710, w_053_2713, w_053_2715, w_053_2717, w_053_2719, w_053_2720, w_053_2721, w_053_2722, w_053_2723, w_053_2728, w_053_2729, w_053_2730, w_053_2731, w_053_2733, w_053_2734, w_053_2736, w_053_2737, w_053_2738, w_053_2739, w_053_2740, w_053_2741, w_053_2745, w_053_2746, w_053_2747, w_053_2748, w_053_2749, w_053_2750, w_053_2751, w_053_2753, w_053_2754, w_053_2755, w_053_2756, w_053_2757, w_053_2758, w_053_2759, w_053_2760, w_053_2762, w_053_2763, w_053_2766, w_053_2767, w_053_2769, w_053_2770, w_053_2772, w_053_2774, w_053_2776, w_053_2778, w_053_2780, w_053_2781, w_053_2785, w_053_2787, w_053_2788, w_053_2789, w_053_2790, w_053_2792, w_053_2793, w_053_2794, w_053_2795, w_053_2799, w_053_2803, w_053_2804, w_053_2805, w_053_2807, w_053_2808, w_053_2809, w_053_2810, w_053_2811, w_053_2812, w_053_2813, w_053_2815, w_053_2818, w_053_2819, w_053_2820, w_053_2821, w_053_2822, w_053_2823, w_053_2825, w_053_2826, w_053_2827, w_053_2828, w_053_2829, w_053_2832, w_053_2833, w_053_2834, w_053_2835, w_053_2838, w_053_2839, w_053_2840, w_053_2842, w_053_2845, w_053_2848, w_053_2849, w_053_2851, w_053_2852, w_053_2853, w_053_2855, w_053_2856, w_053_2857, w_053_2860, w_053_2862, w_053_2864, w_053_2865, w_053_2866, w_053_2867, w_053_2868, w_053_2870, w_053_2871, w_053_2872, w_053_2873, w_053_2874, w_053_2875, w_053_2877, w_053_2878, w_053_2879, w_053_2880, w_053_2882, w_053_2884, w_053_2885, w_053_2886, w_053_2887, w_053_2888, w_053_2889, w_053_2890, w_053_2891, w_053_2894, w_053_2895, w_053_2896, w_053_2897, w_053_2898, w_053_2899, w_053_2900, w_053_2901, w_053_2902, w_053_2904, w_053_2906, w_053_2907, w_053_2908, w_053_2910, w_053_2914, w_053_2915, w_053_2916, w_053_2917, w_053_2919, w_053_2922, w_053_2923, w_053_2924, w_053_2925, w_053_2927, w_053_2928, w_053_2929, w_053_2930, w_053_2932, w_053_2934, w_053_2936, w_053_2937, w_053_2938, w_053_2941, w_053_2942, w_053_2944, w_053_2947, w_053_2948, w_053_2949, w_053_2950, w_053_2953, w_053_2954, w_053_2955, w_053_2956, w_053_2958, w_053_2960, w_053_2961, w_053_2964, w_053_2970, w_053_2972, w_053_2973, w_053_2974, w_053_2976, w_053_2977, w_053_2982, w_053_2984, w_053_2985, w_053_2986, w_053_2987, w_053_2989, w_053_2990, w_053_2991, w_053_2993, w_053_2995, w_053_2996, w_053_2997, w_053_2998, w_053_3000, w_053_3001, w_053_3003, w_053_3006, w_053_3010, w_053_3011, w_053_3014, w_053_3015, w_053_3016, w_053_3017, w_053_3018, w_053_3020, w_053_3022, w_053_3024, w_053_3025, w_053_3026, w_053_3027, w_053_3031, w_053_3032, w_053_3033, w_053_3035, w_053_3036, w_053_3041, w_053_3042, w_053_3044, w_053_3045, w_053_3048, w_053_3049, w_053_3053, w_053_3054, w_053_3055, w_053_3056, w_053_3058, w_053_3060, w_053_3061, w_053_3062, w_053_3063, w_053_3064, w_053_3065, w_053_3066, w_053_3068, w_053_3069, w_053_3070, w_053_3071, w_053_3072, w_053_3073, w_053_3075, w_053_3077, w_053_3079, w_053_3080, w_053_3081, w_053_3082, w_053_3083, w_053_3084, w_053_3085, w_053_3086, w_053_3088, w_053_3089, w_053_3091, w_053_3093, w_053_3095, w_053_3097, w_053_3098, w_053_3099, w_053_3100, w_053_3101, w_053_3102, w_053_3103, w_053_3104, w_053_3105, w_053_3109, w_053_3110, w_053_3113, w_053_3114, w_053_3116, w_053_3118, w_053_3120, w_053_3124, w_053_3125, w_053_3126, w_053_3127, w_053_3128, w_053_3129, w_053_3130, w_053_3133, w_053_3134, w_053_3135, w_053_3136, w_053_3138, w_053_3139, w_053_3140, w_053_3141, w_053_3142, w_053_3143, w_053_3144, w_053_3145, w_053_3146, w_053_3147, w_053_3148, w_053_3150, w_053_3151, w_053_3153, w_053_3155, w_053_3157, w_053_3160, w_053_3161, w_053_3163, w_053_3164, w_053_3166, w_053_3167, w_053_3168, w_053_3169, w_053_3172, w_053_3173, w_053_3174, w_053_3175, w_053_3177, w_053_3180, w_053_3181, w_053_3183, w_053_3185, w_053_3186, w_053_3187, w_053_3188, w_053_3189, w_053_3190, w_053_3192, w_053_3193, w_053_3194, w_053_3195, w_053_3198, w_053_3202, w_053_3204, w_053_3207, w_053_3208, w_053_3209, w_053_3210, w_053_3214, w_053_3215, w_053_3217, w_053_3219, w_053_3220, w_053_3221, w_053_3222, w_053_3224, w_053_3226, w_053_3227, w_053_3228, w_053_3229, w_053_3230, w_053_3232, w_053_3233, w_053_3234, w_053_3235, w_053_3239, w_053_3240, w_053_3241, w_053_3242, w_053_3244, w_053_3248, w_053_3250, w_053_3251, w_053_3252, w_053_3253, w_053_3254, w_053_3255, w_053_3256, w_053_3257, w_053_3258, w_053_3260, w_053_3263, w_053_3266, w_053_3268, w_053_3269, w_053_3270, w_053_3271, w_053_3273, w_053_3275, w_053_3276, w_053_3277, w_053_3278, w_053_3280, w_053_3281, w_053_3285, w_053_3287, w_053_3289, w_053_3291, w_053_3292, w_053_3293, w_053_3294, w_053_3296, w_053_3297, w_053_3298, w_053_3299, w_053_3300, w_053_3302, w_053_3303, w_053_3304, w_053_3309, w_053_3310, w_053_3315, w_053_3316, w_053_3318, w_053_3319, w_053_3320, w_053_3322, w_053_3326, w_053_3328, w_053_3329, w_053_3334, w_053_3336, w_053_3337, w_053_3338, w_053_3339, w_053_3340, w_053_3341, w_053_3342, w_053_3343, w_053_3344, w_053_3346, w_053_3347, w_053_3348, w_053_3349, w_053_3354, w_053_3355, w_053_3357, w_053_3358, w_053_3359, w_053_3360, w_053_3361, w_053_3362, w_053_3363, w_053_3364, w_053_3365, w_053_3367, w_053_3369, w_053_3371, w_053_3372, w_053_3373, w_053_3375, w_053_3379, w_053_3380, w_053_3382, w_053_3383, w_053_3385, w_053_3388, w_053_3389, w_053_3390, w_053_3392, w_053_3393, w_053_3395, w_053_3396, w_053_3397, w_053_3398, w_053_3401, w_053_3402, w_053_3403, w_053_3404, w_053_3408, w_053_3409, w_053_3411, w_053_3413, w_053_3417, w_053_3418, w_053_3420, w_053_3422, w_053_3423, w_053_3425, w_053_3426, w_053_3427, w_053_3430, w_053_3431, w_053_3435, w_053_3437, w_053_3438, w_053_3440, w_053_3441, w_053_3442, w_053_3443, w_053_3445, w_053_3447, w_053_3448, w_053_3449, w_053_3450, w_053_3454, w_053_3456, w_053_3457, w_053_3459, w_053_3460, w_053_3461, w_053_3465, w_053_3466, w_053_3468, w_053_3470, w_053_3471, w_053_3472, w_053_3473, w_053_3474, w_053_3476, w_053_3478, w_053_3479, w_053_3481, w_053_3482, w_053_3483, w_053_3484, w_053_3486, w_053_3487, w_053_3492, w_053_3493, w_053_3494, w_053_3496, w_053_3497, w_053_3498, w_053_3499, w_053_3500, w_053_3502, w_053_3504, w_053_3505, w_053_3507, w_053_3508, w_053_3509, w_053_3510, w_053_3511, w_053_3512, w_053_3514, w_053_3516, w_053_3517, w_053_3518, w_053_3521, w_053_3522, w_053_3523, w_053_3524, w_053_3526, w_053_3527, w_053_3528, w_053_3529, w_053_3530, w_053_3531, w_053_3532, w_053_3533, w_053_3537, w_053_3538, w_053_3539, w_053_3541, w_053_3543, w_053_3544, w_053_3546, w_053_3547, w_053_3548, w_053_3549, w_053_3550, w_053_3551, w_053_3552, w_053_3553, w_053_3554, w_053_3555, w_053_3557, w_053_3559, w_053_3560, w_053_3562, w_053_3563, w_053_3564, w_053_3565, w_053_3570, w_053_3571, w_053_3572, w_053_3575, w_053_3576, w_053_3578, w_053_3579, w_053_3580, w_053_3581, w_053_3583, w_053_3584, w_053_3587, w_053_3588, w_053_3589, w_053_3590, w_053_3591, w_053_3595, w_053_3596, w_053_3597, w_053_3598, w_053_3599, w_053_3601, w_053_3602, w_053_3603, w_053_3606, w_053_3607, w_053_3610, w_053_3612, w_053_3615, w_053_3616, w_053_3619, w_053_3621, w_053_3623, w_053_3624, w_053_3626, w_053_3628, w_053_3630, w_053_3631, w_053_3632, w_053_3633, w_053_3634, w_053_3635, w_053_3636, w_053_3639, w_053_3640, w_053_3642, w_053_3645, w_053_3648, w_053_3649, w_053_3650, w_053_3651, w_053_3654, w_053_3655, w_053_3656, w_053_3659, w_053_3660, w_053_3661, w_053_3662, w_053_3663, w_053_3664, w_053_3666, w_053_3667, w_053_3668, w_053_3669, w_053_3670, w_053_3671, w_053_3672, w_053_3673, w_053_3675, w_053_3677, w_053_3678, w_053_3679, w_053_3680, w_053_3682, w_053_3683, w_053_3684, w_053_3685, w_053_3686, w_053_3687, w_053_3688, w_053_3690, w_053_3691, w_053_3692, w_053_3693, w_053_3696, w_053_3697, w_053_3698, w_053_3699, w_053_3700, w_053_3702, w_053_3703, w_053_3704, w_053_3706, w_053_3707, w_053_3708, w_053_3709, w_053_3711, w_053_3712, w_053_3715, w_053_3717, w_053_3718, w_053_3721, w_053_3722, w_053_3724, w_053_3726, w_053_3727, w_053_3729, w_053_3730, w_053_3731, w_053_3732, w_053_3734, w_053_3738, w_053_3745, w_053_3746, w_053_3748, w_053_3749, w_053_3750, w_053_3751, w_053_3752, w_053_3753, w_053_3754, w_053_3755, w_053_3756, w_053_3758, w_053_3759, w_053_3760, w_053_3761, w_053_3764, w_053_3765, w_053_3768, w_053_3769, w_053_3770, w_053_3772, w_053_3775, w_053_3776, w_053_3777, w_053_3778, w_053_3779, w_053_3780, w_053_3781, w_053_3782, w_053_3783, w_053_3784, w_053_3786, w_053_3787, w_053_3788, w_053_3790, w_053_3791, w_053_3792, w_053_3793, w_053_3794, w_053_3795, w_053_3798, w_053_3799, w_053_3800, w_053_3801, w_053_3802, w_053_3803, w_053_3804, w_053_3808, w_053_3813, w_053_3814, w_053_3816, w_053_3817, w_053_3820, w_053_3821, w_053_3822, w_053_3824, w_053_3825, w_053_3827, w_053_3828, w_053_3829, w_053_3830, w_053_3832, w_053_3833, w_053_3835, w_053_3836, w_053_3837, w_053_3838, w_053_3839, w_053_3840, w_053_3841, w_053_3842, w_053_3843, w_053_3844, w_053_3845, w_053_3848, w_053_3850, w_053_3852, w_053_3853, w_053_3854, w_053_3856, w_053_3858, w_053_3859, w_053_3861, w_053_3862, w_053_3863, w_053_3864, w_053_3865, w_053_3867, w_053_3868, w_053_3869, w_053_3871, w_053_3874, w_053_3875, w_053_3876, w_053_3877, w_053_3880, w_053_3882, w_053_3884, w_053_3885, w_053_3886, w_053_3888, w_053_3889, w_053_3893, w_053_3894, w_053_3896, w_053_3897, w_053_3901, w_053_3904, w_053_3905, w_053_3906, w_053_3908, w_053_3910, w_053_3911, w_053_3913, w_053_3914, w_053_3915, w_053_3916, w_053_3917, w_053_3918, w_053_3920, w_053_3921, w_053_3922, w_053_3923, w_053_3925, w_053_3926, w_053_3927, w_053_3928, w_053_3930, w_053_3931, w_053_3932, w_053_3933, w_053_3934, w_053_3935, w_053_3936, w_053_3939, w_053_3941, w_053_3942, w_053_3943, w_053_3944, w_053_3946, w_053_3948, w_053_3952, w_053_3953, w_053_3954, w_053_3956, w_053_3958, w_053_3960, w_053_3964, w_053_3965, w_053_3966, w_053_3968, w_053_3969, w_053_3970, w_053_3971, w_053_3972, w_053_3973, w_053_3974, w_053_3975, w_053_3977, w_053_3978, w_053_3979, w_053_3980, w_053_3981, w_053_3982, w_053_3984, w_053_3985, w_053_3986, w_053_3987, w_053_3988, w_053_3989, w_053_3990, w_053_3992, w_053_3993, w_053_3994, w_053_3995, w_053_3997, w_053_3998, w_053_4000, w_053_4001, w_053_4003, w_053_4004, w_053_4005, w_053_4006, w_053_4007, w_053_4010, w_053_4011, w_053_4012, w_053_4013, w_053_4014, w_053_4015, w_053_4016, w_053_4017, w_053_4018, w_053_4019, w_053_4021, w_053_4023, w_053_4024, w_053_4025, w_053_4026, w_053_4029, w_053_4030, w_053_4031, w_053_4033, w_053_4034, w_053_4037, w_053_4038, w_053_4039, w_053_4040, w_053_4042, w_053_4043, w_053_4045, w_053_4046, w_053_4048, w_053_4050, w_053_4051, w_053_4052, w_053_4053, w_053_4055, w_053_4057, w_053_4058, w_053_4059, w_053_4060, w_053_4062, w_053_4063, w_053_4064, w_053_4067, w_053_4069, w_053_4071, w_053_4072, w_053_4073, w_053_4074, w_053_4075, w_053_4076, w_053_4078, w_053_4079, w_053_4081, w_053_4082, w_053_4084, w_053_4086, w_053_4088, w_053_4089, w_053_4090, w_053_4091, w_053_4093, w_053_4094, w_053_4095, w_053_4096, w_053_4100, w_053_4101, w_053_4102, w_053_4103, w_053_4105, w_053_4106, w_053_4108, w_053_4110, w_053_4114, w_053_4118, w_053_4120, w_053_4123, w_053_4124, w_053_4127, w_053_4130, w_053_4131, w_053_4132, w_053_4134, w_053_4135, w_053_4136, w_053_4137, w_053_4138, w_053_4141, w_053_4144, w_053_4145, w_053_4147, w_053_4148, w_053_4150, w_053_4151, w_053_4153, w_053_4155, w_053_4157, w_053_4158, w_053_4159, w_053_4160, w_053_4161, w_053_4162, w_053_4163, w_053_4164, w_053_4166, w_053_4167, w_053_4169, w_053_4171, w_053_4174, w_053_4175, w_053_4176, w_053_4177, w_053_4178, w_053_4180, w_053_4182, w_053_4183, w_053_4184, w_053_4185, w_053_4186, w_053_4187, w_053_4188, w_053_4191, w_053_4192, w_053_4193, w_053_4194, w_053_4195, w_053_4196, w_053_4198, w_053_4199, w_053_4201, w_053_4202, w_053_4205, w_053_4206, w_053_4207, w_053_4208, w_053_4209, w_053_4212, w_053_4213, w_053_4214, w_053_4216, w_053_4217, w_053_4218, w_053_4221, w_053_4222, w_053_4223, w_053_4224, w_053_4225, w_053_4226, w_053_4227, w_053_4229, w_053_4230, w_053_4234, w_053_4235, w_053_4236, w_053_4237, w_053_4238, w_053_4239, w_053_4240, w_053_4241, w_053_4242, w_053_4243, w_053_4244, w_053_4245, w_053_4246, w_053_4248, w_053_4249, w_053_4250, w_053_4251, w_053_4252, w_053_4255, w_053_4256, w_053_4258, w_053_4261, w_053_4262, w_053_4263, w_053_4266, w_053_4267, w_053_4268, w_053_4270, w_053_4272, w_053_4274, w_053_4275, w_053_4276, w_053_4277, w_053_4278, w_053_4279, w_053_4280, w_053_4281, w_053_4283, w_053_4284, w_053_4287, w_053_4288, w_053_4289, w_053_4290, w_053_4291, w_053_4292, w_053_4293, w_053_4296, w_053_4297, w_053_4298, w_053_4299, w_053_4301, w_053_4302, w_053_4303, w_053_4305, w_053_4306, w_053_4307, w_053_4309, w_053_4310, w_053_4312, w_053_4313, w_053_4315, w_053_4316, w_053_4318, w_053_4319, w_053_4322, w_053_4323, w_053_4324, w_053_4326, w_053_4327, w_053_4330, w_053_4331, w_053_4334, w_053_4335, w_053_4336, w_053_4339, w_053_4340, w_053_4341, w_053_4342, w_053_4344, w_053_4345, w_053_4346, w_053_4348, w_053_4351, w_053_4353, w_053_4355, w_053_4356, w_053_4358, w_053_4359, w_053_4361, w_053_4362, w_053_4364, w_053_4365, w_053_4366, w_053_4367, w_053_4369, w_053_4370, w_053_4371, w_053_4372, w_053_4373, w_053_4374, w_053_4376, w_053_4378, w_053_4381, w_053_4382, w_053_4383, w_053_4384, w_053_4385, w_053_4387, w_053_4388, w_053_4389, w_053_4390, w_053_4392, w_053_4395, w_053_4396, w_053_4397, w_053_4398, w_053_4400, w_053_4401, w_053_4402, w_053_4404, w_053_4406, w_053_4409, w_053_4411, w_053_4412, w_053_4413, w_053_4414, w_053_4415, w_053_4419, w_053_4420, w_053_4422, w_053_4423, w_053_4424, w_053_4425, w_053_4426, w_053_4428, w_053_4429, w_053_4431, w_053_4433, w_053_4434, w_053_4435, w_053_4436, w_053_4437, w_053_4438, w_053_4439, w_053_4440, w_053_4441, w_053_4442, w_053_4443, w_053_4445, w_053_4447, w_053_4450, w_053_4451, w_053_4452, w_053_4453, w_053_4458, w_053_4460, w_053_4461, w_053_4462, w_053_4463, w_053_4464, w_053_4465, w_053_4466, w_053_4468, w_053_4469, w_053_4470, w_053_4471, w_053_4472, w_053_4474, w_053_4476, w_053_4477, w_053_4478, w_053_4480, w_053_4481, w_053_4482, w_053_4494, w_053_4495, w_053_4503, w_053_4505, w_053_4506, w_053_4509, w_053_4517, w_053_4518, w_053_4519, w_053_4520, w_053_4521, w_053_4522, w_053_4523, w_053_4524, w_053_4528, w_053_4532, w_053_4535, w_053_4536, w_053_4537, w_053_4542, w_053_4544, w_053_4550, w_053_4557, w_053_4558, w_053_4560, w_053_4561, w_053_4563, w_053_4566, w_053_4567, w_053_4571, w_053_4573, w_053_4579, w_053_4582, w_053_4588, w_053_4589, w_053_4591, w_053_4593, w_053_4594, w_053_4597, w_053_4598, w_053_4605, w_053_4609, w_053_4610, w_053_4614, w_053_4616, w_053_4617, w_053_4622, w_053_4624, w_053_4626, w_053_4629, w_053_4632, w_053_4633, w_053_4634, w_053_4636, w_053_4637, w_053_4638, w_053_4639, w_053_4641, w_053_4643, w_053_4651, w_053_4662, w_053_4664, w_053_4665, w_053_4670, w_053_4676, w_053_4677, w_053_4678, w_053_4679, w_053_4684, w_053_4685, w_053_4686, w_053_4689, w_053_4691, w_053_4695, w_053_4696, w_053_4698, w_053_4700, w_053_4702, w_053_4705, w_053_4707, w_053_4716, w_053_4719, w_053_4720, w_053_4721, w_053_4723, w_053_4724, w_053_4732, w_053_4733, w_053_4734, w_053_4736, w_053_4737, w_053_4739, w_053_4741, w_053_4742, w_053_4754, w_053_4755, w_053_4758, w_053_4759, w_053_4762, w_053_4763, w_053_4766, w_053_4772, w_053_4779, w_053_4781, w_053_4794, w_053_4796, w_053_4797, w_053_4801, w_053_4803, w_053_4808, w_053_4811, w_053_4813, w_053_4814, w_053_4815, w_053_4817, w_053_4818, w_053_4822, w_053_4824, w_053_4829, w_053_4830, w_053_4831, w_053_4832, w_053_4834, w_053_4837, w_053_4839, w_053_4844, w_053_4845, w_053_4846, w_053_4847, w_053_4849, w_053_4854, w_053_4856, w_053_4858, w_053_4862, w_053_4863, w_053_4866, w_053_4867, w_053_4868, w_053_4870, w_053_4871, w_053_4875, w_053_4877, w_053_4878, w_053_4880, w_053_4882, w_053_4883, w_053_4887, w_053_4888, w_053_4894, w_053_4896, w_053_4897, w_053_4899, w_053_4900, w_053_4902, w_053_4906, w_053_4907, w_053_4910, w_053_4912, w_053_4914, w_053_4918, w_053_4921, w_053_4928, w_053_4930, w_053_4933, w_053_4934, w_053_4935, w_053_4936, w_053_4937, w_053_4939, w_053_4940, w_053_4942, w_053_4943, w_053_4944, w_053_4945, w_053_4946, w_053_4948, w_053_4952, w_053_4953, w_053_4960, w_053_4968, w_053_4970, w_053_4972, w_053_4973, w_053_4974, w_053_4976, w_053_4979, w_053_4980, w_053_4982, w_053_4983, w_053_4984, w_053_4985, w_053_4988, w_053_4990, w_053_4991, w_053_4992, w_053_4999, w_053_5000, w_053_5004, w_053_5005, w_053_5008, w_053_5009, w_053_5010, w_053_5011, w_053_5012, w_053_5015, w_053_5016, w_053_5017, w_053_5019, w_053_5023, w_053_5024, w_053_5025, w_053_5026, w_053_5029, w_053_5032, w_053_5034, w_053_5035, w_053_5036, w_053_5040, w_053_5042, w_053_5051, w_053_5052, w_053_5054, w_053_5055, w_053_5057, w_053_5060, w_053_5067, w_053_5069, w_053_5071, w_053_5072, w_053_5074, w_053_5076, w_053_5082, w_053_5084, w_053_5085, w_053_5087, w_053_5091, w_053_5094, w_053_5095, w_053_5096, w_053_5097, w_053_5098, w_053_5099, w_053_5103, w_053_5109, w_053_5110, w_053_5111, w_053_5116, w_053_5124, w_053_5127, w_053_5129, w_053_5130, w_053_5131, w_053_5140, w_053_5145, w_053_5146, w_053_5148, w_053_5155, w_053_5162, w_053_5165, w_053_5168, w_053_5171, w_053_5173, w_053_5176, w_053_5179, w_053_5180, w_053_5181, w_053_5183, w_053_5185, w_053_5188, w_053_5189, w_053_5191, w_053_5192, w_053_5199, w_053_5201, w_053_5204, w_053_5206, w_053_5207, w_053_5209, w_053_5210, w_053_5212, w_053_5216, w_053_5219, w_053_5223, w_053_5228, w_053_5229, w_053_5230, w_053_5231, w_053_5232, w_053_5236, w_053_5237, w_053_5239, w_053_5240, w_053_5243, w_053_5249, w_053_5250, w_053_5251, w_053_5261, w_053_5262, w_053_5264, w_053_5265, w_053_5271, w_053_5274, w_053_5275, w_053_5277, w_053_5278, w_053_5287, w_053_5288, w_053_5291, w_053_5294, w_053_5305, w_053_5314, w_053_5316, w_053_5328, w_053_5334, w_053_5337, w_053_5338, w_053_5342, w_053_5343, w_053_5348, w_053_5349, w_053_5350, w_053_5351, w_053_5355, w_053_5358, w_053_5360, w_053_5362, w_053_5363, w_053_5367, w_053_5368, w_053_5375, w_053_5376, w_053_5378, w_053_5379, w_053_5380, w_053_5382, w_053_5385, w_053_5386, w_053_5388, w_053_5393, w_053_5395, w_053_5396, w_053_5399, w_053_5400, w_053_5401, w_053_5402, w_053_5406, w_053_5408, w_053_5409, w_053_5417, w_053_5421, w_053_5425, w_053_5426, w_053_5432, w_053_5434, w_053_5435, w_053_5436, w_053_5440, w_053_5443, w_053_5447, w_053_5451, w_053_5452, w_053_5453, w_053_5454, w_053_5457, w_053_5458, w_053_5459, w_053_5470, w_053_5474, w_053_5479, w_053_5480, w_053_5482, w_053_5483, w_053_5484, w_053_5485, w_053_5489, w_053_5492, w_053_5495, w_053_5506, w_053_5511, w_053_5512;
  wire w_054_000, w_054_002, w_054_003, w_054_004, w_054_007, w_054_008, w_054_009, w_054_010, w_054_013, w_054_014, w_054_015, w_054_017, w_054_019, w_054_020, w_054_021, w_054_022, w_054_023, w_054_027, w_054_028, w_054_029, w_054_030, w_054_031, w_054_032, w_054_035, w_054_037, w_054_038, w_054_040, w_054_046, w_054_047, w_054_049, w_054_050, w_054_051, w_054_052, w_054_053, w_054_055, w_054_056, w_054_057, w_054_059, w_054_061, w_054_063, w_054_064, w_054_066, w_054_070, w_054_071, w_054_072, w_054_073, w_054_074, w_054_075, w_054_076, w_054_078, w_054_080, w_054_081, w_054_084, w_054_085, w_054_087, w_054_088, w_054_089, w_054_092, w_054_093, w_054_096, w_054_097, w_054_098, w_054_099, w_054_100, w_054_102, w_054_105, w_054_106, w_054_107, w_054_108, w_054_109, w_054_111, w_054_117, w_054_121, w_054_122, w_054_123, w_054_126, w_054_129, w_054_131, w_054_132, w_054_137, w_054_139, w_054_143, w_054_144, w_054_146, w_054_147, w_054_148, w_054_150, w_054_151, w_054_152, w_054_155, w_054_156, w_054_157, w_054_159, w_054_160, w_054_164, w_054_165, w_054_169, w_054_170, w_054_171, w_054_172, w_054_175, w_054_176, w_054_178, w_054_179, w_054_180, w_054_183, w_054_185, w_054_187, w_054_189, w_054_191, w_054_192, w_054_193, w_054_194, w_054_195, w_054_196, w_054_198, w_054_200, w_054_202, w_054_204, w_054_206, w_054_210, w_054_211, w_054_212, w_054_213, w_054_215, w_054_216, w_054_217, w_054_220, w_054_221, w_054_223, w_054_224, w_054_225, w_054_226, w_054_227, w_054_230, w_054_232, w_054_233, w_054_235, w_054_237, w_054_238, w_054_239, w_054_242, w_054_243, w_054_244, w_054_245, w_054_246, w_054_247, w_054_251, w_054_252, w_054_253, w_054_255, w_054_258, w_054_260, w_054_262, w_054_264, w_054_268, w_054_269, w_054_275, w_054_277, w_054_278, w_054_280, w_054_282, w_054_284, w_054_286, w_054_289, w_054_290, w_054_296, w_054_297, w_054_298, w_054_299, w_054_300, w_054_301, w_054_302, w_054_303, w_054_304, w_054_307, w_054_308, w_054_310, w_054_311, w_054_312, w_054_313, w_054_315, w_054_322, w_054_324, w_054_325, w_054_326, w_054_327, w_054_330, w_054_332, w_054_333, w_054_337, w_054_338, w_054_339, w_054_341, w_054_342, w_054_343, w_054_344, w_054_345, w_054_346, w_054_349, w_054_350, w_054_351, w_054_352, w_054_353, w_054_354, w_054_355, w_054_356, w_054_359, w_054_362, w_054_363, w_054_366, w_054_367, w_054_369, w_054_370, w_054_371, w_054_373, w_054_375, w_054_377, w_054_379, w_054_381, w_054_384, w_054_385, w_054_390, w_054_391, w_054_393, w_054_394, w_054_395, w_054_398, w_054_400, w_054_402, w_054_403, w_054_405, w_054_408, w_054_410, w_054_412, w_054_414, w_054_416, w_054_417, w_054_418, w_054_419, w_054_421, w_054_422, w_054_424, w_054_428, w_054_432, w_054_433, w_054_434, w_054_436, w_054_437, w_054_439, w_054_442, w_054_443, w_054_444, w_054_446, w_054_447, w_054_449, w_054_453, w_054_455, w_054_456, w_054_457, w_054_460, w_054_461, w_054_462, w_054_463, w_054_464, w_054_465, w_054_467, w_054_468, w_054_470, w_054_471, w_054_472, w_054_473, w_054_475, w_054_476, w_054_477, w_054_478, w_054_480, w_054_482, w_054_483, w_054_484, w_054_485, w_054_489, w_054_490, w_054_492, w_054_493, w_054_494, w_054_498, w_054_499, w_054_500, w_054_502, w_054_505, w_054_506, w_054_507, w_054_510, w_054_511, w_054_512, w_054_514, w_054_519, w_054_520, w_054_522, w_054_525, w_054_527, w_054_528, w_054_530, w_054_531, w_054_532, w_054_534, w_054_535, w_054_537, w_054_539, w_054_541, w_054_543, w_054_545, w_054_546, w_054_547, w_054_549, w_054_552, w_054_553, w_054_555, w_054_556, w_054_560, w_054_561, w_054_563, w_054_564, w_054_565, w_054_566, w_054_568, w_054_569, w_054_570, w_054_571, w_054_572, w_054_573, w_054_576, w_054_577, w_054_578, w_054_579, w_054_580, w_054_581, w_054_582, w_054_584, w_054_587, w_054_588, w_054_589, w_054_591, w_054_592, w_054_593, w_054_595, w_054_596, w_054_597, w_054_598, w_054_599, w_054_601, w_054_602, w_054_604, w_054_605, w_054_609, w_054_611, w_054_612, w_054_615, w_054_616, w_054_617, w_054_618, w_054_620, w_054_622, w_054_624, w_054_628, w_054_629, w_054_630, w_054_631, w_054_632, w_054_633, w_054_634, w_054_636, w_054_637, w_054_640, w_054_641, w_054_642, w_054_643, w_054_644, w_054_646, w_054_647, w_054_648, w_054_650, w_054_653, w_054_654, w_054_655, w_054_656, w_054_657, w_054_658, w_054_659, w_054_660, w_054_664, w_054_665, w_054_666, w_054_667, w_054_672, w_054_673, w_054_674, w_054_675, w_054_676, w_054_678, w_054_679, w_054_681, w_054_682, w_054_683, w_054_684, w_054_686, w_054_687, w_054_688, w_054_689, w_054_690, w_054_691, w_054_694, w_054_695, w_054_699, w_054_700, w_054_701, w_054_706, w_054_709, w_054_710, w_054_711, w_054_715, w_054_716, w_054_717, w_054_718, w_054_719, w_054_720, w_054_721, w_054_726, w_054_727, w_054_728, w_054_729, w_054_730, w_054_732, w_054_733, w_054_736, w_054_737, w_054_739, w_054_744, w_054_745, w_054_746, w_054_747, w_054_749, w_054_751, w_054_752, w_054_754, w_054_755, w_054_757, w_054_758, w_054_759, w_054_760, w_054_761, w_054_764, w_054_767, w_054_769, w_054_771, w_054_772, w_054_775, w_054_776, w_054_779, w_054_780, w_054_782, w_054_783, w_054_785, w_054_786, w_054_787, w_054_788, w_054_789, w_054_793, w_054_797, w_054_799, w_054_800, w_054_801, w_054_802, w_054_803, w_054_804, w_054_806, w_054_807, w_054_810, w_054_813, w_054_814, w_054_815, w_054_816, w_054_819, w_054_820, w_054_821, w_054_823, w_054_824, w_054_825, w_054_826, w_054_827, w_054_828, w_054_829, w_054_831, w_054_834, w_054_835, w_054_838, w_054_839, w_054_840, w_054_842, w_054_843, w_054_844, w_054_846, w_054_847, w_054_848, w_054_849, w_054_850, w_054_851, w_054_853, w_054_854, w_054_856, w_054_857, w_054_859, w_054_860, w_054_861, w_054_862, w_054_866, w_054_869, w_054_870, w_054_872, w_054_873, w_054_875, w_054_876, w_054_877, w_054_878, w_054_879, w_054_881, w_054_883, w_054_884, w_054_885, w_054_886, w_054_887, w_054_890, w_054_891, w_054_892, w_054_893, w_054_894, w_054_896, w_054_898, w_054_903, w_054_904, w_054_906, w_054_909, w_054_910, w_054_911, w_054_913, w_054_914, w_054_916, w_054_920, w_054_921, w_054_923, w_054_924, w_054_926, w_054_927, w_054_929, w_054_932, w_054_933, w_054_934, w_054_935, w_054_936, w_054_940, w_054_941, w_054_943, w_054_944, w_054_945, w_054_946, w_054_950, w_054_951, w_054_952, w_054_953, w_054_954, w_054_955, w_054_958, w_054_961, w_054_964, w_054_966, w_054_967, w_054_968, w_054_969, w_054_970, w_054_972, w_054_974, w_054_975, w_054_976, w_054_977, w_054_978, w_054_979, w_054_981, w_054_983, w_054_984, w_054_985, w_054_986, w_054_987, w_054_988, w_054_990, w_054_993, w_054_994, w_054_997, w_054_998, w_054_1000, w_054_1001, w_054_1002, w_054_1003, w_054_1004, w_054_1006, w_054_1008, w_054_1009, w_054_1010, w_054_1012, w_054_1014, w_054_1015, w_054_1017, w_054_1019, w_054_1022, w_054_1023, w_054_1024, w_054_1025, w_054_1027, w_054_1028, w_054_1029, w_054_1031, w_054_1032, w_054_1033, w_054_1038, w_054_1039, w_054_1042, w_054_1043, w_054_1044, w_054_1045, w_054_1046, w_054_1047, w_054_1048, w_054_1049, w_054_1050, w_054_1052, w_054_1053, w_054_1054, w_054_1055, w_054_1056, w_054_1057, w_054_1058, w_054_1059, w_054_1060, w_054_1061, w_054_1063, w_054_1064, w_054_1065, w_054_1066, w_054_1067, w_054_1068, w_054_1069, w_054_1070, w_054_1072, w_054_1074, w_054_1075, w_054_1076, w_054_1077, w_054_1078, w_054_1081, w_054_1082, w_054_1085, w_054_1086, w_054_1087, w_054_1088, w_054_1089, w_054_1090, w_054_1092, w_054_1094, w_054_1095, w_054_1096, w_054_1099, w_054_1102, w_054_1104, w_054_1105, w_054_1109, w_054_1110, w_054_1114, w_054_1115, w_054_1120, w_054_1121, w_054_1122, w_054_1123, w_054_1126, w_054_1127, w_054_1129, w_054_1130, w_054_1131, w_054_1132, w_054_1134, w_054_1136, w_054_1140, w_054_1141, w_054_1142, w_054_1145, w_054_1147, w_054_1149, w_054_1151, w_054_1152, w_054_1154, w_054_1155, w_054_1156, w_054_1157, w_054_1158, w_054_1159, w_054_1161, w_054_1162, w_054_1163, w_054_1164, w_054_1167, w_054_1168, w_054_1170, w_054_1171, w_054_1172, w_054_1173, w_054_1175, w_054_1176, w_054_1177, w_054_1179, w_054_1180, w_054_1182, w_054_1183, w_054_1186, w_054_1188, w_054_1189, w_054_1190, w_054_1191, w_054_1192, w_054_1193, w_054_1195, w_054_1196, w_054_1197, w_054_1198, w_054_1204, w_054_1205, w_054_1206, w_054_1207, w_054_1208, w_054_1211, w_054_1212, w_054_1216, w_054_1217, w_054_1220, w_054_1221, w_054_1226, w_054_1230, w_054_1232, w_054_1236, w_054_1238, w_054_1240, w_054_1243, w_054_1244, w_054_1245, w_054_1246, w_054_1248, w_054_1249, w_054_1251, w_054_1252, w_054_1253, w_054_1254, w_054_1255, w_054_1259, w_054_1262, w_054_1263, w_054_1266, w_054_1269, w_054_1270, w_054_1272, w_054_1274, w_054_1275, w_054_1276, w_054_1277, w_054_1279, w_054_1280, w_054_1281, w_054_1283, w_054_1287, w_054_1289, w_054_1292, w_054_1294, w_054_1296, w_054_1297, w_054_1298, w_054_1299, w_054_1300, w_054_1301, w_054_1302, w_054_1304, w_054_1307, w_054_1309, w_054_1310, w_054_1312, w_054_1314, w_054_1317, w_054_1318, w_054_1319, w_054_1321, w_054_1324, w_054_1326, w_054_1328, w_054_1329, w_054_1330, w_054_1331, w_054_1332, w_054_1333, w_054_1335, w_054_1338, w_054_1339, w_054_1340, w_054_1341, w_054_1343, w_054_1344, w_054_1345, w_054_1346, w_054_1347, w_054_1350, w_054_1352, w_054_1354, w_054_1355, w_054_1356, w_054_1357, w_054_1358, w_054_1359, w_054_1361, w_054_1363, w_054_1364, w_054_1366, w_054_1368, w_054_1370, w_054_1371, w_054_1372, w_054_1373, w_054_1375, w_054_1377, w_054_1379, w_054_1380, w_054_1381, w_054_1383, w_054_1384, w_054_1387, w_054_1388, w_054_1389, w_054_1393, w_054_1394, w_054_1395, w_054_1396, w_054_1399, w_054_1400, w_054_1401, w_054_1403, w_054_1405, w_054_1406, w_054_1409, w_054_1410, w_054_1412, w_054_1413, w_054_1414, w_054_1415, w_054_1417, w_054_1418, w_054_1420, w_054_1422, w_054_1423, w_054_1424, w_054_1425, w_054_1426, w_054_1427, w_054_1428, w_054_1429, w_054_1430, w_054_1431, w_054_1433, w_054_1434, w_054_1436, w_054_1437, w_054_1438, w_054_1439, w_054_1440, w_054_1441, w_054_1443, w_054_1444, w_054_1446, w_054_1448, w_054_1450, w_054_1451, w_054_1452, w_054_1456, w_054_1458, w_054_1463, w_054_1468, w_054_1470, w_054_1471, w_054_1473, w_054_1474, w_054_1475, w_054_1476, w_054_1478, w_054_1480, w_054_1482, w_054_1483, w_054_1484, w_054_1485, w_054_1487, w_054_1489, w_054_1490, w_054_1493, w_054_1494, w_054_1496, w_054_1498, w_054_1501, w_054_1502, w_054_1504, w_054_1505, w_054_1506, w_054_1507, w_054_1513, w_054_1516, w_054_1518, w_054_1521, w_054_1522, w_054_1523, w_054_1528, w_054_1529, w_054_1531, w_054_1533, w_054_1537, w_054_1539, w_054_1542, w_054_1544, w_054_1545, w_054_1547, w_054_1549, w_054_1551, w_054_1552, w_054_1553, w_054_1554, w_054_1555, w_054_1556, w_054_1557, w_054_1558, w_054_1559, w_054_1561, w_054_1562, w_054_1563, w_054_1564, w_054_1565, w_054_1567, w_054_1569, w_054_1570, w_054_1571, w_054_1572, w_054_1574, w_054_1576, w_054_1579, w_054_1580, w_054_1581, w_054_1582, w_054_1583, w_054_1584, w_054_1586, w_054_1587, w_054_1588, w_054_1589, w_054_1590, w_054_1591, w_054_1592, w_054_1593, w_054_1596, w_054_1597, w_054_1599, w_054_1600, w_054_1603, w_054_1604, w_054_1605, w_054_1606, w_054_1607, w_054_1614, w_054_1615, w_054_1616, w_054_1617, w_054_1618, w_054_1619, w_054_1620, w_054_1621, w_054_1622, w_054_1624, w_054_1626, w_054_1627, w_054_1628, w_054_1629, w_054_1630, w_054_1633, w_054_1637, w_054_1639, w_054_1640, w_054_1641, w_054_1642, w_054_1643, w_054_1644, w_054_1645, w_054_1647, w_054_1650, w_054_1651, w_054_1652, w_054_1653, w_054_1654, w_054_1655, w_054_1656, w_054_1657, w_054_1658, w_054_1659, w_054_1661, w_054_1662, w_054_1663, w_054_1664, w_054_1666, w_054_1668, w_054_1672, w_054_1673, w_054_1674, w_054_1677, w_054_1678, w_054_1684, w_054_1686, w_054_1691, w_054_1692, w_054_1696, w_054_1698, w_054_1700, w_054_1701, w_054_1702, w_054_1703, w_054_1705, w_054_1706, w_054_1707, w_054_1711, w_054_1712, w_054_1714, w_054_1717, w_054_1718, w_054_1720, w_054_1721, w_054_1722, w_054_1723, w_054_1725, w_054_1727, w_054_1728, w_054_1729, w_054_1731, w_054_1734, w_054_1735, w_054_1739, w_054_1740, w_054_1741, w_054_1743, w_054_1745, w_054_1746, w_054_1750, w_054_1751, w_054_1752, w_054_1753, w_054_1754, w_054_1757, w_054_1758, w_054_1760, w_054_1762, w_054_1764, w_054_1765, w_054_1767, w_054_1771, w_054_1774, w_054_1775, w_054_1776, w_054_1777, w_054_1778, w_054_1779, w_054_1780, w_054_1781, w_054_1788, w_054_1790, w_054_1792, w_054_1793, w_054_1795, w_054_1797, w_054_1798, w_054_1799, w_054_1801, w_054_1803, w_054_1804, w_054_1805, w_054_1806, w_054_1807, w_054_1808, w_054_1809, w_054_1810, w_054_1813, w_054_1814, w_054_1815, w_054_1816, w_054_1817, w_054_1819, w_054_1820, w_054_1821, w_054_1822, w_054_1823, w_054_1824, w_054_1825, w_054_1827, w_054_1828, w_054_1829, w_054_1830, w_054_1831, w_054_1832, w_054_1833, w_054_1838, w_054_1839, w_054_1840, w_054_1841, w_054_1842, w_054_1844, w_054_1845, w_054_1846, w_054_1847, w_054_1849, w_054_1852, w_054_1854, w_054_1855, w_054_1859, w_054_1860, w_054_1861, w_054_1863, w_054_1864, w_054_1865, w_054_1866, w_054_1868, w_054_1869, w_054_1870, w_054_1871, w_054_1872, w_054_1873, w_054_1880, w_054_1881, w_054_1883, w_054_1885, w_054_1886, w_054_1888, w_054_1889, w_054_1891, w_054_1893, w_054_1900, w_054_1901, w_054_1905, w_054_1907, w_054_1909, w_054_1912, w_054_1916, w_054_1918, w_054_1919, w_054_1920, w_054_1922, w_054_1923, w_054_1925, w_054_1926, w_054_1927, w_054_1928, w_054_1930, w_054_1931, w_054_1932, w_054_1934, w_054_1935, w_054_1937, w_054_1938, w_054_1939, w_054_1940, w_054_1941, w_054_1942, w_054_1944, w_054_1946, w_054_1947, w_054_1949, w_054_1950, w_054_1951, w_054_1952, w_054_1954, w_054_1955, w_054_1959, w_054_1962, w_054_1963, w_054_1966, w_054_1969, w_054_1970, w_054_1971, w_054_1974, w_054_1975, w_054_1976, w_054_1979, w_054_1982, w_054_1984, w_054_1985, w_054_1986, w_054_1987, w_054_1988, w_054_1989, w_054_1990, w_054_1992, w_054_1994, w_054_1996, w_054_1997, w_054_2000, w_054_2002, w_054_2003, w_054_2004, w_054_2006, w_054_2010, w_054_2011, w_054_2012, w_054_2013, w_054_2014, w_054_2015, w_054_2017, w_054_2019, w_054_2020, w_054_2021, w_054_2023, w_054_2024, w_054_2025, w_054_2026, w_054_2028, w_054_2030, w_054_2032, w_054_2034, w_054_2036, w_054_2038, w_054_2039, w_054_2040, w_054_2041, w_054_2043, w_054_2046, w_054_2047, w_054_2048, w_054_2050, w_054_2051, w_054_2053, w_054_2054, w_054_2056, w_054_2057, w_054_2058, w_054_2060, w_054_2061, w_054_2065, w_054_2067, w_054_2068, w_054_2069, w_054_2072, w_054_2073, w_054_2074, w_054_2075, w_054_2076, w_054_2080, w_054_2081, w_054_2083, w_054_2084, w_054_2088, w_054_2090, w_054_2092, w_054_2093, w_054_2095, w_054_2096, w_054_2097, w_054_2098, w_054_2101, w_054_2102, w_054_2104, w_054_2106, w_054_2107, w_054_2108, w_054_2109, w_054_2110, w_054_2111, w_054_2112, w_054_2114, w_054_2115, w_054_2116, w_054_2117, w_054_2118, w_054_2119, w_054_2122, w_054_2123, w_054_2124, w_054_2126, w_054_2127, w_054_2128, w_054_2129, w_054_2130, w_054_2133, w_054_2134, w_054_2135, w_054_2136, w_054_2140, w_054_2141, w_054_2143, w_054_2144, w_054_2146, w_054_2147, w_054_2148, w_054_2149, w_054_2150, w_054_2154, w_054_2155, w_054_2156, w_054_2158, w_054_2159, w_054_2160, w_054_2161, w_054_2162, w_054_2163, w_054_2164, w_054_2165, w_054_2166, w_054_2167, w_054_2168, w_054_2170, w_054_2171, w_054_2174, w_054_2175, w_054_2177, w_054_2179, w_054_2181, w_054_2186, w_054_2192, w_054_2193, w_054_2194, w_054_2195, w_054_2200, w_054_2202, w_054_2203, w_054_2205, w_054_2206, w_054_2209, w_054_2210, w_054_2213, w_054_2215, w_054_2216, w_054_2220, w_054_2222, w_054_2223, w_054_2224, w_054_2227, w_054_2228, w_054_2231, w_054_2234, w_054_2235, w_054_2237, w_054_2240, w_054_2241, w_054_2242, w_054_2244, w_054_2245, w_054_2246, w_054_2247, w_054_2249, w_054_2251, w_054_2252, w_054_2253, w_054_2255, w_054_2258, w_054_2259, w_054_2260, w_054_2261, w_054_2263, w_054_2264, w_054_2266, w_054_2267, w_054_2268, w_054_2272, w_054_2276, w_054_2277, w_054_2278, w_054_2279, w_054_2280, w_054_2281, w_054_2282, w_054_2283, w_054_2284, w_054_2285, w_054_2286, w_054_2290, w_054_2292, w_054_2294, w_054_2295, w_054_2296, w_054_2297, w_054_2298, w_054_2304, w_054_2305, w_054_2307, w_054_2309, w_054_2311, w_054_2313, w_054_2314, w_054_2317, w_054_2321, w_054_2322, w_054_2323, w_054_2324, w_054_2325, w_054_2327, w_054_2330, w_054_2331, w_054_2332, w_054_2333, w_054_2334, w_054_2335, w_054_2336, w_054_2338, w_054_2339, w_054_2340, w_054_2341, w_054_2342, w_054_2343, w_054_2344, w_054_2345, w_054_2346, w_054_2348, w_054_2355, w_054_2357, w_054_2360, w_054_2361, w_054_2362, w_054_2365, w_054_2366, w_054_2367, w_054_2368, w_054_2371, w_054_2372, w_054_2374, w_054_2375, w_054_2376, w_054_2378, w_054_2379, w_054_2381, w_054_2383, w_054_2386, w_054_2387, w_054_2389, w_054_2390, w_054_2391, w_054_2393, w_054_2394, w_054_2395, w_054_2398, w_054_2399, w_054_2400, w_054_2402, w_054_2403, w_054_2404, w_054_2405, w_054_2408, w_054_2410, w_054_2411, w_054_2413, w_054_2416, w_054_2418, w_054_2419, w_054_2422, w_054_2423, w_054_2424, w_054_2425, w_054_2427, w_054_2428, w_054_2431, w_054_2432, w_054_2433, w_054_2434, w_054_2436, w_054_2440, w_054_2441, w_054_2443, w_054_2444, w_054_2446, w_054_2448, w_054_2449, w_054_2450, w_054_2452, w_054_2454, w_054_2455, w_054_2457, w_054_2458, w_054_2460, w_054_2461, w_054_2463, w_054_2466, w_054_2467, w_054_2468, w_054_2469, w_054_2470, w_054_2472, w_054_2473, w_054_2474, w_054_2477, w_054_2478, w_054_2479, w_054_2480, w_054_2481, w_054_2482, w_054_2484, w_054_2487, w_054_2488, w_054_2490, w_054_2491, w_054_2492, w_054_2493, w_054_2494, w_054_2495, w_054_2497, w_054_2499, w_054_2503, w_054_2505, w_054_2506, w_054_2507, w_054_2512, w_054_2513, w_054_2519, w_054_2520, w_054_2521, w_054_2523, w_054_2524, w_054_2525, w_054_2526, w_054_2527, w_054_2528, w_054_2529, w_054_2531, w_054_2532, w_054_2533, w_054_2534, w_054_2535, w_054_2536, w_054_2538, w_054_2540, w_054_2541, w_054_2543, w_054_2544, w_054_2545, w_054_2546, w_054_2548, w_054_2549, w_054_2551, w_054_2552, w_054_2554, w_054_2556, w_054_2557, w_054_2559, w_054_2562, w_054_2563, w_054_2564, w_054_2566, w_054_2569, w_054_2570, w_054_2573, w_054_2579, w_054_2580, w_054_2583, w_054_2585, w_054_2586, w_054_2590, w_054_2591, w_054_2592, w_054_2593, w_054_2594, w_054_2595, w_054_2596, w_054_2598, w_054_2600, w_054_2601, w_054_2602, w_054_2604, w_054_2605, w_054_2606, w_054_2608, w_054_2609, w_054_2610, w_054_2612, w_054_2614, w_054_2615, w_054_2616, w_054_2619, w_054_2621, w_054_2623, w_054_2626, w_054_2628, w_054_2630, w_054_2631, w_054_2632, w_054_2634, w_054_2636, w_054_2637, w_054_2639, w_054_2640, w_054_2641, w_054_2643, w_054_2644, w_054_2645, w_054_2647, w_054_2648, w_054_2649, w_054_2650, w_054_2651, w_054_2652, w_054_2653, w_054_2654, w_054_2655, w_054_2658, w_054_2660, w_054_2662, w_054_2663, w_054_2664, w_054_2665, w_054_2668, w_054_2672, w_054_2674, w_054_2675, w_054_2677, w_054_2678, w_054_2681, w_054_2683, w_054_2686, w_054_2687, w_054_2688, w_054_2689, w_054_2691, w_054_2692, w_054_2695, w_054_2696, w_054_2700, w_054_2701, w_054_2702, w_054_2704, w_054_2707, w_054_2708, w_054_2710, w_054_2711, w_054_2712, w_054_2713, w_054_2716, w_054_2717, w_054_2718, w_054_2719, w_054_2720, w_054_2721, w_054_2722, w_054_2724, w_054_2725, w_054_2726, w_054_2728, w_054_2729, w_054_2730, w_054_2734, w_054_2736, w_054_2741, w_054_2742, w_054_2743, w_054_2745, w_054_2746, w_054_2749, w_054_2750, w_054_2751, w_054_2753, w_054_2756, w_054_2760, w_054_2761, w_054_2762, w_054_2764, w_054_2765, w_054_2766, w_054_2767, w_054_2768, w_054_2770, w_054_2771, w_054_2773, w_054_2775, w_054_2777, w_054_2778, w_054_2779, w_054_2781, w_054_2784, w_054_2786, w_054_2788, w_054_2789, w_054_2791, w_054_2792, w_054_2793, w_054_2794, w_054_2795, w_054_2797, w_054_2798, w_054_2799, w_054_2800, w_054_2801, w_054_2802, w_054_2803, w_054_2804, w_054_2805, w_054_2806, w_054_2808, w_054_2809, w_054_2810, w_054_2811, w_054_2812, w_054_2813, w_054_2815, w_054_2816, w_054_2817, w_054_2818, w_054_2820, w_054_2821, w_054_2822, w_054_2825, w_054_2826, w_054_2827, w_054_2828, w_054_2830, w_054_2831, w_054_2832, w_054_2833, w_054_2834, w_054_2836, w_054_2838, w_054_2840, w_054_2842, w_054_2845, w_054_2848, w_054_2852, w_054_2853, w_054_2854, w_054_2855, w_054_2857, w_054_2859, w_054_2860, w_054_2864, w_054_2865, w_054_2866, w_054_2868, w_054_2869, w_054_2870, w_054_2871, w_054_2873, w_054_2875, w_054_2878, w_054_2880, w_054_2883, w_054_2884, w_054_2885, w_054_2887, w_054_2888, w_054_2889, w_054_2890, w_054_2891, w_054_2893, w_054_2894, w_054_2895, w_054_2896, w_054_2897, w_054_2898, w_054_2903, w_054_2904, w_054_2905, w_054_2907, w_054_2908, w_054_2909, w_054_2910, w_054_2911, w_054_2913, w_054_2914, w_054_2915, w_054_2916, w_054_2917, w_054_2918, w_054_2919, w_054_2920, w_054_2921, w_054_2924, w_054_2925, w_054_2926, w_054_2927, w_054_2931, w_054_2935, w_054_2937, w_054_2939, w_054_2940, w_054_2941, w_054_2942, w_054_2943, w_054_2944, w_054_2947, w_054_2948, w_054_2949, w_054_2950, w_054_2951, w_054_2954, w_054_2955, w_054_2956, w_054_2959, w_054_2963, w_054_2965, w_054_2966, w_054_2967, w_054_2968, w_054_2970, w_054_2971, w_054_2973, w_054_2974, w_054_2975, w_054_2978, w_054_2979, w_054_2980, w_054_2981, w_054_2982, w_054_2983, w_054_2984, w_054_2986, w_054_2991, w_054_2992, w_054_2993, w_054_2994, w_054_2995, w_054_2996, w_054_2998, w_054_3000, w_054_3001, w_054_3002, w_054_3003, w_054_3005, w_054_3007, w_054_3009, w_054_3010, w_054_3011, w_054_3013, w_054_3014, w_054_3018, w_054_3019, w_054_3020, w_054_3021, w_054_3022, w_054_3023, w_054_3024, w_054_3025, w_054_3026, w_054_3028, w_054_3033, w_054_3034, w_054_3035, w_054_3036, w_054_3038, w_054_3040, w_054_3042, w_054_3043, w_054_3044, w_054_3046, w_054_3049, w_054_3050, w_054_3051, w_054_3052, w_054_3053, w_054_3054, w_054_3056, w_054_3057, w_054_3060, w_054_3061, w_054_3062, w_054_3063, w_054_3064, w_054_3065, w_054_3066, w_054_3067, w_054_3068, w_054_3071, w_054_3073, w_054_3078, w_054_3079, w_054_3080, w_054_3084, w_054_3085, w_054_3086, w_054_3087, w_054_3088, w_054_3091, w_054_3092, w_054_3093, w_054_3094, w_054_3097, w_054_3098, w_054_3099, w_054_3100, w_054_3101, w_054_3102, w_054_3105, w_054_3106, w_054_3107, w_054_3108, w_054_3109, w_054_3110, w_054_3113, w_054_3114, w_054_3115, w_054_3117, w_054_3118, w_054_3119, w_054_3120, w_054_3122, w_054_3123, w_054_3126, w_054_3127, w_054_3128, w_054_3132, w_054_3135, w_054_3136, w_054_3137, w_054_3138, w_054_3139, w_054_3140, w_054_3143, w_054_3144, w_054_3145, w_054_3146, w_054_3147, w_054_3149, w_054_3150, w_054_3153, w_054_3154, w_054_3155, w_054_3156, w_054_3157, w_054_3158, w_054_3163, w_054_3165, w_054_3166, w_054_3167, w_054_3168, w_054_3169, w_054_3170, w_054_3172, w_054_3173, w_054_3174, w_054_3177, w_054_3180, w_054_3184, w_054_3185, w_054_3186, w_054_3187, w_054_3190, w_054_3191, w_054_3193, w_054_3195, w_054_3196, w_054_3197, w_054_3198, w_054_3199, w_054_3201, w_054_3202, w_054_3203, w_054_3204, w_054_3205, w_054_3206, w_054_3208, w_054_3209, w_054_3210, w_054_3213, w_054_3214, w_054_3215, w_054_3216, w_054_3217, w_054_3218, w_054_3219, w_054_3221, w_054_3223, w_054_3224, w_054_3225, w_054_3226, w_054_3227, w_054_3228, w_054_3230, w_054_3231, w_054_3233, w_054_3234, w_054_3237, w_054_3242, w_054_3246, w_054_3247, w_054_3248, w_054_3249, w_054_3252, w_054_3254, w_054_3255, w_054_3256, w_054_3258, w_054_3259, w_054_3260, w_054_3263, w_054_3264, w_054_3266, w_054_3267, w_054_3268, w_054_3269, w_054_3270, w_054_3271, w_054_3273, w_054_3274, w_054_3277, w_054_3278, w_054_3279, w_054_3281, w_054_3283, w_054_3286, w_054_3287, w_054_3289, w_054_3290, w_054_3294, w_054_3297, w_054_3299, w_054_3302, w_054_3305, w_054_3307, w_054_3310, w_054_3311, w_054_3313, w_054_3314, w_054_3315, w_054_3316, w_054_3317, w_054_3318, w_054_3319, w_054_3321, w_054_3322, w_054_3323, w_054_3324, w_054_3325, w_054_3326, w_054_3331, w_054_3333, w_054_3334, w_054_3337, w_054_3340, w_054_3342, w_054_3343, w_054_3344, w_054_3345, w_054_3346, w_054_3347, w_054_3348, w_054_3351, w_054_3352, w_054_3354, w_054_3355, w_054_3356, w_054_3357, w_054_3358, w_054_3360, w_054_3364, w_054_3365, w_054_3366, w_054_3367, w_054_3368, w_054_3371, w_054_3372, w_054_3373, w_054_3375, w_054_3376, w_054_3377, w_054_3380, w_054_3381, w_054_3382, w_054_3385, w_054_3387, w_054_3389, w_054_3390, w_054_3391, w_054_3392, w_054_3393, w_054_3394, w_054_3395, w_054_3396, w_054_3398, w_054_3399, w_054_3400, w_054_3401, w_054_3402, w_054_3405, w_054_3407, w_054_3409, w_054_3410, w_054_3411, w_054_3412, w_054_3413, w_054_3415, w_054_3417, w_054_3418, w_054_3420, w_054_3422, w_054_3423, w_054_3424, w_054_3426, w_054_3427, w_054_3429, w_054_3431, w_054_3432, w_054_3433, w_054_3434, w_054_3435, w_054_3436, w_054_3439, w_054_3440, w_054_3442, w_054_3443, w_054_3444, w_054_3450, w_054_3451, w_054_3452, w_054_3453, w_054_3454, w_054_3455, w_054_3457, w_054_3460, w_054_3463, w_054_3465, w_054_3466, w_054_3467, w_054_3468, w_054_3469, w_054_3470, w_054_3472, w_054_3474, w_054_3475, w_054_3477, w_054_3479, w_054_3480, w_054_3481, w_054_3482, w_054_3485, w_054_3487, w_054_3488, w_054_3492, w_054_3494, w_054_3495, w_054_3496, w_054_3497, w_054_3499, w_054_3500, w_054_3501, w_054_3505, w_054_3506, w_054_3508, w_054_3509, w_054_3510, w_054_3511, w_054_3512, w_054_3513, w_054_3515, w_054_3518, w_054_3520, w_054_3521, w_054_3522, w_054_3524, w_054_3525, w_054_3526, w_054_3529, w_054_3532, w_054_3533, w_054_3534, w_054_3535, w_054_3538, w_054_3539, w_054_3540, w_054_3541, w_054_3542, w_054_3544, w_054_3545, w_054_3546, w_054_3547, w_054_3548, w_054_3553, w_054_3555, w_054_3556, w_054_3557, w_054_3560, w_054_3565, w_054_3566, w_054_3567, w_054_3568, w_054_3570, w_054_3571, w_054_3572, w_054_3574, w_054_3575, w_054_3576, w_054_3577, w_054_3578, w_054_3580, w_054_3581, w_054_3582, w_054_3587, w_054_3588, w_054_3589, w_054_3591, w_054_3594, w_054_3599, w_054_3600, w_054_3601, w_054_3602, w_054_3605, w_054_3606, w_054_3607, w_054_3608, w_054_3609, w_054_3610, w_054_3611, w_054_3614, w_054_3615, w_054_3616, w_054_3619, w_054_3620, w_054_3621, w_054_3622, w_054_3623, w_054_3626, w_054_3630, w_054_3631, w_054_3635, w_054_3636, w_054_3638, w_054_3639, w_054_3642, w_054_3645, w_054_3651, w_054_3652, w_054_3653, w_054_3656, w_054_3657, w_054_3658, w_054_3659, w_054_3660, w_054_3661, w_054_3662, w_054_3664, w_054_3665, w_054_3666, w_054_3667, w_054_3668, w_054_3669, w_054_3670, w_054_3671, w_054_3672, w_054_3673, w_054_3674, w_054_3676, w_054_3677, w_054_3678, w_054_3680, w_054_3681, w_054_3682, w_054_3683, w_054_3684, w_054_3685, w_054_3689, w_054_3690, w_054_3691, w_054_3693, w_054_3695, w_054_3697, w_054_3698, w_054_3700, w_054_3703, w_054_3705, w_054_3707, w_054_3712, w_054_3714, w_054_3715, w_054_3717, w_054_3718, w_054_3720, w_054_3721, w_054_3722, w_054_3724, w_054_3725, w_054_3728, w_054_3729, w_054_3731, w_054_3732, w_054_3734, w_054_3737, w_054_3739, w_054_3740, w_054_3741, w_054_3744, w_054_3748, w_054_3750, w_054_3752, w_054_3753, w_054_3754, w_054_3755, w_054_3756, w_054_3757, w_054_3759, w_054_3761, w_054_3763, w_054_3764, w_054_3766, w_054_3769, w_054_3770, w_054_3772, w_054_3773, w_054_3774, w_054_3775, w_054_3777, w_054_3780, w_054_3788, w_054_3790, w_054_3792, w_054_3793, w_054_3794, w_054_3795, w_054_3796, w_054_3799, w_054_3801, w_054_3802, w_054_3803, w_054_3804, w_054_3805, w_054_3808, w_054_3809, w_054_3810, w_054_3811, w_054_3815, w_054_3817, w_054_3818, w_054_3819, w_054_3820, w_054_3822, w_054_3823, w_054_3824, w_054_3828, w_054_3829, w_054_3830, w_054_3831, w_054_3832, w_054_3833, w_054_3834, w_054_3835, w_054_3840, w_054_3842, w_054_3843, w_054_3845, w_054_3847, w_054_3849, w_054_3852, w_054_3853, w_054_3854, w_054_3855, w_054_3857, w_054_3860, w_054_3861, w_054_3865, w_054_3867, w_054_3868, w_054_3870, w_054_3871, w_054_3873, w_054_3874, w_054_3875, w_054_3876, w_054_3880, w_054_3882, w_054_3883, w_054_3885, w_054_3886, w_054_3887, w_054_3888, w_054_3890, w_054_3891, w_054_3892, w_054_3894, w_054_3895, w_054_3896, w_054_3897, w_054_3899, w_054_3900, w_054_3903, w_054_3905, w_054_3906, w_054_3908, w_054_3909, w_054_3910, w_054_3911, w_054_3912, w_054_3913, w_054_3915, w_054_3920, w_054_3921, w_054_3922, w_054_3923, w_054_3924, w_054_3925, w_054_3928, w_054_3929, w_054_3931, w_054_3932, w_054_3935, w_054_3936, w_054_3938, w_054_3940, w_054_3942, w_054_3943, w_054_3944, w_054_3946, w_054_3948, w_054_3949, w_054_3953, w_054_3955, w_054_3958, w_054_3961, w_054_3964, w_054_3966, w_054_3968, w_054_3969, w_054_3970, w_054_3974, w_054_3975, w_054_3980, w_054_3981, w_054_3982, w_054_3984, w_054_3987, w_054_3991, w_054_3992, w_054_3994, w_054_3996, w_054_3997, w_054_3998, w_054_3999, w_054_4000, w_054_4001, w_054_4003, w_054_4004, w_054_4005, w_054_4006, w_054_4007, w_054_4009, w_054_4010, w_054_4012, w_054_4014, w_054_4018, w_054_4019, w_054_4020, w_054_4021, w_054_4022, w_054_4023, w_054_4024, w_054_4028, w_054_4030, w_054_4031, w_054_4032, w_054_4033, w_054_4034, w_054_4036, w_054_4037, w_054_4038, w_054_4039, w_054_4040, w_054_4041, w_054_4042, w_054_4045, w_054_4046, w_054_4047, w_054_4048, w_054_4051, w_054_4053, w_054_4055, w_054_4059, w_054_4060, w_054_4063, w_054_4064, w_054_4065, w_054_4067, w_054_4069, w_054_4071, w_054_4072, w_054_4073, w_054_4074, w_054_4075, w_054_4076, w_054_4078, w_054_4079, w_054_4083, w_054_4084, w_054_4085, w_054_4086, w_054_4088, w_054_4091, w_054_4093, w_054_4094, w_054_4095, w_054_4097, w_054_4099, w_054_4100, w_054_4101, w_054_4103, w_054_4104, w_054_4107, w_054_4108, w_054_4110, w_054_4111, w_054_4112, w_054_4115, w_054_4116, w_054_4118, w_054_4120, w_054_4121, w_054_4122, w_054_4125, w_054_4127, w_054_4129, w_054_4130, w_054_4131, w_054_4132, w_054_4133, w_054_4134, w_054_4135, w_054_4136, w_054_4137, w_054_4138, w_054_4139, w_054_4140, w_054_4141, w_054_4143, w_054_4144, w_054_4146, w_054_4148, w_054_4150, w_054_4151, w_054_4152, w_054_4153, w_054_4154, w_054_4155, w_054_4156, w_054_4158, w_054_4160, w_054_4163, w_054_4164, w_054_4165, w_054_4166, w_054_4167, w_054_4170, w_054_4171, w_054_4172, w_054_4173, w_054_4175, w_054_4176, w_054_4179, w_054_4183, w_054_4185, w_054_4186, w_054_4190, w_054_4191, w_054_4192, w_054_4193, w_054_4194, w_054_4196, w_054_4198, w_054_4202, w_054_4203, w_054_4204, w_054_4205, w_054_4207, w_054_4209, w_054_4211, w_054_4212, w_054_4213, w_054_4214, w_054_4215, w_054_4216, w_054_4218, w_054_4220, w_054_4223, w_054_4227, w_054_4229, w_054_4230, w_054_4232, w_054_4233, w_054_4234, w_054_4236, w_054_4237, w_054_4238, w_054_4239, w_054_4241, w_054_4242, w_054_4243, w_054_4244, w_054_4246, w_054_4248, w_054_4249, w_054_4250, w_054_4251, w_054_4252, w_054_4254, w_054_4256, w_054_4257, w_054_4258, w_054_4259, w_054_4260, w_054_4261, w_054_4263, w_054_4264, w_054_4265, w_054_4266, w_054_4268, w_054_4269, w_054_4270, w_054_4271, w_054_4272, w_054_4274, w_054_4275, w_054_4276, w_054_4277, w_054_4278, w_054_4279, w_054_4280, w_054_4282, w_054_4284, w_054_4285, w_054_4286, w_054_4287, w_054_4288, w_054_4289, w_054_4291, w_054_4292, w_054_4293, w_054_4294, w_054_4296, w_054_4298, w_054_4301, w_054_4302, w_054_4303, w_054_4304, w_054_4305, w_054_4306, w_054_4307, w_054_4308, w_054_4310, w_054_4311, w_054_4312, w_054_4313, w_054_4314, w_054_4315, w_054_4316, w_054_4319, w_054_4320, w_054_4321, w_054_4322, w_054_4325, w_054_4326, w_054_4328, w_054_4329, w_054_4332, w_054_4333, w_054_4335, w_054_4336, w_054_4337, w_054_4338, w_054_4339, w_054_4340, w_054_4341, w_054_4345, w_054_4346, w_054_4347, w_054_4348, w_054_4349, w_054_4350, w_054_4351, w_054_4353, w_054_4354, w_054_4355, w_054_4356, w_054_4357, w_054_4358, w_054_4359, w_054_4360, w_054_4361, w_054_4364, w_054_4365, w_054_4366, w_054_4371, w_054_4372, w_054_4373, w_054_4374, w_054_4376, w_054_4377, w_054_4378, w_054_4379, w_054_4382, w_054_4384, w_054_4385, w_054_4386, w_054_4387, w_054_4388, w_054_4389, w_054_4393, w_054_4394, w_054_4400, w_054_4401, w_054_4402, w_054_4404, w_054_4406, w_054_4408, w_054_4409, w_054_4411, w_054_4414, w_054_4415, w_054_4416, w_054_4419, w_054_4421, w_054_4422, w_054_4423, w_054_4424, w_054_4425, w_054_4426, w_054_4427, w_054_4430, w_054_4434, w_054_4435, w_054_4436, w_054_4437, w_054_4438, w_054_4439, w_054_4442, w_054_4444, w_054_4445, w_054_4446, w_054_4450, w_054_4451, w_054_4456, w_054_4457, w_054_4458, w_054_4459, w_054_4461, w_054_4462, w_054_4463, w_054_4464, w_054_4465, w_054_4466, w_054_4467, w_054_4468, w_054_4469, w_054_4470, w_054_4471, w_054_4473, w_054_4475, w_054_4476, w_054_4479, w_054_4480, w_054_4481, w_054_4482, w_054_4484, w_054_4486, w_054_4488, w_054_4495, w_054_4496, w_054_4498, w_054_4499, w_054_4500, w_054_4501, w_054_4502, w_054_4503, w_054_4504, w_054_4505, w_054_4506, w_054_4509, w_054_4510, w_054_4512, w_054_4513, w_054_4514, w_054_4515, w_054_4516, w_054_4517, w_054_4520, w_054_4522, w_054_4523, w_054_4525, w_054_4526, w_054_4527, w_054_4531, w_054_4532, w_054_4533, w_054_4535, w_054_4539, w_054_4541, w_054_4543, w_054_4544, w_054_4545, w_054_4546, w_054_4548, w_054_4550, w_054_4551, w_054_4553, w_054_4554, w_054_4555, w_054_4556, w_054_4559, w_054_4560, w_054_4561, w_054_4564, w_054_4566, w_054_4568, w_054_4569, w_054_4570, w_054_4571, w_054_4572, w_054_4575, w_054_4578, w_054_4579, w_054_4580, w_054_4581, w_054_4583, w_054_4584, w_054_4585, w_054_4586, w_054_4587, w_054_4588, w_054_4589, w_054_4591, w_054_4592, w_054_4593, w_054_4594, w_054_4597, w_054_4598, w_054_4599, w_054_4600, w_054_4602, w_054_4605, w_054_4606, w_054_4610, w_054_4616, w_054_4618, w_054_4627, w_054_4628, w_054_4629, w_054_4630, w_054_4631, w_054_4633, w_054_4637, w_054_4638, w_054_4639, w_054_4643, w_054_4645, w_054_4649, w_054_4651, w_054_4652, w_054_4653, w_054_4654, w_054_4655, w_054_4660, w_054_4661, w_054_4662, w_054_4666, w_054_4669, w_054_4670, w_054_4674, w_054_4675, w_054_4678, w_054_4684, w_054_4688, w_054_4690, w_054_4691, w_054_4693, w_054_4695, w_054_4697, w_054_4698, w_054_4715, w_054_4717, w_054_4721, w_054_4726, w_054_4730, w_054_4731, w_054_4732, w_054_4737, w_054_4739, w_054_4740, w_054_4741, w_054_4743, w_054_4744, w_054_4749, w_054_4751, w_054_4752, w_054_4755, w_054_4756, w_054_4759, w_054_4760, w_054_4762, w_054_4764, w_054_4766, w_054_4768, w_054_4769, w_054_4771, w_054_4772, w_054_4778, w_054_4782, w_054_4783, w_054_4784, w_054_4788, w_054_4792, w_054_4793, w_054_4797, w_054_4798, w_054_4800, w_054_4801, w_054_4802, w_054_4804, w_054_4808, w_054_4809, w_054_4811, w_054_4813, w_054_4814, w_054_4815, w_054_4816, w_054_4818, w_054_4822, w_054_4824, w_054_4825, w_054_4826, w_054_4832, w_054_4833, w_054_4834, w_054_4837, w_054_4840, w_054_4843, w_054_4847, w_054_4850, w_054_4852, w_054_4854, w_054_4856, w_054_4860, w_054_4862, w_054_4868, w_054_4871, w_054_4872, w_054_4882, w_054_4885, w_054_4890, w_054_4895, w_054_4896, w_054_4897, w_054_4900, w_054_4902, w_054_4903, w_054_4909, w_054_4910, w_054_4911, w_054_4913, w_054_4914, w_054_4918, w_054_4924, w_054_4925, w_054_4927, w_054_4928, w_054_4929, w_054_4930, w_054_4931, w_054_4936, w_054_4940, w_054_4941, w_054_4942, w_054_4943, w_054_4945, w_054_4946, w_054_4952, w_054_4953, w_054_4958, w_054_4962, w_054_4964, w_054_4970, w_054_4972, w_054_4974, w_054_4977, w_054_4978, w_054_4984, w_054_4986, w_054_4990, w_054_4992, w_054_4999, w_054_5000, w_054_5002, w_054_5004, w_054_5005, w_054_5006, w_054_5008, w_054_5009, w_054_5011, w_054_5013, w_054_5014, w_054_5016, w_054_5021, w_054_5023, w_054_5024, w_054_5026, w_054_5029, w_054_5030, w_054_5032, w_054_5035, w_054_5036, w_054_5039, w_054_5040, w_054_5044, w_054_5045, w_054_5047, w_054_5051, w_054_5056, w_054_5057, w_054_5058, w_054_5066, w_054_5068, w_054_5070, w_054_5072, w_054_5073, w_054_5077, w_054_5079, w_054_5081, w_054_5085, w_054_5089, w_054_5092, w_054_5093, w_054_5097, w_054_5099, w_054_5100, w_054_5102, w_054_5103, w_054_5104, w_054_5109, w_054_5111, w_054_5114, w_054_5116, w_054_5117, w_054_5118, w_054_5119, w_054_5121, w_054_5124, w_054_5128, w_054_5129, w_054_5132, w_054_5135, w_054_5136, w_054_5137, w_054_5138, w_054_5139, w_054_5148, w_054_5150, w_054_5156, w_054_5159, w_054_5163, w_054_5166, w_054_5167, w_054_5169, w_054_5172, w_054_5173, w_054_5174, w_054_5175, w_054_5179, w_054_5183, w_054_5184, w_054_5192, w_054_5193, w_054_5194, w_054_5196, w_054_5197, w_054_5198, w_054_5200, w_054_5204, w_054_5206, w_054_5208, w_054_5209, w_054_5211, w_054_5216, w_054_5221, w_054_5222, w_054_5223, w_054_5230, w_054_5233, w_054_5235, w_054_5236, w_054_5237, w_054_5239, w_054_5240, w_054_5242, w_054_5244, w_054_5249, w_054_5250, w_054_5252, w_054_5255, w_054_5258, w_054_5259, w_054_5262, w_054_5266, w_054_5268, w_054_5270, w_054_5271, w_054_5272, w_054_5273, w_054_5278, w_054_5282, w_054_5288, w_054_5289, w_054_5291, w_054_5292, w_054_5294, w_054_5295, w_054_5300, w_054_5302, w_054_5303, w_054_5309, w_054_5311, w_054_5314, w_054_5319, w_054_5320, w_054_5324, w_054_5325, w_054_5328, w_054_5329, w_054_5330, w_054_5333, w_054_5336, w_054_5339, w_054_5343, w_054_5344, w_054_5347;
  wire w_055_001, w_055_003, w_055_004, w_055_005, w_055_007, w_055_009, w_055_010, w_055_011, w_055_012, w_055_013, w_055_015, w_055_016, w_055_018, w_055_019, w_055_020, w_055_022, w_055_024, w_055_025, w_055_026, w_055_027, w_055_028, w_055_029, w_055_030, w_055_031, w_055_033, w_055_034, w_055_035, w_055_036, w_055_037, w_055_038, w_055_039, w_055_040, w_055_042, w_055_043, w_055_045, w_055_046, w_055_047, w_055_048, w_055_049, w_055_050, w_055_051, w_055_052, w_055_053, w_055_054, w_055_055, w_055_056, w_055_059, w_055_061, w_055_063, w_055_064, w_055_065, w_055_067, w_055_069, w_055_070, w_055_071, w_055_073, w_055_074, w_055_075, w_055_077, w_055_078, w_055_079, w_055_080, w_055_083, w_055_084, w_055_085, w_055_086, w_055_088, w_055_090, w_055_091, w_055_095, w_055_098, w_055_099, w_055_104, w_055_105, w_055_106, w_055_107, w_055_108, w_055_110, w_055_112, w_055_114, w_055_115, w_055_116, w_055_117, w_055_119, w_055_120, w_055_121, w_055_122, w_055_123, w_055_126, w_055_127, w_055_128, w_055_130, w_055_131, w_055_133, w_055_134, w_055_137, w_055_138, w_055_142, w_055_144, w_055_145, w_055_147, w_055_148, w_055_149, w_055_150, w_055_151, w_055_152, w_055_153, w_055_154, w_055_156, w_055_159, w_055_162, w_055_164, w_055_167, w_055_168, w_055_171, w_055_172, w_055_173, w_055_175, w_055_180, w_055_182, w_055_184, w_055_185, w_055_187, w_055_188, w_055_189, w_055_190, w_055_191, w_055_192, w_055_201, w_055_203, w_055_204, w_055_207, w_055_208, w_055_211, w_055_215, w_055_218, w_055_220, w_055_221, w_055_222, w_055_226, w_055_227, w_055_228, w_055_229, w_055_230, w_055_232, w_055_233, w_055_234, w_055_235, w_055_237, w_055_238, w_055_240, w_055_241, w_055_251, w_055_252, w_055_254, w_055_255, w_055_259, w_055_261, w_055_262, w_055_263, w_055_265, w_055_266, w_055_267, w_055_271, w_055_272, w_055_275, w_055_276, w_055_277, w_055_278, w_055_281, w_055_282, w_055_283, w_055_284, w_055_286, w_055_287, w_055_288, w_055_289, w_055_291, w_055_292, w_055_295, w_055_296, w_055_297, w_055_298, w_055_299, w_055_302, w_055_303, w_055_304, w_055_305, w_055_306, w_055_307, w_055_310, w_055_311, w_055_312, w_055_313, w_055_314, w_055_315, w_055_316, w_055_319, w_055_320, w_055_321, w_055_322, w_055_323, w_055_324, w_055_325, w_055_326, w_055_327, w_055_328, w_055_330, w_055_333, w_055_339, w_055_341, w_055_343, w_055_344, w_055_345, w_055_346, w_055_347, w_055_348, w_055_351, w_055_354, w_055_355, w_055_357, w_055_358, w_055_359, w_055_360, w_055_361, w_055_362, w_055_363, w_055_364, w_055_366, w_055_367, w_055_368, w_055_370, w_055_372, w_055_376, w_055_378, w_055_379, w_055_382, w_055_383, w_055_384, w_055_389, w_055_390, w_055_391, w_055_392, w_055_393, w_055_394, w_055_398, w_055_400, w_055_401, w_055_403, w_055_407, w_055_409, w_055_410, w_055_412, w_055_413, w_055_414, w_055_415, w_055_417, w_055_418, w_055_419, w_055_420, w_055_421, w_055_422, w_055_423, w_055_424, w_055_426, w_055_428, w_055_429, w_055_431, w_055_432, w_055_433, w_055_434, w_055_436, w_055_437, w_055_438, w_055_439, w_055_441, w_055_442, w_055_443, w_055_444, w_055_445, w_055_446, w_055_447, w_055_450, w_055_451, w_055_452, w_055_453, w_055_454, w_055_457, w_055_462, w_055_463, w_055_466, w_055_467, w_055_468, w_055_469, w_055_471, w_055_474, w_055_477, w_055_478, w_055_479, w_055_480, w_055_483, w_055_486, w_055_487, w_055_489, w_055_492, w_055_493, w_055_494, w_055_497, w_055_498, w_055_499, w_055_500, w_055_501, w_055_502, w_055_503, w_055_504, w_055_505, w_055_506, w_055_508, w_055_509, w_055_511, w_055_513, w_055_514, w_055_516, w_055_517, w_055_519, w_055_520, w_055_521, w_055_522, w_055_524, w_055_526, w_055_528, w_055_529, w_055_532, w_055_533, w_055_536, w_055_537, w_055_538, w_055_539, w_055_541, w_055_542, w_055_543, w_055_544, w_055_546, w_055_547, w_055_548, w_055_549, w_055_551, w_055_552, w_055_555, w_055_556, w_055_557, w_055_560, w_055_561, w_055_563, w_055_567, w_055_569, w_055_570, w_055_571, w_055_573, w_055_574, w_055_575, w_055_576, w_055_577, w_055_578, w_055_579, w_055_583, w_055_584, w_055_585, w_055_586, w_055_587, w_055_588, w_055_589, w_055_592, w_055_593, w_055_594, w_055_595, w_055_596, w_055_597, w_055_598, w_055_600, w_055_605, w_055_606, w_055_607, w_055_608, w_055_609, w_055_611, w_055_612, w_055_614, w_055_616, w_055_619, w_055_621, w_055_623, w_055_624, w_055_625, w_055_627, w_055_628, w_055_630, w_055_631, w_055_632, w_055_636, w_055_637, w_055_638, w_055_639, w_055_640, w_055_641, w_055_642, w_055_643, w_055_645, w_055_649, w_055_650, w_055_651, w_055_652, w_055_653, w_055_654, w_055_655, w_055_656, w_055_659, w_055_661, w_055_663, w_055_664, w_055_665, w_055_666, w_055_669, w_055_670, w_055_671, w_055_674, w_055_676, w_055_677, w_055_678, w_055_680, w_055_682, w_055_683, w_055_684, w_055_686, w_055_687, w_055_689, w_055_690, w_055_691, w_055_694, w_055_695, w_055_696, w_055_697, w_055_698, w_055_700, w_055_704, w_055_705, w_055_706, w_055_708, w_055_709, w_055_713, w_055_715, w_055_716, w_055_717, w_055_719, w_055_725, w_055_726, w_055_727, w_055_728, w_055_729, w_055_730, w_055_731, w_055_732, w_055_733, w_055_734, w_055_737, w_055_738, w_055_741, w_055_743, w_055_745, w_055_746, w_055_747, w_055_748, w_055_750, w_055_751, w_055_752, w_055_754, w_055_756, w_055_758, w_055_761, w_055_763, w_055_765, w_055_767, w_055_769, w_055_770, w_055_772, w_055_775, w_055_776, w_055_777, w_055_779, w_055_781, w_055_783, w_055_785, w_055_787, w_055_790, w_055_791, w_055_792, w_055_793, w_055_794, w_055_796, w_055_797, w_055_798, w_055_800, w_055_802, w_055_804, w_055_805, w_055_806, w_055_808, w_055_811, w_055_812, w_055_813, w_055_815, w_055_816, w_055_817, w_055_818, w_055_819, w_055_820, w_055_821, w_055_822, w_055_824, w_055_828, w_055_829, w_055_830, w_055_831, w_055_832, w_055_833, w_055_834, w_055_835, w_055_836, w_055_839, w_055_840, w_055_841, w_055_843, w_055_848, w_055_849, w_055_853, w_055_854, w_055_855, w_055_857, w_055_860, w_055_861, w_055_863, w_055_864, w_055_865, w_055_866, w_055_867, w_055_869, w_055_870, w_055_871, w_055_872, w_055_875, w_055_877, w_055_879, w_055_880, w_055_885, w_055_886, w_055_889, w_055_890, w_055_891, w_055_892, w_055_893, w_055_896, w_055_897, w_055_898, w_055_900, w_055_901, w_055_902, w_055_903, w_055_906, w_055_907, w_055_908, w_055_910, w_055_911, w_055_913, w_055_914, w_055_915, w_055_917, w_055_919, w_055_926, w_055_927, w_055_928, w_055_930, w_055_931, w_055_934, w_055_935, w_055_936, w_055_937, w_055_938, w_055_939, w_055_942, w_055_944, w_055_945, w_055_946, w_055_948, w_055_949, w_055_952, w_055_955, w_055_956, w_055_958, w_055_960, w_055_961, w_055_962, w_055_965, w_055_968, w_055_969, w_055_973, w_055_975, w_055_978, w_055_979, w_055_980, w_055_984, w_055_985, w_055_987, w_055_988, w_055_989, w_055_991, w_055_994, w_055_995, w_055_997, w_055_999, w_055_1000, w_055_1003, w_055_1004, w_055_1005, w_055_1006, w_055_1007, w_055_1008, w_055_1009, w_055_1010, w_055_1012, w_055_1013, w_055_1014, w_055_1015, w_055_1016, w_055_1017, w_055_1019, w_055_1020, w_055_1022, w_055_1023, w_055_1024, w_055_1025, w_055_1027, w_055_1028, w_055_1030, w_055_1031, w_055_1032, w_055_1033, w_055_1034, w_055_1035, w_055_1037, w_055_1038, w_055_1039, w_055_1040, w_055_1042, w_055_1043, w_055_1045, w_055_1049, w_055_1050, w_055_1051, w_055_1052, w_055_1053, w_055_1054, w_055_1056, w_055_1057, w_055_1059, w_055_1060, w_055_1061, w_055_1062, w_055_1063, w_055_1065, w_055_1067, w_055_1068, w_055_1069, w_055_1070, w_055_1071, w_055_1074, w_055_1075, w_055_1076, w_055_1077, w_055_1078, w_055_1079, w_055_1080, w_055_1083, w_055_1085, w_055_1086, w_055_1087, w_055_1088, w_055_1089, w_055_1090, w_055_1091, w_055_1094, w_055_1096, w_055_1097, w_055_1098, w_055_1100, w_055_1102, w_055_1103, w_055_1104, w_055_1105, w_055_1107, w_055_1109, w_055_1110, w_055_1111, w_055_1116, w_055_1118, w_055_1119, w_055_1120, w_055_1122, w_055_1124, w_055_1125, w_055_1126, w_055_1127, w_055_1128, w_055_1135, w_055_1137, w_055_1138, w_055_1140, w_055_1141, w_055_1143, w_055_1144, w_055_1145, w_055_1147, w_055_1149, w_055_1151, w_055_1152, w_055_1153, w_055_1155, w_055_1156, w_055_1157, w_055_1158, w_055_1159, w_055_1160, w_055_1161, w_055_1162, w_055_1163, w_055_1165, w_055_1166, w_055_1167, w_055_1170, w_055_1173, w_055_1177, w_055_1178, w_055_1180, w_055_1182, w_055_1183, w_055_1185, w_055_1186, w_055_1187, w_055_1188, w_055_1190, w_055_1191, w_055_1192, w_055_1193, w_055_1195, w_055_1196, w_055_1197, w_055_1198, w_055_1199, w_055_1200, w_055_1202, w_055_1203, w_055_1204, w_055_1207, w_055_1208, w_055_1209, w_055_1210, w_055_1211, w_055_1212, w_055_1213, w_055_1214, w_055_1216, w_055_1217, w_055_1219, w_055_1221, w_055_1222, w_055_1225, w_055_1226, w_055_1227, w_055_1228, w_055_1230, w_055_1231, w_055_1232, w_055_1233, w_055_1234, w_055_1237, w_055_1238, w_055_1239, w_055_1240, w_055_1241, w_055_1242, w_055_1243, w_055_1244, w_055_1245, w_055_1246, w_055_1248, w_055_1249, w_055_1253, w_055_1255, w_055_1256, w_055_1257, w_055_1258, w_055_1260, w_055_1264, w_055_1265, w_055_1266, w_055_1267, w_055_1271, w_055_1272, w_055_1274, w_055_1276, w_055_1279, w_055_1281, w_055_1282, w_055_1283, w_055_1285, w_055_1286, w_055_1288, w_055_1289, w_055_1291, w_055_1294, w_055_1295, w_055_1298, w_055_1305, w_055_1308, w_055_1309, w_055_1310, w_055_1311, w_055_1312, w_055_1316, w_055_1317, w_055_1318, w_055_1321, w_055_1322, w_055_1323, w_055_1324, w_055_1325, w_055_1326, w_055_1327, w_055_1329, w_055_1330, w_055_1332, w_055_1333, w_055_1334, w_055_1335, w_055_1336, w_055_1337, w_055_1338, w_055_1342, w_055_1343, w_055_1344, w_055_1345, w_055_1346, w_055_1348, w_055_1350, w_055_1353, w_055_1354, w_055_1356, w_055_1357, w_055_1359, w_055_1360, w_055_1361, w_055_1365, w_055_1366, w_055_1368, w_055_1370, w_055_1372, w_055_1374, w_055_1375, w_055_1377, w_055_1378, w_055_1379, w_055_1380, w_055_1381, w_055_1384, w_055_1386, w_055_1387, w_055_1388, w_055_1389, w_055_1393, w_055_1396, w_055_1398, w_055_1400, w_055_1404, w_055_1405, w_055_1406, w_055_1407, w_055_1408, w_055_1409, w_055_1410, w_055_1411, w_055_1412, w_055_1414, w_055_1416, w_055_1417, w_055_1418, w_055_1419, w_055_1420, w_055_1422, w_055_1424, w_055_1425, w_055_1426, w_055_1427, w_055_1429, w_055_1430, w_055_1431, w_055_1432, w_055_1433, w_055_1435, w_055_1436, w_055_1437, w_055_1438, w_055_1439, w_055_1440, w_055_1441, w_055_1442, w_055_1445, w_055_1446, w_055_1447, w_055_1449, w_055_1450, w_055_1452, w_055_1454, w_055_1455, w_055_1457, w_055_1459, w_055_1460, w_055_1461, w_055_1465, w_055_1466, w_055_1468, w_055_1471, w_055_1474, w_055_1478, w_055_1479, w_055_1480, w_055_1481, w_055_1482, w_055_1484, w_055_1486, w_055_1487, w_055_1488, w_055_1489, w_055_1490, w_055_1493, w_055_1495, w_055_1498, w_055_1503, w_055_1504, w_055_1505, w_055_1507, w_055_1508, w_055_1509, w_055_1510, w_055_1511, w_055_1512, w_055_1513, w_055_1515, w_055_1516, w_055_1517, w_055_1519, w_055_1521, w_055_1522, w_055_1524, w_055_1525, w_055_1527, w_055_1529, w_055_1530, w_055_1531, w_055_1534, w_055_1536, w_055_1541, w_055_1544, w_055_1545, w_055_1546, w_055_1548, w_055_1551, w_055_1552, w_055_1554, w_055_1555, w_055_1556, w_055_1557, w_055_1558, w_055_1561, w_055_1562, w_055_1563, w_055_1566, w_055_1567, w_055_1568, w_055_1569, w_055_1572, w_055_1573, w_055_1575, w_055_1576, w_055_1577, w_055_1578, w_055_1582, w_055_1586, w_055_1589, w_055_1590, w_055_1591, w_055_1593, w_055_1594, w_055_1596, w_055_1597, w_055_1598, w_055_1599, w_055_1601, w_055_1604, w_055_1605, w_055_1607, w_055_1609, w_055_1610, w_055_1611, w_055_1613, w_055_1615, w_055_1619, w_055_1622, w_055_1623, w_055_1624, w_055_1625, w_055_1627, w_055_1631, w_055_1633, w_055_1634, w_055_1636, w_055_1638, w_055_1641, w_055_1642, w_055_1644, w_055_1645, w_055_1647, w_055_1648, w_055_1649, w_055_1650, w_055_1651, w_055_1657, w_055_1659, w_055_1660, w_055_1661, w_055_1662, w_055_1663, w_055_1664, w_055_1668, w_055_1669, w_055_1670, w_055_1671, w_055_1673, w_055_1675, w_055_1676, w_055_1677, w_055_1679, w_055_1680, w_055_1681, w_055_1684, w_055_1687, w_055_1689, w_055_1690, w_055_1691, w_055_1692, w_055_1693, w_055_1694, w_055_1696, w_055_1700, w_055_1702, w_055_1704, w_055_1705, w_055_1710, w_055_1711, w_055_1712, w_055_1716, w_055_1718, w_055_1719, w_055_1720, w_055_1722, w_055_1723, w_055_1724, w_055_1725, w_055_1729, w_055_1731, w_055_1732, w_055_1733, w_055_1734, w_055_1736, w_055_1738, w_055_1740, w_055_1742, w_055_1743, w_055_1744, w_055_1745, w_055_1747, w_055_1748, w_055_1749, w_055_1750, w_055_1753, w_055_1754, w_055_1755, w_055_1756, w_055_1758, w_055_1759, w_055_1760, w_055_1761, w_055_1762, w_055_1763, w_055_1764, w_055_1765, w_055_1767, w_055_1768, w_055_1770, w_055_1771, w_055_1773, w_055_1774, w_055_1775, w_055_1778, w_055_1781, w_055_1782, w_055_1783, w_055_1784, w_055_1785, w_055_1786, w_055_1787, w_055_1792, w_055_1793, w_055_1794, w_055_1796, w_055_1797, w_055_1798, w_055_1799, w_055_1801, w_055_1803, w_055_1804, w_055_1805, w_055_1807, w_055_1808, w_055_1809, w_055_1811, w_055_1812, w_055_1816, w_055_1819, w_055_1820, w_055_1822, w_055_1824, w_055_1827, w_055_1830, w_055_1832, w_055_1834, w_055_1835, w_055_1836, w_055_1837, w_055_1839, w_055_1841, w_055_1842, w_055_1844, w_055_1847, w_055_1849, w_055_1851, w_055_1852, w_055_1853, w_055_1854, w_055_1855, w_055_1856, w_055_1857, w_055_1858, w_055_1863, w_055_1864, w_055_1865, w_055_1866, w_055_1867, w_055_1868, w_055_1870, w_055_1871, w_055_1872, w_055_1874, w_055_1875, w_055_1877, w_055_1878, w_055_1879, w_055_1883, w_055_1885, w_055_1886, w_055_1887, w_055_1888, w_055_1889, w_055_1890, w_055_1891, w_055_1893, w_055_1896, w_055_1897, w_055_1898, w_055_1899, w_055_1900, w_055_1903, w_055_1904, w_055_1906, w_055_1907, w_055_1908, w_055_1911, w_055_1912, w_055_1913, w_055_1914, w_055_1915, w_055_1916, w_055_1918, w_055_1919, w_055_1922, w_055_1923, w_055_1924, w_055_1927, w_055_1929, w_055_1930, w_055_1934, w_055_1935, w_055_1936, w_055_1937, w_055_1938, w_055_1939, w_055_1940, w_055_1941, w_055_1942, w_055_1945, w_055_1947, w_055_1949, w_055_1950, w_055_1952, w_055_1954, w_055_1955, w_055_1957, w_055_1958, w_055_1959, w_055_1961, w_055_1962, w_055_1964, w_055_1968, w_055_1969, w_055_1970, w_055_1971, w_055_1972, w_055_1973, w_055_1974, w_055_1975, w_055_1976, w_055_1977, w_055_1979, w_055_1980, w_055_1981, w_055_1982, w_055_1983, w_055_1984, w_055_1986, w_055_1992, w_055_1994, w_055_1995, w_055_1996, w_055_1998, w_055_2002, w_055_2003, w_055_2004, w_055_2006, w_055_2007, w_055_2008, w_055_2009, w_055_2013, w_055_2014, w_055_2015, w_055_2016, w_055_2017, w_055_2018, w_055_2020, w_055_2021, w_055_2022, w_055_2024, w_055_2025, w_055_2026, w_055_2028, w_055_2032, w_055_2033, w_055_2034, w_055_2035, w_055_2037, w_055_2038, w_055_2039, w_055_2041, w_055_2042, w_055_2043, w_055_2044, w_055_2045, w_055_2047, w_055_2049, w_055_2051, w_055_2052, w_055_2053, w_055_2054, w_055_2058, w_055_2059, w_055_2060, w_055_2062, w_055_2064, w_055_2065, w_055_2066, w_055_2068, w_055_2069, w_055_2070, w_055_2072, w_055_2075, w_055_2077, w_055_2078, w_055_2079, w_055_2080, w_055_2081, w_055_2082, w_055_2083, w_055_2084, w_055_2085, w_055_2086, w_055_2087, w_055_2088, w_055_2092, w_055_2095, w_055_2096, w_055_2097, w_055_2099, w_055_2100, w_055_2101, w_055_2102, w_055_2103, w_055_2104, w_055_2105, w_055_2107, w_055_2109, w_055_2110, w_055_2113, w_055_2114, w_055_2115, w_055_2117, w_055_2118, w_055_2119, w_055_2120, w_055_2121, w_055_2122, w_055_2123, w_055_2124, w_055_2127, w_055_2128, w_055_2130, w_055_2132, w_055_2133, w_055_2134, w_055_2135, w_055_2136, w_055_2139, w_055_2140, w_055_2142, w_055_2143, w_055_2144, w_055_2146, w_055_2152, w_055_2153, w_055_2154, w_055_2156, w_055_2157, w_055_2158, w_055_2159, w_055_2160, w_055_2162, w_055_2163, w_055_2164, w_055_2166, w_055_2167, w_055_2169, w_055_2170, w_055_2171, w_055_2172, w_055_2173, w_055_2175, w_055_2176, w_055_2177, w_055_2179, w_055_2180, w_055_2181, w_055_2182, w_055_2183, w_055_2184, w_055_2185, w_055_2186, w_055_2189, w_055_2190, w_055_2191, w_055_2192, w_055_2193, w_055_2194, w_055_2196, w_055_2197, w_055_2199, w_055_2200, w_055_2201, w_055_2203, w_055_2204, w_055_2205, w_055_2206, w_055_2210, w_055_2211, w_055_2213, w_055_2214, w_055_2215, w_055_2216, w_055_2218, w_055_2219, w_055_2220, w_055_2222, w_055_2223, w_055_2224, w_055_2225, w_055_2226, w_055_2227, w_055_2228, w_055_2230, w_055_2232, w_055_2233, w_055_2234, w_055_2235, w_055_2236, w_055_2238, w_055_2242, w_055_2246, w_055_2250, w_055_2251, w_055_2253, w_055_2254, w_055_2255, w_055_2256, w_055_2259, w_055_2260, w_055_2261, w_055_2262, w_055_2264, w_055_2266, w_055_2268, w_055_2269, w_055_2271, w_055_2272, w_055_2274, w_055_2275, w_055_2277, w_055_2278, w_055_2279, w_055_2281, w_055_2282, w_055_2283, w_055_2284, w_055_2286, w_055_2287, w_055_2288, w_055_2290, w_055_2291, w_055_2292, w_055_2293, w_055_2295, w_055_2297, w_055_2301, w_055_2304, w_055_2306, w_055_2307, w_055_2311, w_055_2313, w_055_2314, w_055_2315, w_055_2316, w_055_2317, w_055_2320, w_055_2323, w_055_2325, w_055_2326, w_055_2329, w_055_2331, w_055_2332, w_055_2333, w_055_2334, w_055_2335, w_055_2337, w_055_2338, w_055_2339, w_055_2342, w_055_2343, w_055_2345, w_055_2346, w_055_2349, w_055_2350, w_055_2352, w_055_2353, w_055_2354, w_055_2356, w_055_2359, w_055_2360, w_055_2361, w_055_2362, w_055_2363, w_055_2365, w_055_2367, w_055_2369, w_055_2370, w_055_2372, w_055_2373, w_055_2375, w_055_2378, w_055_2379, w_055_2382, w_055_2384, w_055_2386, w_055_2390, w_055_2391, w_055_2392, w_055_2394, w_055_2395, w_055_2396, w_055_2397, w_055_2398, w_055_2400, w_055_2403, w_055_2404, w_055_2405, w_055_2407, w_055_2408, w_055_2409, w_055_2411, w_055_2412, w_055_2413, w_055_2415, w_055_2417, w_055_2418, w_055_2419, w_055_2422, w_055_2425, w_055_2427, w_055_2430, w_055_2431, w_055_2432, w_055_2437, w_055_2438, w_055_2439, w_055_2440, w_055_2441, w_055_2442, w_055_2443, w_055_2444, w_055_2446, w_055_2447, w_055_2448, w_055_2456, w_055_2462, w_055_2465, w_055_2466, w_055_2471, w_055_2472, w_055_2474, w_055_2475, w_055_2476, w_055_2479, w_055_2481, w_055_2482, w_055_2484, w_055_2487, w_055_2489, w_055_2490, w_055_2491, w_055_2493, w_055_2494, w_055_2495, w_055_2496, w_055_2498, w_055_2502, w_055_2504, w_055_2505, w_055_2506, w_055_2507, w_055_2508, w_055_2510, w_055_2511, w_055_2513, w_055_2514, w_055_2515, w_055_2516, w_055_2519, w_055_2520, w_055_2521, w_055_2522, w_055_2523, w_055_2524, w_055_2528, w_055_2530, w_055_2531, w_055_2532, w_055_2533, w_055_2534, w_055_2536, w_055_2537, w_055_2538, w_055_2539, w_055_2540, w_055_2543, w_055_2544, w_055_2545, w_055_2546, w_055_2547, w_055_2549, w_055_2551, w_055_2552, w_055_2554, w_055_2555, w_055_2556, w_055_2557, w_055_2558, w_055_2559, w_055_2560, w_055_2562, w_055_2563, w_055_2564, w_055_2566, w_055_2570, w_055_2571, w_055_2573, w_055_2574, w_055_2575, w_055_2576, w_055_2577, w_055_2579, w_055_2580, w_055_2581, w_055_2582, w_055_2584, w_055_2587, w_055_2588, w_055_2591, w_055_2593, w_055_2594, w_055_2596, w_055_2597, w_055_2598, w_055_2599, w_055_2600, w_055_2601, w_055_2603, w_055_2604, w_055_2605, w_055_2606, w_055_2607, w_055_2609, w_055_2610, w_055_2611, w_055_2612, w_055_2613, w_055_2615, w_055_2616, w_055_2617, w_055_2619, w_055_2620, w_055_2621, w_055_2622, w_055_2624, w_055_2625, w_055_2626, w_055_2627, w_055_2629, w_055_2630, w_055_2631, w_055_2633, w_055_2634, w_055_2635, w_055_2636, w_055_2637, w_055_2638, w_055_2639, w_055_2640, w_055_2641, w_055_2645, w_055_2649, w_055_2653, w_055_2654, w_055_2656, w_055_2661, w_055_2662, w_055_2664, w_055_2667, w_055_2670, w_055_2671, w_055_2673, w_055_2674, w_055_2675, w_055_2677, w_055_2679, w_055_2681, w_055_2682, w_055_2683, w_055_2684, w_055_2689, w_055_2690, w_055_2691, w_055_2692, w_055_2693, w_055_2696, w_055_2697, w_055_2701, w_055_2702, w_055_2705, w_055_2707, w_055_2709, w_055_2710, w_055_2712, w_055_2714, w_055_2715, w_055_2716, w_055_2718, w_055_2719, w_055_2720, w_055_2721, w_055_2722, w_055_2724, w_055_2725, w_055_2726, w_055_2727, w_055_2733, w_055_2734, w_055_2735, w_055_2736, w_055_2737, w_055_2738, w_055_2739, w_055_2740, w_055_2741, w_055_2743, w_055_2744, w_055_2746, w_055_2747, w_055_2748, w_055_2750, w_055_2751, w_055_2753, w_055_2754, w_055_2756, w_055_2758, w_055_2759, w_055_2760, w_055_2762, w_055_2763, w_055_2765, w_055_2766, w_055_2767, w_055_2773, w_055_2774, w_055_2776, w_055_2778, w_055_2779, w_055_2781, w_055_2782, w_055_2784, w_055_2788, w_055_2790, w_055_2791, w_055_2792, w_055_2793, w_055_2795, w_055_2797, w_055_2800, w_055_2804, w_055_2805, w_055_2808, w_055_2811, w_055_2812, w_055_2813, w_055_2818, w_055_2820, w_055_2821, w_055_2822, w_055_2824, w_055_2826, w_055_2828, w_055_2831, w_055_2833, w_055_2834, w_055_2838, w_055_2840, w_055_2841, w_055_2842, w_055_2843, w_055_2848, w_055_2851, w_055_2852, w_055_2854, w_055_2855, w_055_2856, w_055_2857, w_055_2858, w_055_2860, w_055_2861, w_055_2862, w_055_2863, w_055_2865, w_055_2866, w_055_2867, w_055_2870, w_055_2875, w_055_2876, w_055_2878, w_055_2879, w_055_2880, w_055_2881, w_055_2884, w_055_2886, w_055_2887, w_055_2888, w_055_2890, w_055_2891, w_055_2893, w_055_2894, w_055_2896, w_055_2898, w_055_2899, w_055_2900, w_055_2902, w_055_2903, w_055_2906, w_055_2907, w_055_2908, w_055_2911, w_055_2912, w_055_2914, w_055_2915, w_055_2916, w_055_2917, w_055_2918, w_055_2919, w_055_2921, w_055_2922, w_055_2923, w_055_2924, w_055_2926, w_055_2927, w_055_2928, w_055_2929, w_055_2931, w_055_2933, w_055_2934, w_055_2937, w_055_2940, w_055_2941, w_055_2942, w_055_2945, w_055_2946, w_055_2947, w_055_2948, w_055_2950, w_055_2952, w_055_2953, w_055_2954, w_055_2955, w_055_2956, w_055_2958, w_055_2960, w_055_2961, w_055_2962, w_055_2963, w_055_2964, w_055_2966, w_055_2967, w_055_2968, w_055_2969, w_055_2970, w_055_2974, w_055_2975, w_055_2978, w_055_2979, w_055_2980, w_055_2981, w_055_2982, w_055_2984, w_055_2985, w_055_2989, w_055_2992, w_055_2995, w_055_2997, w_055_2999, w_055_3000, w_055_3003, w_055_3005, w_055_3007, w_055_3008, w_055_3010, w_055_3011, w_055_3012, w_055_3013, w_055_3014, w_055_3015, w_055_3016, w_055_3018, w_055_3019, w_055_3020, w_055_3022, w_055_3023, w_055_3024, w_055_3025, w_055_3026, w_055_3028, w_055_3029, w_055_3034, w_055_3037, w_055_3038, w_055_3041, w_055_3043, w_055_3044, w_055_3045, w_055_3046, w_055_3048, w_055_3050, w_055_3052, w_055_3053, w_055_3056, w_055_3058, w_055_3059, w_055_3061, w_055_3062, w_055_3063, w_055_3065, w_055_3067, w_055_3069, w_055_3074, w_055_3075, w_055_3076, w_055_3077, w_055_3078, w_055_3081, w_055_3084, w_055_3085, w_055_3087, w_055_3089, w_055_3090, w_055_3091, w_055_3092, w_055_3094, w_055_3098, w_055_3099, w_055_3100, w_055_3101, w_055_3102, w_055_3103, w_055_3104, w_055_3105, w_055_3106, w_055_3107, w_055_3109, w_055_3111, w_055_3112, w_055_3113, w_055_3115, w_055_3119, w_055_3121, w_055_3122, w_055_3124, w_055_3126, w_055_3128, w_055_3129, w_055_3131, w_055_3132, w_055_3133, w_055_3134, w_055_3135, w_055_3136, w_055_3138, w_055_3141, w_055_3142, w_055_3143, w_055_3144, w_055_3145, w_055_3150, w_055_3153, w_055_3154, w_055_3156, w_055_3157, w_055_3159, w_055_3161, w_055_3164, w_055_3168, w_055_3170, w_055_3171, w_055_3172, w_055_3173, w_055_3174, w_055_3175, w_055_3176, w_055_3177, w_055_3179, w_055_3183, w_055_3186, w_055_3188, w_055_3189, w_055_3190, w_055_3191, w_055_3194, w_055_3196, w_055_3198, w_055_3200, w_055_3204, w_055_3208, w_055_3209, w_055_3210, w_055_3213, w_055_3215, w_055_3216, w_055_3217, w_055_3218, w_055_3219, w_055_3220, w_055_3223, w_055_3224, w_055_3226, w_055_3227, w_055_3228, w_055_3229, w_055_3230, w_055_3231, w_055_3232, w_055_3233, w_055_3234, w_055_3235, w_055_3236, w_055_3238, w_055_3240, w_055_3241, w_055_3245, w_055_3246, w_055_3247, w_055_3248, w_055_3249, w_055_3250, w_055_3251, w_055_3252, w_055_3253, w_055_3254, w_055_3255, w_055_3257, w_055_3258, w_055_3259, w_055_3260, w_055_3261, w_055_3262, w_055_3265, w_055_3267, w_055_3268, w_055_3269, w_055_3270, w_055_3271, w_055_3272, w_055_3274, w_055_3275, w_055_3276, w_055_3277, w_055_3278, w_055_3279, w_055_3283, w_055_3284, w_055_3286, w_055_3289, w_055_3291, w_055_3292, w_055_3294, w_055_3297, w_055_3299, w_055_3300, w_055_3301, w_055_3302, w_055_3303, w_055_3306, w_055_3307, w_055_3308, w_055_3311, w_055_3313, w_055_3314, w_055_3315, w_055_3318, w_055_3319, w_055_3321, w_055_3323, w_055_3325, w_055_3328, w_055_3329, w_055_3330, w_055_3331, w_055_3332, w_055_3333, w_055_3334, w_055_3335, w_055_3336, w_055_3338, w_055_3339, w_055_3340, w_055_3341, w_055_3345, w_055_3347, w_055_3350, w_055_3351, w_055_3352, w_055_3353, w_055_3356, w_055_3357, w_055_3359, w_055_3360, w_055_3361, w_055_3363, w_055_3365, w_055_3368, w_055_3369, w_055_3370, w_055_3371, w_055_3373, w_055_3374, w_055_3375, w_055_3376, w_055_3377, w_055_3379, w_055_3381, w_055_3382, w_055_3383, w_055_3384, w_055_3386, w_055_3387, w_055_3388, w_055_3389, w_055_3390, w_055_3392, w_055_3393, w_055_3394, w_055_3395, w_055_3396, w_055_3398, w_055_3399, w_055_3400, w_055_3401, w_055_3403, w_055_3404, w_055_3409, w_055_3410, w_055_3411, w_055_3413, w_055_3414, w_055_3415, w_055_3416, w_055_3417, w_055_3419, w_055_3420, w_055_3421, w_055_3422, w_055_3423, w_055_3424, w_055_3425, w_055_3426, w_055_3427, w_055_3428, w_055_3429, w_055_3430, w_055_3431, w_055_3432, w_055_3439, w_055_3440, w_055_3442, w_055_3443, w_055_3444, w_055_3445, w_055_3447, w_055_3449, w_055_3450, w_055_3452, w_055_3453, w_055_3454, w_055_3459, w_055_3461, w_055_3466, w_055_3468, w_055_3471, w_055_3474, w_055_3476, w_055_3477, w_055_3479, w_055_3480, w_055_3481, w_055_3482, w_055_3483, w_055_3484, w_055_3485, w_055_3486, w_055_3488, w_055_3490, w_055_3491, w_055_3493, w_055_3494, w_055_3496, w_055_3498, w_055_3499, w_055_3502, w_055_3503, w_055_3504, w_055_3507, w_055_3510, w_055_3513, w_055_3514, w_055_3515, w_055_3516, w_055_3521, w_055_3522, w_055_3524, w_055_3526, w_055_3527, w_055_3528, w_055_3529, w_055_3531, w_055_3532, w_055_3533, w_055_3534, w_055_3535, w_055_3536, w_055_3537, w_055_3542, w_055_3543, w_055_3544, w_055_3546, w_055_3547, w_055_3551, w_055_3552, w_055_3553, w_055_3554, w_055_3555, w_055_3556, w_055_3557, w_055_3560, w_055_3562, w_055_3563, w_055_3564, w_055_3567, w_055_3568, w_055_3570, w_055_3573, w_055_3575, w_055_3576, w_055_3577, w_055_3579, w_055_3580, w_055_3581, w_055_3584, w_055_3585, w_055_3587, w_055_3588, w_055_3590, w_055_3591, w_055_3592, w_055_3593, w_055_3596, w_055_3597, w_055_3599, w_055_3601, w_055_3603, w_055_3604, w_055_3605, w_055_3606, w_055_3614, w_055_3616, w_055_3617, w_055_3618, w_055_3619, w_055_3620, w_055_3621, w_055_3622, w_055_3624, w_055_3625, w_055_3626, w_055_3627, w_055_3630, w_055_3631, w_055_3632, w_055_3633, w_055_3634, w_055_3635, w_055_3637, w_055_3641, w_055_3642, w_055_3644, w_055_3646, w_055_3649, w_055_3650, w_055_3651, w_055_3652, w_055_3654, w_055_3656, w_055_3657, w_055_3659, w_055_3660, w_055_3661, w_055_3662, w_055_3663, w_055_3665, w_055_3666, w_055_3667, w_055_3668, w_055_3669, w_055_3670, w_055_3671, w_055_3672, w_055_3674, w_055_3675, w_055_3676, w_055_3678, w_055_3679, w_055_3680, w_055_3684, w_055_3686, w_055_3687, w_055_3688, w_055_3692, w_055_3693, w_055_3694, w_055_3695, w_055_3697, w_055_3699, w_055_3701, w_055_3702, w_055_3703, w_055_3704, w_055_3705, w_055_3706, w_055_3708, w_055_3709, w_055_3710, w_055_3711, w_055_3712, w_055_3714, w_055_3716, w_055_3717, w_055_3718, w_055_3719, w_055_3720, w_055_3721, w_055_3722, w_055_3723, w_055_3725, w_055_3726, w_055_3727, w_055_3728, w_055_3730, w_055_3732, w_055_3735, w_055_3736, w_055_3739, w_055_3740, w_055_3742, w_055_3743, w_055_3744, w_055_3745, w_055_3749, w_055_3750, w_055_3751, w_055_3753, w_055_3754, w_055_3755, w_055_3756, w_055_3757, w_055_3758, w_055_3759, w_055_3760, w_055_3761, w_055_3763, w_055_3764, w_055_3766, w_055_3767, w_055_3769, w_055_3771, w_055_3773, w_055_3774, w_055_3775, w_055_3777, w_055_3778, w_055_3779, w_055_3780, w_055_3783, w_055_3785, w_055_3786, w_055_3787, w_055_3790, w_055_3793, w_055_3795, w_055_3798, w_055_3799, w_055_3800, w_055_3803, w_055_3805, w_055_3806, w_055_3807, w_055_3808, w_055_3809, w_055_3810, w_055_3811, w_055_3812, w_055_3813, w_055_3814, w_055_3815, w_055_3816, w_055_3817, w_055_3822, w_055_3823, w_055_3824, w_055_3825, w_055_3829, w_055_3830, w_055_3832, w_055_3833, w_055_3835, w_055_3836, w_055_3837, w_055_3838, w_055_3839, w_055_3840, w_055_3841, w_055_3842, w_055_3843, w_055_3845, w_055_3847, w_055_3848, w_055_3850, w_055_3851, w_055_3852, w_055_3853, w_055_3854, w_055_3855, w_055_3857, w_055_3859, w_055_3860, w_055_3862, w_055_3863, w_055_3865, w_055_3867, w_055_3869, w_055_3870, w_055_3873, w_055_3874, w_055_3875, w_055_3876, w_055_3877, w_055_3878, w_055_3879, w_055_3880, w_055_3881, w_055_3882, w_055_3886, w_055_3887, w_055_3889, w_055_3890, w_055_3893, w_055_3895, w_055_3896, w_055_3898, w_055_3899, w_055_3901, w_055_3902, w_055_3903, w_055_3905, w_055_3908, w_055_3909, w_055_3910, w_055_3911, w_055_3913, w_055_3914, w_055_3915, w_055_3916, w_055_3918, w_055_3920, w_055_3922, w_055_3923, w_055_3924, w_055_3925, w_055_3926, w_055_3927, w_055_3928, w_055_3929, w_055_3930, w_055_3932, w_055_3933, w_055_3934, w_055_3935, w_055_3937, w_055_3938, w_055_3941, w_055_3945, w_055_3947, w_055_3948, w_055_3952, w_055_3953, w_055_3955, w_055_3957, w_055_3958, w_055_3960, w_055_3961, w_055_3962, w_055_3963, w_055_3964, w_055_3965, w_055_3966, w_055_3967, w_055_3969, w_055_3970, w_055_3971, w_055_3972, w_055_3973, w_055_3974, w_055_3975, w_055_3976, w_055_3977, w_055_3978, w_055_3981, w_055_3982, w_055_3983, w_055_3985, w_055_3986, w_055_3987, w_055_3988, w_055_3989, w_055_3990, w_055_3992, w_055_3993, w_055_3994, w_055_3995, w_055_3996, w_055_3998, w_055_4000, w_055_4001, w_055_4002, w_055_4006, w_055_4008, w_055_4010, w_055_4011, w_055_4012, w_055_4013, w_055_4016, w_055_4017, w_055_4018, w_055_4019, w_055_4020, w_055_4023, w_055_4025, w_055_4026, w_055_4027, w_055_4028, w_055_4029, w_055_4030, w_055_4031, w_055_4032, w_055_4034, w_055_4035, w_055_4036, w_055_4037, w_055_4039, w_055_4040, w_055_4043, w_055_4046, w_055_4049, w_055_4050, w_055_4052, w_055_4055, w_055_4056, w_055_4057, w_055_4058, w_055_4059, w_055_4060, w_055_4064, w_055_4065, w_055_4067, w_055_4068, w_055_4069, w_055_4071, w_055_4072, w_055_4073, w_055_4074, w_055_4075, w_055_4076, w_055_4077, w_055_4078, w_055_4079, w_055_4080, w_055_4081, w_055_4083, w_055_4085, w_055_4087, w_055_4089, w_055_4091, w_055_4092, w_055_4094, w_055_4095, w_055_4096, w_055_4097, w_055_4098, w_055_4099, w_055_4100, w_055_4101, w_055_4103, w_055_4104, w_055_4105, w_055_4106, w_055_4107, w_055_4110, w_055_4111, w_055_4112, w_055_4113, w_055_4114, w_055_4115, w_055_4116, w_055_4118, w_055_4119, w_055_4120, w_055_4122, w_055_4123, w_055_4124, w_055_4125, w_055_4126, w_055_4127, w_055_4128, w_055_4130, w_055_4131, w_055_4132, w_055_4133, w_055_4134, w_055_4135, w_055_4136, w_055_4137, w_055_4138, w_055_4139, w_055_4140, w_055_4142, w_055_4144, w_055_4146, w_055_4147, w_055_4148, w_055_4151, w_055_4152, w_055_4154, w_055_4156, w_055_4160, w_055_4161, w_055_4162, w_055_4165, w_055_4168, w_055_4169, w_055_4170, w_055_4171, w_055_4173, w_055_4174, w_055_4175, w_055_4176, w_055_4178, w_055_4179, w_055_4181, w_055_4182, w_055_4183, w_055_4184, w_055_4185, w_055_4186, w_055_4188, w_055_4190, w_055_4193, w_055_4194, w_055_4196, w_055_4200, w_055_4201, w_055_4202, w_055_4203, w_055_4204, w_055_4205, w_055_4206, w_055_4207, w_055_4209, w_055_4210, w_055_4212, w_055_4214, w_055_4217, w_055_4218, w_055_4219, w_055_4221, w_055_4222, w_055_4224, w_055_4227, w_055_4229, w_055_4230, w_055_4231, w_055_4232, w_055_4233, w_055_4237, w_055_4238, w_055_4239, w_055_4240, w_055_4241, w_055_4242, w_055_4243, w_055_4244, w_055_4245, w_055_4246, w_055_4248, w_055_4249, w_055_4250, w_055_4255, w_055_4256, w_055_4257, w_055_4258, w_055_4259, w_055_4260, w_055_4261, w_055_4262, w_055_4264, w_055_4267, w_055_4268, w_055_4269, w_055_4270, w_055_4272, w_055_4273, w_055_4276, w_055_4277, w_055_4278, w_055_4280, w_055_4281, w_055_4283, w_055_4286, w_055_4287, w_055_4293, w_055_4295, w_055_4297, w_055_4298, w_055_4300, w_055_4302, w_055_4304, w_055_4305, w_055_4307, w_055_4308, w_055_4309, w_055_4310, w_055_4313, w_055_4315, w_055_4317, w_055_4318, w_055_4320, w_055_4322, w_055_4323, w_055_4327, w_055_4328, w_055_4330, w_055_4332, w_055_4333, w_055_4335, w_055_4336, w_055_4337, w_055_4338, w_055_4340, w_055_4341, w_055_4342, w_055_4344, w_055_4345, w_055_4346, w_055_4348, w_055_4349, w_055_4351, w_055_4355, w_055_4356, w_055_4357, w_055_4358, w_055_4359, w_055_4360, w_055_4361, w_055_4362, w_055_4363, w_055_4364, w_055_4365, w_055_4366, w_055_4367, w_055_4369, w_055_4372, w_055_4373, w_055_4374, w_055_4375, w_055_4376, w_055_4378, w_055_4380, w_055_4383, w_055_4385, w_055_4386, w_055_4387, w_055_4393, w_055_4394, w_055_4396, w_055_4397, w_055_4401, w_055_4403, w_055_4404, w_055_4405, w_055_4406, w_055_4407, w_055_4408, w_055_4409, w_055_4411, w_055_4412, w_055_4414, w_055_4416, w_055_4418, w_055_4419, w_055_4421, w_055_4422, w_055_4423, w_055_4424, w_055_4426, w_055_4427, w_055_4428, w_055_4431, w_055_4436, w_055_4438, w_055_4441, w_055_4443, w_055_4444, w_055_4445, w_055_4449, w_055_4450, w_055_4452, w_055_4454, w_055_4455, w_055_4457, w_055_4460, w_055_4461, w_055_4462, w_055_4463, w_055_4466, w_055_4467, w_055_4471, w_055_4473, w_055_4474, w_055_4475, w_055_4476, w_055_4478, w_055_4479, w_055_4480, w_055_4483, w_055_4484, w_055_4485, w_055_4486, w_055_4487, w_055_4488, w_055_4489, w_055_4490, w_055_4491, w_055_4492, w_055_4493, w_055_4494, w_055_4495, w_055_4496, w_055_4497, w_055_4499, w_055_4500, w_055_4501, w_055_4502, w_055_4503, w_055_4504, w_055_4506, w_055_4508, w_055_4510, w_055_4511, w_055_4513, w_055_4515, w_055_4516, w_055_4518, w_055_4521, w_055_4522, w_055_4523, w_055_4524, w_055_4525, w_055_4526, w_055_4527, w_055_4528, w_055_4531, w_055_4533, w_055_4534, w_055_4538, w_055_4540, w_055_4541, w_055_4543, w_055_4545, w_055_4546, w_055_4548, w_055_4553, w_055_4555, w_055_4556, w_055_4557, w_055_4559, w_055_4560, w_055_4561, w_055_4562, w_055_4564, w_055_4569, w_055_4571, w_055_4572, w_055_4573, w_055_4575, w_055_4577, w_055_4578, w_055_4579, w_055_4581, w_055_4582, w_055_4585, w_055_4586, w_055_4587, w_055_4588, w_055_4589, w_055_4590, w_055_4591, w_055_4592, w_055_4595, w_055_4600, w_055_4605, w_055_4606, w_055_4607, w_055_4608, w_055_4609, w_055_4610, w_055_4611, w_055_4612, w_055_4613, w_055_4615, w_055_4617, w_055_4619, w_055_4620, w_055_4621, w_055_4623, w_055_4624, w_055_4625, w_055_4626, w_055_4627, w_055_4632, w_055_4633, w_055_4636, w_055_4637, w_055_4638, w_055_4639, w_055_4640, w_055_4641, w_055_4642, w_055_4643, w_055_4644, w_055_4647, w_055_4648, w_055_4650, w_055_4651, w_055_4652, w_055_4653, w_055_4654, w_055_4656, w_055_4657, w_055_4659, w_055_4660, w_055_4663, w_055_4666, w_055_4669, w_055_4670, w_055_4673, w_055_4676, w_055_4680, w_055_4682, w_055_4684, w_055_4686, w_055_4687, w_055_4690, w_055_4692, w_055_4693, w_055_4694, w_055_4696, w_055_4697, w_055_4699, w_055_4700, w_055_4701, w_055_4702, w_055_4703, w_055_4707, w_055_4709, w_055_4710, w_055_4711, w_055_4712, w_055_4713, w_055_4714, w_055_4715, w_055_4716, w_055_4718, w_055_4720, w_055_4721, w_055_4722, w_055_4725, w_055_4726, w_055_4727, w_055_4729, w_055_4737, w_055_4738, w_055_4739, w_055_4740, w_055_4741, w_055_4742, w_055_4743, w_055_4744, w_055_4745, w_055_4747, w_055_4748, w_055_4749, w_055_4750, w_055_4751, w_055_4753, w_055_4755, w_055_4756, w_055_4757, w_055_4759, w_055_4760, w_055_4765, w_055_4766, w_055_4771, w_055_4772, w_055_4773, w_055_4776, w_055_4779, w_055_4781, w_055_4782, w_055_4792, w_055_4794, w_055_4795, w_055_4796, w_055_4797, w_055_4798, w_055_4800, w_055_4801, w_055_4803, w_055_4806, w_055_4809, w_055_4813, w_055_4821, w_055_4822, w_055_4825, w_055_4828, w_055_4832, w_055_4833, w_055_4834, w_055_4835, w_055_4840, w_055_4843, w_055_4847, w_055_4849, w_055_4850, w_055_4851, w_055_4852, w_055_4853, w_055_4859, w_055_4860, w_055_4861, w_055_4865, w_055_4868, w_055_4872, w_055_4874, w_055_4875, w_055_4876, w_055_4880, w_055_4882, w_055_4885, w_055_4889, w_055_4893, w_055_4896, w_055_4897, w_055_4899, w_055_4900, w_055_4904, w_055_4905, w_055_4914, w_055_4917, w_055_4923, w_055_4924, w_055_4926, w_055_4927, w_055_4928, w_055_4930, w_055_4933, w_055_4934, w_055_4939, w_055_4941, w_055_4944, w_055_4947, w_055_4948, w_055_4949, w_055_4956, w_055_4958, w_055_4965, w_055_4968, w_055_4969, w_055_4973, w_055_4975, w_055_4986, w_055_4987, w_055_4989, w_055_4990, w_055_4994, w_055_4997, w_055_5000, w_055_5001, w_055_5002, w_055_5004, w_055_5005, w_055_5007, w_055_5010, w_055_5013, w_055_5015, w_055_5016, w_055_5017, w_055_5018, w_055_5019, w_055_5020, w_055_5021, w_055_5023, w_055_5028, w_055_5030, w_055_5031, w_055_5033, w_055_5037, w_055_5039, w_055_5042, w_055_5043, w_055_5047, w_055_5051, w_055_5054, w_055_5059, w_055_5063, w_055_5066, w_055_5068, w_055_5069, w_055_5076, w_055_5078, w_055_5080, w_055_5084, w_055_5087, w_055_5088, w_055_5097, w_055_5099, w_055_5100, w_055_5106, w_055_5107, w_055_5112, w_055_5113, w_055_5114, w_055_5116, w_055_5118, w_055_5123, w_055_5125, w_055_5126, w_055_5128, w_055_5129, w_055_5131, w_055_5135, w_055_5136, w_055_5140, w_055_5142, w_055_5146, w_055_5148, w_055_5149, w_055_5156, w_055_5169, w_055_5172, w_055_5178, w_055_5180, w_055_5181, w_055_5182, w_055_5184, w_055_5185, w_055_5189, w_055_5190, w_055_5191, w_055_5192, w_055_5194, w_055_5195, w_055_5197, w_055_5202, w_055_5206, w_055_5208, w_055_5209, w_055_5211, w_055_5212, w_055_5213, w_055_5214, w_055_5215, w_055_5218, w_055_5219, w_055_5220, w_055_5221, w_055_5222, w_055_5227, w_055_5228, w_055_5229, w_055_5231;
  wire w_056_000, w_056_001, w_056_003, w_056_004, w_056_005, w_056_007, w_056_008, w_056_009, w_056_010, w_056_012, w_056_013, w_056_014, w_056_015, w_056_016, w_056_017, w_056_018, w_056_019, w_056_020, w_056_021, w_056_022, w_056_023, w_056_024, w_056_025, w_056_026, w_056_027, w_056_028, w_056_029, w_056_030, w_056_031, w_056_032, w_056_033, w_056_034, w_056_035, w_056_036, w_056_037, w_056_038, w_056_039, w_056_040, w_056_041, w_056_042, w_056_043, w_056_044, w_056_045, w_056_046, w_056_047, w_056_048, w_056_049, w_056_050, w_056_051, w_056_052, w_056_053, w_056_054, w_056_055, w_056_057, w_056_058, w_056_059, w_056_060, w_056_061, w_056_062, w_056_063, w_056_064, w_056_065, w_056_066, w_056_067, w_056_068, w_056_069, w_056_070, w_056_071, w_056_072, w_056_073, w_056_074, w_056_075, w_056_078, w_056_079, w_056_080, w_056_081, w_056_082, w_056_083, w_056_085, w_056_086, w_056_087, w_056_088, w_056_089, w_056_090, w_056_091, w_056_092, w_056_093, w_056_094, w_056_096, w_056_097, w_056_099, w_056_100, w_056_101, w_056_103, w_056_104, w_056_105, w_056_106, w_056_109, w_056_110, w_056_111, w_056_112, w_056_114, w_056_115, w_056_116, w_056_117, w_056_118, w_056_119, w_056_120, w_056_121, w_056_122, w_056_124, w_056_125, w_056_126, w_056_127, w_056_128, w_056_129, w_056_130, w_056_131, w_056_132, w_056_133, w_056_134, w_056_135, w_056_136, w_056_137, w_056_138, w_056_141, w_056_143, w_056_144, w_056_145, w_056_146, w_056_147, w_056_148, w_056_149, w_056_150, w_056_151, w_056_153, w_056_154, w_056_155, w_056_156, w_056_157, w_056_158, w_056_159, w_056_160, w_056_161, w_056_162, w_056_163, w_056_164, w_056_165, w_056_166, w_056_168, w_056_169, w_056_170, w_056_171, w_056_173, w_056_175, w_056_176, w_056_177, w_056_178, w_056_179, w_056_180, w_056_181, w_056_182, w_056_183, w_056_184, w_056_185, w_056_186, w_056_187, w_056_188, w_056_189, w_056_190, w_056_191, w_056_192, w_056_193, w_056_194, w_056_195, w_056_196, w_056_197, w_056_198, w_056_199, w_056_200, w_056_201, w_056_202, w_056_203, w_056_204, w_056_205, w_056_206, w_056_207, w_056_208, w_056_209, w_056_210, w_056_211, w_056_212, w_056_213, w_056_214, w_056_215, w_056_216, w_056_217, w_056_219, w_056_220, w_056_221, w_056_222, w_056_223, w_056_224, w_056_226, w_056_227, w_056_228, w_056_229, w_056_230, w_056_231, w_056_232, w_056_233, w_056_234, w_056_235, w_056_236, w_056_237, w_056_238, w_056_239, w_056_240, w_056_241, w_056_242, w_056_243, w_056_244, w_056_245, w_056_246, w_056_248, w_056_249, w_056_250, w_056_251, w_056_252, w_056_253, w_056_254, w_056_255, w_056_256, w_056_257, w_056_258, w_056_259, w_056_260, w_056_261, w_056_263, w_056_264, w_056_265, w_056_266, w_056_267, w_056_268, w_056_269, w_056_270, w_056_271, w_056_272, w_056_273, w_056_275, w_056_276, w_056_277, w_056_278, w_056_279, w_056_280, w_056_281, w_056_282, w_056_283, w_056_284, w_056_285, w_056_286, w_056_287, w_056_288, w_056_289, w_056_290, w_056_291, w_056_292, w_056_293, w_056_294, w_056_295, w_056_296, w_056_297, w_056_298, w_056_299, w_056_300, w_056_301, w_056_302, w_056_303, w_056_304, w_056_305, w_056_306, w_056_307, w_056_308, w_056_309, w_056_310, w_056_311, w_056_312, w_056_314, w_056_315, w_056_316, w_056_317, w_056_318, w_056_319, w_056_320, w_056_322, w_056_323, w_056_324, w_056_325, w_056_326, w_056_327, w_056_328, w_056_329, w_056_330, w_056_331, w_056_332, w_056_334, w_056_335, w_056_336, w_056_338, w_056_339, w_056_340, w_056_341, w_056_342, w_056_343, w_056_345, w_056_346, w_056_347, w_056_349, w_056_350, w_056_351, w_056_352, w_056_353, w_056_354, w_056_355, w_056_356, w_056_357, w_056_358, w_056_359, w_056_362, w_056_363, w_056_365, w_056_366, w_056_367, w_056_368, w_056_370, w_056_371, w_056_372, w_056_373, w_056_374, w_056_377, w_056_378, w_056_379, w_056_380, w_056_381, w_056_383, w_056_384, w_056_385, w_056_386, w_056_387, w_056_388, w_056_390, w_056_391, w_056_392, w_056_393, w_056_394, w_056_395, w_056_396, w_056_397, w_056_398, w_056_399, w_056_400, w_056_401, w_056_402, w_056_403, w_056_405, w_056_406, w_056_407, w_056_410, w_056_411, w_056_412, w_056_413, w_056_414, w_056_415, w_056_416, w_056_417, w_056_418, w_056_419, w_056_420, w_056_421, w_056_422, w_056_423, w_056_424, w_056_425, w_056_426, w_056_427, w_056_430, w_056_431, w_056_432, w_056_433, w_056_434, w_056_435, w_056_436, w_056_437, w_056_438, w_056_439, w_056_440, w_056_441, w_056_442, w_056_443, w_056_444, w_056_445, w_056_446, w_056_447, w_056_448, w_056_449, w_056_450, w_056_451, w_056_452, w_056_453, w_056_454, w_056_455, w_056_456, w_056_457, w_056_458, w_056_459, w_056_460, w_056_461, w_056_462, w_056_463, w_056_464, w_056_465, w_056_466, w_056_467, w_056_468, w_056_469, w_056_470, w_056_471, w_056_472, w_056_473, w_056_474, w_056_475, w_056_476, w_056_477, w_056_478, w_056_479, w_056_480, w_056_481, w_056_483, w_056_484, w_056_485, w_056_486, w_056_487, w_056_488, w_056_489, w_056_490, w_056_491, w_056_492, w_056_493, w_056_494, w_056_495, w_056_496, w_056_497, w_056_498, w_056_499, w_056_500, w_056_501, w_056_502, w_056_503, w_056_504, w_056_505, w_056_506, w_056_507, w_056_508, w_056_509, w_056_510, w_056_511, w_056_512, w_056_513, w_056_514, w_056_516, w_056_517, w_056_518, w_056_519, w_056_520, w_056_521, w_056_522, w_056_523, w_056_524, w_056_525, w_056_526, w_056_527, w_056_528, w_056_530, w_056_531, w_056_532, w_056_533, w_056_534, w_056_535, w_056_536, w_056_538, w_056_539, w_056_540, w_056_541, w_056_542, w_056_543, w_056_545, w_056_547, w_056_548, w_056_549, w_056_550, w_056_551, w_056_552, w_056_553, w_056_555, w_056_556, w_056_557, w_056_558, w_056_559, w_056_560, w_056_561, w_056_562, w_056_563, w_056_564, w_056_565, w_056_566, w_056_567, w_056_569, w_056_570, w_056_571, w_056_572, w_056_573, w_056_574, w_056_575, w_056_576, w_056_579, w_056_580, w_056_581, w_056_582, w_056_583, w_056_584, w_056_585, w_056_586, w_056_587, w_056_588, w_056_589, w_056_590, w_056_591, w_056_592, w_056_593, w_056_594, w_056_595, w_056_596, w_056_597, w_056_598, w_056_600, w_056_601, w_056_602, w_056_603, w_056_604, w_056_605, w_056_606, w_056_607, w_056_608, w_056_609, w_056_610, w_056_611, w_056_612, w_056_613, w_056_614, w_056_615, w_056_616, w_056_617, w_056_618, w_056_619, w_056_620, w_056_621, w_056_622, w_056_623, w_056_624, w_056_625, w_056_628, w_056_629, w_056_630, w_056_631, w_056_632, w_056_633, w_056_634, w_056_635, w_056_636, w_056_637, w_056_638, w_056_639, w_056_640, w_056_641, w_056_642, w_056_644, w_056_645, w_056_646, w_056_647, w_056_648, w_056_649, w_056_650, w_056_651, w_056_652, w_056_653, w_056_654, w_056_655, w_056_656, w_056_657, w_056_659, w_056_661, w_056_662, w_056_663, w_056_666, w_056_667, w_056_668, w_056_669, w_056_670, w_056_671, w_056_672, w_056_673, w_056_677, w_056_678, w_056_679, w_056_680, w_056_681, w_056_682, w_056_684, w_056_685, w_056_686, w_056_687, w_056_688, w_056_689, w_056_690, w_056_692, w_056_693, w_056_694, w_056_696, w_056_697, w_056_698, w_056_699, w_056_700, w_056_701, w_056_703, w_056_704, w_056_705, w_056_706, w_056_707, w_056_709, w_056_711, w_056_712, w_056_713, w_056_714, w_056_715, w_056_716, w_056_717, w_056_719, w_056_720, w_056_721, w_056_722, w_056_723, w_056_724, w_056_725, w_056_726, w_056_727, w_056_728, w_056_729, w_056_730, w_056_731, w_056_732, w_056_733, w_056_735, w_056_736, w_056_737, w_056_740, w_056_741, w_056_742, w_056_743, w_056_744, w_056_745, w_056_746, w_056_747, w_056_748, w_056_749, w_056_750, w_056_751, w_056_752, w_056_753, w_056_754, w_056_755, w_056_757, w_056_758, w_056_760, w_056_761, w_056_762, w_056_763, w_056_765, w_056_767, w_056_769, w_056_770, w_056_771, w_056_772, w_056_773, w_056_774, w_056_775, w_056_776, w_056_777, w_056_778, w_056_779, w_056_780, w_056_781, w_056_784, w_056_785, w_056_786, w_056_787, w_056_788, w_056_791, w_056_792, w_056_793, w_056_794, w_056_796, w_056_797, w_056_798, w_056_799, w_056_800, w_056_802, w_056_804, w_056_805, w_056_806, w_056_807, w_056_809, w_056_810, w_056_811, w_056_812, w_056_813, w_056_814, w_056_815, w_056_816, w_056_817, w_056_818, w_056_819, w_056_820, w_056_821, w_056_822, w_056_824, w_056_825, w_056_826, w_056_827, w_056_830, w_056_831, w_056_834, w_056_835, w_056_836, w_056_837, w_056_838, w_056_839, w_056_840, w_056_841, w_056_842, w_056_843, w_056_844, w_056_845, w_056_846, w_056_847, w_056_848, w_056_849, w_056_850, w_056_851, w_056_853, w_056_854, w_056_855, w_056_856, w_056_857, w_056_858, w_056_859, w_056_860, w_056_861, w_056_862, w_056_863, w_056_864, w_056_865, w_056_866, w_056_867, w_056_868, w_056_869, w_056_870, w_056_871, w_056_872, w_056_873, w_056_874, w_056_875, w_056_877, w_056_878, w_056_880, w_056_881, w_056_882, w_056_883, w_056_884, w_056_885, w_056_886, w_056_888, w_056_891, w_056_892, w_056_893, w_056_895, w_056_897, w_056_898, w_056_899, w_056_900, w_056_901, w_056_902, w_056_903, w_056_905, w_056_906, w_056_907, w_056_911, w_056_912, w_056_914, w_056_915, w_056_916, w_056_917, w_056_918, w_056_920, w_056_921, w_056_922, w_056_923, w_056_925, w_056_926, w_056_927, w_056_928, w_056_929, w_056_930, w_056_931, w_056_932, w_056_933, w_056_934, w_056_935, w_056_936, w_056_937, w_056_938, w_056_939, w_056_940, w_056_941, w_056_942, w_056_943, w_056_944, w_056_946, w_056_947, w_056_948, w_056_949, w_056_950, w_056_952, w_056_953, w_056_954, w_056_955, w_056_956, w_056_957, w_056_958, w_056_959, w_056_960, w_056_962, w_056_963, w_056_964, w_056_965, w_056_967, w_056_968, w_056_969, w_056_970, w_056_971, w_056_972, w_056_973, w_056_975, w_056_976, w_056_977, w_056_978, w_056_979, w_056_980, w_056_982, w_056_983, w_056_985, w_056_986, w_056_987, w_056_988, w_056_989, w_056_990, w_056_991, w_056_992, w_056_993, w_056_994, w_056_995, w_056_996, w_056_997, w_056_998, w_056_1000, w_056_1002, w_056_1003, w_056_1004, w_056_1005, w_056_1006, w_056_1008, w_056_1009, w_056_1010, w_056_1011, w_056_1012, w_056_1013, w_056_1014, w_056_1015, w_056_1016, w_056_1017, w_056_1018, w_056_1019, w_056_1020, w_056_1021, w_056_1022, w_056_1023, w_056_1025, w_056_1026, w_056_1027, w_056_1028, w_056_1030, w_056_1033, w_056_1034, w_056_1035, w_056_1037, w_056_1038, w_056_1039, w_056_1040, w_056_1041, w_056_1042, w_056_1043, w_056_1044, w_056_1045, w_056_1046, w_056_1047, w_056_1048, w_056_1049, w_056_1050, w_056_1051, w_056_1052, w_056_1053, w_056_1055, w_056_1056, w_056_1057, w_056_1058, w_056_1059, w_056_1060, w_056_1061, w_056_1062, w_056_1063, w_056_1064, w_056_1065, w_056_1066, w_056_1067, w_056_1068, w_056_1069, w_056_1070, w_056_1071, w_056_1072, w_056_1073, w_056_1074, w_056_1075, w_056_1078, w_056_1079, w_056_1080, w_056_1081, w_056_1082, w_056_1083, w_056_1084, w_056_1085, w_056_1086, w_056_1087, w_056_1088, w_056_1089, w_056_1090, w_056_1091, w_056_1093, w_056_1094, w_056_1095, w_056_1096, w_056_1097, w_056_1098, w_056_1099, w_056_1100, w_056_1101, w_056_1102, w_056_1103, w_056_1104, w_056_1105, w_056_1106, w_056_1107, w_056_1108, w_056_1109, w_056_1110, w_056_1111, w_056_1112, w_056_1113, w_056_1114, w_056_1115, w_056_1116, w_056_1117, w_056_1118, w_056_1119, w_056_1120, w_056_1121, w_056_1122, w_056_1123, w_056_1124, w_056_1127, w_056_1128, w_056_1129, w_056_1130, w_056_1131, w_056_1132, w_056_1133, w_056_1134, w_056_1135, w_056_1136, w_056_1137, w_056_1138, w_056_1139, w_056_1140, w_056_1141, w_056_1142, w_056_1143, w_056_1145, w_056_1146, w_056_1147, w_056_1148, w_056_1150, w_056_1151, w_056_1152, w_056_1153, w_056_1154, w_056_1156, w_056_1157, w_056_1158, w_056_1159, w_056_1160, w_056_1161, w_056_1163, w_056_1164, w_056_1165, w_056_1166, w_056_1167, w_056_1168, w_056_1169, w_056_1170, w_056_1171, w_056_1172, w_056_1174, w_056_1175, w_056_1176, w_056_1178, w_056_1179, w_056_1180, w_056_1182, w_056_1183, w_056_1185, w_056_1187, w_056_1188, w_056_1189, w_056_1190, w_056_1191, w_056_1192, w_056_1193, w_056_1194, w_056_1195, w_056_1196, w_056_1197, w_056_1198, w_056_1199, w_056_1200, w_056_1201, w_056_1202, w_056_1203, w_056_1204, w_056_1205, w_056_1206, w_056_1207, w_056_1208, w_056_1209, w_056_1211, w_056_1212, w_056_1214, w_056_1216, w_056_1217, w_056_1219, w_056_1220, w_056_1221, w_056_1223, w_056_1224, w_056_1225, w_056_1226, w_056_1228, w_056_1229, w_056_1231, w_056_1232, w_056_1233, w_056_1234, w_056_1235, w_056_1236, w_056_1237, w_056_1238, w_056_1239, w_056_1240, w_056_1241, w_056_1243, w_056_1244, w_056_1245, w_056_1247, w_056_1248, w_056_1249, w_056_1250, w_056_1251, w_056_1252, w_056_1253, w_056_1254, w_056_1255, w_056_1256, w_056_1257, w_056_1258, w_056_1259, w_056_1261, w_056_1262, w_056_1263, w_056_1264, w_056_1265, w_056_1266, w_056_1267, w_056_1268, w_056_1269, w_056_1270, w_056_1271, w_056_1273, w_056_1274, w_056_1275, w_056_1276, w_056_1277, w_056_1278, w_056_1279, w_056_1281, w_056_1282, w_056_1284, w_056_1287, w_056_1289, w_056_1290, w_056_1294, w_056_1297, w_056_1298, w_056_1299, w_056_1300, w_056_1301, w_056_1302, w_056_1304, w_056_1305, w_056_1306, w_056_1307, w_056_1309, w_056_1310, w_056_1311, w_056_1312, w_056_1313, w_056_1315, w_056_1317, w_056_1318, w_056_1319, w_056_1320, w_056_1321, w_056_1322, w_056_1323, w_056_1324, w_056_1326, w_056_1327, w_056_1328, w_056_1329, w_056_1332, w_056_1333, w_056_1334, w_056_1335, w_056_1336, w_056_1337, w_056_1338, w_056_1339, w_056_1340, w_056_1342, w_056_1343, w_056_1345, w_056_1346, w_056_1348, w_056_1349, w_056_1350, w_056_1351, w_056_1353, w_056_1354, w_056_1355, w_056_1356, w_056_1358, w_056_1359, w_056_1360, w_056_1361, w_056_1362, w_056_1364, w_056_1366, w_056_1367, w_056_1368, w_056_1369, w_056_1370, w_056_1371, w_056_1372, w_056_1373, w_056_1374, w_056_1375, w_056_1376, w_056_1377, w_056_1378, w_056_1380, w_056_1382, w_056_1383, w_056_1384, w_056_1385, w_056_1386, w_056_1387, w_056_1388, w_056_1389, w_056_1390, w_056_1391, w_056_1392, w_056_1395, w_056_1396, w_056_1398, w_056_1399, w_056_1400, w_056_1401, w_056_1402, w_056_1403, w_056_1404, w_056_1405, w_056_1406, w_056_1407, w_056_1408, w_056_1409, w_056_1410, w_056_1411, w_056_1412, w_056_1413, w_056_1414, w_056_1415, w_056_1416, w_056_1417, w_056_1418, w_056_1419, w_056_1420, w_056_1422, w_056_1423, w_056_1424, w_056_1425, w_056_1426, w_056_1427, w_056_1429, w_056_1430, w_056_1431, w_056_1432, w_056_1433, w_056_1435, w_056_1436, w_056_1437, w_056_1438, w_056_1439, w_056_1442, w_056_1443, w_056_1444, w_056_1446, w_056_1447, w_056_1448, w_056_1449, w_056_1450, w_056_1451, w_056_1453, w_056_1456, w_056_1458, w_056_1459, w_056_1460, w_056_1461, w_056_1462, w_056_1463, w_056_1464, w_056_1465, w_056_1467, w_056_1468, w_056_1469, w_056_1470, w_056_1471, w_056_1472, w_056_1473, w_056_1474, w_056_1475, w_056_1476, w_056_1477, w_056_1478, w_056_1479, w_056_1480, w_056_1481, w_056_1482, w_056_1483, w_056_1484, w_056_1485, w_056_1486, w_056_1487, w_056_1488, w_056_1489, w_056_1490, w_056_1491, w_056_1493, w_056_1494, w_056_1495, w_056_1496, w_056_1497, w_056_1499, w_056_1500, w_056_1502, w_056_1503, w_056_1504, w_056_1505, w_056_1507, w_056_1508, w_056_1509, w_056_1510, w_056_1514, w_056_1516, w_056_1519, w_056_1520, w_056_1521, w_056_1524, w_056_1525, w_056_1526, w_056_1527, w_056_1529, w_056_1530, w_056_1531, w_056_1533, w_056_1534, w_056_1535, w_056_1536, w_056_1537, w_056_1538, w_056_1539, w_056_1542, w_056_1543, w_056_1544, w_056_1545, w_056_1546, w_056_1547, w_056_1548, w_056_1549, w_056_1550, w_056_1552, w_056_1553, w_056_1555, w_056_1556, w_056_1557, w_056_1559, w_056_1560, w_056_1561, w_056_1562, w_056_1563, w_056_1564, w_056_1566, w_056_1567, w_056_1568, w_056_1569, w_056_1570, w_056_1573, w_056_1574, w_056_1575, w_056_1576, w_056_1577, w_056_1578, w_056_1579, w_056_1582, w_056_1583, w_056_1584, w_056_1585, w_056_1586, w_056_1587, w_056_1588, w_056_1589, w_056_1590, w_056_1591, w_056_1594, w_056_1595, w_056_1596, w_056_1597, w_056_1598, w_056_1599, w_056_1601, w_056_1603, w_056_1604, w_056_1605, w_056_1606, w_056_1607, w_056_1608, w_056_1609, w_056_1610, w_056_1611, w_056_1612, w_056_1613, w_056_1614, w_056_1616, w_056_1617, w_056_1618, w_056_1619, w_056_1620, w_056_1621, w_056_1622, w_056_1623, w_056_1624, w_056_1625, w_056_1627, w_056_1628, w_056_1630, w_056_1632, w_056_1633, w_056_1634, w_056_1635, w_056_1636, w_056_1637, w_056_1638, w_056_1639, w_056_1640, w_056_1641, w_056_1642, w_056_1643, w_056_1644, w_056_1645, w_056_1646, w_056_1647, w_056_1648, w_056_1649, w_056_1650, w_056_1651, w_056_1652, w_056_1653, w_056_1654, w_056_1655, w_056_1656, w_056_1657, w_056_1659, w_056_1660, w_056_1661, w_056_1662, w_056_1663, w_056_1665, w_056_1666, w_056_1669, w_056_1670, w_056_1672, w_056_1673, w_056_1674, w_056_1675, w_056_1677, w_056_1678, w_056_1679, w_056_1680, w_056_1681, w_056_1682, w_056_1683, w_056_1686, w_056_1687, w_056_1690, w_056_1691, w_056_1692, w_056_1693, w_056_1694, w_056_1695, w_056_1696, w_056_1697, w_056_1698, w_056_1699, w_056_1700, w_056_1701, w_056_1702, w_056_1703, w_056_1704, w_056_1705, w_056_1706, w_056_1707, w_056_1708, w_056_1710, w_056_1711, w_056_1712, w_056_1713, w_056_1714, w_056_1716, w_056_1717, w_056_1719, w_056_1720, w_056_1721, w_056_1722, w_056_1723, w_056_1724, w_056_1725, w_056_1728, w_056_1729, w_056_1730, w_056_1731, w_056_1732, w_056_1733, w_056_1734, w_056_1735, w_056_1736, w_056_1737, w_056_1738, w_056_1739, w_056_1740, w_056_1741, w_056_1742, w_056_1743, w_056_1744, w_056_1746, w_056_1747, w_056_1748, w_056_1749, w_056_1750, w_056_1751, w_056_1752, w_056_1753, w_056_1754, w_056_1755, w_056_1756, w_056_1758, w_056_1760, w_056_1761, w_056_1762, w_056_1763, w_056_1764, w_056_1765, w_056_1766, w_056_1767, w_056_1768, w_056_1770, w_056_1771, w_056_1772, w_056_1773, w_056_1774, w_056_1775, w_056_1776, w_056_1777, w_056_1779, w_056_1780, w_056_1781, w_056_1783, w_056_1784, w_056_1785, w_056_1786, w_056_1787, w_056_1788, w_056_1789, w_056_1790, w_056_1791, w_056_1793, w_056_1794, w_056_1795, w_056_1796, w_056_1797, w_056_1798, w_056_1799, w_056_1800, w_056_1801, w_056_1802, w_056_1803, w_056_1804, w_056_1805, w_056_1806, w_056_1807, w_056_1808, w_056_1809, w_056_1810, w_056_1811, w_056_1814, w_056_1815, w_056_1816, w_056_1817, w_056_1820, w_056_1822, w_056_1824, w_056_1825, w_056_1826, w_056_1827, w_056_1828, w_056_1829, w_056_1830, w_056_1832, w_056_1833, w_056_1834, w_056_1835, w_056_1838, w_056_1839, w_056_1840, w_056_1842, w_056_1843, w_056_1844, w_056_1846, w_056_1847, w_056_1848, w_056_1849, w_056_1850, w_056_1851, w_056_1852, w_056_1854, w_056_1856, w_056_1857, w_056_1858, w_056_1859, w_056_1860, w_056_1861, w_056_1862, w_056_1863, w_056_1864, w_056_1865, w_056_1866, w_056_1867, w_056_1868, w_056_1872, w_056_1873, w_056_1874, w_056_1875, w_056_1876, w_056_1877, w_056_1881, w_056_1882, w_056_1883, w_056_1884, w_056_1885, w_056_1887, w_056_1888, w_056_1889, w_056_1890, w_056_1891, w_056_1892, w_056_1893, w_056_1894, w_056_1895, w_056_1896, w_056_1898, w_056_1899, w_056_1900, w_056_1901, w_056_1902, w_056_1903, w_056_1905, w_056_1907, w_056_1908, w_056_1909, w_056_1910, w_056_1911, w_056_1912, w_056_1913, w_056_1914, w_056_1915, w_056_1916, w_056_1917, w_056_1918, w_056_1919, w_056_1920, w_056_1921, w_056_1924, w_056_1925, w_056_1928, w_056_1929, w_056_1930, w_056_1931, w_056_1932, w_056_1933, w_056_1935, w_056_1939, w_056_1940, w_056_1941, w_056_1942, w_056_1943, w_056_1944, w_056_1945, w_056_1946, w_056_1947, w_056_1949, w_056_1950, w_056_1951, w_056_1953, w_056_1955, w_056_1956, w_056_1957, w_056_1958, w_056_1959, w_056_1960, w_056_1961, w_056_1962, w_056_1963, w_056_1964, w_056_1965, w_056_1966, w_056_1967, w_056_1968, w_056_1969, w_056_1971, w_056_1972, w_056_1974, w_056_1976, w_056_1977, w_056_1978, w_056_1980, w_056_1981, w_056_1982, w_056_1983, w_056_1984, w_056_1985, w_056_1986, w_056_1987, w_056_1988, w_056_1989, w_056_1990, w_056_1991, w_056_1992, w_056_1993, w_056_1994, w_056_1995, w_056_1996, w_056_1997, w_056_1999, w_056_2000, w_056_2001, w_056_2003, w_056_2004, w_056_2005, w_056_2006, w_056_2007, w_056_2009, w_056_2010, w_056_2012, w_056_2014, w_056_2015, w_056_2016, w_056_2017, w_056_2018, w_056_2019, w_056_2020, w_056_2021, w_056_2022, w_056_2023, w_056_2024, w_056_2025, w_056_2026, w_056_2027, w_056_2028, w_056_2029, w_056_2030, w_056_2031, w_056_2032, w_056_2033, w_056_2034, w_056_2035, w_056_2036, w_056_2037, w_056_2039, w_056_2041, w_056_2042, w_056_2043, w_056_2044, w_056_2047, w_056_2048, w_056_2050, w_056_2052, w_056_2053, w_056_2054, w_056_2055, w_056_2056, w_056_2057, w_056_2058, w_056_2059, w_056_2060, w_056_2061, w_056_2062, w_056_2063, w_056_2064, w_056_2065, w_056_2066, w_056_2067, w_056_2068, w_056_2069, w_056_2070, w_056_2071, w_056_2072, w_056_2073, w_056_2074, w_056_2075, w_056_2076, w_056_2077, w_056_2078, w_056_2079, w_056_2080, w_056_2081, w_056_2082, w_056_2083, w_056_2084, w_056_2085, w_056_2086, w_056_2087, w_056_2090, w_056_2091, w_056_2092, w_056_2093, w_056_2095, w_056_2096, w_056_2097, w_056_2098, w_056_2099, w_056_2100, w_056_2101, w_056_2102, w_056_2103, w_056_2104, w_056_2105, w_056_2107, w_056_2108, w_056_2109, w_056_2110, w_056_2112, w_056_2113, w_056_2114, w_056_2115, w_056_2117, w_056_2118, w_056_2119, w_056_2121, w_056_2122, w_056_2123, w_056_2124, w_056_2125, w_056_2126, w_056_2130, w_056_2131, w_056_2132, w_056_2133, w_056_2134, w_056_2135, w_056_2136, w_056_2137, w_056_2138, w_056_2139, w_056_2140, w_056_2141, w_056_2142, w_056_2143, w_056_2144, w_056_2145, w_056_2146, w_056_2147, w_056_2148, w_056_2149, w_056_2150, w_056_2151, w_056_2152, w_056_2153, w_056_2154, w_056_2155, w_056_2156, w_056_2158, w_056_2160, w_056_2161, w_056_2162, w_056_2163, w_056_2164, w_056_2166, w_056_2167, w_056_2168, w_056_2170, w_056_2173, w_056_2174, w_056_2175, w_056_2176, w_056_2177, w_056_2178, w_056_2179, w_056_2180, w_056_2181, w_056_2182, w_056_2183, w_056_2184, w_056_2185, w_056_2186, w_056_2187, w_056_2188, w_056_2189, w_056_2190, w_056_2192, w_056_2193, w_056_2194, w_056_2195, w_056_2196, w_056_2197, w_056_2199, w_056_2200, w_056_2201, w_056_2202, w_056_2203, w_056_2204, w_056_2205, w_056_2206, w_056_2207, w_056_2208, w_056_2209, w_056_2210, w_056_2211, w_056_2212, w_056_2213, w_056_2215, w_056_2217, w_056_2218, w_056_2219, w_056_2220, w_056_2221, w_056_2222, w_056_2223, w_056_2224, w_056_2225, w_056_2226, w_056_2227, w_056_2229, w_056_2230, w_056_2232, w_056_2233, w_056_2234, w_056_2236, w_056_2237, w_056_2238, w_056_2241, w_056_2242, w_056_2243, w_056_2244, w_056_2245, w_056_2246, w_056_2247, w_056_2248, w_056_2249, w_056_2250, w_056_2251, w_056_2252, w_056_2254, w_056_2255, w_056_2256, w_056_2257, w_056_2259, w_056_2260, w_056_2261, w_056_2262, w_056_2263, w_056_2264, w_056_2265, w_056_2266, w_056_2267, w_056_2268, w_056_2270, w_056_2271, w_056_2274, w_056_2275, w_056_2276, w_056_2277, w_056_2278, w_056_2279, w_056_2280, w_056_2281, w_056_2282, w_056_2283, w_056_2284, w_056_2286, w_056_2287, w_056_2288, w_056_2289, w_056_2290, w_056_2291, w_056_2292, w_056_2293, w_056_2294, w_056_2295, w_056_2297, w_056_2298, w_056_2299, w_056_2300, w_056_2301, w_056_2302, w_056_2303, w_056_2304, w_056_2305, w_056_2306, w_056_2307, w_056_2308, w_056_2309, w_056_2310, w_056_2311, w_056_2312, w_056_2313, w_056_2315, w_056_2316, w_056_2317, w_056_2318, w_056_2319, w_056_2320, w_056_2321, w_056_2322, w_056_2323, w_056_2324, w_056_2325, w_056_2327, w_056_2328, w_056_2329, w_056_2332, w_056_2333, w_056_2334, w_056_2336, w_056_2338, w_056_2339, w_056_2340, w_056_2342, w_056_2345, w_056_2346, w_056_2347, w_056_2348, w_056_2349, w_056_2350, w_056_2351, w_056_2352, w_056_2353, w_056_2354, w_056_2355, w_056_2356, w_056_2357, w_056_2358, w_056_2359, w_056_2360, w_056_2361, w_056_2362, w_056_2364, w_056_2367, w_056_2368, w_056_2369, w_056_2370, w_056_2371;
  wire w_057_001, w_057_002, w_057_004, w_057_006, w_057_007, w_057_009, w_057_010, w_057_011, w_057_012, w_057_014, w_057_015, w_057_016, w_057_021, w_057_022, w_057_023, w_057_024, w_057_025, w_057_026, w_057_027, w_057_029, w_057_030, w_057_032, w_057_033, w_057_035, w_057_036, w_057_038, w_057_039, w_057_040, w_057_041, w_057_043, w_057_044, w_057_045, w_057_048, w_057_049, w_057_050, w_057_051, w_057_052, w_057_053, w_057_054, w_057_056, w_057_057, w_057_058, w_057_059, w_057_060, w_057_062, w_057_063, w_057_064, w_057_065, w_057_066, w_057_067, w_057_068, w_057_069, w_057_070, w_057_071, w_057_072, w_057_074, w_057_075, w_057_076, w_057_077, w_057_078, w_057_079, w_057_081, w_057_082, w_057_084, w_057_085, w_057_087, w_057_088, w_057_089, w_057_090, w_057_091, w_057_092, w_057_093, w_057_094, w_057_095, w_057_096, w_057_098, w_057_100, w_057_101, w_057_102, w_057_105, w_057_107, w_057_108, w_057_111, w_057_113, w_057_114, w_057_115, w_057_116, w_057_117, w_057_118, w_057_119, w_057_121, w_057_122, w_057_123, w_057_124, w_057_125, w_057_126, w_057_127, w_057_128, w_057_129, w_057_130, w_057_131, w_057_132, w_057_133, w_057_134, w_057_136, w_057_137, w_057_139, w_057_140, w_057_141, w_057_142, w_057_143, w_057_144, w_057_147, w_057_148, w_057_149, w_057_150, w_057_151, w_057_152, w_057_154, w_057_156, w_057_157, w_057_159, w_057_160, w_057_161, w_057_162, w_057_163, w_057_164, w_057_165, w_057_166, w_057_167, w_057_168, w_057_170, w_057_171, w_057_172, w_057_173, w_057_174, w_057_176, w_057_177, w_057_178, w_057_179, w_057_181, w_057_182, w_057_183, w_057_184, w_057_188, w_057_189, w_057_190, w_057_191, w_057_192, w_057_193, w_057_194, w_057_195, w_057_196, w_057_197, w_057_198, w_057_199, w_057_200, w_057_201, w_057_202, w_057_206, w_057_207, w_057_208, w_057_209, w_057_210, w_057_211, w_057_212, w_057_214, w_057_215, w_057_216, w_057_217, w_057_218, w_057_219, w_057_220, w_057_222, w_057_224, w_057_225, w_057_226, w_057_228, w_057_230, w_057_231, w_057_234, w_057_235, w_057_237, w_057_240, w_057_243, w_057_244, w_057_245, w_057_246, w_057_247, w_057_249, w_057_251, w_057_252, w_057_253, w_057_256, w_057_258, w_057_260, w_057_261, w_057_262, w_057_265, w_057_266, w_057_269, w_057_270, w_057_271, w_057_272, w_057_273, w_057_274, w_057_276, w_057_277, w_057_278, w_057_279, w_057_280, w_057_281, w_057_282, w_057_283, w_057_284, w_057_285, w_057_286, w_057_287, w_057_288, w_057_289, w_057_291, w_057_293, w_057_294, w_057_295, w_057_296, w_057_297, w_057_298, w_057_300, w_057_302, w_057_303, w_057_304, w_057_305, w_057_306, w_057_309, w_057_311, w_057_312, w_057_313, w_057_314, w_057_315, w_057_316, w_057_317, w_057_318, w_057_319, w_057_320, w_057_321, w_057_324, w_057_325, w_057_326, w_057_327, w_057_329, w_057_330, w_057_331, w_057_332, w_057_336, w_057_337, w_057_338, w_057_339, w_057_340, w_057_341, w_057_344, w_057_345, w_057_346, w_057_347, w_057_348, w_057_349, w_057_351, w_057_352, w_057_353, w_057_356, w_057_357, w_057_358, w_057_359, w_057_361, w_057_363, w_057_364, w_057_365, w_057_366, w_057_367, w_057_368, w_057_369, w_057_370, w_057_372, w_057_374, w_057_375, w_057_376, w_057_378, w_057_379, w_057_380, w_057_381, w_057_382, w_057_383, w_057_384, w_057_385, w_057_386, w_057_388, w_057_389, w_057_390, w_057_392, w_057_393, w_057_394, w_057_395, w_057_396, w_057_397, w_057_399, w_057_401, w_057_402, w_057_407, w_057_408, w_057_409, w_057_410, w_057_411, w_057_412, w_057_413, w_057_414, w_057_416, w_057_417, w_057_419, w_057_420, w_057_421, w_057_422, w_057_423, w_057_424, w_057_425, w_057_426, w_057_427, w_057_428, w_057_429, w_057_430, w_057_431, w_057_432, w_057_433, w_057_435, w_057_436, w_057_437, w_057_438, w_057_439, w_057_440, w_057_442, w_057_443, w_057_444, w_057_446, w_057_447, w_057_448, w_057_449, w_057_450, w_057_452, w_057_453, w_057_454, w_057_455, w_057_456, w_057_457, w_057_458, w_057_459, w_057_461, w_057_462, w_057_463, w_057_465, w_057_468, w_057_469, w_057_470, w_057_471, w_057_472, w_057_473, w_057_474, w_057_475, w_057_476, w_057_477, w_057_478, w_057_479, w_057_480, w_057_481, w_057_482, w_057_483, w_057_484, w_057_486, w_057_487, w_057_488, w_057_489, w_057_491, w_057_492, w_057_493, w_057_494, w_057_495, w_057_496, w_057_497, w_057_498, w_057_501, w_057_502, w_057_503, w_057_504, w_057_506, w_057_508, w_057_510, w_057_511, w_057_512, w_057_514, w_057_516, w_057_517, w_057_518, w_057_519, w_057_520, w_057_521, w_057_525, w_057_527, w_057_528, w_057_529, w_057_531, w_057_532, w_057_533, w_057_535, w_057_536, w_057_537, w_057_538, w_057_539, w_057_540, w_057_542, w_057_543, w_057_544, w_057_545, w_057_546, w_057_547, w_057_549, w_057_550, w_057_551, w_057_553, w_057_554, w_057_555, w_057_556, w_057_557, w_057_560, w_057_561, w_057_563, w_057_564, w_057_567, w_057_568, w_057_569, w_057_570, w_057_571, w_057_573, w_057_575, w_057_576, w_057_577, w_057_578, w_057_579, w_057_580, w_057_581, w_057_582, w_057_583, w_057_584, w_057_585, w_057_587, w_057_588, w_057_589, w_057_591, w_057_597, w_057_599, w_057_601, w_057_602, w_057_603, w_057_608, w_057_609, w_057_610, w_057_611, w_057_612, w_057_614, w_057_615, w_057_616, w_057_618, w_057_619, w_057_621, w_057_622, w_057_623, w_057_624, w_057_625, w_057_627, w_057_628, w_057_631, w_057_632, w_057_633, w_057_635, w_057_636, w_057_637, w_057_638, w_057_639, w_057_640, w_057_641, w_057_642, w_057_646, w_057_647, w_057_649, w_057_650, w_057_651, w_057_652, w_057_653, w_057_654, w_057_655, w_057_656, w_057_657, w_057_658, w_057_660, w_057_661, w_057_662, w_057_664, w_057_665, w_057_667, w_057_668, w_057_670, w_057_671, w_057_672, w_057_673, w_057_674, w_057_675, w_057_676, w_057_677, w_057_678, w_057_680, w_057_682, w_057_684, w_057_687, w_057_688, w_057_689, w_057_692, w_057_693, w_057_694, w_057_695, w_057_696, w_057_697, w_057_698, w_057_699, w_057_702, w_057_703, w_057_705, w_057_706, w_057_707, w_057_709, w_057_710, w_057_711, w_057_712, w_057_713, w_057_714, w_057_715, w_057_717, w_057_718, w_057_720, w_057_721, w_057_722, w_057_723, w_057_724, w_057_725, w_057_726, w_057_727, w_057_728, w_057_730, w_057_731, w_057_733, w_057_734, w_057_735, w_057_736, w_057_737, w_057_738, w_057_739, w_057_740, w_057_741, w_057_743, w_057_744, w_057_745, w_057_746, w_057_747, w_057_748, w_057_749, w_057_750, w_057_753, w_057_755, w_057_756, w_057_759, w_057_760, w_057_763, w_057_764, w_057_765, w_057_766, w_057_767, w_057_769, w_057_771, w_057_773, w_057_774, w_057_775, w_057_776, w_057_777, w_057_778, w_057_779, w_057_780, w_057_781, w_057_782, w_057_783, w_057_785, w_057_786, w_057_788, w_057_789, w_057_790, w_057_791, w_057_792, w_057_793, w_057_794, w_057_795, w_057_797, w_057_798, w_057_799, w_057_800, w_057_801, w_057_802, w_057_803, w_057_804, w_057_805, w_057_806, w_057_807, w_057_808, w_057_809, w_057_810, w_057_811, w_057_812, w_057_814, w_057_816, w_057_818, w_057_819, w_057_820, w_057_821, w_057_822, w_057_826, w_057_829, w_057_830, w_057_831, w_057_832, w_057_833, w_057_834, w_057_835, w_057_836, w_057_837, w_057_838, w_057_839, w_057_842, w_057_843, w_057_845, w_057_846, w_057_848, w_057_849, w_057_850, w_057_851, w_057_853, w_057_854, w_057_855, w_057_859, w_057_860, w_057_863, w_057_865, w_057_866, w_057_867, w_057_868, w_057_869, w_057_870, w_057_871, w_057_873, w_057_874, w_057_875, w_057_876, w_057_877, w_057_879, w_057_880, w_057_881, w_057_883, w_057_888, w_057_889, w_057_892, w_057_893, w_057_895, w_057_896, w_057_897, w_057_899, w_057_900, w_057_902, w_057_903, w_057_906, w_057_907, w_057_909, w_057_910, w_057_911, w_057_913, w_057_914, w_057_916, w_057_917, w_057_919, w_057_920, w_057_921, w_057_922, w_057_923, w_057_924, w_057_925, w_057_926, w_057_927, w_057_928, w_057_929, w_057_930, w_057_932, w_057_934, w_057_935, w_057_936, w_057_937, w_057_938, w_057_939, w_057_940, w_057_941, w_057_942, w_057_943, w_057_945, w_057_946, w_057_948, w_057_949, w_057_953, w_057_954, w_057_956, w_057_957, w_057_958, w_057_959, w_057_961, w_057_962, w_057_963, w_057_964, w_057_965, w_057_966, w_057_967, w_057_968, w_057_969, w_057_971, w_057_972, w_057_973, w_057_976, w_057_979, w_057_980, w_057_981, w_057_982, w_057_984, w_057_985, w_057_986, w_057_987, w_057_988, w_057_989, w_057_990, w_057_991, w_057_993, w_057_994, w_057_995, w_057_997, w_057_1000, w_057_1001, w_057_1002, w_057_1004, w_057_1005, w_057_1007, w_057_1008, w_057_1009, w_057_1010, w_057_1011, w_057_1012, w_057_1013, w_057_1014, w_057_1017, w_057_1018, w_057_1019, w_057_1020, w_057_1021, w_057_1022, w_057_1023, w_057_1024, w_057_1025, w_057_1026, w_057_1027, w_057_1030, w_057_1032, w_057_1033, w_057_1034, w_057_1036, w_057_1037, w_057_1038, w_057_1039, w_057_1040, w_057_1041, w_057_1042, w_057_1043, w_057_1044, w_057_1045, w_057_1046, w_057_1047, w_057_1049, w_057_1051, w_057_1052, w_057_1053, w_057_1055, w_057_1056, w_057_1057, w_057_1060, w_057_1062, w_057_1063, w_057_1066, w_057_1067, w_057_1068, w_057_1069, w_057_1071, w_057_1073, w_057_1074, w_057_1075, w_057_1076, w_057_1077, w_057_1078, w_057_1079, w_057_1080, w_057_1081, w_057_1082, w_057_1083, w_057_1084, w_057_1085, w_057_1086, w_057_1087, w_057_1088, w_057_1089, w_057_1091, w_057_1093, w_057_1094, w_057_1095, w_057_1096, w_057_1098, w_057_1099, w_057_1100, w_057_1101, w_057_1102, w_057_1104, w_057_1107, w_057_1108, w_057_1110, w_057_1113, w_057_1115, w_057_1117, w_057_1119, w_057_1120, w_057_1121, w_057_1122, w_057_1123, w_057_1124, w_057_1126, w_057_1127, w_057_1130, w_057_1132, w_057_1133, w_057_1137, w_057_1138, w_057_1139, w_057_1142, w_057_1144, w_057_1145, w_057_1146, w_057_1148, w_057_1149, w_057_1152, w_057_1155, w_057_1156, w_057_1158, w_057_1159, w_057_1161, w_057_1163, w_057_1165, w_057_1166, w_057_1171, w_057_1172, w_057_1173, w_057_1174, w_057_1175, w_057_1177, w_057_1178, w_057_1179, w_057_1182, w_057_1183, w_057_1184, w_057_1185, w_057_1186, w_057_1187, w_057_1188, w_057_1190, w_057_1193, w_057_1194, w_057_1195, w_057_1197, w_057_1200, w_057_1202, w_057_1203, w_057_1205, w_057_1206, w_057_1207, w_057_1209, w_057_1211, w_057_1212, w_057_1221, w_057_1222, w_057_1223, w_057_1224, w_057_1225, w_057_1226, w_057_1227, w_057_1228, w_057_1229, w_057_1231, w_057_1232, w_057_1233, w_057_1234, w_057_1235, w_057_1236, w_057_1239, w_057_1240, w_057_1241, w_057_1242, w_057_1243, w_057_1244, w_057_1248, w_057_1249, w_057_1250, w_057_1251, w_057_1252, w_057_1254, w_057_1255, w_057_1257, w_057_1259, w_057_1260, w_057_1261, w_057_1262, w_057_1264, w_057_1265, w_057_1271, w_057_1272, w_057_1273, w_057_1277, w_057_1278, w_057_1280, w_057_1283, w_057_1286, w_057_1288, w_057_1289, w_057_1291, w_057_1294, w_057_1296, w_057_1297, w_057_1298, w_057_1299, w_057_1300, w_057_1301, w_057_1303, w_057_1306, w_057_1307, w_057_1308, w_057_1313, w_057_1314, w_057_1316, w_057_1317, w_057_1318, w_057_1319, w_057_1321, w_057_1322, w_057_1323, w_057_1324, w_057_1325, w_057_1326, w_057_1327, w_057_1331, w_057_1333, w_057_1334, w_057_1335, w_057_1338, w_057_1340, w_057_1341, w_057_1342, w_057_1343, w_057_1344, w_057_1347, w_057_1350, w_057_1352, w_057_1353, w_057_1354, w_057_1355, w_057_1357, w_057_1359, w_057_1360, w_057_1361, w_057_1362, w_057_1363, w_057_1364, w_057_1367, w_057_1368, w_057_1369, w_057_1370, w_057_1371, w_057_1373, w_057_1374, w_057_1376, w_057_1377, w_057_1379, w_057_1381, w_057_1382, w_057_1388, w_057_1389, w_057_1391, w_057_1393, w_057_1394, w_057_1395, w_057_1396, w_057_1398, w_057_1403, w_057_1405, w_057_1407, w_057_1408, w_057_1413, w_057_1415, w_057_1416, w_057_1418, w_057_1419, w_057_1421, w_057_1422, w_057_1423, w_057_1425, w_057_1426, w_057_1427, w_057_1428, w_057_1431, w_057_1432, w_057_1433, w_057_1434, w_057_1435, w_057_1439, w_057_1440, w_057_1441, w_057_1442, w_057_1443, w_057_1444, w_057_1446, w_057_1447, w_057_1449, w_057_1450, w_057_1451, w_057_1455, w_057_1457, w_057_1458, w_057_1459, w_057_1461, w_057_1463, w_057_1464, w_057_1466, w_057_1467, w_057_1470, w_057_1471, w_057_1472, w_057_1475, w_057_1477, w_057_1478, w_057_1479, w_057_1481, w_057_1482, w_057_1483, w_057_1484, w_057_1485, w_057_1486, w_057_1488, w_057_1489, w_057_1493, w_057_1497, w_057_1499, w_057_1502, w_057_1503, w_057_1504, w_057_1505, w_057_1506, w_057_1507, w_057_1508, w_057_1509, w_057_1510, w_057_1511, w_057_1512, w_057_1513, w_057_1514, w_057_1516, w_057_1518, w_057_1519, w_057_1520, w_057_1522, w_057_1524, w_057_1525, w_057_1527, w_057_1529, w_057_1531, w_057_1532, w_057_1533, w_057_1534, w_057_1538, w_057_1539, w_057_1542, w_057_1549, w_057_1552, w_057_1554, w_057_1555, w_057_1558, w_057_1560, w_057_1561, w_057_1562, w_057_1563, w_057_1565, w_057_1566, w_057_1567, w_057_1568, w_057_1569, w_057_1571, w_057_1572, w_057_1573, w_057_1574, w_057_1575, w_057_1577, w_057_1578, w_057_1580, w_057_1581, w_057_1582, w_057_1585, w_057_1588, w_057_1590, w_057_1591, w_057_1592, w_057_1593, w_057_1594, w_057_1595, w_057_1597, w_057_1598, w_057_1600, w_057_1601, w_057_1602, w_057_1605, w_057_1606, w_057_1607, w_057_1608, w_057_1610, w_057_1613, w_057_1615, w_057_1616, w_057_1619, w_057_1620, w_057_1622, w_057_1623, w_057_1624, w_057_1625, w_057_1628, w_057_1629, w_057_1630, w_057_1631, w_057_1632, w_057_1633, w_057_1634, w_057_1635, w_057_1637, w_057_1638, w_057_1642, w_057_1643, w_057_1645, w_057_1646, w_057_1648, w_057_1651, w_057_1653, w_057_1654, w_057_1655, w_057_1656, w_057_1660, w_057_1661, w_057_1662, w_057_1665, w_057_1668, w_057_1669, w_057_1672, w_057_1674, w_057_1677, w_057_1679, w_057_1680, w_057_1682, w_057_1683, w_057_1685, w_057_1686, w_057_1688, w_057_1689, w_057_1690, w_057_1691, w_057_1692, w_057_1694, w_057_1695, w_057_1696, w_057_1697, w_057_1698, w_057_1699, w_057_1701, w_057_1702, w_057_1703, w_057_1704, w_057_1706, w_057_1707, w_057_1711, w_057_1712, w_057_1713, w_057_1714, w_057_1715, w_057_1716, w_057_1717, w_057_1718, w_057_1720, w_057_1721, w_057_1725, w_057_1726, w_057_1727, w_057_1728, w_057_1730, w_057_1731, w_057_1733, w_057_1735, w_057_1737, w_057_1738, w_057_1739, w_057_1740, w_057_1741, w_057_1742, w_057_1743, w_057_1744, w_057_1745, w_057_1746, w_057_1747, w_057_1748, w_057_1749, w_057_1750, w_057_1751, w_057_1752, w_057_1754, w_057_1755, w_057_1757, w_057_1758, w_057_1759, w_057_1760, w_057_1761, w_057_1762, w_057_1763, w_057_1765, w_057_1766, w_057_1768, w_057_1771, w_057_1772, w_057_1773, w_057_1774, w_057_1776, w_057_1777, w_057_1779, w_057_1780, w_057_1781, w_057_1789, w_057_1791, w_057_1792, w_057_1793, w_057_1794, w_057_1795, w_057_1796, w_057_1798, w_057_1800, w_057_1801, w_057_1802, w_057_1805, w_057_1809, w_057_1811, w_057_1812, w_057_1814, w_057_1818, w_057_1820, w_057_1821, w_057_1823, w_057_1826, w_057_1827, w_057_1828, w_057_1829, w_057_1830, w_057_1831, w_057_1832, w_057_1833, w_057_1834, w_057_1836, w_057_1838, w_057_1839, w_057_1840, w_057_1841, w_057_1844, w_057_1845, w_057_1846, w_057_1849, w_057_1851, w_057_1854, w_057_1855, w_057_1856, w_057_1859, w_057_1861, w_057_1862, w_057_1863, w_057_1865, w_057_1866, w_057_1868, w_057_1870, w_057_1871, w_057_1874, w_057_1875, w_057_1876, w_057_1878, w_057_1880, w_057_1881, w_057_1883, w_057_1885, w_057_1887, w_057_1889, w_057_1890, w_057_1891, w_057_1895, w_057_1896, w_057_1897, w_057_1898, w_057_1899, w_057_1900, w_057_1902, w_057_1903, w_057_1905, w_057_1908, w_057_1909, w_057_1910, w_057_1912, w_057_1915, w_057_1916, w_057_1917, w_057_1918, w_057_1919, w_057_1923, w_057_1925, w_057_1927, w_057_1929, w_057_1931, w_057_1933, w_057_1934, w_057_1935, w_057_1936, w_057_1937, w_057_1938, w_057_1941, w_057_1942, w_057_1943, w_057_1944, w_057_1945, w_057_1946, w_057_1947, w_057_1948, w_057_1951, w_057_1954, w_057_1955, w_057_1957, w_057_1958, w_057_1960, w_057_1963, w_057_1965, w_057_1966, w_057_1967, w_057_1968, w_057_1969, w_057_1970, w_057_1976, w_057_1978, w_057_1979, w_057_1982, w_057_1983, w_057_1984, w_057_1985, w_057_1987, w_057_1988, w_057_1989, w_057_1991, w_057_1992, w_057_1993, w_057_1994, w_057_1997, w_057_1998, w_057_1999, w_057_2001, w_057_2004, w_057_2005, w_057_2006, w_057_2007, w_057_2008, w_057_2010, w_057_2012, w_057_2013, w_057_2014, w_057_2015, w_057_2016, w_057_2017, w_057_2019, w_057_2020, w_057_2021, w_057_2022, w_057_2025, w_057_2026, w_057_2027, w_057_2028, w_057_2029, w_057_2030, w_057_2031, w_057_2032, w_057_2033, w_057_2034, w_057_2035, w_057_2036, w_057_2037, w_057_2038, w_057_2039, w_057_2040, w_057_2041, w_057_2043, w_057_2044, w_057_2045, w_057_2050, w_057_2051, w_057_2053, w_057_2054, w_057_2058, w_057_2060, w_057_2061, w_057_2063, w_057_2064, w_057_2066, w_057_2068, w_057_2069, w_057_2070, w_057_2071, w_057_2072, w_057_2073, w_057_2075, w_057_2077, w_057_2078, w_057_2079, w_057_2081, w_057_2084, w_057_2086, w_057_2087, w_057_2088, w_057_2090, w_057_2091, w_057_2094, w_057_2095, w_057_2096, w_057_2098, w_057_2100, w_057_2101, w_057_2106, w_057_2107, w_057_2108, w_057_2109, w_057_2114, w_057_2117, w_057_2118, w_057_2121, w_057_2123, w_057_2124, w_057_2126, w_057_2127, w_057_2128, w_057_2136, w_057_2137, w_057_2138, w_057_2139, w_057_2140, w_057_2143, w_057_2144, w_057_2145, w_057_2146, w_057_2147, w_057_2148, w_057_2149, w_057_2150, w_057_2151, w_057_2155, w_057_2157, w_057_2158, w_057_2159, w_057_2160, w_057_2161, w_057_2162, w_057_2163, w_057_2166, w_057_2167, w_057_2168, w_057_2169, w_057_2170, w_057_2171, w_057_2172, w_057_2173, w_057_2174, w_057_2175, w_057_2176, w_057_2177, w_057_2178, w_057_2179, w_057_2180, w_057_2182, w_057_2185, w_057_2186, w_057_2187, w_057_2188, w_057_2189, w_057_2192, w_057_2193, w_057_2194, w_057_2196, w_057_2197, w_057_2200, w_057_2201, w_057_2202, w_057_2203, w_057_2204, w_057_2205, w_057_2206, w_057_2207, w_057_2209, w_057_2210, w_057_2211, w_057_2212, w_057_2217, w_057_2219, w_057_2220, w_057_2222, w_057_2223, w_057_2224, w_057_2225, w_057_2226, w_057_2228, w_057_2230, w_057_2231, w_057_2233, w_057_2235, w_057_2237, w_057_2238, w_057_2239, w_057_2240, w_057_2243, w_057_2244, w_057_2245, w_057_2246, w_057_2247, w_057_2250, w_057_2253, w_057_2254, w_057_2255, w_057_2256, w_057_2258, w_057_2260, w_057_2261, w_057_2263, w_057_2265, w_057_2266, w_057_2268, w_057_2269, w_057_2270, w_057_2271, w_057_2274, w_057_2275, w_057_2276, w_057_2277, w_057_2278, w_057_2279, w_057_2280, w_057_2281, w_057_2282, w_057_2284, w_057_2289, w_057_2290, w_057_2291, w_057_2292, w_057_2294, w_057_2296, w_057_2298, w_057_2301, w_057_2302, w_057_2304, w_057_2305, w_057_2306, w_057_2307, w_057_2309, w_057_2310, w_057_2311, w_057_2316, w_057_2317, w_057_2321, w_057_2322, w_057_2326, w_057_2327, w_057_2329, w_057_2330, w_057_2331, w_057_2332, w_057_2333, w_057_2334, w_057_2335, w_057_2336, w_057_2337, w_057_2338, w_057_2339, w_057_2340, w_057_2342, w_057_2344, w_057_2345, w_057_2348, w_057_2351, w_057_2352, w_057_2354, w_057_2355, w_057_2356, w_057_2359, w_057_2360, w_057_2363, w_057_2364, w_057_2365, w_057_2368, w_057_2369, w_057_2372, w_057_2373, w_057_2376, w_057_2377, w_057_2378, w_057_2379, w_057_2381, w_057_2382, w_057_2383, w_057_2385, w_057_2386, w_057_2387, w_057_2388, w_057_2389, w_057_2390, w_057_2391, w_057_2392, w_057_2393, w_057_2395, w_057_2397, w_057_2398, w_057_2399, w_057_2400, w_057_2404, w_057_2405, w_057_2407, w_057_2409, w_057_2411, w_057_2412, w_057_2414, w_057_2415, w_057_2416, w_057_2417, w_057_2418, w_057_2420, w_057_2421, w_057_2424, w_057_2425, w_057_2426, w_057_2427, w_057_2430, w_057_2431, w_057_2432, w_057_2433, w_057_2435, w_057_2436, w_057_2438, w_057_2439, w_057_2440, w_057_2441, w_057_2442, w_057_2444, w_057_2445, w_057_2446, w_057_2447, w_057_2449, w_057_2454, w_057_2456, w_057_2457, w_057_2461, w_057_2462, w_057_2464, w_057_2465, w_057_2467, w_057_2469, w_057_2473, w_057_2475, w_057_2476, w_057_2478, w_057_2479, w_057_2480, w_057_2481, w_057_2482, w_057_2483, w_057_2484, w_057_2485, w_057_2486, w_057_2488, w_057_2491, w_057_2492, w_057_2493, w_057_2494, w_057_2499, w_057_2500, w_057_2502, w_057_2503, w_057_2504, w_057_2505, w_057_2506, w_057_2508, w_057_2509, w_057_2512, w_057_2513, w_057_2514, w_057_2515, w_057_2516, w_057_2520, w_057_2522, w_057_2525, w_057_2526, w_057_2527, w_057_2528, w_057_2529, w_057_2530, w_057_2533, w_057_2534, w_057_2537, w_057_2538, w_057_2539, w_057_2540, w_057_2541, w_057_2542, w_057_2543, w_057_2544, w_057_2545, w_057_2546, w_057_2548, w_057_2549, w_057_2550, w_057_2558, w_057_2561, w_057_2562, w_057_2563, w_057_2564, w_057_2567, w_057_2568, w_057_2569, w_057_2571, w_057_2572, w_057_2573, w_057_2574, w_057_2575, w_057_2576, w_057_2577, w_057_2578, w_057_2579, w_057_2582, w_057_2583, w_057_2584, w_057_2587, w_057_2589, w_057_2590, w_057_2591, w_057_2592, w_057_2594, w_057_2596, w_057_2597, w_057_2598, w_057_2600, w_057_2602, w_057_2605, w_057_2607, w_057_2608, w_057_2609, w_057_2613, w_057_2615, w_057_2617, w_057_2619, w_057_2620, w_057_2621, w_057_2622, w_057_2626, w_057_2627, w_057_2628, w_057_2630, w_057_2631, w_057_2636, w_057_2637, w_057_2638, w_057_2639, w_057_2640, w_057_2641, w_057_2643, w_057_2644, w_057_2645, w_057_2646, w_057_2647, w_057_2655, w_057_2658, w_057_2659, w_057_2660, w_057_2661, w_057_2662, w_057_2663, w_057_2665, w_057_2666, w_057_2668, w_057_2669, w_057_2671, w_057_2672, w_057_2674, w_057_2676, w_057_2679, w_057_2680, w_057_2682, w_057_2683, w_057_2685, w_057_2686, w_057_2689, w_057_2693, w_057_2695, w_057_2698, w_057_2703, w_057_2704, w_057_2705, w_057_2706, w_057_2707, w_057_2711, w_057_2712, w_057_2716, w_057_2719, w_057_2720, w_057_2721, w_057_2723, w_057_2724, w_057_2725, w_057_2726, w_057_2727, w_057_2728, w_057_2730, w_057_2734, w_057_2735, w_057_2737, w_057_2738, w_057_2740, w_057_2741, w_057_2742, w_057_2743, w_057_2744, w_057_2745, w_057_2746, w_057_2747, w_057_2748, w_057_2749, w_057_2752, w_057_2755, w_057_2756, w_057_2757, w_057_2759, w_057_2761, w_057_2763, w_057_2764, w_057_2765, w_057_2766, w_057_2767, w_057_2768, w_057_2771, w_057_2772, w_057_2774, w_057_2778, w_057_2782, w_057_2783, w_057_2784, w_057_2785, w_057_2786, w_057_2787, w_057_2794, w_057_2795, w_057_2799, w_057_2800, w_057_2801, w_057_2802, w_057_2806, w_057_2807, w_057_2808, w_057_2809, w_057_2810, w_057_2814, w_057_2815, w_057_2817, w_057_2818, w_057_2821, w_057_2822, w_057_2825, w_057_2828, w_057_2831, w_057_2833, w_057_2836, w_057_2838, w_057_2839, w_057_2843, w_057_2844, w_057_2845, w_057_2849, w_057_2850, w_057_2851, w_057_2852, w_057_2853, w_057_2854, w_057_2855, w_057_2856, w_057_2857, w_057_2860, w_057_2861, w_057_2865, w_057_2868, w_057_2869, w_057_2870, w_057_2872, w_057_2873, w_057_2874, w_057_2875, w_057_2876, w_057_2880, w_057_2883, w_057_2885, w_057_2887, w_057_2889, w_057_2890, w_057_2893, w_057_2894, w_057_2895, w_057_2897, w_057_2898, w_057_2900, w_057_2901, w_057_2902, w_057_2903, w_057_2905, w_057_2908, w_057_2915, w_057_2916, w_057_2917, w_057_2918, w_057_2921, w_057_2922, w_057_2923, w_057_2924, w_057_2925, w_057_2926, w_057_2927, w_057_2928, w_057_2929, w_057_2930, w_057_2931, w_057_2932, w_057_2935, w_057_2936, w_057_2938, w_057_2941, w_057_2943, w_057_2945, w_057_2946, w_057_2947, w_057_2948, w_057_2951, w_057_2952, w_057_2954, w_057_2956, w_057_2958, w_057_2959, w_057_2960, w_057_2961, w_057_2963, w_057_2964, w_057_2966, w_057_2967, w_057_2968, w_057_2971, w_057_2972, w_057_2973, w_057_2978, w_057_2979, w_057_2983, w_057_2985, w_057_2986, w_057_2989, w_057_2990, w_057_2991, w_057_2992, w_057_2993, w_057_2994, w_057_2995, w_057_2998, w_057_2999, w_057_3001, w_057_3002, w_057_3003, w_057_3005, w_057_3007, w_057_3008, w_057_3010, w_057_3012, w_057_3013, w_057_3014, w_057_3015, w_057_3016, w_057_3017, w_057_3018, w_057_3019, w_057_3022, w_057_3024, w_057_3025, w_057_3026, w_057_3027, w_057_3029, w_057_3030, w_057_3031, w_057_3035, w_057_3037, w_057_3038, w_057_3039, w_057_3044, w_057_3047, w_057_3048, w_057_3051, w_057_3052, w_057_3054, w_057_3057, w_057_3058, w_057_3059, w_057_3061, w_057_3062, w_057_3063, w_057_3064, w_057_3065, w_057_3066, w_057_3068, w_057_3071, w_057_3075, w_057_3076, w_057_3077, w_057_3080, w_057_3083, w_057_3084, w_057_3086, w_057_3087, w_057_3089, w_057_3090, w_057_3092, w_057_3094, w_057_3095, w_057_3096, w_057_3097, w_057_3098, w_057_3099, w_057_3100, w_057_3101, w_057_3103, w_057_3104, w_057_3106, w_057_3110, w_057_3111, w_057_3112, w_057_3113, w_057_3116, w_057_3118, w_057_3119, w_057_3123, w_057_3124, w_057_3125, w_057_3126, w_057_3128, w_057_3129, w_057_3130, w_057_3131, w_057_3132, w_057_3134, w_057_3136, w_057_3140, w_057_3143, w_057_3148, w_057_3149, w_057_3150, w_057_3151, w_057_3152, w_057_3154, w_057_3156, w_057_3157, w_057_3158, w_057_3160, w_057_3161, w_057_3162, w_057_3163, w_057_3166, w_057_3169, w_057_3170, w_057_3172, w_057_3174, w_057_3176, w_057_3177, w_057_3178, w_057_3184, w_057_3185, w_057_3187, w_057_3191, w_057_3192, w_057_3193, w_057_3194, w_057_3195, w_057_3196, w_057_3197, w_057_3201, w_057_3202, w_057_3204, w_057_3205, w_057_3206, w_057_3208, w_057_3209, w_057_3210, w_057_3211, w_057_3214, w_057_3215, w_057_3216, w_057_3217, w_057_3219, w_057_3222, w_057_3224, w_057_3226, w_057_3227, w_057_3230, w_057_3231, w_057_3232, w_057_3233, w_057_3235, w_057_3237, w_057_3239, w_057_3240, w_057_3242, w_057_3245, w_057_3246, w_057_3247, w_057_3248, w_057_3249, w_057_3253, w_057_3255, w_057_3256, w_057_3257, w_057_3258, w_057_3259, w_057_3261, w_057_3262, w_057_3263, w_057_3264, w_057_3266, w_057_3268, w_057_3271, w_057_3272, w_057_3273, w_057_3275, w_057_3276, w_057_3277, w_057_3278, w_057_3279, w_057_3280, w_057_3281, w_057_3283, w_057_3284, w_057_3285, w_057_3286, w_057_3288, w_057_3289, w_057_3291, w_057_3292, w_057_3293, w_057_3295, w_057_3296, w_057_3297, w_057_3298, w_057_3302, w_057_3303, w_057_3305, w_057_3306, w_057_3307, w_057_3308, w_057_3311, w_057_3314, w_057_3315, w_057_3318, w_057_3319, w_057_3322, w_057_3324, w_057_3325, w_057_3326, w_057_3328, w_057_3329, w_057_3330, w_057_3331, w_057_3332, w_057_3334, w_057_3335, w_057_3336, w_057_3337, w_057_3339, w_057_3341, w_057_3342, w_057_3343, w_057_3346, w_057_3348, w_057_3349, w_057_3350, w_057_3353, w_057_3357, w_057_3358, w_057_3360, w_057_3361, w_057_3363, w_057_3364, w_057_3365, w_057_3366, w_057_3368, w_057_3369, w_057_3370, w_057_3371, w_057_3372, w_057_3373, w_057_3375, w_057_3378, w_057_3380, w_057_3381, w_057_3384, w_057_3385, w_057_3387, w_057_3388, w_057_3390, w_057_3392, w_057_3393, w_057_3394, w_057_3396, w_057_3397, w_057_3398, w_057_3401, w_057_3402, w_057_3403, w_057_3405, w_057_3407, w_057_3408, w_057_3409, w_057_3413, w_057_3416, w_057_3417, w_057_3418, w_057_3419, w_057_3420, w_057_3421, w_057_3423, w_057_3424, w_057_3425, w_057_3427, w_057_3428, w_057_3429, w_057_3430, w_057_3431, w_057_3435, w_057_3438, w_057_3439, w_057_3440, w_057_3442, w_057_3445, w_057_3446, w_057_3447, w_057_3449, w_057_3453, w_057_3454, w_057_3455, w_057_3456, w_057_3457, w_057_3458, w_057_3459, w_057_3460, w_057_3461, w_057_3462, w_057_3464, w_057_3466, w_057_3467, w_057_3468, w_057_3469, w_057_3470, w_057_3471, w_057_3472, w_057_3473, w_057_3474, w_057_3475, w_057_3477, w_057_3479, w_057_3480, w_057_3482, w_057_3483, w_057_3484, w_057_3485, w_057_3487, w_057_3490, w_057_3491, w_057_3492, w_057_3493, w_057_3494, w_057_3495, w_057_3496, w_057_3499, w_057_3501, w_057_3502, w_057_3503, w_057_3504, w_057_3505, w_057_3506, w_057_3507, w_057_3509, w_057_3512, w_057_3514, w_057_3515, w_057_3521, w_057_3522, w_057_3523, w_057_3525, w_057_3528, w_057_3529, w_057_3530, w_057_3531, w_057_3536, w_057_3538, w_057_3539, w_057_3540, w_057_3541, w_057_3542, w_057_3544, w_057_3546, w_057_3548, w_057_3549, w_057_3550, w_057_3551, w_057_3554, w_057_3555, w_057_3557, w_057_3559, w_057_3562, w_057_3564, w_057_3567, w_057_3569, w_057_3572, w_057_3573, w_057_3574, w_057_3576, w_057_3577, w_057_3578, w_057_3580, w_057_3581, w_057_3582, w_057_3583, w_057_3584, w_057_3586, w_057_3588, w_057_3589, w_057_3592, w_057_3593, w_057_3594, w_057_3595, w_057_3598, w_057_3600, w_057_3601, w_057_3602, w_057_3603, w_057_3605, w_057_3606, w_057_3607, w_057_3609, w_057_3611, w_057_3613, w_057_3614, w_057_3617, w_057_3618, w_057_3620, w_057_3621, w_057_3622, w_057_3623, w_057_3624, w_057_3625, w_057_3626, w_057_3627, w_057_3628, w_057_3630, w_057_3631, w_057_3632, w_057_3634, w_057_3635, w_057_3637, w_057_3639, w_057_3643, w_057_3645, w_057_3646, w_057_3647, w_057_3649, w_057_3651, w_057_3652, w_057_3653, w_057_3655, w_057_3656, w_057_3657, w_057_3658, w_057_3662, w_057_3664, w_057_3665, w_057_3667, w_057_3668, w_057_3669, w_057_3670, w_057_3672, w_057_3673, w_057_3674, w_057_3677, w_057_3678, w_057_3679, w_057_3680, w_057_3683, w_057_3686, w_057_3689, w_057_3690, w_057_3691, w_057_3692, w_057_3695, w_057_3696, w_057_3697, w_057_3698, w_057_3700, w_057_3702, w_057_3703, w_057_3704, w_057_3705, w_057_3706, w_057_3708, w_057_3709, w_057_3710, w_057_3713, w_057_3716, w_057_3718, w_057_3719, w_057_3720, w_057_3721, w_057_3724, w_057_3726, w_057_3727, w_057_3728, w_057_3729, w_057_3730, w_057_3732, w_057_3733, w_057_3734, w_057_3735, w_057_3736, w_057_3739, w_057_3742, w_057_3743, w_057_3744, w_057_3747, w_057_3748, w_057_3749, w_057_3751, w_057_3755, w_057_3756, w_057_3757, w_057_3758, w_057_3761, w_057_3766, w_057_3767, w_057_3768, w_057_3769, w_057_3770, w_057_3771, w_057_3772, w_057_3773, w_057_3775, w_057_3776, w_057_3777, w_057_3778, w_057_3779, w_057_3780, w_057_3781, w_057_3783, w_057_3790, w_057_3792, w_057_3793, w_057_3794, w_057_3795, w_057_3796, w_057_3799, w_057_3801, w_057_3803, w_057_3804, w_057_3805, w_057_3807, w_057_3808, w_057_3809, w_057_3810, w_057_3812, w_057_3815, w_057_3816, w_057_3817, w_057_3818, w_057_3820, w_057_3821, w_057_3822, w_057_3823, w_057_3827, w_057_3828, w_057_3830, w_057_3831, w_057_3835, w_057_3836, w_057_3838, w_057_3839, w_057_3840, w_057_3842, w_057_3843, w_057_3845, w_057_3846, w_057_3847, w_057_3849, w_057_3852, w_057_3853, w_057_3855, w_057_3856, w_057_3857, w_057_3858, w_057_3859, w_057_3860, w_057_3862, w_057_3863, w_057_3864, w_057_3865, w_057_3867, w_057_3869, w_057_3871, w_057_3872, w_057_3874, w_057_3875, w_057_3877, w_057_3878, w_057_3879, w_057_3880, w_057_3882, w_057_3883, w_057_3884, w_057_3885, w_057_3886, w_057_3889, w_057_3896, w_057_3900, w_057_3901, w_057_3902, w_057_3903, w_057_3904, w_057_3905, w_057_3907, w_057_3908, w_057_3910, w_057_3911, w_057_3913, w_057_3915, w_057_3917, w_057_3918, w_057_3920, w_057_3922, w_057_3923, w_057_3925, w_057_3926, w_057_3931, w_057_3933, w_057_3934, w_057_3935, w_057_3936, w_057_3937, w_057_3938, w_057_3939, w_057_3940, w_057_3942, w_057_3943, w_057_3944, w_057_3946, w_057_3947, w_057_3949, w_057_3952, w_057_3956, w_057_3957, w_057_3958, w_057_3959, w_057_3960, w_057_3961, w_057_3962, w_057_3965, w_057_3966, w_057_3967, w_057_3968, w_057_3970, w_057_3971, w_057_3972, w_057_3973, w_057_3974, w_057_3977, w_057_3979, w_057_3980, w_057_3981, w_057_3982, w_057_3983, w_057_3984, w_057_3987, w_057_3990, w_057_3991, w_057_3993, w_057_3996, w_057_3997, w_057_3998, w_057_3999, w_057_4000, w_057_4001, w_057_4002, w_057_4004, w_057_4005, w_057_4007, w_057_4008, w_057_4009, w_057_4016, w_057_4021, w_057_4028, w_057_4030, w_057_4031, w_057_4032, w_057_4033, w_057_4034, w_057_4035, w_057_4038, w_057_4040, w_057_4042, w_057_4044, w_057_4046, w_057_4047, w_057_4048, w_057_4050, w_057_4053, w_057_4055, w_057_4056, w_057_4057, w_057_4058, w_057_4060, w_057_4061, w_057_4062, w_057_4063, w_057_4064, w_057_4065, w_057_4066, w_057_4067, w_057_4068, w_057_4069, w_057_4073, w_057_4074, w_057_4078, w_057_4079, w_057_4080, w_057_4082, w_057_4084, w_057_4086, w_057_4087, w_057_4089, w_057_4090, w_057_4091, w_057_4092, w_057_4093, w_057_4096, w_057_4097, w_057_4103, w_057_4105, w_057_4106, w_057_4107, w_057_4110, w_057_4112, w_057_4113, w_057_4114, w_057_4115, w_057_4116, w_057_4117, w_057_4118, w_057_4119, w_057_4120, w_057_4121, w_057_4122, w_057_4124, w_057_4126, w_057_4127, w_057_4129, w_057_4130, w_057_4131, w_057_4133, w_057_4134, w_057_4135, w_057_4138, w_057_4139, w_057_4141, w_057_4142, w_057_4143, w_057_4144, w_057_4145, w_057_4147, w_057_4148, w_057_4150, w_057_4151, w_057_4153, w_057_4155, w_057_4156, w_057_4157, w_057_4158, w_057_4160, w_057_4161, w_057_4166, w_057_4169, w_057_4171, w_057_4172, w_057_4175, w_057_4178, w_057_4180, w_057_4185, w_057_4186, w_057_4187, w_057_4188, w_057_4189, w_057_4190, w_057_4191, w_057_4192, w_057_4193, w_057_4199, w_057_4200, w_057_4201, w_057_4205, w_057_4206, w_057_4207, w_057_4209, w_057_4210, w_057_4211, w_057_4212, w_057_4214, w_057_4215, w_057_4218, w_057_4219, w_057_4220, w_057_4221, w_057_4222, w_057_4223, w_057_4224, w_057_4225, w_057_4226, w_057_4230, w_057_4231, w_057_4232, w_057_4233, w_057_4234, w_057_4235, w_057_4237, w_057_4238, w_057_4240, w_057_4243, w_057_4245, w_057_4247, w_057_4250, w_057_4252, w_057_4255, w_057_4257, w_057_4258, w_057_4259, w_057_4260, w_057_4262, w_057_4264, w_057_4265, w_057_4266, w_057_4267, w_057_4273, w_057_4274, w_057_4279, w_057_4280, w_057_4282, w_057_4283, w_057_4284, w_057_4287, w_057_4288, w_057_4289, w_057_4290, w_057_4296, w_057_4297, w_057_4300, w_057_4302, w_057_4303, w_057_4305, w_057_4306, w_057_4307, w_057_4308, w_057_4309, w_057_4310, w_057_4311, w_057_4312, w_057_4313, w_057_4315, w_057_4317, w_057_4318, w_057_4319, w_057_4322, w_057_4325, w_057_4326, w_057_4328, w_057_4329, w_057_4330, w_057_4343, w_057_4344, w_057_4348, w_057_4349, w_057_4351, w_057_4352, w_057_4353, w_057_4354, w_057_4356, w_057_4357, w_057_4358, w_057_4359, w_057_4361, w_057_4362, w_057_4365, w_057_4370, w_057_4371, w_057_4372, w_057_4373, w_057_4374, w_057_4375, w_057_4376, w_057_4377, w_057_4378, w_057_4379, w_057_4380, w_057_4381, w_057_4383, w_057_4385, w_057_4386, w_057_4387, w_057_4389, w_057_4391, w_057_4393, w_057_4396, w_057_4397, w_057_4398, w_057_4400, w_057_4401, w_057_4402, w_057_4404, w_057_4405, w_057_4407, w_057_4408, w_057_4410, w_057_4411, w_057_4412, w_057_4414, w_057_4415, w_057_4417, w_057_4419, w_057_4420, w_057_4423, w_057_4427, w_057_4428, w_057_4429, w_057_4430, w_057_4431, w_057_4432, w_057_4434, w_057_4435, w_057_4436, w_057_4437;
  wire w_058_000, w_058_002, w_058_003, w_058_005, w_058_007, w_058_009, w_058_010, w_058_011, w_058_012, w_058_013, w_058_014, w_058_015, w_058_016, w_058_017, w_058_018, w_058_019, w_058_020, w_058_022, w_058_024, w_058_025, w_058_027, w_058_028, w_058_029, w_058_030, w_058_031, w_058_032, w_058_033, w_058_034, w_058_036, w_058_037, w_058_039, w_058_040, w_058_041, w_058_042, w_058_044, w_058_045, w_058_047, w_058_048, w_058_049, w_058_050, w_058_051, w_058_055, w_058_057, w_058_058, w_058_059, w_058_060, w_058_062, w_058_063, w_058_064, w_058_066, w_058_067, w_058_069, w_058_071, w_058_072, w_058_073, w_058_074, w_058_075, w_058_076, w_058_077, w_058_078, w_058_079, w_058_080, w_058_081, w_058_082, w_058_083, w_058_084, w_058_085, w_058_086, w_058_087, w_058_088, w_058_090, w_058_091, w_058_092, w_058_093, w_058_094, w_058_095, w_058_096, w_058_097, w_058_098, w_058_099, w_058_100, w_058_101, w_058_102, w_058_103, w_058_105, w_058_106, w_058_107, w_058_108, w_058_111, w_058_113, w_058_114, w_058_115, w_058_116, w_058_117, w_058_118, w_058_120, w_058_122, w_058_124, w_058_125, w_058_126, w_058_128, w_058_130, w_058_131, w_058_133, w_058_134, w_058_135, w_058_136, w_058_137, w_058_138, w_058_140, w_058_141, w_058_143, w_058_144, w_058_145, w_058_149, w_058_150, w_058_151, w_058_153, w_058_154, w_058_155, w_058_156, w_058_157, w_058_158, w_058_159, w_058_160, w_058_161, w_058_162, w_058_163, w_058_164, w_058_165, w_058_166, w_058_167, w_058_168, w_058_169, w_058_170, w_058_172, w_058_173, w_058_174, w_058_175, w_058_177, w_058_178, w_058_179, w_058_180, w_058_181, w_058_182, w_058_183, w_058_185, w_058_188, w_058_190, w_058_192, w_058_195, w_058_196, w_058_197, w_058_198, w_058_200, w_058_202, w_058_203, w_058_204, w_058_205, w_058_206, w_058_207, w_058_209, w_058_210, w_058_212, w_058_213, w_058_214, w_058_215, w_058_216, w_058_218, w_058_220, w_058_221, w_058_222, w_058_223, w_058_224, w_058_225, w_058_226, w_058_227, w_058_228, w_058_230, w_058_231, w_058_233, w_058_234, w_058_235, w_058_236, w_058_237, w_058_238, w_058_240, w_058_241, w_058_243, w_058_245, w_058_246, w_058_247, w_058_248, w_058_249, w_058_250, w_058_251, w_058_252, w_058_254, w_058_256, w_058_257, w_058_258, w_058_260, w_058_261, w_058_262, w_058_263, w_058_265, w_058_267, w_058_270, w_058_271, w_058_272, w_058_273, w_058_274, w_058_276, w_058_277, w_058_279, w_058_280, w_058_281, w_058_282, w_058_284, w_058_285, w_058_286, w_058_287, w_058_290, w_058_291, w_058_296, w_058_297, w_058_298, w_058_299, w_058_301, w_058_303, w_058_305, w_058_307, w_058_308, w_058_309, w_058_310, w_058_311, w_058_312, w_058_314, w_058_315, w_058_316, w_058_318, w_058_319, w_058_320, w_058_321, w_058_324, w_058_325, w_058_326, w_058_327, w_058_328, w_058_329, w_058_330, w_058_331, w_058_334, w_058_335, w_058_339, w_058_340, w_058_341, w_058_342, w_058_343, w_058_344, w_058_345, w_058_346, w_058_348, w_058_349, w_058_350, w_058_351, w_058_352, w_058_353, w_058_354, w_058_355, w_058_356, w_058_358, w_058_359, w_058_360, w_058_362, w_058_365, w_058_367, w_058_368, w_058_370, w_058_371, w_058_373, w_058_374, w_058_375, w_058_378, w_058_379, w_058_380, w_058_381, w_058_382, w_058_384, w_058_385, w_058_390, w_058_391, w_058_392, w_058_393, w_058_396, w_058_397, w_058_400, w_058_402, w_058_403, w_058_406, w_058_407, w_058_408, w_058_409, w_058_411, w_058_412, w_058_415, w_058_416, w_058_417, w_058_419, w_058_420, w_058_421, w_058_422, w_058_423, w_058_424, w_058_425, w_058_427, w_058_428, w_058_429, w_058_430, w_058_433, w_058_434, w_058_435, w_058_436, w_058_438, w_058_439, w_058_440, w_058_442, w_058_443, w_058_444, w_058_445, w_058_446, w_058_447, w_058_448, w_058_449, w_058_450, w_058_451, w_058_453, w_058_455, w_058_456, w_058_457, w_058_458, w_058_460, w_058_461, w_058_462, w_058_463, w_058_465, w_058_467, w_058_468, w_058_469, w_058_470, w_058_471, w_058_472, w_058_473, w_058_474, w_058_475, w_058_476, w_058_477, w_058_478, w_058_479, w_058_480, w_058_481, w_058_482, w_058_483, w_058_484, w_058_486, w_058_487, w_058_489, w_058_490, w_058_491, w_058_492, w_058_493, w_058_494, w_058_495, w_058_497, w_058_498, w_058_499, w_058_500, w_058_501, w_058_503, w_058_504, w_058_507, w_058_508, w_058_509, w_058_512, w_058_514, w_058_515, w_058_518, w_058_519, w_058_520, w_058_523, w_058_524, w_058_525, w_058_526, w_058_527, w_058_528, w_058_529, w_058_532, w_058_536, w_058_538, w_058_539, w_058_541, w_058_543, w_058_545, w_058_546, w_058_548, w_058_549, w_058_551, w_058_552, w_058_553, w_058_554, w_058_556, w_058_557, w_058_559, w_058_560, w_058_561, w_058_562, w_058_563, w_058_564, w_058_567, w_058_568, w_058_569, w_058_570, w_058_571, w_058_573, w_058_574, w_058_575, w_058_576, w_058_577, w_058_578, w_058_579, w_058_580, w_058_581, w_058_582, w_058_583, w_058_584, w_058_585, w_058_586, w_058_587, w_058_588, w_058_589, w_058_590, w_058_591, w_058_593, w_058_594, w_058_596, w_058_597, w_058_598, w_058_600, w_058_601, w_058_602, w_058_603, w_058_604, w_058_605, w_058_606, w_058_607, w_058_608, w_058_609, w_058_610, w_058_611, w_058_613, w_058_615, w_058_618, w_058_620, w_058_621, w_058_622, w_058_623, w_058_624, w_058_625, w_058_626, w_058_627, w_058_628, w_058_630, w_058_631, w_058_632, w_058_633, w_058_634, w_058_635, w_058_637, w_058_638, w_058_639, w_058_640, w_058_641, w_058_642, w_058_643, w_058_644, w_058_645, w_058_646, w_058_647, w_058_648, w_058_649, w_058_650, w_058_651, w_058_652, w_058_653, w_058_654, w_058_655, w_058_656, w_058_657, w_058_658, w_058_659, w_058_661, w_058_662, w_058_663, w_058_664, w_058_665, w_058_668, w_058_669, w_058_670, w_058_671, w_058_672, w_058_673, w_058_675, w_058_676, w_058_678, w_058_680, w_058_681, w_058_684, w_058_685, w_058_686, w_058_688, w_058_689, w_058_691, w_058_692, w_058_693, w_058_694, w_058_697, w_058_698, w_058_699, w_058_700, w_058_701, w_058_702, w_058_703, w_058_704, w_058_705, w_058_706, w_058_707, w_058_708, w_058_710, w_058_711, w_058_712, w_058_714, w_058_715, w_058_716, w_058_717, w_058_718, w_058_720, w_058_721, w_058_723, w_058_724, w_058_725, w_058_726, w_058_727, w_058_729, w_058_730, w_058_731, w_058_734, w_058_736, w_058_737, w_058_738, w_058_741, w_058_744, w_058_747, w_058_748, w_058_749, w_058_750, w_058_751, w_058_752, w_058_753, w_058_757, w_058_760, w_058_761, w_058_763, w_058_764, w_058_766, w_058_768, w_058_770, w_058_771, w_058_772, w_058_773, w_058_776, w_058_777, w_058_778, w_058_779, w_058_780, w_058_781, w_058_783, w_058_785, w_058_786, w_058_787, w_058_789, w_058_790, w_058_791, w_058_793, w_058_797, w_058_798, w_058_799, w_058_800, w_058_802, w_058_803, w_058_804, w_058_805, w_058_808, w_058_809, w_058_810, w_058_811, w_058_812, w_058_813, w_058_814, w_058_815, w_058_817, w_058_818, w_058_819, w_058_823, w_058_824, w_058_825, w_058_826, w_058_828, w_058_829, w_058_830, w_058_831, w_058_832, w_058_833, w_058_834, w_058_835, w_058_836, w_058_837, w_058_838, w_058_840, w_058_841, w_058_842, w_058_843, w_058_845, w_058_846, w_058_847, w_058_848, w_058_849, w_058_850, w_058_851, w_058_855, w_058_857, w_058_858, w_058_859, w_058_860, w_058_861, w_058_862, w_058_863, w_058_864, w_058_866, w_058_869, w_058_870, w_058_871, w_058_872, w_058_873, w_058_874, w_058_875, w_058_876, w_058_877, w_058_878, w_058_879, w_058_880, w_058_881, w_058_882, w_058_883, w_058_884, w_058_885, w_058_888, w_058_889, w_058_890, w_058_891, w_058_892, w_058_893, w_058_894, w_058_895, w_058_896, w_058_897, w_058_898, w_058_899, w_058_900, w_058_901, w_058_902, w_058_905, w_058_906, w_058_907, w_058_908, w_058_909, w_058_910, w_058_911, w_058_912, w_058_913, w_058_914, w_058_916, w_058_917, w_058_919, w_058_920, w_058_921, w_058_922, w_058_923, w_058_924, w_058_926, w_058_927, w_058_928, w_058_930, w_058_931, w_058_932, w_058_933, w_058_936, w_058_937, w_058_938, w_058_939, w_058_940, w_058_941, w_058_942, w_058_943, w_058_945, w_058_946, w_058_947, w_058_949, w_058_950, w_058_951, w_058_952, w_058_954, w_058_955, w_058_956, w_058_957, w_058_958, w_058_959, w_058_960, w_058_961, w_058_964, w_058_965, w_058_966, w_058_968, w_058_969, w_058_970, w_058_971, w_058_972, w_058_974, w_058_975, w_058_977, w_058_980, w_058_981, w_058_982, w_058_985, w_058_990, w_058_991, w_058_993, w_058_995, w_058_996, w_058_997, w_058_1000, w_058_1002, w_058_1003, w_058_1004, w_058_1008, w_058_1009, w_058_1010, w_058_1011, w_058_1012, w_058_1013, w_058_1014, w_058_1016, w_058_1017, w_058_1018, w_058_1019, w_058_1020, w_058_1021, w_058_1022, w_058_1023, w_058_1024, w_058_1025, w_058_1027, w_058_1028, w_058_1029, w_058_1030, w_058_1031, w_058_1032, w_058_1033, w_058_1034, w_058_1035, w_058_1036, w_058_1037, w_058_1038, w_058_1039, w_058_1040, w_058_1041, w_058_1042, w_058_1043, w_058_1045, w_058_1048, w_058_1049, w_058_1050, w_058_1051, w_058_1053, w_058_1054, w_058_1055, w_058_1056, w_058_1059, w_058_1061, w_058_1062, w_058_1063, w_058_1064, w_058_1065, w_058_1066, w_058_1068, w_058_1070, w_058_1071, w_058_1072, w_058_1073, w_058_1074, w_058_1076, w_058_1077, w_058_1078, w_058_1079, w_058_1082, w_058_1084, w_058_1086, w_058_1087, w_058_1089, w_058_1090, w_058_1091, w_058_1092, w_058_1093, w_058_1094, w_058_1096, w_058_1098, w_058_1099, w_058_1101, w_058_1102, w_058_1103, w_058_1104, w_058_1105, w_058_1110, w_058_1111, w_058_1112, w_058_1113, w_058_1114, w_058_1115, w_058_1116, w_058_1117, w_058_1118, w_058_1120, w_058_1122, w_058_1123, w_058_1124, w_058_1125, w_058_1126, w_058_1128, w_058_1129, w_058_1130, w_058_1131, w_058_1132, w_058_1134, w_058_1135, w_058_1137, w_058_1139, w_058_1140, w_058_1141, w_058_1143, w_058_1144, w_058_1146, w_058_1147, w_058_1148, w_058_1149, w_058_1150, w_058_1151, w_058_1153, w_058_1154, w_058_1155, w_058_1156, w_058_1157, w_058_1158, w_058_1159, w_058_1160, w_058_1161, w_058_1162, w_058_1163, w_058_1165, w_058_1166, w_058_1167, w_058_1168, w_058_1169, w_058_1172, w_058_1173, w_058_1174, w_058_1175, w_058_1178, w_058_1179, w_058_1180, w_058_1181, w_058_1182, w_058_1185, w_058_1186, w_058_1187, w_058_1188, w_058_1189, w_058_1190, w_058_1191, w_058_1192, w_058_1196, w_058_1197, w_058_1198, w_058_1200, w_058_1201, w_058_1203, w_058_1204, w_058_1205, w_058_1206, w_058_1207, w_058_1208, w_058_1209, w_058_1211, w_058_1212, w_058_1213, w_058_1215, w_058_1216, w_058_1217, w_058_1218, w_058_1219, w_058_1222, w_058_1223, w_058_1224, w_058_1225, w_058_1226, w_058_1227, w_058_1228, w_058_1229, w_058_1230, w_058_1231, w_058_1232, w_058_1233, w_058_1234, w_058_1236, w_058_1238, w_058_1241, w_058_1242, w_058_1243, w_058_1244, w_058_1245, w_058_1246, w_058_1247, w_058_1249, w_058_1250, w_058_1252, w_058_1253, w_058_1254, w_058_1255, w_058_1257, w_058_1258, w_058_1259, w_058_1261, w_058_1262, w_058_1264, w_058_1265, w_058_1266, w_058_1267, w_058_1268, w_058_1269, w_058_1271, w_058_1272, w_058_1275, w_058_1277, w_058_1279, w_058_1280, w_058_1282, w_058_1283, w_058_1284, w_058_1285, w_058_1286, w_058_1287, w_058_1288, w_058_1290, w_058_1293, w_058_1294, w_058_1295, w_058_1296, w_058_1297, w_058_1298, w_058_1300, w_058_1301, w_058_1303, w_058_1304, w_058_1305, w_058_1306, w_058_1307, w_058_1308, w_058_1309, w_058_1313, w_058_1314, w_058_1315, w_058_1318, w_058_1319, w_058_1321, w_058_1322, w_058_1323, w_058_1326, w_058_1327, w_058_1329, w_058_1331, w_058_1334, w_058_1335, w_058_1336, w_058_1338, w_058_1339, w_058_1341, w_058_1342, w_058_1343, w_058_1344, w_058_1345, w_058_1346, w_058_1348, w_058_1349, w_058_1350, w_058_1353, w_058_1354, w_058_1356, w_058_1357, w_058_1358, w_058_1360, w_058_1361, w_058_1362, w_058_1364, w_058_1365, w_058_1366, w_058_1368, w_058_1369, w_058_1370, w_058_1371, w_058_1375, w_058_1376, w_058_1377, w_058_1378, w_058_1379, w_058_1380, w_058_1381, w_058_1384, w_058_1385, w_058_1387, w_058_1388, w_058_1389, w_058_1390, w_058_1392, w_058_1393, w_058_1394, w_058_1395, w_058_1396, w_058_1398, w_058_1400, w_058_1401, w_058_1403, w_058_1404, w_058_1405, w_058_1407, w_058_1408, w_058_1409, w_058_1410, w_058_1412, w_058_1413, w_058_1414, w_058_1415, w_058_1418, w_058_1419, w_058_1420, w_058_1421, w_058_1422, w_058_1423, w_058_1424, w_058_1426, w_058_1428, w_058_1429, w_058_1430, w_058_1435, w_058_1436, w_058_1437, w_058_1438, w_058_1439, w_058_1440, w_058_1441, w_058_1442, w_058_1444, w_058_1447, w_058_1448, w_058_1451, w_058_1452, w_058_1454, w_058_1456, w_058_1458, w_058_1459, w_058_1460, w_058_1461, w_058_1462, w_058_1463, w_058_1464, w_058_1465, w_058_1466, w_058_1469, w_058_1471, w_058_1472, w_058_1473, w_058_1475, w_058_1476, w_058_1477, w_058_1478, w_058_1479, w_058_1480, w_058_1481, w_058_1482, w_058_1483, w_058_1484, w_058_1485, w_058_1486, w_058_1487, w_058_1488, w_058_1491, w_058_1492, w_058_1494, w_058_1495, w_058_1496, w_058_1500, w_058_1501, w_058_1502, w_058_1504, w_058_1505, w_058_1506, w_058_1507, w_058_1509, w_058_1511, w_058_1512, w_058_1516, w_058_1517, w_058_1518, w_058_1521, w_058_1522, w_058_1523, w_058_1525, w_058_1526, w_058_1527, w_058_1529, w_058_1531, w_058_1532, w_058_1533, w_058_1534, w_058_1536, w_058_1537, w_058_1538, w_058_1539, w_058_1543, w_058_1544, w_058_1545, w_058_1546, w_058_1547, w_058_1548, w_058_1550, w_058_1552, w_058_1553, w_058_1554, w_058_1555, w_058_1556, w_058_1559, w_058_1560, w_058_1561, w_058_1563, w_058_1564, w_058_1565, w_058_1567, w_058_1569, w_058_1570, w_058_1573, w_058_1574, w_058_1575, w_058_1576, w_058_1577, w_058_1578, w_058_1579, w_058_1581, w_058_1582, w_058_1583, w_058_1584, w_058_1585, w_058_1587, w_058_1588, w_058_1589, w_058_1591, w_058_1592, w_058_1593, w_058_1594, w_058_1595, w_058_1596, w_058_1597, w_058_1598, w_058_1599, w_058_1601, w_058_1602, w_058_1603, w_058_1604, w_058_1605, w_058_1606, w_058_1608, w_058_1609, w_058_1610, w_058_1612, w_058_1613, w_058_1614, w_058_1615, w_058_1616, w_058_1617, w_058_1618, w_058_1619, w_058_1620, w_058_1621, w_058_1622, w_058_1623, w_058_1624, w_058_1625, w_058_1626, w_058_1627, w_058_1628, w_058_1629, w_058_1631, w_058_1633, w_058_1634, w_058_1635, w_058_1636, w_058_1637, w_058_1638, w_058_1640, w_058_1641, w_058_1642, w_058_1643, w_058_1645, w_058_1646, w_058_1647, w_058_1649, w_058_1650, w_058_1651, w_058_1652, w_058_1653, w_058_1655, w_058_1657, w_058_1658, w_058_1659, w_058_1660, w_058_1661, w_058_1662, w_058_1663, w_058_1664, w_058_1665, w_058_1666, w_058_1667, w_058_1669, w_058_1671, w_058_1677, w_058_1678, w_058_1680, w_058_1681, w_058_1683, w_058_1684, w_058_1685, w_058_1686, w_058_1688, w_058_1690, w_058_1691, w_058_1692, w_058_1695, w_058_1696, w_058_1699, w_058_1700, w_058_1702, w_058_1703, w_058_1704, w_058_1705, w_058_1707, w_058_1708, w_058_1710, w_058_1711, w_058_1712, w_058_1713, w_058_1714, w_058_1715, w_058_1716, w_058_1717, w_058_1718, w_058_1721, w_058_1722, w_058_1723, w_058_1726, w_058_1727, w_058_1729, w_058_1730, w_058_1731, w_058_1732, w_058_1733, w_058_1734, w_058_1735, w_058_1736, w_058_1738, w_058_1740, w_058_1742, w_058_1743, w_058_1745, w_058_1746, w_058_1747, w_058_1748, w_058_1749, w_058_1751, w_058_1755, w_058_1757, w_058_1758, w_058_1760, w_058_1761, w_058_1762, w_058_1763, w_058_1766, w_058_1767, w_058_1768, w_058_1772, w_058_1773, w_058_1774, w_058_1775, w_058_1776, w_058_1777, w_058_1778, w_058_1780, w_058_1782, w_058_1783, w_058_1784, w_058_1785, w_058_1787, w_058_1788, w_058_1789, w_058_1790, w_058_1791, w_058_1792, w_058_1793, w_058_1794, w_058_1797, w_058_1798, w_058_1799, w_058_1805, w_058_1806, w_058_1807, w_058_1808, w_058_1809, w_058_1810, w_058_1811, w_058_1812, w_058_1813, w_058_1814, w_058_1815, w_058_1817, w_058_1818, w_058_1819, w_058_1820, w_058_1822, w_058_1823, w_058_1824, w_058_1825, w_058_1826, w_058_1827, w_058_1828, w_058_1829, w_058_1830, w_058_1832, w_058_1834, w_058_1835, w_058_1838, w_058_1839, w_058_1841, w_058_1843, w_058_1845, w_058_1848, w_058_1852, w_058_1853, w_058_1854, w_058_1856, w_058_1857, w_058_1858, w_058_1859, w_058_1860, w_058_1861, w_058_1862, w_058_1863, w_058_1864, w_058_1865, w_058_1867, w_058_1868, w_058_1871, w_058_1872, w_058_1873, w_058_1875, w_058_1876, w_058_1877, w_058_1878, w_058_1879, w_058_1880, w_058_1881, w_058_1882, w_058_1883, w_058_1885, w_058_1887, w_058_1889, w_058_1891, w_058_1893, w_058_1894, w_058_1895, w_058_1896, w_058_1897, w_058_1900, w_058_1901, w_058_1902, w_058_1903, w_058_1904, w_058_1905, w_058_1906, w_058_1907, w_058_1908, w_058_1910, w_058_1911, w_058_1912, w_058_1916, w_058_1917, w_058_1918, w_058_1919, w_058_1920, w_058_1921, w_058_1922, w_058_1923, w_058_1924, w_058_1926, w_058_1928, w_058_1929, w_058_1931, w_058_1932, w_058_1934, w_058_1935, w_058_1936, w_058_1938, w_058_1939, w_058_1943, w_058_1944, w_058_1945, w_058_1946, w_058_1947, w_058_1948, w_058_1950, w_058_1951, w_058_1953, w_058_1954, w_058_1955, w_058_1956, w_058_1957, w_058_1959, w_058_1960, w_058_1962, w_058_1963, w_058_1964, w_058_1965, w_058_1967, w_058_1968, w_058_1969, w_058_1972, w_058_1973, w_058_1974, w_058_1975, w_058_1977, w_058_1978, w_058_1979, w_058_1980, w_058_1981, w_058_1982, w_058_1983, w_058_1985, w_058_1986, w_058_1987, w_058_1989, w_058_1990, w_058_1991, w_058_1992, w_058_1993, w_058_1994, w_058_1995, w_058_1996, w_058_1997, w_058_1998, w_058_1999, w_058_2000, w_058_2001, w_058_2002, w_058_2003, w_058_2006, w_058_2008, w_058_2010, w_058_2011, w_058_2012, w_058_2014, w_058_2015, w_058_2016, w_058_2017, w_058_2018, w_058_2019, w_058_2020, w_058_2021, w_058_2023, w_058_2024, w_058_2026, w_058_2027, w_058_2028, w_058_2030, w_058_2031, w_058_2033, w_058_2034, w_058_2035, w_058_2036, w_058_2037, w_058_2038, w_058_2039, w_058_2040, w_058_2041, w_058_2042, w_058_2043, w_058_2044, w_058_2045, w_058_2046, w_058_2047, w_058_2048, w_058_2051, w_058_2054, w_058_2055, w_058_2056, w_058_2057, w_058_2059, w_058_2060, w_058_2062, w_058_2063, w_058_2064, w_058_2065, w_058_2068, w_058_2070, w_058_2072, w_058_2073, w_058_2075, w_058_2076, w_058_2077, w_058_2079, w_058_2080, w_058_2083, w_058_2084, w_058_2085, w_058_2086, w_058_2088, w_058_2089, w_058_2090, w_058_2091, w_058_2092, w_058_2094, w_058_2095, w_058_2096, w_058_2099, w_058_2100, w_058_2102, w_058_2103, w_058_2105, w_058_2106, w_058_2107, w_058_2108, w_058_2109, w_058_2110, w_058_2111, w_058_2112, w_058_2113, w_058_2114, w_058_2115, w_058_2116, w_058_2117, w_058_2119, w_058_2120, w_058_2123, w_058_2124, w_058_2126, w_058_2127, w_058_2128, w_058_2129, w_058_2130, w_058_2131, w_058_2132, w_058_2133, w_058_2135, w_058_2139, w_058_2141, w_058_2142, w_058_2143, w_058_2144, w_058_2145, w_058_2146, w_058_2147, w_058_2148, w_058_2150, w_058_2151, w_058_2152, w_058_2154, w_058_2155, w_058_2156, w_058_2158, w_058_2160, w_058_2161, w_058_2162, w_058_2163, w_058_2164, w_058_2166, w_058_2167, w_058_2169, w_058_2172, w_058_2173, w_058_2174, w_058_2175, w_058_2176, w_058_2177, w_058_2178, w_058_2180, w_058_2181, w_058_2182, w_058_2183, w_058_2185, w_058_2186, w_058_2187, w_058_2188, w_058_2190, w_058_2192, w_058_2194, w_058_2195, w_058_2196, w_058_2198, w_058_2199, w_058_2200, w_058_2201, w_058_2202, w_058_2203, w_058_2204, w_058_2205, w_058_2206, w_058_2207, w_058_2208, w_058_2209, w_058_2210, w_058_2211, w_058_2212, w_058_2214, w_058_2215, w_058_2217, w_058_2219, w_058_2220, w_058_2221, w_058_2222, w_058_2223, w_058_2224, w_058_2225, w_058_2226, w_058_2227, w_058_2228, w_058_2229, w_058_2230, w_058_2231, w_058_2233, w_058_2236, w_058_2238, w_058_2239, w_058_2240, w_058_2241, w_058_2243, w_058_2244, w_058_2245, w_058_2246, w_058_2247, w_058_2248, w_058_2249, w_058_2251, w_058_2253, w_058_2254, w_058_2255, w_058_2256, w_058_2258, w_058_2259, w_058_2260, w_058_2261, w_058_2262, w_058_2264, w_058_2265, w_058_2267, w_058_2268, w_058_2270, w_058_2271, w_058_2273, w_058_2274, w_058_2275, w_058_2276, w_058_2277, w_058_2278, w_058_2280, w_058_2281, w_058_2282, w_058_2283, w_058_2284, w_058_2285, w_058_2287, w_058_2290, w_058_2291, w_058_2292, w_058_2293, w_058_2294, w_058_2295, w_058_2296, w_058_2297, w_058_2298, w_058_2299, w_058_2300, w_058_2301, w_058_2303, w_058_2305, w_058_2306, w_058_2307, w_058_2308, w_058_2310, w_058_2311, w_058_2312, w_058_2313, w_058_2314, w_058_2316, w_058_2317, w_058_2318, w_058_2321, w_058_2323, w_058_2324, w_058_2325, w_058_2326, w_058_2327, w_058_2330, w_058_2331, w_058_2332, w_058_2334, w_058_2335, w_058_2336, w_058_2338, w_058_2340, w_058_2341, w_058_2343, w_058_2345, w_058_2346, w_058_2347, w_058_2348, w_058_2349, w_058_2350, w_058_2352, w_058_2353, w_058_2354, w_058_2356, w_058_2357, w_058_2358, w_058_2359, w_058_2361, w_058_2363, w_058_2364, w_058_2365, w_058_2366, w_058_2367, w_058_2368, w_058_2369, w_058_2371, w_058_2372, w_058_2375, w_058_2377, w_058_2378, w_058_2382, w_058_2383, w_058_2384, w_058_2385, w_058_2386, w_058_2387, w_058_2388, w_058_2389, w_058_2390, w_058_2391, w_058_2393, w_058_2394, w_058_2395, w_058_2396, w_058_2397, w_058_2399, w_058_2400, w_058_2402, w_058_2403, w_058_2406, w_058_2407, w_058_2408, w_058_2411, w_058_2412, w_058_2413, w_058_2415, w_058_2417, w_058_2418, w_058_2419, w_058_2420, w_058_2421, w_058_2422, w_058_2423, w_058_2424, w_058_2426, w_058_2428, w_058_2429, w_058_2430, w_058_2431, w_058_2432, w_058_2433, w_058_2434, w_058_2435, w_058_2437, w_058_2439, w_058_2440, w_058_2441, w_058_2444, w_058_2445, w_058_2446, w_058_2449, w_058_2450, w_058_2451, w_058_2452, w_058_2453, w_058_2454, w_058_2455, w_058_2457, w_058_2459, w_058_2460, w_058_2461, w_058_2462, w_058_2463, w_058_2464, w_058_2465, w_058_2466, w_058_2467, w_058_2469, w_058_2470, w_058_2471, w_058_2472, w_058_2473, w_058_2474, w_058_2475, w_058_2477, w_058_2479, w_058_2482, w_058_2483, w_058_2484, w_058_2485, w_058_2487, w_058_2488, w_058_2489, w_058_2490, w_058_2491, w_058_2492, w_058_2494, w_058_2495, w_058_2496, w_058_2497, w_058_2498, w_058_2500, w_058_2501, w_058_2502, w_058_2505, w_058_2507, w_058_2508, w_058_2509, w_058_2510, w_058_2511, w_058_2512, w_058_2513, w_058_2514, w_058_2515, w_058_2517, w_058_2518, w_058_2519, w_058_2520, w_058_2522, w_058_2523, w_058_2526, w_058_2528, w_058_2529, w_058_2530, w_058_2531, w_058_2533, w_058_2535, w_058_2536, w_058_2538, w_058_2540, w_058_2542, w_058_2543, w_058_2545, w_058_2546, w_058_2547, w_058_2550, w_058_2551, w_058_2552, w_058_2553, w_058_2554, w_058_2556, w_058_2557, w_058_2558, w_058_2559, w_058_2560, w_058_2561, w_058_2564, w_058_2568, w_058_2571, w_058_2572, w_058_2573, w_058_2574, w_058_2575, w_058_2577, w_058_2581, w_058_2582, w_058_2586, w_058_2587, w_058_2588, w_058_2589, w_058_2590, w_058_2591, w_058_2595, w_058_2596, w_058_2597, w_058_2598, w_058_2600, w_058_2601, w_058_2602, w_058_2603, w_058_2604, w_058_2606, w_058_2607, w_058_2608, w_058_2609, w_058_2610, w_058_2611, w_058_2612, w_058_2613, w_058_2614, w_058_2615, w_058_2616, w_058_2617, w_058_2619, w_058_2620, w_058_2621, w_058_2622, w_058_2623, w_058_2624, w_058_2625, w_058_2626, w_058_2627, w_058_2628, w_058_2630, w_058_2632, w_058_2633, w_058_2634, w_058_2635, w_058_2636, w_058_2637, w_058_2638, w_058_2639, w_058_2642, w_058_2643, w_058_2645, w_058_2646, w_058_2647, w_058_2648, w_058_2650, w_058_2651, w_058_2652, w_058_2654, w_058_2655, w_058_2656, w_058_2659, w_058_2660, w_058_2661, w_058_2662, w_058_2663, w_058_2664, w_058_2665, w_058_2666, w_058_2667, w_058_2670, w_058_2671, w_058_2672, w_058_2673, w_058_2674, w_058_2675, w_058_2676, w_058_2677, w_058_2678, w_058_2679, w_058_2681, w_058_2683, w_058_2684, w_058_2685, w_058_2686, w_058_2687, w_058_2688, w_058_2690, w_058_2692, w_058_2693, w_058_2697, w_058_2698, w_058_2699, w_058_2700, w_058_2701, w_058_2702, w_058_2703, w_058_2705, w_058_2706, w_058_2707, w_058_2708, w_058_2709, w_058_2710, w_058_2711, w_058_2712, w_058_2713, w_058_2714, w_058_2715, w_058_2717, w_058_2718, w_058_2719, w_058_2720, w_058_2721, w_058_2723, w_058_2724, w_058_2725, w_058_2727, w_058_2728, w_058_2729, w_058_2730, w_058_2732, w_058_2734, w_058_2735, w_058_2736, w_058_2738, w_058_2739, w_058_2741, w_058_2742, w_058_2743, w_058_2744, w_058_2745, w_058_2746, w_058_2747, w_058_2749, w_058_2750, w_058_2751, w_058_2752, w_058_2753, w_058_2754, w_058_2755, w_058_2756, w_058_2757, w_058_2758, w_058_2759, w_058_2760, w_058_2761, w_058_2762, w_058_2763, w_058_2766, w_058_2767, w_058_2768, w_058_2770, w_058_2771, w_058_2772, w_058_2773, w_058_2774, w_058_2775, w_058_2778, w_058_2779, w_058_2780, w_058_2781, w_058_2782, w_058_2783, w_058_2784, w_058_2785, w_058_2786, w_058_2788, w_058_2789, w_058_2790, w_058_2791, w_058_2793, w_058_2794, w_058_2797, w_058_2799, w_058_2800, w_058_2801, w_058_2802, w_058_2804, w_058_2805, w_058_2806, w_058_2807, w_058_2808, w_058_2809, w_058_2810, w_058_2811, w_058_2812, w_058_2813, w_058_2814, w_058_2815, w_058_2816, w_058_2818, w_058_2820, w_058_2821, w_058_2822, w_058_2824, w_058_2825, w_058_2826, w_058_2828, w_058_2829, w_058_2831, w_058_2834, w_058_2835, w_058_2836, w_058_2837, w_058_2838, w_058_2840, w_058_2841, w_058_2842, w_058_2843, w_058_2844, w_058_2845, w_058_2846, w_058_2849, w_058_2850, w_058_2851, w_058_2853, w_058_2854, w_058_2855, w_058_2856, w_058_2857, w_058_2858, w_058_2859, w_058_2860, w_058_2861, w_058_2862, w_058_2863, w_058_2864, w_058_2865, w_058_2866, w_058_2867, w_058_2869, w_058_2871, w_058_2872, w_058_2873, w_058_2874, w_058_2875, w_058_2876, w_058_2877, w_058_2878, w_058_2879, w_058_2880, w_058_2881, w_058_2885, w_058_2886, w_058_2887, w_058_2888, w_058_2889, w_058_2890, w_058_2891, w_058_2892, w_058_2893, w_058_2895, w_058_2896, w_058_2897, w_058_2899, w_058_2900, w_058_2901, w_058_2902, w_058_2908, w_058_2910, w_058_2911, w_058_2913, w_058_2914, w_058_2916, w_058_2917, w_058_2918, w_058_2919, w_058_2920, w_058_2921, w_058_2922, w_058_2926, w_058_2927, w_058_2929, w_058_2930, w_058_2934, w_058_2935, w_058_2936, w_058_2937, w_058_2938, w_058_2939, w_058_2940, w_058_2941, w_058_2944, w_058_2945, w_058_2946, w_058_2947, w_058_2948, w_058_2950, w_058_2952, w_058_2953, w_058_2955, w_058_2956, w_058_2957, w_058_2958, w_058_2959, w_058_2960, w_058_2962, w_058_2963, w_058_2964, w_058_2965, w_058_2966, w_058_2967, w_058_2968, w_058_2969, w_058_2970, w_058_2971, w_058_2976, w_058_2978, w_058_2979, w_058_2980, w_058_2981, w_058_2982, w_058_2983, w_058_2984, w_058_2985, w_058_2986, w_058_2987, w_058_2990, w_058_2991, w_058_2993, w_058_2994, w_058_2995, w_058_2996, w_058_2997, w_058_2998, w_058_2999, w_058_3000, w_058_3001, w_058_3002, w_058_3006, w_058_3008, w_058_3010, w_058_3012, w_058_3013, w_058_3014, w_058_3015, w_058_3016, w_058_3017, w_058_3018, w_058_3019, w_058_3022, w_058_3023, w_058_3024, w_058_3025, w_058_3026, w_058_3031, w_058_3032, w_058_3039, w_058_3040, w_058_3042, w_058_3044, w_058_3045, w_058_3047, w_058_3051, w_058_3052, w_058_3053, w_058_3054, w_058_3057, w_058_3058, w_058_3059, w_058_3060, w_058_3061, w_058_3063, w_058_3064, w_058_3067, w_058_3069, w_058_3072, w_058_3074, w_058_3077, w_058_3078, w_058_3079, w_058_3080, w_058_3082, w_058_3083, w_058_3085, w_058_3091, w_058_3095, w_058_3096, w_058_3097, w_058_3099, w_058_3100, w_058_3101, w_058_3102, w_058_3103, w_058_3104, w_058_3105, w_058_3106, w_058_3108, w_058_3109, w_058_3110, w_058_3111, w_058_3112, w_058_3113, w_058_3116, w_058_3118, w_058_3119, w_058_3120, w_058_3123, w_058_3125, w_058_3126, w_058_3127, w_058_3129, w_058_3132, w_058_3135, w_058_3137, w_058_3138, w_058_3142, w_058_3143, w_058_3146, w_058_3148, w_058_3149, w_058_3150, w_058_3152, w_058_3153, w_058_3154, w_058_3155, w_058_3157, w_058_3159, w_058_3160, w_058_3162, w_058_3163, w_058_3166, w_058_3167, w_058_3169, w_058_3171, w_058_3172, w_058_3174, w_058_3176, w_058_3179, w_058_3180, w_058_3183, w_058_3184, w_058_3189, w_058_3190, w_058_3191, w_058_3192, w_058_3193, w_058_3198, w_058_3200, w_058_3201, w_058_3203, w_058_3205, w_058_3206, w_058_3207, w_058_3208, w_058_3209, w_058_3213, w_058_3214, w_058_3219, w_058_3220, w_058_3221, w_058_3222, w_058_3223, w_058_3224, w_058_3225, w_058_3226, w_058_3227, w_058_3228, w_058_3230, w_058_3233, w_058_3234, w_058_3236, w_058_3237, w_058_3238, w_058_3239, w_058_3240, w_058_3241, w_058_3242, w_058_3243, w_058_3244, w_058_3246, w_058_3248, w_058_3249, w_058_3250, w_058_3254, w_058_3255, w_058_3258, w_058_3262, w_058_3263, w_058_3265, w_058_3266, w_058_3270, w_058_3273, w_058_3274, w_058_3275, w_058_3276, w_058_3278, w_058_3279, w_058_3280, w_058_3281, w_058_3282, w_058_3283, w_058_3286, w_058_3287, w_058_3288, w_058_3289, w_058_3290, w_058_3291, w_058_3293, w_058_3295, w_058_3296, w_058_3297, w_058_3298, w_058_3299, w_058_3302, w_058_3303, w_058_3304, w_058_3305, w_058_3307, w_058_3308, w_058_3313, w_058_3314, w_058_3318, w_058_3319, w_058_3322, w_058_3323, w_058_3324, w_058_3325, w_058_3326, w_058_3327, w_058_3328, w_058_3329, w_058_3331, w_058_3332, w_058_3334, w_058_3335, w_058_3336, w_058_3337, w_058_3338, w_058_3339, w_058_3341, w_058_3345, w_058_3348, w_058_3349, w_058_3350, w_058_3354, w_058_3357, w_058_3360, w_058_3361, w_058_3362, w_058_3363, w_058_3364, w_058_3365, w_058_3368, w_058_3369, w_058_3371, w_058_3373, w_058_3376, w_058_3378, w_058_3379, w_058_3380, w_058_3381, w_058_3382, w_058_3383, w_058_3384, w_058_3385, w_058_3388, w_058_3389, w_058_3390, w_058_3392, w_058_3394, w_058_3395, w_058_3396, w_058_3397, w_058_3398, w_058_3399, w_058_3400, w_058_3401, w_058_3403, w_058_3404, w_058_3406, w_058_3407, w_058_3412, w_058_3414, w_058_3416, w_058_3418, w_058_3419, w_058_3421, w_058_3422, w_058_3424, w_058_3428, w_058_3429, w_058_3430, w_058_3431, w_058_3434, w_058_3436, w_058_3437, w_058_3438, w_058_3440, w_058_3442, w_058_3444, w_058_3445, w_058_3447, w_058_3448, w_058_3451, w_058_3452, w_058_3454, w_058_3455, w_058_3456, w_058_3457, w_058_3461, w_058_3463, w_058_3466, w_058_3467, w_058_3469, w_058_3470, w_058_3471, w_058_3472, w_058_3473, w_058_3474, w_058_3475, w_058_3476, w_058_3477, w_058_3478, w_058_3480, w_058_3482, w_058_3483, w_058_3484, w_058_3485;
  wire w_059_000, w_059_001, w_059_002, w_059_003, w_059_004, w_059_005, w_059_006, w_059_007, w_059_008, w_059_009, w_059_010, w_059_011, w_059_012, w_059_013, w_059_014, w_059_015, w_059_016, w_059_017, w_059_018, w_059_019, w_059_021, w_059_022, w_059_023, w_059_024, w_059_025, w_059_026, w_059_027, w_059_028, w_059_029, w_059_030, w_059_031, w_059_032, w_059_033, w_059_034, w_059_035, w_059_036, w_059_037, w_059_038, w_059_039, w_059_040, w_059_041, w_059_042, w_059_043, w_059_044, w_059_045, w_059_046, w_059_047, w_059_048, w_059_049, w_059_050, w_059_051, w_059_052, w_059_053, w_059_054, w_059_055, w_059_056, w_059_057, w_059_058, w_059_059, w_059_060, w_059_061, w_059_062, w_059_063, w_059_064, w_059_065, w_059_066, w_059_067, w_059_068, w_059_069, w_059_070, w_059_071, w_059_072, w_059_073, w_059_074, w_059_075, w_059_076, w_059_077, w_059_078, w_059_079, w_059_080, w_059_081, w_059_082, w_059_083, w_059_084, w_059_085, w_059_086, w_059_087, w_059_088, w_059_089, w_059_090, w_059_091, w_059_092, w_059_093, w_059_094, w_059_095, w_059_096, w_059_097, w_059_098, w_059_099, w_059_100, w_059_101, w_059_102, w_059_103, w_059_104, w_059_105, w_059_106, w_059_107, w_059_108, w_059_109, w_059_110, w_059_111, w_059_112, w_059_113, w_059_114, w_059_115, w_059_116, w_059_117, w_059_118, w_059_119, w_059_120, w_059_121, w_059_122, w_059_123, w_059_124, w_059_125, w_059_126, w_059_127, w_059_128, w_059_129, w_059_130, w_059_131, w_059_132, w_059_133, w_059_134, w_059_135, w_059_136, w_059_137, w_059_138, w_059_139, w_059_140, w_059_141, w_059_142, w_059_143, w_059_144, w_059_145, w_059_146, w_059_147, w_059_148, w_059_149, w_059_150, w_059_151, w_059_152, w_059_153, w_059_154, w_059_155, w_059_156, w_059_157, w_059_158, w_059_159, w_059_160, w_059_161, w_059_162, w_059_163, w_059_164, w_059_165, w_059_166, w_059_167, w_059_168, w_059_169, w_059_170, w_059_171, w_059_172, w_059_173, w_059_174, w_059_175, w_059_176, w_059_177, w_059_178, w_059_179, w_059_180, w_059_181, w_059_182, w_059_183, w_059_184, w_059_185, w_059_186, w_059_188, w_059_189, w_059_190, w_059_191, w_059_192, w_059_193, w_059_194, w_059_195, w_059_196, w_059_197, w_059_198, w_059_199, w_059_200, w_059_201, w_059_202, w_059_203, w_059_204, w_059_205, w_059_206, w_059_207, w_059_208, w_059_209, w_059_210, w_059_211, w_059_212, w_059_213, w_059_214, w_059_215, w_059_216, w_059_217, w_059_218, w_059_219, w_059_220, w_059_221, w_059_222, w_059_223, w_059_224, w_059_225, w_059_226, w_059_227, w_059_228, w_059_229, w_059_230, w_059_231, w_059_232, w_059_233, w_059_234, w_059_235, w_059_236, w_059_237, w_059_238, w_059_239, w_059_240, w_059_241, w_059_242, w_059_243, w_059_244, w_059_245, w_059_246, w_059_247, w_059_248, w_059_249, w_059_250, w_059_251, w_059_252, w_059_253, w_059_254, w_059_255, w_059_256, w_059_257, w_059_258, w_059_259, w_059_260, w_059_261, w_059_262, w_059_263, w_059_264, w_059_265, w_059_266, w_059_267, w_059_268, w_059_269, w_059_270, w_059_271, w_059_272, w_059_273, w_059_274, w_059_275, w_059_276, w_059_277, w_059_278, w_059_279, w_059_280, w_059_281, w_059_282, w_059_283, w_059_284, w_059_285, w_059_286, w_059_287, w_059_288, w_059_289, w_059_290, w_059_291, w_059_292, w_059_293, w_059_294, w_059_296, w_059_297, w_059_298, w_059_299, w_059_300, w_059_301, w_059_302, w_059_303, w_059_304, w_059_305, w_059_306, w_059_307, w_059_308, w_059_309, w_059_310, w_059_311, w_059_312, w_059_313, w_059_314, w_059_315, w_059_316, w_059_317, w_059_318, w_059_319, w_059_320, w_059_321, w_059_322, w_059_323, w_059_324, w_059_325, w_059_326, w_059_327, w_059_329, w_059_330, w_059_331, w_059_332, w_059_333, w_059_334, w_059_336, w_059_337, w_059_338, w_059_339, w_059_340, w_059_341, w_059_342, w_059_343, w_059_344, w_059_345, w_059_346, w_059_347, w_059_348, w_059_349, w_059_350, w_059_351, w_059_352, w_059_353, w_059_354, w_059_355, w_059_356, w_059_357, w_059_358, w_059_359, w_059_360, w_059_361, w_059_362, w_059_363, w_059_364, w_059_365, w_059_366, w_059_367, w_059_368, w_059_369, w_059_370, w_059_371, w_059_372, w_059_373, w_059_374, w_059_375, w_059_376, w_059_377, w_059_378, w_059_379, w_059_380, w_059_381, w_059_382, w_059_383, w_059_384, w_059_385, w_059_386, w_059_387, w_059_388, w_059_389, w_059_390, w_059_391, w_059_392, w_059_393, w_059_394, w_059_395, w_059_396, w_059_397, w_059_398, w_059_399, w_059_400, w_059_401, w_059_402, w_059_403, w_059_404, w_059_405, w_059_406, w_059_407, w_059_408, w_059_409, w_059_410, w_059_411, w_059_412, w_059_413, w_059_414, w_059_415, w_059_416, w_059_417, w_059_418, w_059_419, w_059_420, w_059_421, w_059_422, w_059_423, w_059_424, w_059_425, w_059_426, w_059_427, w_059_428, w_059_429, w_059_430, w_059_431, w_059_432, w_059_433, w_059_434, w_059_435, w_059_437, w_059_438, w_059_439, w_059_440, w_059_441, w_059_442, w_059_443, w_059_444, w_059_445, w_059_446, w_059_447, w_059_448, w_059_449, w_059_450, w_059_451, w_059_452, w_059_453, w_059_454, w_059_455, w_059_457, w_059_458, w_059_459, w_059_460, w_059_461, w_059_462, w_059_463, w_059_464, w_059_465, w_059_467, w_059_468, w_059_469, w_059_470, w_059_471, w_059_472, w_059_473, w_059_474, w_059_475, w_059_476, w_059_477, w_059_478, w_059_479, w_059_480, w_059_481, w_059_482, w_059_484, w_059_485, w_059_486, w_059_487, w_059_488, w_059_489, w_059_490, w_059_491, w_059_492, w_059_493, w_059_494, w_059_495, w_059_496, w_059_497, w_059_498, w_059_500, w_059_501, w_059_502, w_059_503, w_059_504, w_059_505, w_059_506, w_059_507, w_059_508, w_059_509, w_059_510, w_059_512, w_059_513, w_059_514, w_059_515, w_059_516, w_059_517, w_059_518, w_059_520, w_059_521, w_059_522, w_059_523, w_059_524, w_059_525, w_059_526, w_059_527, w_059_528, w_059_529, w_059_530, w_059_531, w_059_532, w_059_533, w_059_534, w_059_535, w_059_536, w_059_537, w_059_538, w_059_539, w_059_540, w_059_541, w_059_542, w_059_543, w_059_544, w_059_545, w_059_546, w_059_547, w_059_548, w_059_549, w_059_550, w_059_551, w_059_552, w_059_553, w_059_554, w_059_555, w_059_556, w_059_557, w_059_558, w_059_559, w_059_560, w_059_561, w_059_562, w_059_563, w_059_565, w_059_566, w_059_567, w_059_568, w_059_569, w_059_570, w_059_571, w_059_572, w_059_573, w_059_574, w_059_575, w_059_576, w_059_577, w_059_578, w_059_579, w_059_580, w_059_581, w_059_582, w_059_583, w_059_584, w_059_585, w_059_586, w_059_587, w_059_588, w_059_589, w_059_590, w_059_591, w_059_593, w_059_594, w_059_595, w_059_596, w_059_597, w_059_598, w_059_599, w_059_600, w_059_601, w_059_602, w_059_603, w_059_604, w_059_605, w_059_606, w_059_607, w_059_608, w_059_609, w_059_610, w_059_611, w_059_612, w_059_613, w_059_614, w_059_615, w_059_616, w_059_617, w_059_618, w_059_619, w_059_620, w_059_621, w_059_622, w_059_623, w_059_624, w_059_625, w_059_626, w_059_627, w_059_628, w_059_629, w_059_630, w_059_631, w_059_632, w_059_633, w_059_634, w_059_635, w_059_636, w_059_637, w_059_638, w_059_639, w_059_640, w_059_641, w_059_642, w_059_643, w_059_644, w_059_645, w_059_646, w_059_647, w_059_648, w_059_649, w_059_650, w_059_651, w_059_652, w_059_653, w_059_654, w_059_655, w_059_656, w_059_657, w_059_658, w_059_659, w_059_660, w_059_661, w_059_662, w_059_663, w_059_664, w_059_665, w_059_666, w_059_667, w_059_668, w_059_669, w_059_670, w_059_671, w_059_672, w_059_673, w_059_674, w_059_675, w_059_676, w_059_677, w_059_678, w_059_679, w_059_680, w_059_681, w_059_682, w_059_683, w_059_684, w_059_685, w_059_686, w_059_687, w_059_688, w_059_689, w_059_690, w_059_691, w_059_692, w_059_693, w_059_694, w_059_695, w_059_696, w_059_697, w_059_698, w_059_699, w_059_700, w_059_701, w_059_702, w_059_703, w_059_704, w_059_705, w_059_706, w_059_707, w_059_708, w_059_709, w_059_710, w_059_711, w_059_712, w_059_713, w_059_714, w_059_715, w_059_716, w_059_717, w_059_718, w_059_719, w_059_720, w_059_721, w_059_722, w_059_723, w_059_724, w_059_725, w_059_726, w_059_727, w_059_728, w_059_729, w_059_730, w_059_731, w_059_732, w_059_733, w_059_734, w_059_736, w_059_737, w_059_738, w_059_739, w_059_740, w_059_741, w_059_742, w_059_743, w_059_744, w_059_745, w_059_746, w_059_747, w_059_748, w_059_749, w_059_750, w_059_751, w_059_752, w_059_755, w_059_756, w_059_758, w_059_759, w_059_760, w_059_761, w_059_762, w_059_763, w_059_764, w_059_765, w_059_766, w_059_767, w_059_768, w_059_769, w_059_770, w_059_771, w_059_773, w_059_774, w_059_775, w_059_776, w_059_777, w_059_778, w_059_779, w_059_781, w_059_782, w_059_783, w_059_784, w_059_785, w_059_786, w_059_787, w_059_788, w_059_789, w_059_790, w_059_791, w_059_792, w_059_793, w_059_794, w_059_795, w_059_796, w_059_797, w_059_798, w_059_799, w_059_800, w_059_801, w_059_802, w_059_803, w_059_804, w_059_805, w_059_806, w_059_807, w_059_808, w_059_809, w_059_811, w_059_812, w_059_813, w_059_814, w_059_815, w_059_816, w_059_817, w_059_818, w_059_819, w_059_820, w_059_821, w_059_822, w_059_823, w_059_824, w_059_825, w_059_826, w_059_827, w_059_828, w_059_829, w_059_830, w_059_831, w_059_832, w_059_833, w_059_835, w_059_836, w_059_837, w_059_838, w_059_839, w_059_840, w_059_841, w_059_842, w_059_843, w_059_844, w_059_845, w_059_846, w_059_847, w_059_848, w_059_849, w_059_850, w_059_851, w_059_852, w_059_853, w_059_854, w_059_855, w_059_856, w_059_857, w_059_858, w_059_859, w_059_860, w_059_861, w_059_862, w_059_863, w_059_864, w_059_865, w_059_866, w_059_867, w_059_868, w_059_869, w_059_870, w_059_871, w_059_872, w_059_873, w_059_874, w_059_875, w_059_876, w_059_877, w_059_878, w_059_879, w_059_880, w_059_881, w_059_882, w_059_883, w_059_884, w_059_885, w_059_886, w_059_887, w_059_888, w_059_889, w_059_890, w_059_891, w_059_892, w_059_893, w_059_894, w_059_895, w_059_896, w_059_898, w_059_899, w_059_900, w_059_901, w_059_902, w_059_903, w_059_904, w_059_905, w_059_906, w_059_907, w_059_908, w_059_909, w_059_910, w_059_911, w_059_912, w_059_913, w_059_914, w_059_915, w_059_916, w_059_917, w_059_918, w_059_919, w_059_920, w_059_921, w_059_922, w_059_923, w_059_924, w_059_925, w_059_926, w_059_927, w_059_928, w_059_929, w_059_930, w_059_931, w_059_932, w_059_933, w_059_934, w_059_935, w_059_936, w_059_937, w_059_938, w_059_939, w_059_940, w_059_941, w_059_942, w_059_943, w_059_944, w_059_945, w_059_946, w_059_947, w_059_948, w_059_949, w_059_950, w_059_951, w_059_952, w_059_953, w_059_954, w_059_955, w_059_956, w_059_958, w_059_959, w_059_960, w_059_961, w_059_962, w_059_963, w_059_964, w_059_965, w_059_966, w_059_967, w_059_968, w_059_969, w_059_970, w_059_971, w_059_972, w_059_973, w_059_974, w_059_975, w_059_976, w_059_977, w_059_978, w_059_979, w_059_980, w_059_981, w_059_982, w_059_983, w_059_984, w_059_985, w_059_986, w_059_987, w_059_988, w_059_989, w_059_990, w_059_991, w_059_992, w_059_993, w_059_994, w_059_995, w_059_996, w_059_997, w_059_998, w_059_999, w_059_1000, w_059_1001, w_059_1003, w_059_1004, w_059_1005, w_059_1006, w_059_1007, w_059_1008, w_059_1009, w_059_1010, w_059_1011, w_059_1012, w_059_1013, w_059_1014, w_059_1016, w_059_1017, w_059_1018, w_059_1019, w_059_1020, w_059_1021, w_059_1022, w_059_1023, w_059_1024, w_059_1025, w_059_1026, w_059_1027, w_059_1028, w_059_1029, w_059_1030, w_059_1031, w_059_1032, w_059_1033, w_059_1034, w_059_1035, w_059_1036, w_059_1037, w_059_1038, w_059_1039, w_059_1040, w_059_1041, w_059_1042, w_059_1043, w_059_1044, w_059_1045, w_059_1046, w_059_1047, w_059_1048, w_059_1049, w_059_1050, w_059_1051, w_059_1052, w_059_1053, w_059_1054, w_059_1055, w_059_1056, w_059_1057, w_059_1058, w_059_1059, w_059_1060, w_059_1061, w_059_1062, w_059_1063, w_059_1064, w_059_1065, w_059_1066, w_059_1067, w_059_1068, w_059_1069, w_059_1070, w_059_1071, w_059_1072, w_059_1073, w_059_1074, w_059_1075, w_059_1076, w_059_1077, w_059_1078, w_059_1079, w_059_1080, w_059_1081, w_059_1082, w_059_1083, w_059_1084, w_059_1085, w_059_1086, w_059_1087, w_059_1089, w_059_1091, w_059_1092, w_059_1094, w_059_1095, w_059_1096, w_059_1097, w_059_1098, w_059_1099, w_059_1100, w_059_1101, w_059_1102, w_059_1103, w_059_1104, w_059_1105, w_059_1106, w_059_1107, w_059_1108, w_059_1109, w_059_1111, w_059_1112, w_059_1113, w_059_1115, w_059_1116, w_059_1117, w_059_1118, w_059_1119, w_059_1120, w_059_1121, w_059_1122, w_059_1123, w_059_1124, w_059_1125, w_059_1127, w_059_1128, w_059_1129, w_059_1130, w_059_1131, w_059_1132, w_059_1133, w_059_1134, w_059_1135, w_059_1136, w_059_1137, w_059_1138, w_059_1140, w_059_1141, w_059_1142, w_059_1143, w_059_1144, w_059_1145, w_059_1146, w_059_1148, w_059_1149, w_059_1150, w_059_1151, w_059_1152, w_059_1153, w_059_1154, w_059_1155, w_059_1156, w_059_1157, w_059_1158, w_059_1159, w_059_1160, w_059_1161, w_059_1163, w_059_1164, w_059_1165, w_059_1166, w_059_1167, w_059_1168, w_059_1169, w_059_1170, w_059_1171, w_059_1172, w_059_1173, w_059_1174, w_059_1177, w_059_1178, w_059_1179, w_059_1180, w_059_1181, w_059_1182, w_059_1183, w_059_1184, w_059_1185, w_059_1186, w_059_1189, w_059_1190, w_059_1191, w_059_1192, w_059_1193, w_059_1195, w_059_1196, w_059_1197, w_059_1198, w_059_1199, w_059_1200, w_059_1201, w_059_1202, w_059_1203, w_059_1204, w_059_1205, w_059_1206, w_059_1207, w_059_1208, w_059_1209, w_059_1210, w_059_1211, w_059_1212, w_059_1213, w_059_1214, w_059_1215, w_059_1216, w_059_1217, w_059_1218, w_059_1219, w_059_1220, w_059_1221, w_059_1222, w_059_1223, w_059_1224, w_059_1225, w_059_1226, w_059_1227, w_059_1228, w_059_1230, w_059_1231, w_059_1232, w_059_1233, w_059_1234, w_059_1235, w_059_1236, w_059_1237, w_059_1238, w_059_1239, w_059_1240, w_059_1241, w_059_1242, w_059_1243, w_059_1244, w_059_1245, w_059_1246, w_059_1247, w_059_1248, w_059_1249, w_059_1250, w_059_1251, w_059_1252, w_059_1253, w_059_1254, w_059_1255, w_059_1256, w_059_1257, w_059_1258, w_059_1259, w_059_1260, w_059_1261, w_059_1262, w_059_1263, w_059_1264, w_059_1265, w_059_1266, w_059_1267, w_059_1268, w_059_1269, w_059_1270, w_059_1271, w_059_1272, w_059_1273, w_059_1274, w_059_1275, w_059_1276;
  wire w_060_000, w_060_002, w_060_003, w_060_004, w_060_007, w_060_009, w_060_011, w_060_013, w_060_017, w_060_018, w_060_019, w_060_020, w_060_021, w_060_023, w_060_024, w_060_025, w_060_026, w_060_027, w_060_029, w_060_030, w_060_031, w_060_032, w_060_033, w_060_034, w_060_035, w_060_036, w_060_040, w_060_041, w_060_042, w_060_043, w_060_044, w_060_045, w_060_046, w_060_048, w_060_049, w_060_050, w_060_051, w_060_052, w_060_053, w_060_054, w_060_056, w_060_057, w_060_058, w_060_059, w_060_060, w_060_061, w_060_062, w_060_063, w_060_064, w_060_065, w_060_066, w_060_067, w_060_070, w_060_073, w_060_074, w_060_075, w_060_076, w_060_077, w_060_078, w_060_079, w_060_080, w_060_081, w_060_082, w_060_083, w_060_084, w_060_086, w_060_087, w_060_088, w_060_089, w_060_090, w_060_091, w_060_092, w_060_093, w_060_094, w_060_095, w_060_096, w_060_097, w_060_098, w_060_099, w_060_100, w_060_101, w_060_102, w_060_103, w_060_104, w_060_105, w_060_106, w_060_107, w_060_108, w_060_109, w_060_110, w_060_111, w_060_112, w_060_113, w_060_114, w_060_115, w_060_116, w_060_117, w_060_118, w_060_119, w_060_120, w_060_121, w_060_122, w_060_123, w_060_125, w_060_127, w_060_128, w_060_129, w_060_130, w_060_132, w_060_133, w_060_134, w_060_135, w_060_137, w_060_138, w_060_139, w_060_140, w_060_141, w_060_142, w_060_145, w_060_146, w_060_147, w_060_148, w_060_149, w_060_150, w_060_151, w_060_152, w_060_153, w_060_154, w_060_155, w_060_156, w_060_158, w_060_159, w_060_160, w_060_161, w_060_163, w_060_164, w_060_165, w_060_166, w_060_167, w_060_168, w_060_169, w_060_170, w_060_171, w_060_172, w_060_173, w_060_174, w_060_175, w_060_176, w_060_177, w_060_180, w_060_181, w_060_182, w_060_183, w_060_184, w_060_185, w_060_187, w_060_189, w_060_190, w_060_191, w_060_192, w_060_193, w_060_195, w_060_196, w_060_197, w_060_198, w_060_199, w_060_200, w_060_201, w_060_202, w_060_203, w_060_204, w_060_205, w_060_206, w_060_207, w_060_208, w_060_209, w_060_210, w_060_211, w_060_213, w_060_214, w_060_215, w_060_216, w_060_217, w_060_218, w_060_219, w_060_220, w_060_221, w_060_222, w_060_223, w_060_224, w_060_225, w_060_226, w_060_227, w_060_228, w_060_229, w_060_230, w_060_231, w_060_232, w_060_235, w_060_236, w_060_237, w_060_238, w_060_239, w_060_240, w_060_241, w_060_242, w_060_244, w_060_245, w_060_246, w_060_249, w_060_251, w_060_253, w_060_254, w_060_256, w_060_257, w_060_258, w_060_259, w_060_260, w_060_261, w_060_262, w_060_263, w_060_264, w_060_265, w_060_266, w_060_267, w_060_268, w_060_269, w_060_270, w_060_271, w_060_272, w_060_273, w_060_276, w_060_277, w_060_279, w_060_280, w_060_281, w_060_283, w_060_284, w_060_285, w_060_286, w_060_287, w_060_288, w_060_289, w_060_290, w_060_291, w_060_292, w_060_294, w_060_295, w_060_296, w_060_297, w_060_298, w_060_299, w_060_300, w_060_301, w_060_302, w_060_304, w_060_306, w_060_307, w_060_308, w_060_309, w_060_310, w_060_311, w_060_313, w_060_314, w_060_315, w_060_316, w_060_317, w_060_318, w_060_319, w_060_321, w_060_322, w_060_324, w_060_325, w_060_326, w_060_327, w_060_328, w_060_329, w_060_331, w_060_332, w_060_333, w_060_334, w_060_335, w_060_336, w_060_337, w_060_339, w_060_340, w_060_341, w_060_342, w_060_343, w_060_344, w_060_345, w_060_346, w_060_347, w_060_348, w_060_349, w_060_350, w_060_351, w_060_352, w_060_353, w_060_354, w_060_355, w_060_356, w_060_357, w_060_358, w_060_359, w_060_360, w_060_361, w_060_362, w_060_363, w_060_364, w_060_366, w_060_367, w_060_368, w_060_369, w_060_370, w_060_371, w_060_372, w_060_373, w_060_375, w_060_377, w_060_378, w_060_379, w_060_380, w_060_381, w_060_382, w_060_383, w_060_384, w_060_385, w_060_386, w_060_387, w_060_388, w_060_389, w_060_390, w_060_392, w_060_393, w_060_394, w_060_396, w_060_398, w_060_399, w_060_400, w_060_401, w_060_402, w_060_403, w_060_404, w_060_405, w_060_406, w_060_407, w_060_408, w_060_409, w_060_410, w_060_411, w_060_412, w_060_413, w_060_414, w_060_416, w_060_417, w_060_418, w_060_420, w_060_422, w_060_423, w_060_424, w_060_426, w_060_427, w_060_428, w_060_429, w_060_430, w_060_431, w_060_432, w_060_434, w_060_435, w_060_436, w_060_438, w_060_439, w_060_440, w_060_441, w_060_442, w_060_443, w_060_444, w_060_445, w_060_446, w_060_447, w_060_449, w_060_450, w_060_451, w_060_453, w_060_454, w_060_455, w_060_456, w_060_457, w_060_458, w_060_459, w_060_460, w_060_462, w_060_463, w_060_464, w_060_465, w_060_466, w_060_467, w_060_468, w_060_469, w_060_470, w_060_471, w_060_472, w_060_474, w_060_476, w_060_477, w_060_478, w_060_479, w_060_480, w_060_481, w_060_482, w_060_483, w_060_484, w_060_485, w_060_486, w_060_488, w_060_489, w_060_490, w_060_491, w_060_492, w_060_493, w_060_494, w_060_495, w_060_497, w_060_498, w_060_499, w_060_501, w_060_502, w_060_503, w_060_504, w_060_505, w_060_506, w_060_507, w_060_508, w_060_509, w_060_510, w_060_511, w_060_512, w_060_513, w_060_514, w_060_515, w_060_516, w_060_517, w_060_518, w_060_519, w_060_521, w_060_522, w_060_523, w_060_525, w_060_526, w_060_527, w_060_528, w_060_530, w_060_531, w_060_532, w_060_533, w_060_534, w_060_535, w_060_536, w_060_537, w_060_539, w_060_540, w_060_541, w_060_542, w_060_543, w_060_545, w_060_546, w_060_547, w_060_548, w_060_551, w_060_552, w_060_553, w_060_554, w_060_555, w_060_556, w_060_557, w_060_558, w_060_559, w_060_560, w_060_561, w_060_562, w_060_563, w_060_564, w_060_565, w_060_566, w_060_567, w_060_568, w_060_569, w_060_571, w_060_572, w_060_573, w_060_574, w_060_575, w_060_576, w_060_577, w_060_580, w_060_581, w_060_582, w_060_583, w_060_584, w_060_585, w_060_586, w_060_587, w_060_588, w_060_590, w_060_591, w_060_592, w_060_593, w_060_594, w_060_595, w_060_597, w_060_598, w_060_600, w_060_601, w_060_602, w_060_603, w_060_604, w_060_605, w_060_606, w_060_608, w_060_609, w_060_611, w_060_613, w_060_614, w_060_615, w_060_616, w_060_617, w_060_618, w_060_619, w_060_620, w_060_621, w_060_622, w_060_623, w_060_624, w_060_625, w_060_626, w_060_627, w_060_628, w_060_629, w_060_630, w_060_632, w_060_633, w_060_634, w_060_635, w_060_636, w_060_637, w_060_638, w_060_639, w_060_640, w_060_641, w_060_642, w_060_643, w_060_645, w_060_647, w_060_648, w_060_650, w_060_651, w_060_652, w_060_653, w_060_654, w_060_655, w_060_656, w_060_657, w_060_658, w_060_659, w_060_660, w_060_663, w_060_664, w_060_665, w_060_666, w_060_667, w_060_669, w_060_670, w_060_671, w_060_672, w_060_673, w_060_674, w_060_675, w_060_676, w_060_677, w_060_678, w_060_679, w_060_680, w_060_681, w_060_682, w_060_683, w_060_684, w_060_686, w_060_688, w_060_689, w_060_690, w_060_692, w_060_693, w_060_694, w_060_696, w_060_697, w_060_698, w_060_700, w_060_701, w_060_704, w_060_705, w_060_706, w_060_707, w_060_709, w_060_711, w_060_712, w_060_713, w_060_714, w_060_715, w_060_716, w_060_718, w_060_720, w_060_721, w_060_722, w_060_724, w_060_725, w_060_726, w_060_727, w_060_728, w_060_729, w_060_730, w_060_731, w_060_733, w_060_734, w_060_736, w_060_737, w_060_738, w_060_739, w_060_741, w_060_742, w_060_743, w_060_744, w_060_745, w_060_746, w_060_747, w_060_749, w_060_750, w_060_751, w_060_753, w_060_754, w_060_755, w_060_756, w_060_757, w_060_758, w_060_759, w_060_760, w_060_761, w_060_762, w_060_763, w_060_764, w_060_766, w_060_767, w_060_768, w_060_769, w_060_770, w_060_771, w_060_772, w_060_775, w_060_776, w_060_777, w_060_778, w_060_779, w_060_780, w_060_781, w_060_782, w_060_783, w_060_784, w_060_785, w_060_786, w_060_787, w_060_788, w_060_789, w_060_790, w_060_791, w_060_793, w_060_794, w_060_795, w_060_796, w_060_797, w_060_798, w_060_799, w_060_800, w_060_802, w_060_804, w_060_805, w_060_806, w_060_807, w_060_808, w_060_809, w_060_810, w_060_811, w_060_812, w_060_813, w_060_814, w_060_815, w_060_816, w_060_817, w_060_818, w_060_819, w_060_820, w_060_821, w_060_822, w_060_823, w_060_828, w_060_830, w_060_831, w_060_832, w_060_833, w_060_834, w_060_835, w_060_836, w_060_837, w_060_838, w_060_839, w_060_841, w_060_842, w_060_843, w_060_844, w_060_845, w_060_846, w_060_847, w_060_848, w_060_849, w_060_850, w_060_851, w_060_854, w_060_855, w_060_856, w_060_857, w_060_860, w_060_861, w_060_863, w_060_864, w_060_865, w_060_866, w_060_868, w_060_869, w_060_870, w_060_872, w_060_873, w_060_874, w_060_875, w_060_877, w_060_878, w_060_879, w_060_880, w_060_881, w_060_882, w_060_883, w_060_884, w_060_885, w_060_886, w_060_887, w_060_888, w_060_889, w_060_891, w_060_893, w_060_894, w_060_895, w_060_896, w_060_897, w_060_898, w_060_899, w_060_900, w_060_901, w_060_902, w_060_905, w_060_906, w_060_907, w_060_908, w_060_909, w_060_910, w_060_911, w_060_912, w_060_913, w_060_914, w_060_915, w_060_916, w_060_917, w_060_918, w_060_919, w_060_920, w_060_921, w_060_922, w_060_923, w_060_924, w_060_925, w_060_927, w_060_929, w_060_930, w_060_931, w_060_932, w_060_933, w_060_934, w_060_935, w_060_936, w_060_940, w_060_941, w_060_942, w_060_943, w_060_944, w_060_945, w_060_946, w_060_947, w_060_948, w_060_950, w_060_951, w_060_952, w_060_953, w_060_954, w_060_955, w_060_956, w_060_957, w_060_958, w_060_959, w_060_960, w_060_961, w_060_962, w_060_964, w_060_965, w_060_966, w_060_967, w_060_968, w_060_970, w_060_971, w_060_972, w_060_973, w_060_974, w_060_975, w_060_977, w_060_978, w_060_979, w_060_981, w_060_982, w_060_983, w_060_984, w_060_985, w_060_986, w_060_987, w_060_988, w_060_989, w_060_990, w_060_991, w_060_992, w_060_993, w_060_994, w_060_995, w_060_996, w_060_997, w_060_998, w_060_999, w_060_1000, w_060_1001, w_060_1002, w_060_1003, w_060_1004, w_060_1005, w_060_1006, w_060_1007, w_060_1008, w_060_1009, w_060_1010, w_060_1011, w_060_1012, w_060_1013, w_060_1014, w_060_1015, w_060_1016, w_060_1017, w_060_1018, w_060_1019, w_060_1020, w_060_1021, w_060_1022, w_060_1023, w_060_1024, w_060_1025, w_060_1027, w_060_1028, w_060_1029, w_060_1030, w_060_1031, w_060_1032, w_060_1034, w_060_1035, w_060_1036, w_060_1037, w_060_1038, w_060_1039, w_060_1040, w_060_1041, w_060_1043, w_060_1044, w_060_1045, w_060_1046, w_060_1047, w_060_1050, w_060_1051, w_060_1053, w_060_1054, w_060_1055, w_060_1056, w_060_1057, w_060_1058, w_060_1059, w_060_1060, w_060_1062, w_060_1064, w_060_1065, w_060_1066, w_060_1067, w_060_1068, w_060_1069, w_060_1070, w_060_1072, w_060_1073, w_060_1074, w_060_1075, w_060_1076, w_060_1077, w_060_1078, w_060_1079, w_060_1080, w_060_1081, w_060_1082, w_060_1083, w_060_1085, w_060_1086, w_060_1087, w_060_1088, w_060_1089, w_060_1090, w_060_1091, w_060_1092, w_060_1093, w_060_1095, w_060_1096, w_060_1099, w_060_1100, w_060_1101, w_060_1102, w_060_1103, w_060_1104, w_060_1105, w_060_1106, w_060_1108, w_060_1109, w_060_1112, w_060_1113, w_060_1115, w_060_1116, w_060_1117, w_060_1118, w_060_1120, w_060_1121, w_060_1122, w_060_1123, w_060_1124, w_060_1125, w_060_1126, w_060_1127, w_060_1128, w_060_1129, w_060_1130, w_060_1131, w_060_1132, w_060_1134, w_060_1135, w_060_1136, w_060_1137, w_060_1138, w_060_1139, w_060_1140, w_060_1141, w_060_1142, w_060_1143, w_060_1144, w_060_1145, w_060_1146, w_060_1148, w_060_1150, w_060_1151, w_060_1152, w_060_1153, w_060_1154, w_060_1156, w_060_1157, w_060_1158, w_060_1159, w_060_1160, w_060_1162, w_060_1164, w_060_1165, w_060_1166, w_060_1167, w_060_1169, w_060_1170, w_060_1173, w_060_1174, w_060_1175, w_060_1176, w_060_1177, w_060_1178, w_060_1180, w_060_1181, w_060_1182, w_060_1183, w_060_1185, w_060_1186, w_060_1187, w_060_1188, w_060_1190, w_060_1191, w_060_1192, w_060_1193, w_060_1194, w_060_1195, w_060_1196, w_060_1197, w_060_1198, w_060_1199, w_060_1201, w_060_1203, w_060_1204, w_060_1205, w_060_1206, w_060_1207, w_060_1208, w_060_1209, w_060_1210, w_060_1211, w_060_1212, w_060_1213, w_060_1214, w_060_1215, w_060_1217, w_060_1218, w_060_1219, w_060_1220, w_060_1221, w_060_1222, w_060_1223, w_060_1224, w_060_1226, w_060_1227, w_060_1228, w_060_1230, w_060_1231, w_060_1232, w_060_1233, w_060_1234, w_060_1235, w_060_1236, w_060_1237, w_060_1238, w_060_1240, w_060_1241, w_060_1242, w_060_1243, w_060_1244, w_060_1245, w_060_1246, w_060_1247, w_060_1248, w_060_1249, w_060_1250, w_060_1251, w_060_1252, w_060_1253, w_060_1254, w_060_1255, w_060_1257, w_060_1258, w_060_1259, w_060_1260, w_060_1262, w_060_1264, w_060_1266, w_060_1268, w_060_1269, w_060_1272, w_060_1273, w_060_1274, w_060_1276, w_060_1277, w_060_1278, w_060_1279, w_060_1281, w_060_1282, w_060_1283, w_060_1284, w_060_1285, w_060_1287, w_060_1289, w_060_1292, w_060_1293, w_060_1294, w_060_1295, w_060_1296, w_060_1297, w_060_1298, w_060_1300, w_060_1302, w_060_1304, w_060_1305, w_060_1306, w_060_1308, w_060_1309, w_060_1311, w_060_1313, w_060_1314, w_060_1315, w_060_1318, w_060_1319, w_060_1320, w_060_1321, w_060_1322, w_060_1324, w_060_1325, w_060_1326, w_060_1328, w_060_1330, w_060_1332, w_060_1333, w_060_1334, w_060_1336, w_060_1337, w_060_1338, w_060_1339, w_060_1341, w_060_1342, w_060_1343, w_060_1344, w_060_1346, w_060_1347, w_060_1349, w_060_1350, w_060_1351, w_060_1352, w_060_1355, w_060_1356, w_060_1357, w_060_1359, w_060_1360, w_060_1361, w_060_1362, w_060_1363, w_060_1365, w_060_1366, w_060_1368, w_060_1369, w_060_1370, w_060_1371, w_060_1373, w_060_1375, w_060_1376, w_060_1377, w_060_1378, w_060_1379, w_060_1380, w_060_1383, w_060_1386, w_060_1387, w_060_1388, w_060_1390, w_060_1391, w_060_1392, w_060_1393, w_060_1394, w_060_1395, w_060_1396, w_060_1397, w_060_1398, w_060_1400, w_060_1401, w_060_1403, w_060_1409, w_060_1410, w_060_1411, w_060_1412, w_060_1413, w_060_1414, w_060_1415, w_060_1417, w_060_1418, w_060_1419, w_060_1421, w_060_1423, w_060_1424, w_060_1426, w_060_1427, w_060_1428, w_060_1429, w_060_1430, w_060_1431, w_060_1432, w_060_1433, w_060_1434, w_060_1435, w_060_1437, w_060_1438, w_060_1441, w_060_1443, w_060_1445, w_060_1446, w_060_1448, w_060_1449, w_060_1451, w_060_1452, w_060_1454, w_060_1455, w_060_1457, w_060_1459, w_060_1460, w_060_1462, w_060_1463, w_060_1465, w_060_1467, w_060_1468, w_060_1469, w_060_1471, w_060_1472, w_060_1473, w_060_1474, w_060_1477, w_060_1478, w_060_1479, w_060_1482, w_060_1483, w_060_1484, w_060_1485, w_060_1487, w_060_1488, w_060_1489, w_060_1490, w_060_1491, w_060_1492, w_060_1493, w_060_1495, w_060_1496, w_060_1497, w_060_1498, w_060_1499, w_060_1500, w_060_1502, w_060_1504, w_060_1505, w_060_1506, w_060_1507, w_060_1509, w_060_1511, w_060_1512, w_060_1513, w_060_1514, w_060_1516, w_060_1517, w_060_1518, w_060_1519, w_060_1521, w_060_1522, w_060_1523, w_060_1524, w_060_1525, w_060_1527, w_060_1529, w_060_1534, w_060_1535, w_060_1537, w_060_1538, w_060_1540, w_060_1541, w_060_1542, w_060_1544, w_060_1545, w_060_1547, w_060_1548, w_060_1550, w_060_1551, w_060_1552, w_060_1553, w_060_1554, w_060_1555, w_060_1556, w_060_1558, w_060_1559, w_060_1560, w_060_1561, w_060_1563, w_060_1564, w_060_1565, w_060_1567, w_060_1568, w_060_1572, w_060_1579, w_060_1581, w_060_1582, w_060_1583, w_060_1585, w_060_1586, w_060_1587, w_060_1588, w_060_1589, w_060_1592, w_060_1594, w_060_1596, w_060_1597, w_060_1598, w_060_1599, w_060_1601, w_060_1602, w_060_1604, w_060_1605, w_060_1606, w_060_1608, w_060_1609, w_060_1610, w_060_1611, w_060_1612, w_060_1615, w_060_1616, w_060_1618, w_060_1620, w_060_1621, w_060_1622, w_060_1623, w_060_1624, w_060_1625, w_060_1627, w_060_1629, w_060_1630, w_060_1632, w_060_1633, w_060_1634, w_060_1635, w_060_1636, w_060_1637, w_060_1640, w_060_1641, w_060_1642, w_060_1643, w_060_1644, w_060_1646, w_060_1647, w_060_1650, w_060_1651, w_060_1652, w_060_1653, w_060_1654, w_060_1655, w_060_1658, w_060_1660, w_060_1661, w_060_1662, w_060_1663, w_060_1664, w_060_1665, w_060_1666, w_060_1667, w_060_1668, w_060_1669, w_060_1670, w_060_1671, w_060_1672, w_060_1673, w_060_1674, w_060_1676, w_060_1677, w_060_1679, w_060_1680, w_060_1681, w_060_1682, w_060_1683, w_060_1685, w_060_1687, w_060_1690, w_060_1692, w_060_1694, w_060_1695, w_060_1696, w_060_1697, w_060_1699, w_060_1701, w_060_1702, w_060_1704, w_060_1705, w_060_1706, w_060_1708, w_060_1709, w_060_1710, w_060_1711, w_060_1712, w_060_1714, w_060_1716, w_060_1717, w_060_1718, w_060_1719, w_060_1720, w_060_1721, w_060_1722, w_060_1723, w_060_1724, w_060_1725, w_060_1726, w_060_1728, w_060_1729, w_060_1733, w_060_1734, w_060_1735, w_060_1736, w_060_1737, w_060_1738, w_060_1739, w_060_1740, w_060_1741, w_060_1742, w_060_1744, w_060_1745, w_060_1746, w_060_1747, w_060_1750, w_060_1751, w_060_1752, w_060_1753, w_060_1754, w_060_1755, w_060_1757, w_060_1759, w_060_1762, w_060_1763, w_060_1765, w_060_1767, w_060_1768, w_060_1770, w_060_1771, w_060_1772, w_060_1773, w_060_1774, w_060_1776, w_060_1778, w_060_1779, w_060_1780, w_060_1781, w_060_1782, w_060_1783, w_060_1784, w_060_1785, w_060_1786, w_060_1787, w_060_1790, w_060_1792, w_060_1793, w_060_1795, w_060_1796, w_060_1797, w_060_1798, w_060_1800, w_060_1801, w_060_1802, w_060_1803, w_060_1804, w_060_1805, w_060_1806, w_060_1807, w_060_1808, w_060_1809, w_060_1810, w_060_1812, w_060_1813, w_060_1814, w_060_1815, w_060_1816, w_060_1817, w_060_1820, w_060_1821, w_060_1822, w_060_1824, w_060_1825, w_060_1826, w_060_1827, w_060_1828, w_060_1829, w_060_1830, w_060_1832, w_060_1833, w_060_1834, w_060_1835, w_060_1836, w_060_1837, w_060_1838, w_060_1839, w_060_1840, w_060_1841, w_060_1845, w_060_1846, w_060_1847, w_060_1849, w_060_1851, w_060_1853, w_060_1854, w_060_1855, w_060_1857, w_060_1858, w_060_1860, w_060_1861, w_060_1862, w_060_1864, w_060_1865, w_060_1866, w_060_1867, w_060_1868, w_060_1872, w_060_1874, w_060_1876, w_060_1877, w_060_1878, w_060_1879, w_060_1880, w_060_1882, w_060_1883, w_060_1884, w_060_1885, w_060_1886, w_060_1891, w_060_1892, w_060_1894, w_060_1895, w_060_1896, w_060_1898, w_060_1900, w_060_1902, w_060_1903, w_060_1904, w_060_1905, w_060_1907, w_060_1908, w_060_1910, w_060_1911, w_060_1912, w_060_1913, w_060_1916, w_060_1917, w_060_1918, w_060_1919, w_060_1920, w_060_1921, w_060_1922, w_060_1923, w_060_1925, w_060_1926, w_060_1927, w_060_1928, w_060_1929, w_060_1930, w_060_1931, w_060_1932, w_060_1934, w_060_1935, w_060_1936, w_060_1937, w_060_1938, w_060_1939, w_060_1941, w_060_1942, w_060_1945, w_060_1947, w_060_1948, w_060_1949, w_060_1951, w_060_1952, w_060_1953, w_060_1954, w_060_1956, w_060_1957, w_060_1959, w_060_1960, w_060_1961, w_060_1963, w_060_1964, w_060_1965, w_060_1966, w_060_1969, w_060_1970, w_060_1971, w_060_1972, w_060_1974, w_060_1978, w_060_1979, w_060_1980, w_060_1981, w_060_1983, w_060_1986, w_060_1987, w_060_1989, w_060_1990, w_060_1991, w_060_1992, w_060_1993, w_060_1994, w_060_1995, w_060_1996, w_060_1997, w_060_1999, w_060_2000, w_060_2001, w_060_2003, w_060_2004, w_060_2005, w_060_2006, w_060_2007, w_060_2009, w_060_2010, w_060_2011, w_060_2012, w_060_2013, w_060_2015, w_060_2016, w_060_2017, w_060_2018, w_060_2021, w_060_2026, w_060_2027, w_060_2028, w_060_2029, w_060_2030, w_060_2031, w_060_2032, w_060_2033, w_060_2034, w_060_2035, w_060_2038, w_060_2039, w_060_2041, w_060_2043, w_060_2044, w_060_2045, w_060_2046, w_060_2047, w_060_2048, w_060_2049, w_060_2050, w_060_2051, w_060_2052, w_060_2053, w_060_2055, w_060_2056, w_060_2058, w_060_2059, w_060_2060, w_060_2062, w_060_2063, w_060_2064, w_060_2068, w_060_2069, w_060_2070, w_060_2071, w_060_2072, w_060_2074, w_060_2075, w_060_2076, w_060_2077, w_060_2078, w_060_2079, w_060_2080, w_060_2081, w_060_2082, w_060_2084, w_060_2085, w_060_2086, w_060_2087, w_060_2089, w_060_2090, w_060_2091, w_060_2092, w_060_2093, w_060_2095, w_060_2096, w_060_2097, w_060_2098, w_060_2099, w_060_2100, w_060_2101, w_060_2102, w_060_2103, w_060_2104, w_060_2105, w_060_2106, w_060_2107, w_060_2109, w_060_2110, w_060_2112, w_060_2114, w_060_2115, w_060_2116, w_060_2119, w_060_2120, w_060_2122, w_060_2123, w_060_2124, w_060_2125, w_060_2126, w_060_2129, w_060_2132, w_060_2133, w_060_2134, w_060_2135, w_060_2137, w_060_2138, w_060_2139, w_060_2140, w_060_2141, w_060_2142, w_060_2143, w_060_2145, w_060_2147, w_060_2148, w_060_2149, w_060_2151, w_060_2152, w_060_2155, w_060_2157, w_060_2159, w_060_2160, w_060_2162, w_060_2163, w_060_2164, w_060_2165, w_060_2167, w_060_2168, w_060_2169, w_060_2170, w_060_2171, w_060_2172, w_060_2173, w_060_2174, w_060_2175, w_060_2176, w_060_2177, w_060_2178, w_060_2179, w_060_2181, w_060_2182, w_060_2183, w_060_2184, w_060_2185, w_060_2188, w_060_2189, w_060_2190, w_060_2191, w_060_2193, w_060_2195, w_060_2196, w_060_2197, w_060_2199, w_060_2200, w_060_2201, w_060_2202, w_060_2203, w_060_2205, w_060_2206, w_060_2208, w_060_2209, w_060_2210, w_060_2211, w_060_2212, w_060_2213, w_060_2214, w_060_2215, w_060_2217, w_060_2219, w_060_2220, w_060_2221, w_060_2222, w_060_2223, w_060_2226, w_060_2227, w_060_2228, w_060_2229, w_060_2230, w_060_2231, w_060_2233, w_060_2234, w_060_2235, w_060_2236, w_060_2237, w_060_2238, w_060_2241, w_060_2242, w_060_2243, w_060_2245, w_060_2246, w_060_2247, w_060_2248, w_060_2249, w_060_2250, w_060_2251, w_060_2252, w_060_2253, w_060_2254, w_060_2255, w_060_2257, w_060_2258, w_060_2259, w_060_2261, w_060_2262, w_060_2263, w_060_2264, w_060_2266, w_060_2267, w_060_2269, w_060_2270, w_060_2271, w_060_2273, w_060_2275, w_060_2276, w_060_2277, w_060_2278, w_060_2279, w_060_2280, w_060_2282, w_060_2286, w_060_2287, w_060_2288, w_060_2289, w_060_2290, w_060_2291, w_060_2295, w_060_2297, w_060_2301, w_060_2302, w_060_2303, w_060_2304, w_060_2305, w_060_2306, w_060_2307, w_060_2308, w_060_2309, w_060_2310, w_060_2311, w_060_2314, w_060_2316, w_060_2317, w_060_2319, w_060_2321, w_060_2322, w_060_2323, w_060_2325, w_060_2326, w_060_2327, w_060_2328, w_060_2329, w_060_2331, w_060_2332, w_060_2333, w_060_2336, w_060_2337, w_060_2338, w_060_2339, w_060_2341, w_060_2344, w_060_2345, w_060_2346, w_060_2347, w_060_2348, w_060_2349, w_060_2350, w_060_2351, w_060_2352, w_060_2353, w_060_2354, w_060_2355, w_060_2357, w_060_2360, w_060_2361, w_060_2363, w_060_2365, w_060_2371, w_060_2372, w_060_2373, w_060_2374, w_060_2376, w_060_2377, w_060_2378, w_060_2379, w_060_2381, w_060_2384, w_060_2385, w_060_2387, w_060_2390, w_060_2393, w_060_2394, w_060_2396, w_060_2398, w_060_2399, w_060_2403, w_060_2404, w_060_2405, w_060_2406, w_060_2407, w_060_2408, w_060_2409, w_060_2410, w_060_2411, w_060_2412, w_060_2413, w_060_2414, w_060_2415, w_060_2417, w_060_2418, w_060_2419, w_060_2420, w_060_2424, w_060_2425, w_060_2426, w_060_2427, w_060_2429, w_060_2431, w_060_2432, w_060_2433, w_060_2434, w_060_2435, w_060_2436, w_060_2438, w_060_2439, w_060_2441, w_060_2443, w_060_2444, w_060_2445, w_060_2447, w_060_2448, w_060_2451, w_060_2452, w_060_2453, w_060_2455, w_060_2456, w_060_2457, w_060_2460, w_060_2461, w_060_2462, w_060_2464, w_060_2465, w_060_2466, w_060_2467, w_060_2468, w_060_2469, w_060_2470, w_060_2471, w_060_2472, w_060_2473, w_060_2474, w_060_2475, w_060_2477, w_060_2478, w_060_2479, w_060_2480, w_060_2481, w_060_2483, w_060_2484, w_060_2485, w_060_2486, w_060_2487, w_060_2488, w_060_2489, w_060_2490, w_060_2493, w_060_2494, w_060_2495, w_060_2496, w_060_2497, w_060_2498, w_060_2499, w_060_2501, w_060_2502, w_060_2503, w_060_2504, w_060_2505, w_060_2506, w_060_2508, w_060_2509, w_060_2510, w_060_2511, w_060_2512, w_060_2513, w_060_2517, w_060_2518, w_060_2519, w_060_2522, w_060_2524, w_060_2525, w_060_2528, w_060_2529, w_060_2530, w_060_2531, w_060_2532, w_060_2533, w_060_2535, w_060_2536, w_060_2537, w_060_2538, w_060_2539, w_060_2540, w_060_2543, w_060_2544, w_060_2545, w_060_2546, w_060_2547, w_060_2548, w_060_2549, w_060_2550, w_060_2551, w_060_2552, w_060_2553, w_060_2554, w_060_2555, w_060_2556, w_060_2557, w_060_2558, w_060_2559, w_060_2560, w_060_2561, w_060_2563, w_060_2564, w_060_2565, w_060_2567, w_060_2568, w_060_2570, w_060_2572, w_060_2576, w_060_2578, w_060_2579, w_060_2580, w_060_2581, w_060_2582, w_060_2583, w_060_2584, w_060_2586, w_060_2587, w_060_2588, w_060_2592, w_060_2594, w_060_2595, w_060_2596, w_060_2597, w_060_2598, w_060_2601, w_060_2602, w_060_2603, w_060_2605, w_060_2606, w_060_2609, w_060_2611, w_060_2612, w_060_2613, w_060_2616, w_060_2617, w_060_2618, w_060_2619, w_060_2620, w_060_2621, w_060_2623, w_060_2625, w_060_2626, w_060_2629, w_060_2632, w_060_2633, w_060_2634, w_060_2635, w_060_2636, w_060_2637, w_060_2638, w_060_2639, w_060_2640, w_060_2641, w_060_2642, w_060_2643, w_060_2644, w_060_2645, w_060_2646, w_060_2647, w_060_2649, w_060_2650, w_060_2651, w_060_2652, w_060_2653, w_060_2654, w_060_2655, w_060_2658, w_060_2659, w_060_2661, w_060_2662, w_060_2665, w_060_2666, w_060_2668, w_060_2670, w_060_2671, w_060_2672, w_060_2673, w_060_2674, w_060_2675, w_060_2676, w_060_2677, w_060_2678, w_060_2679, w_060_2680, w_060_2683, w_060_2684, w_060_2685, w_060_2686, w_060_2687, w_060_2688, w_060_2689, w_060_2691, w_060_2692, w_060_2694, w_060_2695, w_060_2696, w_060_2697, w_060_2698, w_060_2699, w_060_2701, w_060_2703, w_060_2706, w_060_2707, w_060_2708, w_060_2709, w_060_2710, w_060_2711, w_060_2712, w_060_2713, w_060_2715, w_060_2716, w_060_2717, w_060_2718, w_060_2719, w_060_2720, w_060_2721, w_060_2722, w_060_2723, w_060_2725, w_060_2726, w_060_2730, w_060_2731, w_060_2732, w_060_2733, w_060_2737, w_060_2738, w_060_2739, w_060_2741, w_060_2742, w_060_2743, w_060_2745, w_060_2747, w_060_2748, w_060_2749, w_060_2750, w_060_2751, w_060_2752, w_060_2754, w_060_2755, w_060_2756, w_060_2757, w_060_2758, w_060_2759, w_060_2760, w_060_2761, w_060_2763, w_060_2764, w_060_2765, w_060_2768, w_060_2771, w_060_2772, w_060_2773, w_060_2774, w_060_2775, w_060_2777, w_060_2780, w_060_2781, w_060_2782, w_060_2784, w_060_2785, w_060_2786, w_060_2787, w_060_2788, w_060_2789, w_060_2791, w_060_2792, w_060_2793, w_060_2794, w_060_2797, w_060_2799, w_060_2800, w_060_2802, w_060_2803, w_060_2804, w_060_2805, w_060_2806, w_060_2807, w_060_2809, w_060_2810, w_060_2811, w_060_2812, w_060_2813, w_060_2814, w_060_2815, w_060_2819, w_060_2820, w_060_2821, w_060_2822, w_060_2823, w_060_2825, w_060_2826, w_060_2827, w_060_2828, w_060_2829, w_060_2830, w_060_2831, w_060_2832, w_060_2833, w_060_2834, w_060_2835, w_060_2836, w_060_2837, w_060_2838, w_060_2839, w_060_2840, w_060_2842, w_060_2844, w_060_2846, w_060_2847, w_060_2848, w_060_2849, w_060_2851, w_060_2852, w_060_2853, w_060_2855, w_060_2856, w_060_2857, w_060_2858, w_060_2859, w_060_2861, w_060_2862, w_060_2863, w_060_2864, w_060_2865, w_060_2866, w_060_2868, w_060_2869, w_060_2870, w_060_2871, w_060_2872, w_060_2873, w_060_2874, w_060_2876, w_060_2878, w_060_2879, w_060_2881, w_060_2883, w_060_2884, w_060_2885, w_060_2886, w_060_2888, w_060_2889, w_060_2890, w_060_2891, w_060_2893, w_060_2895, w_060_2896, w_060_2897, w_060_2898, w_060_2899, w_060_2901, w_060_2903, w_060_2907, w_060_2908, w_060_2909, w_060_2910, w_060_2911, w_060_2912;
  wire w_061_001, w_061_002, w_061_003, w_061_004, w_061_005, w_061_006, w_061_007, w_061_009, w_061_010, w_061_011, w_061_012, w_061_013, w_061_014, w_061_015, w_061_016, w_061_017, w_061_018, w_061_019, w_061_020, w_061_021, w_061_022, w_061_023, w_061_024, w_061_025, w_061_026, w_061_027, w_061_028, w_061_029, w_061_030, w_061_031, w_061_032, w_061_033, w_061_034, w_061_035, w_061_036, w_061_037, w_061_038, w_061_039, w_061_040, w_061_041, w_061_043, w_061_044, w_061_045, w_061_047, w_061_048, w_061_049, w_061_050, w_061_051, w_061_052, w_061_053, w_061_054, w_061_055, w_061_056, w_061_057, w_061_058, w_061_059, w_061_060, w_061_061, w_061_062, w_061_063, w_061_064, w_061_065, w_061_066, w_061_067, w_061_068, w_061_069, w_061_070, w_061_071, w_061_072, w_061_073, w_061_074, w_061_075, w_061_076, w_061_077, w_061_078, w_061_079, w_061_080, w_061_081, w_061_082, w_061_083, w_061_084, w_061_085, w_061_086, w_061_087, w_061_088, w_061_089, w_061_090, w_061_091, w_061_092, w_061_093, w_061_094, w_061_095, w_061_096, w_061_097, w_061_098, w_061_099, w_061_100, w_061_101, w_061_102, w_061_103, w_061_104, w_061_105, w_061_106, w_061_107, w_061_108, w_061_109, w_061_110, w_061_111, w_061_112, w_061_113, w_061_114, w_061_115, w_061_116, w_061_117, w_061_118, w_061_119, w_061_120, w_061_121, w_061_122, w_061_123, w_061_124, w_061_125, w_061_126, w_061_127, w_061_128, w_061_129, w_061_130, w_061_131, w_061_132, w_061_133, w_061_134, w_061_135, w_061_136, w_061_137, w_061_138, w_061_139, w_061_140, w_061_141, w_061_142, w_061_143, w_061_144, w_061_145, w_061_146, w_061_147, w_061_148, w_061_149, w_061_150, w_061_151, w_061_152, w_061_153, w_061_154, w_061_155, w_061_156, w_061_157, w_061_158, w_061_159, w_061_160, w_061_161, w_061_162, w_061_163, w_061_164, w_061_165, w_061_166, w_061_167, w_061_168, w_061_169, w_061_170, w_061_171, w_061_172, w_061_173, w_061_174, w_061_175, w_061_176, w_061_177, w_061_178, w_061_179, w_061_180, w_061_181, w_061_182, w_061_183, w_061_184, w_061_185, w_061_186, w_061_187, w_061_188, w_061_189, w_061_190, w_061_191, w_061_192, w_061_193, w_061_194, w_061_195, w_061_196, w_061_197, w_061_198, w_061_199, w_061_200, w_061_201, w_061_202, w_061_204, w_061_205, w_061_206, w_061_207, w_061_208, w_061_209, w_061_210, w_061_211, w_061_212, w_061_213, w_061_214, w_061_215, w_061_216, w_061_217, w_061_218, w_061_219, w_061_220, w_061_221, w_061_222, w_061_223, w_061_224, w_061_225, w_061_226, w_061_227, w_061_228, w_061_229, w_061_231, w_061_232, w_061_233, w_061_234, w_061_235, w_061_236, w_061_237, w_061_238, w_061_239, w_061_241, w_061_242, w_061_243, w_061_244, w_061_245, w_061_246, w_061_247, w_061_248, w_061_249, w_061_250, w_061_251, w_061_252, w_061_253, w_061_254, w_061_255, w_061_256, w_061_257, w_061_258, w_061_259, w_061_260, w_061_261, w_061_263, w_061_264, w_061_265, w_061_266, w_061_267, w_061_268, w_061_269, w_061_270, w_061_271, w_061_272, w_061_273, w_061_274, w_061_275, w_061_276, w_061_277, w_061_278, w_061_279, w_061_280, w_061_281, w_061_282, w_061_283, w_061_284, w_061_285, w_061_287, w_061_288, w_061_289, w_061_290, w_061_291, w_061_292, w_061_293, w_061_294, w_061_295, w_061_296, w_061_297, w_061_298, w_061_299, w_061_300, w_061_301, w_061_302, w_061_303, w_061_304, w_061_305, w_061_306, w_061_307, w_061_308, w_061_309, w_061_310, w_061_311, w_061_312, w_061_313, w_061_314, w_061_315, w_061_316, w_061_317, w_061_318, w_061_319, w_061_320, w_061_321, w_061_322, w_061_323, w_061_324, w_061_325, w_061_326, w_061_327, w_061_328, w_061_329, w_061_330, w_061_331, w_061_332, w_061_333, w_061_334, w_061_335, w_061_336, w_061_337, w_061_338, w_061_339, w_061_340, w_061_341, w_061_342, w_061_343, w_061_344, w_061_345, w_061_347, w_061_348, w_061_349, w_061_350, w_061_351, w_061_352, w_061_353, w_061_354, w_061_355, w_061_356, w_061_357, w_061_358, w_061_359, w_061_360, w_061_361, w_061_362, w_061_363, w_061_364, w_061_365, w_061_366, w_061_367, w_061_368, w_061_369, w_061_370, w_061_372, w_061_373, w_061_374, w_061_375, w_061_376, w_061_377, w_061_378, w_061_379, w_061_380, w_061_381, w_061_382, w_061_383, w_061_384, w_061_385, w_061_386, w_061_387, w_061_388, w_061_389, w_061_390, w_061_391, w_061_392, w_061_393, w_061_395, w_061_396, w_061_397, w_061_398, w_061_399, w_061_400, w_061_401, w_061_402, w_061_403, w_061_404, w_061_405, w_061_406, w_061_407, w_061_408, w_061_409, w_061_410, w_061_411, w_061_412, w_061_413, w_061_414, w_061_415, w_061_417, w_061_418, w_061_419, w_061_420, w_061_423, w_061_424, w_061_425, w_061_426, w_061_427, w_061_429, w_061_430, w_061_431, w_061_432, w_061_433, w_061_434, w_061_435, w_061_436, w_061_437, w_061_438, w_061_439, w_061_440, w_061_441, w_061_442, w_061_443, w_061_444, w_061_445, w_061_446, w_061_447, w_061_448, w_061_449, w_061_450, w_061_451, w_061_452, w_061_453, w_061_454, w_061_455, w_061_456, w_061_457, w_061_458, w_061_459, w_061_460, w_061_461, w_061_462, w_061_463, w_061_464, w_061_465, w_061_466, w_061_467, w_061_468, w_061_469, w_061_470, w_061_471, w_061_472, w_061_473, w_061_474, w_061_476, w_061_477, w_061_478, w_061_479, w_061_480, w_061_481, w_061_482, w_061_484, w_061_485, w_061_486, w_061_487, w_061_488, w_061_489, w_061_490, w_061_491, w_061_492, w_061_493, w_061_494, w_061_495, w_061_496, w_061_497, w_061_498, w_061_499, w_061_500, w_061_501, w_061_502, w_061_504, w_061_505, w_061_506, w_061_507, w_061_509, w_061_510, w_061_511, w_061_512, w_061_513, w_061_514, w_061_515, w_061_516, w_061_517, w_061_518, w_061_519, w_061_520, w_061_521, w_061_522, w_061_523, w_061_524, w_061_525, w_061_526, w_061_527, w_061_528, w_061_529, w_061_530, w_061_531, w_061_532, w_061_533, w_061_534, w_061_535, w_061_536, w_061_537, w_061_538, w_061_539, w_061_540, w_061_541, w_061_542, w_061_543, w_061_544, w_061_545, w_061_546, w_061_547, w_061_548, w_061_549, w_061_550, w_061_552, w_061_553, w_061_554, w_061_555, w_061_556, w_061_557, w_061_558, w_061_559, w_061_560, w_061_561, w_061_562, w_061_563, w_061_564, w_061_565, w_061_566, w_061_567, w_061_568, w_061_569, w_061_570, w_061_571, w_061_572, w_061_573, w_061_574, w_061_575, w_061_576, w_061_577, w_061_578, w_061_579, w_061_580, w_061_581, w_061_582, w_061_583, w_061_584, w_061_585, w_061_586, w_061_587, w_061_588, w_061_589, w_061_590, w_061_591, w_061_592, w_061_593, w_061_594, w_061_595, w_061_596, w_061_597, w_061_598, w_061_599, w_061_601, w_061_602, w_061_603, w_061_604, w_061_605, w_061_606, w_061_607, w_061_608, w_061_609, w_061_610, w_061_611, w_061_612, w_061_613, w_061_615, w_061_616, w_061_617, w_061_618, w_061_619, w_061_620, w_061_621, w_061_622, w_061_623, w_061_624, w_061_625, w_061_626, w_061_627, w_061_628, w_061_629, w_061_630, w_061_631, w_061_633, w_061_634, w_061_635, w_061_636, w_061_637, w_061_638, w_061_639, w_061_640, w_061_641, w_061_642, w_061_643, w_061_644, w_061_645, w_061_646, w_061_647, w_061_648, w_061_649, w_061_650, w_061_651, w_061_652, w_061_653, w_061_654, w_061_655, w_061_656, w_061_657, w_061_658, w_061_659, w_061_660, w_061_661, w_061_662, w_061_663, w_061_665, w_061_666, w_061_667, w_061_668, w_061_669, w_061_670, w_061_671, w_061_672, w_061_673, w_061_674, w_061_675, w_061_676, w_061_677, w_061_679, w_061_680, w_061_681, w_061_682, w_061_683, w_061_684, w_061_685, w_061_686, w_061_687, w_061_688, w_061_690, w_061_691, w_061_692, w_061_693, w_061_694, w_061_695, w_061_696, w_061_698, w_061_699, w_061_700, w_061_701, w_061_702, w_061_703, w_061_704, w_061_705, w_061_706, w_061_707, w_061_708, w_061_709, w_061_710, w_061_711, w_061_712, w_061_713, w_061_714, w_061_715, w_061_716, w_061_717, w_061_718, w_061_719, w_061_720, w_061_721, w_061_722, w_061_723, w_061_724, w_061_725, w_061_726, w_061_727, w_061_728, w_061_729, w_061_730, w_061_731, w_061_732, w_061_733, w_061_734, w_061_735, w_061_736, w_061_737, w_061_738, w_061_739, w_061_740, w_061_741, w_061_742, w_061_743, w_061_744, w_061_745, w_061_746, w_061_747, w_061_748, w_061_749, w_061_750, w_061_751, w_061_752, w_061_753, w_061_754, w_061_755, w_061_757, w_061_758, w_061_759, w_061_760, w_061_761, w_061_762, w_061_763, w_061_764, w_061_765, w_061_766, w_061_767, w_061_768, w_061_769, w_061_770, w_061_771, w_061_772, w_061_773, w_061_774, w_061_775, w_061_776, w_061_777, w_061_779, w_061_780, w_061_781, w_061_782, w_061_783, w_061_784, w_061_785, w_061_786, w_061_787, w_061_788, w_061_790, w_061_791, w_061_792, w_061_793, w_061_794, w_061_795, w_061_796, w_061_797, w_061_798, w_061_799, w_061_800, w_061_801, w_061_802, w_061_803, w_061_804, w_061_805, w_061_806, w_061_807, w_061_808, w_061_809, w_061_810, w_061_811, w_061_812, w_061_813, w_061_814, w_061_815, w_061_816, w_061_817, w_061_818, w_061_819, w_061_820, w_061_821, w_061_822, w_061_823, w_061_824, w_061_825, w_061_826, w_061_827, w_061_828, w_061_829, w_061_830, w_061_831, w_061_832, w_061_833, w_061_834, w_061_835, w_061_836, w_061_837, w_061_838, w_061_839, w_061_840, w_061_841, w_061_842, w_061_843, w_061_845, w_061_846, w_061_847, w_061_848, w_061_849, w_061_850, w_061_851, w_061_854, w_061_855, w_061_856, w_061_857, w_061_858, w_061_859, w_061_860, w_061_861, w_061_862, w_061_863, w_061_864, w_061_865, w_061_866, w_061_867, w_061_869, w_061_870, w_061_871, w_061_872, w_061_873, w_061_874, w_061_875, w_061_876, w_061_877, w_061_878, w_061_879, w_061_880, w_061_881, w_061_882, w_061_883, w_061_884, w_061_885, w_061_886, w_061_887, w_061_888, w_061_889, w_061_890, w_061_891, w_061_892, w_061_893, w_061_894, w_061_895, w_061_896, w_061_897, w_061_898, w_061_899, w_061_900, w_061_901, w_061_902, w_061_903, w_061_904, w_061_905, w_061_906, w_061_907, w_061_908, w_061_909, w_061_911, w_061_912, w_061_914, w_061_915, w_061_916, w_061_917, w_061_918, w_061_919, w_061_920, w_061_921, w_061_922, w_061_923, w_061_924, w_061_925, w_061_926, w_061_927, w_061_928, w_061_929, w_061_930, w_061_931, w_061_932, w_061_933, w_061_934, w_061_935, w_061_936, w_061_937, w_061_938, w_061_939, w_061_940, w_061_941, w_061_942, w_061_943, w_061_944, w_061_945, w_061_946, w_061_947, w_061_948, w_061_949, w_061_950, w_061_951, w_061_952, w_061_953, w_061_954, w_061_955, w_061_956, w_061_957, w_061_958, w_061_959, w_061_960, w_061_961, w_061_962, w_061_963, w_061_964, w_061_965, w_061_966, w_061_967, w_061_968, w_061_969, w_061_970, w_061_971, w_061_972, w_061_973, w_061_975, w_061_976, w_061_977, w_061_978, w_061_979, w_061_980, w_061_981, w_061_982, w_061_983, w_061_984, w_061_985, w_061_986, w_061_987, w_061_988, w_061_991, w_061_992, w_061_993, w_061_994, w_061_996, w_061_997, w_061_998, w_061_999, w_061_1000, w_061_1001, w_061_1002, w_061_1003, w_061_1004, w_061_1005, w_061_1006, w_061_1007, w_061_1008, w_061_1009, w_061_1010, w_061_1011, w_061_1012, w_061_1013, w_061_1014, w_061_1015, w_061_1016, w_061_1017, w_061_1018, w_061_1020, w_061_1021, w_061_1022, w_061_1023, w_061_1024, w_061_1025, w_061_1026, w_061_1027, w_061_1028, w_061_1029, w_061_1030, w_061_1031, w_061_1032, w_061_1033, w_061_1034, w_061_1035, w_061_1036, w_061_1037, w_061_1038, w_061_1039, w_061_1040, w_061_1041, w_061_1042, w_061_1043, w_061_1044, w_061_1045, w_061_1046, w_061_1048, w_061_1049, w_061_1050, w_061_1051, w_061_1052, w_061_1053, w_061_1054, w_061_1055, w_061_1056, w_061_1057, w_061_1058, w_061_1059, w_061_1060, w_061_1061, w_061_1062, w_061_1063, w_061_1064, w_061_1065, w_061_1066, w_061_1067, w_061_1068, w_061_1069, w_061_1070, w_061_1071, w_061_1072, w_061_1073, w_061_1074, w_061_1075, w_061_1076, w_061_1077, w_061_1078, w_061_1079, w_061_1080, w_061_1081, w_061_1082, w_061_1083, w_061_1085, w_061_1086, w_061_1087, w_061_1088, w_061_1090, w_061_1091, w_061_1092, w_061_1093, w_061_1094, w_061_1095, w_061_1096, w_061_1097, w_061_1098, w_061_1099, w_061_1101, w_061_1102, w_061_1103, w_061_1104, w_061_1105, w_061_1106, w_061_1107, w_061_1108, w_061_1109, w_061_1110, w_061_1111, w_061_1112, w_061_1113, w_061_1114, w_061_1115, w_061_1116, w_061_1117, w_061_1118, w_061_1119, w_061_1120, w_061_1121, w_061_1122, w_061_1123, w_061_1125, w_061_1126, w_061_1127, w_061_1128, w_061_1129, w_061_1130, w_061_1131, w_061_1132, w_061_1133, w_061_1134, w_061_1135, w_061_1136, w_061_1137, w_061_1138, w_061_1139, w_061_1140, w_061_1141, w_061_1142, w_061_1143, w_061_1144, w_061_1145, w_061_1146, w_061_1147, w_061_1148, w_061_1149, w_061_1150, w_061_1151, w_061_1152, w_061_1153, w_061_1154, w_061_1155, w_061_1156, w_061_1157, w_061_1158, w_061_1160, w_061_1161, w_061_1162, w_061_1163, w_061_1164, w_061_1165, w_061_1166, w_061_1167, w_061_1168, w_061_1169, w_061_1170, w_061_1171, w_061_1172, w_061_1173, w_061_1174, w_061_1175, w_061_1176, w_061_1177, w_061_1178, w_061_1179, w_061_1180, w_061_1181, w_061_1182, w_061_1183, w_061_1184, w_061_1185, w_061_1186, w_061_1187, w_061_1188, w_061_1189, w_061_1190, w_061_1191, w_061_1192, w_061_1193, w_061_1194, w_061_1196, w_061_1197, w_061_1198, w_061_1199, w_061_1200, w_061_1201, w_061_1202, w_061_1203, w_061_1204, w_061_1205, w_061_1206, w_061_1207, w_061_1208, w_061_1209, w_061_1210, w_061_1211, w_061_1212, w_061_1213, w_061_1214, w_061_1215, w_061_1216, w_061_1217, w_061_1218, w_061_1219, w_061_1220, w_061_1221, w_061_1222, w_061_1223, w_061_1224, w_061_1225, w_061_1226, w_061_1227, w_061_1228, w_061_1229, w_061_1230, w_061_1231, w_061_1232, w_061_1233, w_061_1234, w_061_1235, w_061_1236, w_061_1237, w_061_1238, w_061_1239, w_061_1240, w_061_1241, w_061_1242, w_061_1243, w_061_1244, w_061_1245, w_061_1246, w_061_1247, w_061_1248, w_061_1249, w_061_1250, w_061_1251, w_061_1252, w_061_1253, w_061_1254, w_061_1255, w_061_1256, w_061_1257, w_061_1258, w_061_1259, w_061_1260, w_061_1261, w_061_1262, w_061_1263, w_061_1264, w_061_1265, w_061_1266, w_061_1267, w_061_1268, w_061_1270, w_061_1271, w_061_1272, w_061_1273, w_061_1274, w_061_1275, w_061_1276, w_061_1277, w_061_1278, w_061_1279, w_061_1280, w_061_1281, w_061_1282, w_061_1283, w_061_1284, w_061_1286, w_061_1287, w_061_1288, w_061_1289, w_061_1290, w_061_1291, w_061_1292, w_061_1293, w_061_1294, w_061_1295, w_061_1296, w_061_1297, w_061_1298, w_061_1299, w_061_1300, w_061_1301, w_061_1302, w_061_1303, w_061_1304, w_061_1305, w_061_1306, w_061_1307, w_061_1308, w_061_1309, w_061_1310, w_061_1311, w_061_1312, w_061_1313, w_061_1314, w_061_1315, w_061_1316, w_061_1318, w_061_1319, w_061_1320, w_061_1321, w_061_1322, w_061_1323, w_061_1324, w_061_1325, w_061_1326, w_061_1327, w_061_1328, w_061_1329, w_061_1330, w_061_1331, w_061_1332, w_061_1333, w_061_1334, w_061_1335, w_061_1336, w_061_1337, w_061_1338, w_061_1339, w_061_1340, w_061_1341, w_061_1342, w_061_1343, w_061_1344, w_061_1345, w_061_1346, w_061_1347, w_061_1348, w_061_1349, w_061_1350, w_061_1351, w_061_1352, w_061_1353, w_061_1354, w_061_1355, w_061_1356, w_061_1357, w_061_1358, w_061_1359, w_061_1360, w_061_1361, w_061_1362, w_061_1363, w_061_1364, w_061_1365, w_061_1366, w_061_1367, w_061_1368, w_061_1369, w_061_1371, w_061_1372, w_061_1373, w_061_1374, w_061_1375, w_061_1376, w_061_1377, w_061_1378, w_061_1379, w_061_1380, w_061_1381, w_061_1382, w_061_1383, w_061_1384, w_061_1385, w_061_1386, w_061_1387, w_061_1388, w_061_1389, w_061_1390, w_061_1391, w_061_1392, w_061_1393, w_061_1394, w_061_1396, w_061_1397, w_061_1398, w_061_1399, w_061_1400, w_061_1401;
  wire w_062_004, w_062_005, w_062_012, w_062_014, w_062_015, w_062_016, w_062_017, w_062_018, w_062_020, w_062_022, w_062_023, w_062_024, w_062_026, w_062_027, w_062_032, w_062_033, w_062_036, w_062_037, w_062_038, w_062_039, w_062_042, w_062_045, w_062_047, w_062_049, w_062_050, w_062_051, w_062_052, w_062_053, w_062_054, w_062_056, w_062_057, w_062_059, w_062_060, w_062_061, w_062_062, w_062_064, w_062_066, w_062_067, w_062_068, w_062_071, w_062_072, w_062_075, w_062_077, w_062_079, w_062_080, w_062_081, w_062_083, w_062_084, w_062_085, w_062_088, w_062_090, w_062_092, w_062_093, w_062_096, w_062_098, w_062_099, w_062_100, w_062_101, w_062_102, w_062_103, w_062_107, w_062_108, w_062_109, w_062_110, w_062_112, w_062_114, w_062_115, w_062_116, w_062_119, w_062_121, w_062_123, w_062_124, w_062_125, w_062_126, w_062_127, w_062_128, w_062_130, w_062_131, w_062_132, w_062_134, w_062_137, w_062_138, w_062_139, w_062_140, w_062_143, w_062_144, w_062_147, w_062_148, w_062_149, w_062_151, w_062_152, w_062_154, w_062_157, w_062_158, w_062_159, w_062_160, w_062_162, w_062_163, w_062_165, w_062_166, w_062_168, w_062_173, w_062_174, w_062_176, w_062_177, w_062_178, w_062_180, w_062_182, w_062_184, w_062_186, w_062_188, w_062_189, w_062_191, w_062_192, w_062_195, w_062_199, w_062_200, w_062_201, w_062_203, w_062_204, w_062_205, w_062_207, w_062_210, w_062_211, w_062_212, w_062_214, w_062_215, w_062_216, w_062_217, w_062_218, w_062_220, w_062_223, w_062_225, w_062_226, w_062_228, w_062_234, w_062_235, w_062_237, w_062_242, w_062_243, w_062_244, w_062_246, w_062_248, w_062_249, w_062_250, w_062_251, w_062_252, w_062_254, w_062_255, w_062_256, w_062_257, w_062_258, w_062_259, w_062_260, w_062_261, w_062_264, w_062_265, w_062_266, w_062_268, w_062_269, w_062_270, w_062_271, w_062_275, w_062_276, w_062_277, w_062_278, w_062_281, w_062_282, w_062_283, w_062_284, w_062_285, w_062_286, w_062_289, w_062_290, w_062_291, w_062_292, w_062_293, w_062_294, w_062_295, w_062_298, w_062_299, w_062_304, w_062_305, w_062_306, w_062_307, w_062_308, w_062_309, w_062_313, w_062_316, w_062_320, w_062_321, w_062_322, w_062_323, w_062_324, w_062_325, w_062_329, w_062_330, w_062_331, w_062_332, w_062_333, w_062_335, w_062_336, w_062_337, w_062_338, w_062_339, w_062_341, w_062_344, w_062_348, w_062_349, w_062_351, w_062_353, w_062_355, w_062_358, w_062_361, w_062_364, w_062_365, w_062_367, w_062_368, w_062_372, w_062_375, w_062_377, w_062_382, w_062_388, w_062_389, w_062_390, w_062_393, w_062_394, w_062_395, w_062_397, w_062_399, w_062_400, w_062_402, w_062_403, w_062_404, w_062_408, w_062_409, w_062_410, w_062_412, w_062_413, w_062_417, w_062_418, w_062_419, w_062_421, w_062_422, w_062_423, w_062_424, w_062_426, w_062_427, w_062_429, w_062_430, w_062_432, w_062_434, w_062_435, w_062_436, w_062_439, w_062_440, w_062_441, w_062_443, w_062_445, w_062_450, w_062_451, w_062_452, w_062_454, w_062_455, w_062_457, w_062_458, w_062_459, w_062_461, w_062_462, w_062_463, w_062_464, w_062_465, w_062_466, w_062_468, w_062_469, w_062_470, w_062_471, w_062_473, w_062_474, w_062_475, w_062_476, w_062_477, w_062_478, w_062_479, w_062_480, w_062_482, w_062_483, w_062_484, w_062_486, w_062_487, w_062_488, w_062_489, w_062_490, w_062_491, w_062_492, w_062_493, w_062_495, w_062_496, w_062_497, w_062_498, w_062_499, w_062_500, w_062_501, w_062_503, w_062_507, w_062_508, w_062_509, w_062_511, w_062_513, w_062_515, w_062_520, w_062_521, w_062_522, w_062_523, w_062_526, w_062_527, w_062_528, w_062_530, w_062_531, w_062_533, w_062_535, w_062_539, w_062_542, w_062_543, w_062_544, w_062_546, w_062_551, w_062_554, w_062_555, w_062_556, w_062_558, w_062_559, w_062_561, w_062_562, w_062_563, w_062_564, w_062_567, w_062_571, w_062_572, w_062_573, w_062_574, w_062_575, w_062_576, w_062_578, w_062_579, w_062_584, w_062_586, w_062_589, w_062_590, w_062_591, w_062_593, w_062_594, w_062_595, w_062_598, w_062_599, w_062_601, w_062_603, w_062_604, w_062_605, w_062_606, w_062_608, w_062_609, w_062_610, w_062_611, w_062_614, w_062_616, w_062_618, w_062_619, w_062_620, w_062_623, w_062_625, w_062_626, w_062_629, w_062_632, w_062_633, w_062_636, w_062_638, w_062_639, w_062_642, w_062_643, w_062_649, w_062_650, w_062_652, w_062_657, w_062_658, w_062_661, w_062_664, w_062_666, w_062_667, w_062_668, w_062_669, w_062_670, w_062_672, w_062_674, w_062_676, w_062_679, w_062_683, w_062_687, w_062_689, w_062_692, w_062_694, w_062_696, w_062_697, w_062_699, w_062_703, w_062_704, w_062_706, w_062_708, w_062_709, w_062_712, w_062_713, w_062_714, w_062_715, w_062_716, w_062_717, w_062_718, w_062_719, w_062_721, w_062_722, w_062_724, w_062_725, w_062_726, w_062_730, w_062_731, w_062_732, w_062_733, w_062_735, w_062_737, w_062_740, w_062_741, w_062_743, w_062_744, w_062_745, w_062_748, w_062_749, w_062_751, w_062_752, w_062_754, w_062_757, w_062_758, w_062_759, w_062_760, w_062_764, w_062_767, w_062_768, w_062_769, w_062_772, w_062_774, w_062_776, w_062_777, w_062_778, w_062_781, w_062_782, w_062_785, w_062_786, w_062_787, w_062_788, w_062_789, w_062_792, w_062_793, w_062_794, w_062_796, w_062_798, w_062_799, w_062_800, w_062_802, w_062_803, w_062_804, w_062_806, w_062_807, w_062_808, w_062_810, w_062_811, w_062_812, w_062_818, w_062_820, w_062_821, w_062_822, w_062_824, w_062_827, w_062_829, w_062_830, w_062_831, w_062_832, w_062_834, w_062_835, w_062_836, w_062_837, w_062_839, w_062_841, w_062_842, w_062_843, w_062_845, w_062_846, w_062_847, w_062_848, w_062_849, w_062_850, w_062_851, w_062_852, w_062_853, w_062_854, w_062_859, w_062_860, w_062_861, w_062_862, w_062_863, w_062_867, w_062_868, w_062_869, w_062_873, w_062_874, w_062_875, w_062_876, w_062_877, w_062_878, w_062_879, w_062_880, w_062_883, w_062_885, w_062_886, w_062_888, w_062_890, w_062_893, w_062_894, w_062_897, w_062_898, w_062_899, w_062_900, w_062_901, w_062_905, w_062_906, w_062_909, w_062_911, w_062_912, w_062_913, w_062_915, w_062_920, w_062_921, w_062_922, w_062_924, w_062_926, w_062_928, w_062_929, w_062_930, w_062_933, w_062_934, w_062_935, w_062_937, w_062_938, w_062_939, w_062_940, w_062_942, w_062_943, w_062_944, w_062_946, w_062_948, w_062_949, w_062_951, w_062_952, w_062_953, w_062_955, w_062_956, w_062_961, w_062_962, w_062_963, w_062_965, w_062_966, w_062_968, w_062_971, w_062_973, w_062_974, w_062_975, w_062_977, w_062_978, w_062_983, w_062_984, w_062_985, w_062_986, w_062_988, w_062_991, w_062_992, w_062_993, w_062_994, w_062_995, w_062_996, w_062_997, w_062_998, w_062_1000, w_062_1001, w_062_1002, w_062_1003, w_062_1004, w_062_1006, w_062_1007, w_062_1008, w_062_1010, w_062_1011, w_062_1012, w_062_1014, w_062_1015, w_062_1016, w_062_1018, w_062_1019, w_062_1020, w_062_1022, w_062_1023, w_062_1024, w_062_1025, w_062_1026, w_062_1028, w_062_1030, w_062_1031, w_062_1035, w_062_1036, w_062_1038, w_062_1039, w_062_1040, w_062_1042, w_062_1043, w_062_1044, w_062_1046, w_062_1048, w_062_1053, w_062_1056, w_062_1058, w_062_1059, w_062_1061, w_062_1063, w_062_1064, w_062_1065, w_062_1069, w_062_1070, w_062_1071, w_062_1072, w_062_1077, w_062_1080, w_062_1081, w_062_1084, w_062_1085, w_062_1088, w_062_1090, w_062_1091, w_062_1093, w_062_1094, w_062_1097, w_062_1100, w_062_1101, w_062_1102, w_062_1103, w_062_1105, w_062_1108, w_062_1109, w_062_1110, w_062_1111, w_062_1112, w_062_1113, w_062_1114, w_062_1115, w_062_1116, w_062_1118, w_062_1123, w_062_1124, w_062_1126, w_062_1127, w_062_1129, w_062_1130, w_062_1131, w_062_1135, w_062_1137, w_062_1138, w_062_1140, w_062_1141, w_062_1145, w_062_1146, w_062_1147, w_062_1149, w_062_1151, w_062_1152, w_062_1153, w_062_1154, w_062_1156, w_062_1157, w_062_1158, w_062_1159, w_062_1160, w_062_1165, w_062_1167, w_062_1170, w_062_1171, w_062_1175, w_062_1176, w_062_1178, w_062_1179, w_062_1181, w_062_1183, w_062_1185, w_062_1186, w_062_1187, w_062_1188, w_062_1189, w_062_1191, w_062_1192, w_062_1193, w_062_1194, w_062_1195, w_062_1196, w_062_1197, w_062_1198, w_062_1199, w_062_1200, w_062_1201, w_062_1203, w_062_1205, w_062_1206, w_062_1207, w_062_1208, w_062_1211, w_062_1212, w_062_1214, w_062_1216, w_062_1217, w_062_1218, w_062_1219, w_062_1220, w_062_1221, w_062_1223, w_062_1224, w_062_1226, w_062_1228, w_062_1229, w_062_1232, w_062_1233, w_062_1235, w_062_1236, w_062_1238, w_062_1241, w_062_1242, w_062_1243, w_062_1244, w_062_1245, w_062_1246, w_062_1247, w_062_1248, w_062_1252, w_062_1255, w_062_1259, w_062_1260, w_062_1262, w_062_1264, w_062_1265, w_062_1267, w_062_1268, w_062_1269, w_062_1270, w_062_1271, w_062_1272, w_062_1274, w_062_1277, w_062_1282, w_062_1283, w_062_1284, w_062_1285, w_062_1287, w_062_1288, w_062_1293, w_062_1294, w_062_1296, w_062_1300, w_062_1302, w_062_1303, w_062_1304, w_062_1305, w_062_1307, w_062_1310, w_062_1314, w_062_1315, w_062_1318, w_062_1319, w_062_1320, w_062_1322, w_062_1324, w_062_1326, w_062_1327, w_062_1328, w_062_1331, w_062_1333, w_062_1334, w_062_1336, w_062_1337, w_062_1339, w_062_1340, w_062_1343, w_062_1346, w_062_1347, w_062_1348, w_062_1349, w_062_1351, w_062_1353, w_062_1354, w_062_1355, w_062_1356, w_062_1358, w_062_1359, w_062_1362, w_062_1364, w_062_1366, w_062_1367, w_062_1370, w_062_1373, w_062_1375, w_062_1376, w_062_1377, w_062_1379, w_062_1382, w_062_1385, w_062_1386, w_062_1388, w_062_1389, w_062_1390, w_062_1391, w_062_1392, w_062_1396, w_062_1397, w_062_1398, w_062_1399, w_062_1402, w_062_1403, w_062_1404, w_062_1405, w_062_1407, w_062_1408, w_062_1409, w_062_1412, w_062_1414, w_062_1415, w_062_1416, w_062_1417, w_062_1422, w_062_1423, w_062_1424, w_062_1426, w_062_1427, w_062_1428, w_062_1431, w_062_1434, w_062_1435, w_062_1438, w_062_1439, w_062_1442, w_062_1444, w_062_1445, w_062_1447, w_062_1449, w_062_1452, w_062_1453, w_062_1454, w_062_1456, w_062_1457, w_062_1458, w_062_1459, w_062_1460, w_062_1461, w_062_1464, w_062_1465, w_062_1466, w_062_1468, w_062_1471, w_062_1472, w_062_1474, w_062_1477, w_062_1478, w_062_1479, w_062_1482, w_062_1484, w_062_1487, w_062_1490, w_062_1491, w_062_1495, w_062_1496, w_062_1497, w_062_1498, w_062_1500, w_062_1502, w_062_1504, w_062_1506, w_062_1507, w_062_1508, w_062_1511, w_062_1518, w_062_1519, w_062_1521, w_062_1522, w_062_1524, w_062_1525, w_062_1526, w_062_1527, w_062_1531, w_062_1532, w_062_1533, w_062_1535, w_062_1536, w_062_1537, w_062_1538, w_062_1539, w_062_1541, w_062_1542, w_062_1543, w_062_1545, w_062_1546, w_062_1547, w_062_1548, w_062_1550, w_062_1551, w_062_1552, w_062_1553, w_062_1554, w_062_1556, w_062_1559, w_062_1561, w_062_1562, w_062_1563, w_062_1564, w_062_1565, w_062_1567, w_062_1568, w_062_1571, w_062_1572, w_062_1573, w_062_1574, w_062_1575, w_062_1577, w_062_1582, w_062_1588, w_062_1589, w_062_1595, w_062_1596, w_062_1599, w_062_1601, w_062_1602, w_062_1604, w_062_1607, w_062_1608, w_062_1611, w_062_1613, w_062_1616, w_062_1620, w_062_1621, w_062_1622, w_062_1623, w_062_1625, w_062_1626, w_062_1628, w_062_1629, w_062_1630, w_062_1631, w_062_1632, w_062_1634, w_062_1636, w_062_1637, w_062_1638, w_062_1639, w_062_1640, w_062_1641, w_062_1642, w_062_1643, w_062_1644, w_062_1646, w_062_1647, w_062_1649, w_062_1650, w_062_1651, w_062_1652, w_062_1654, w_062_1655, w_062_1656, w_062_1657, w_062_1659, w_062_1660, w_062_1662, w_062_1664, w_062_1665, w_062_1668, w_062_1669, w_062_1670, w_062_1674, w_062_1675, w_062_1676, w_062_1677, w_062_1678, w_062_1683, w_062_1684, w_062_1685, w_062_1686, w_062_1690, w_062_1691, w_062_1692, w_062_1694, w_062_1695, w_062_1696, w_062_1698, w_062_1699, w_062_1703, w_062_1704, w_062_1705, w_062_1706, w_062_1707, w_062_1708, w_062_1710, w_062_1712, w_062_1713, w_062_1715, w_062_1717, w_062_1718, w_062_1721, w_062_1724, w_062_1726, w_062_1727, w_062_1732, w_062_1734, w_062_1739, w_062_1740, w_062_1741, w_062_1742, w_062_1743, w_062_1744, w_062_1745, w_062_1746, w_062_1747, w_062_1748, w_062_1749, w_062_1750, w_062_1752, w_062_1755, w_062_1757, w_062_1759, w_062_1760, w_062_1761, w_062_1762, w_062_1763, w_062_1764, w_062_1765, w_062_1766, w_062_1767, w_062_1768, w_062_1771, w_062_1775, w_062_1776, w_062_1777, w_062_1778, w_062_1780, w_062_1781, w_062_1784, w_062_1786, w_062_1787, w_062_1788, w_062_1789, w_062_1792, w_062_1794, w_062_1795, w_062_1797, w_062_1800, w_062_1801, w_062_1802, w_062_1803, w_062_1804, w_062_1806, w_062_1807, w_062_1808, w_062_1810, w_062_1811, w_062_1813, w_062_1815, w_062_1816, w_062_1817, w_062_1818, w_062_1819, w_062_1822, w_062_1823, w_062_1824, w_062_1825, w_062_1828, w_062_1829, w_062_1830, w_062_1831, w_062_1832, w_062_1834, w_062_1835, w_062_1836, w_062_1839, w_062_1841, w_062_1843, w_062_1845, w_062_1846, w_062_1847, w_062_1849, w_062_1850, w_062_1851, w_062_1852, w_062_1853, w_062_1854, w_062_1856, w_062_1860, w_062_1861, w_062_1862, w_062_1863, w_062_1864, w_062_1865, w_062_1866, w_062_1868, w_062_1869, w_062_1872, w_062_1873, w_062_1874, w_062_1879, w_062_1880, w_062_1882, w_062_1884, w_062_1885, w_062_1887, w_062_1888, w_062_1890, w_062_1891, w_062_1893, w_062_1894, w_062_1895, w_062_1896, w_062_1897, w_062_1898, w_062_1902, w_062_1906, w_062_1907, w_062_1908, w_062_1909, w_062_1910, w_062_1912, w_062_1913, w_062_1917, w_062_1921, w_062_1922, w_062_1924, w_062_1925, w_062_1926, w_062_1929, w_062_1930, w_062_1937, w_062_1938, w_062_1939, w_062_1941, w_062_1943, w_062_1944, w_062_1946, w_062_1947, w_062_1948, w_062_1949, w_062_1950, w_062_1953, w_062_1955, w_062_1957, w_062_1958, w_062_1963, w_062_1965, w_062_1966, w_062_1967, w_062_1969, w_062_1971, w_062_1972, w_062_1974, w_062_1975, w_062_1976, w_062_1978, w_062_1979, w_062_1980, w_062_1982, w_062_1984, w_062_1985, w_062_1986, w_062_1987, w_062_1988, w_062_1989, w_062_1990, w_062_1993, w_062_1995, w_062_1996, w_062_1998, w_062_2003, w_062_2005, w_062_2008, w_062_2010, w_062_2013, w_062_2014, w_062_2015, w_062_2016, w_062_2017, w_062_2018, w_062_2020, w_062_2025, w_062_2026, w_062_2028, w_062_2029, w_062_2030, w_062_2033, w_062_2034, w_062_2035, w_062_2036, w_062_2042, w_062_2044, w_062_2046, w_062_2049, w_062_2051, w_062_2052, w_062_2054, w_062_2057, w_062_2058, w_062_2059, w_062_2060, w_062_2061, w_062_2063, w_062_2064, w_062_2068, w_062_2069, w_062_2070, w_062_2071, w_062_2074, w_062_2075, w_062_2076, w_062_2077, w_062_2078, w_062_2079, w_062_2080, w_062_2081, w_062_2083, w_062_2084, w_062_2085, w_062_2088, w_062_2089, w_062_2092, w_062_2093, w_062_2094, w_062_2097, w_062_2099, w_062_2100, w_062_2101, w_062_2102, w_062_2103, w_062_2105, w_062_2106, w_062_2108, w_062_2109, w_062_2110, w_062_2112, w_062_2113, w_062_2114, w_062_2115, w_062_2116, w_062_2118, w_062_2119, w_062_2122, w_062_2127, w_062_2129, w_062_2130, w_062_2131, w_062_2132, w_062_2133, w_062_2134, w_062_2136, w_062_2137, w_062_2138, w_062_2140, w_062_2141, w_062_2142, w_062_2144, w_062_2146, w_062_2151, w_062_2152, w_062_2154, w_062_2155, w_062_2156, w_062_2157, w_062_2158, w_062_2159, w_062_2161, w_062_2162, w_062_2164, w_062_2165, w_062_2166, w_062_2169, w_062_2170, w_062_2171, w_062_2174, w_062_2175, w_062_2176, w_062_2177, w_062_2178, w_062_2180, w_062_2181, w_062_2184, w_062_2187, w_062_2189, w_062_2190, w_062_2191, w_062_2192, w_062_2193, w_062_2194, w_062_2195, w_062_2196, w_062_2198, w_062_2199, w_062_2200, w_062_2202, w_062_2203, w_062_2204, w_062_2206, w_062_2207, w_062_2208, w_062_2209, w_062_2210, w_062_2211, w_062_2212, w_062_2214, w_062_2216, w_062_2219, w_062_2220, w_062_2222, w_062_2223, w_062_2228, w_062_2229, w_062_2230, w_062_2231, w_062_2232, w_062_2233, w_062_2234, w_062_2236, w_062_2240, w_062_2241, w_062_2242, w_062_2243, w_062_2245, w_062_2246, w_062_2248, w_062_2250, w_062_2251, w_062_2253, w_062_2254, w_062_2256, w_062_2259, w_062_2262, w_062_2265, w_062_2267, w_062_2268, w_062_2269, w_062_2272, w_062_2274, w_062_2275, w_062_2278, w_062_2280, w_062_2282, w_062_2283, w_062_2284, w_062_2285, w_062_2288, w_062_2289, w_062_2291, w_062_2292, w_062_2293, w_062_2295, w_062_2296, w_062_2297, w_062_2298, w_062_2299, w_062_2300, w_062_2301, w_062_2304, w_062_2306, w_062_2308, w_062_2309, w_062_2310, w_062_2313, w_062_2320, w_062_2321, w_062_2325, w_062_2327, w_062_2328, w_062_2329, w_062_2331, w_062_2333, w_062_2335, w_062_2341, w_062_2343, w_062_2344, w_062_2345, w_062_2347, w_062_2351, w_062_2352, w_062_2353, w_062_2354, w_062_2355, w_062_2356, w_062_2357, w_062_2361, w_062_2363, w_062_2364, w_062_2365, w_062_2367, w_062_2370, w_062_2371, w_062_2373, w_062_2374, w_062_2375, w_062_2376, w_062_2378, w_062_2379, w_062_2380, w_062_2384, w_062_2385, w_062_2386, w_062_2387, w_062_2388, w_062_2391, w_062_2392, w_062_2394, w_062_2395, w_062_2398, w_062_2399, w_062_2400, w_062_2401, w_062_2404, w_062_2406, w_062_2409, w_062_2415, w_062_2416, w_062_2417, w_062_2418, w_062_2419, w_062_2420, w_062_2421, w_062_2424, w_062_2426, w_062_2427, w_062_2430, w_062_2435, w_062_2436, w_062_2437, w_062_2439, w_062_2440, w_062_2443, w_062_2444, w_062_2445, w_062_2446, w_062_2449, w_062_2452, w_062_2453, w_062_2454, w_062_2455, w_062_2456, w_062_2458, w_062_2459, w_062_2460, w_062_2461, w_062_2462, w_062_2464, w_062_2465, w_062_2466, w_062_2467, w_062_2469, w_062_2471, w_062_2472, w_062_2474, w_062_2478, w_062_2479, w_062_2480, w_062_2482, w_062_2486, w_062_2488, w_062_2491, w_062_2495, w_062_2496, w_062_2498, w_062_2501, w_062_2502, w_062_2505, w_062_2508, w_062_2509, w_062_2510, w_062_2511, w_062_2515, w_062_2516, w_062_2517, w_062_2520, w_062_2521, w_062_2523, w_062_2525, w_062_2526, w_062_2527, w_062_2529, w_062_2530, w_062_2531, w_062_2532, w_062_2535, w_062_2537, w_062_2538, w_062_2540, w_062_2541, w_062_2543, w_062_2544, w_062_2546, w_062_2547, w_062_2550, w_062_2551, w_062_2553, w_062_2554, w_062_2555, w_062_2557, w_062_2558, w_062_2560, w_062_2561, w_062_2563, w_062_2564, w_062_2565, w_062_2566, w_062_2568, w_062_2569, w_062_2570, w_062_2571, w_062_2572, w_062_2573, w_062_2574, w_062_2576, w_062_2579, w_062_2580, w_062_2581, w_062_2586, w_062_2587, w_062_2591, w_062_2594, w_062_2595, w_062_2596, w_062_2597, w_062_2598, w_062_2599, w_062_2601, w_062_2602, w_062_2604, w_062_2605, w_062_2606, w_062_2607, w_062_2608, w_062_2609, w_062_2610, w_062_2611, w_062_2616, w_062_2618, w_062_2619, w_062_2622, w_062_2623, w_062_2624, w_062_2625, w_062_2627, w_062_2628, w_062_2629, w_062_2630, w_062_2631, w_062_2632, w_062_2636, w_062_2637, w_062_2638, w_062_2642, w_062_2643, w_062_2644, w_062_2645, w_062_2646, w_062_2647, w_062_2650, w_062_2652, w_062_2654, w_062_2658, w_062_2659, w_062_2660, w_062_2664, w_062_2669, w_062_2670, w_062_2671, w_062_2676, w_062_2678, w_062_2680, w_062_2681, w_062_2682, w_062_2687, w_062_2688, w_062_2689, w_062_2690, w_062_2691, w_062_2700, w_062_2704, w_062_2705, w_062_2707, w_062_2709, w_062_2717, w_062_2719, w_062_2723, w_062_2725, w_062_2728, w_062_2729, w_062_2734, w_062_2736, w_062_2737, w_062_2743, w_062_2745, w_062_2746, w_062_2748, w_062_2749, w_062_2752, w_062_2753, w_062_2754, w_062_2756, w_062_2758, w_062_2760, w_062_2761, w_062_2762, w_062_2768, w_062_2775, w_062_2776, w_062_2785, w_062_2790, w_062_2792, w_062_2795, w_062_2797, w_062_2798, w_062_2801, w_062_2803, w_062_2807, w_062_2811, w_062_2813, w_062_2814, w_062_2820, w_062_2821, w_062_2824, w_062_2825, w_062_2826, w_062_2827, w_062_2831, w_062_2832, w_062_2833, w_062_2835, w_062_2840, w_062_2844, w_062_2848, w_062_2851, w_062_2853, w_062_2859, w_062_2866, w_062_2871, w_062_2872, w_062_2875, w_062_2878, w_062_2879, w_062_2881, w_062_2883, w_062_2884, w_062_2887, w_062_2898, w_062_2899, w_062_2901, w_062_2905, w_062_2906, w_062_2908, w_062_2909, w_062_2910, w_062_2911, w_062_2915, w_062_2920, w_062_2921, w_062_2924, w_062_2925, w_062_2926, w_062_2927, w_062_2928, w_062_2938, w_062_2942, w_062_2946, w_062_2947, w_062_2950, w_062_2953, w_062_2954, w_062_2955, w_062_2956, w_062_2957, w_062_2959, w_062_2960, w_062_2961, w_062_2962, w_062_2963, w_062_2964, w_062_2966, w_062_2968, w_062_2975, w_062_2976, w_062_2980, w_062_2983, w_062_2986, w_062_2987, w_062_2989, w_062_2991, w_062_2994, w_062_2999, w_062_3000, w_062_3003, w_062_3005, w_062_3006, w_062_3009, w_062_3010, w_062_3012, w_062_3014, w_062_3015, w_062_3017, w_062_3019, w_062_3023, w_062_3024, w_062_3025, w_062_3026, w_062_3027, w_062_3028, w_062_3029, w_062_3031, w_062_3032, w_062_3033, w_062_3041, w_062_3042, w_062_3047, w_062_3048, w_062_3053, w_062_3054, w_062_3059, w_062_3060, w_062_3065, w_062_3069, w_062_3070, w_062_3074, w_062_3075, w_062_3087, w_062_3089, w_062_3094, w_062_3096, w_062_3097, w_062_3099, w_062_3106, w_062_3108, w_062_3113, w_062_3116, w_062_3118, w_062_3119, w_062_3123, w_062_3124, w_062_3126, w_062_3129, w_062_3130, w_062_3131, w_062_3132, w_062_3140, w_062_3143, w_062_3144, w_062_3147, w_062_3150, w_062_3152, w_062_3154, w_062_3156, w_062_3157, w_062_3161, w_062_3162, w_062_3165, w_062_3169, w_062_3170, w_062_3171, w_062_3172, w_062_3175, w_062_3176, w_062_3177, w_062_3188, w_062_3189, w_062_3197, w_062_3199, w_062_3210, w_062_3211, w_062_3212, w_062_3215, w_062_3219, w_062_3224, w_062_3228, w_062_3230, w_062_3231, w_062_3235, w_062_3245, w_062_3246, w_062_3252, w_062_3256, w_062_3257, w_062_3258, w_062_3259, w_062_3262, w_062_3269, w_062_3274, w_062_3278, w_062_3280, w_062_3284, w_062_3287, w_062_3292, w_062_3296, w_062_3299, w_062_3301, w_062_3302, w_062_3303, w_062_3308, w_062_3309, w_062_3310, w_062_3313, w_062_3315, w_062_3319, w_062_3322, w_062_3324, w_062_3325, w_062_3326, w_062_3327, w_062_3328, w_062_3330, w_062_3331, w_062_3334, w_062_3335, w_062_3336, w_062_3338, w_062_3339, w_062_3340, w_062_3341, w_062_3344, w_062_3345, w_062_3346, w_062_3349, w_062_3351, w_062_3353, w_062_3354, w_062_3359, w_062_3360, w_062_3362, w_062_3365, w_062_3368, w_062_3370, w_062_3373, w_062_3375, w_062_3376, w_062_3382, w_062_3383, w_062_3384, w_062_3386, w_062_3387, w_062_3396, w_062_3401, w_062_3407, w_062_3412, w_062_3419, w_062_3423, w_062_3424, w_062_3425, w_062_3429, w_062_3433, w_062_3435, w_062_3440, w_062_3441, w_062_3446, w_062_3450, w_062_3451, w_062_3456, w_062_3457, w_062_3463, w_062_3465, w_062_3467, w_062_3468, w_062_3470, w_062_3471, w_062_3476, w_062_3477, w_062_3479, w_062_3482, w_062_3486, w_062_3492, w_062_3498, w_062_3499, w_062_3501, w_062_3502, w_062_3503, w_062_3506, w_062_3508, w_062_3511, w_062_3523, w_062_3524, w_062_3528, w_062_3529, w_062_3530, w_062_3531, w_062_3533, w_062_3539, w_062_3541, w_062_3544, w_062_3548, w_062_3549, w_062_3556, w_062_3557, w_062_3560, w_062_3561, w_062_3562, w_062_3564, w_062_3574, w_062_3576, w_062_3579, w_062_3580, w_062_3582, w_062_3596, w_062_3598, w_062_3599, w_062_3602, w_062_3604, w_062_3607, w_062_3608, w_062_3610, w_062_3612, w_062_3617, w_062_3618, w_062_3620, w_062_3622, w_062_3626, w_062_3627, w_062_3628, w_062_3631, w_062_3635, w_062_3636, w_062_3639, w_062_3642, w_062_3643, w_062_3653, w_062_3655, w_062_3656, w_062_3659, w_062_3661, w_062_3664, w_062_3666, w_062_3668, w_062_3671, w_062_3673, w_062_3676, w_062_3677, w_062_3682, w_062_3686, w_062_3692, w_062_3693, w_062_3694, w_062_3695, w_062_3696, w_062_3697, w_062_3699, w_062_3700, w_062_3706, w_062_3710, w_062_3711, w_062_3712, w_062_3718, w_062_3719, w_062_3724, w_062_3728, w_062_3729, w_062_3732, w_062_3733, w_062_3734, w_062_3735, w_062_3738, w_062_3739, w_062_3754, w_062_3764, w_062_3766, w_062_3769, w_062_3775, w_062_3778, w_062_3785, w_062_3791, w_062_3793, w_062_3796, w_062_3797, w_062_3800, w_062_3801, w_062_3807, w_062_3811, w_062_3814, w_062_3816, w_062_3818, w_062_3820, w_062_3822, w_062_3828, w_062_3830, w_062_3843, w_062_3845, w_062_3846, w_062_3847, w_062_3848, w_062_3849, w_062_3850, w_062_3851, w_062_3852, w_062_3853, w_062_3855, w_062_3858, w_062_3861, w_062_3863, w_062_3869, w_062_3872, w_062_3874, w_062_3879, w_062_3882, w_062_3887, w_062_3888, w_062_3890, w_062_3892, w_062_3893, w_062_3901, w_062_3904, w_062_3906, w_062_3907, w_062_3911, w_062_3912, w_062_3913, w_062_3918, w_062_3921, w_062_3923, w_062_3924, w_062_3928, w_062_3929, w_062_3930, w_062_3932, w_062_3940, w_062_3941, w_062_3945, w_062_3946, w_062_3948, w_062_3954, w_062_3955, w_062_3957, w_062_3958, w_062_3959, w_062_3961, w_062_3971, w_062_3973, w_062_3980, w_062_3982, w_062_3988, w_062_3993, w_062_3994, w_062_3997, w_062_3998, w_062_4001, w_062_4002, w_062_4006, w_062_4012, w_062_4018, w_062_4020, w_062_4022, w_062_4023, w_062_4027, w_062_4030, w_062_4035, w_062_4037, w_062_4038, w_062_4039, w_062_4040, w_062_4043, w_062_4044, w_062_4045, w_062_4047, w_062_4049, w_062_4051, w_062_4055, w_062_4056, w_062_4057, w_062_4059, w_062_4060, w_062_4064, w_062_4071, w_062_4075, w_062_4076, w_062_4077, w_062_4080, w_062_4083, w_062_4084, w_062_4086, w_062_4087, w_062_4088, w_062_4092, w_062_4094, w_062_4095, w_062_4101, w_062_4109, w_062_4113, w_062_4114, w_062_4125, w_062_4127, w_062_4129, w_062_4131, w_062_4133, w_062_4134, w_062_4139, w_062_4144, w_062_4145, w_062_4147, w_062_4149, w_062_4150, w_062_4152, w_062_4154, w_062_4155, w_062_4158, w_062_4160, w_062_4163, w_062_4165, w_062_4167, w_062_4168, w_062_4170, w_062_4175, w_062_4181, w_062_4182, w_062_4183, w_062_4189, w_062_4190, w_062_4194, w_062_4197, w_062_4199, w_062_4208, w_062_4209, w_062_4211, w_062_4212, w_062_4217, w_062_4218, w_062_4222, w_062_4227, w_062_4229, w_062_4230, w_062_4231, w_062_4232, w_062_4235, w_062_4236, w_062_4237, w_062_4240, w_062_4245, w_062_4246, w_062_4249, w_062_4257, w_062_4259, w_062_4263, w_062_4265, w_062_4269, w_062_4271, w_062_4272, w_062_4278, w_062_4281, w_062_4283, w_062_4284, w_062_4291, w_062_4294, w_062_4295, w_062_4297, w_062_4299, w_062_4309, w_062_4315, w_062_4317, w_062_4318, w_062_4319, w_062_4322, w_062_4324, w_062_4326, w_062_4327, w_062_4328, w_062_4330, w_062_4333, w_062_4335, w_062_4338, w_062_4341, w_062_4345, w_062_4347, w_062_4348, w_062_4356, w_062_4359, w_062_4360, w_062_4363, w_062_4366, w_062_4369, w_062_4372, w_062_4373, w_062_4375, w_062_4378, w_062_4380, w_062_4383, w_062_4387, w_062_4389, w_062_4390, w_062_4393, w_062_4394, w_062_4395, w_062_4397, w_062_4398, w_062_4405, w_062_4409, w_062_4410, w_062_4415, w_062_4418, w_062_4419, w_062_4421, w_062_4423, w_062_4428, w_062_4432, w_062_4434, w_062_4438, w_062_4453, w_062_4455, w_062_4456, w_062_4460, w_062_4462, w_062_4471, w_062_4473, w_062_4474, w_062_4476, w_062_4483, w_062_4484, w_062_4487, w_062_4493, w_062_4496, w_062_4501, w_062_4503, w_062_4504, w_062_4505, w_062_4506, w_062_4512, w_062_4513, w_062_4515, w_062_4516, w_062_4518, w_062_4519, w_062_4522, w_062_4525, w_062_4528, w_062_4533, w_062_4536, w_062_4538, w_062_4540, w_062_4541, w_062_4542, w_062_4550, w_062_4551, w_062_4553, w_062_4554, w_062_4558, w_062_4559, w_062_4560, w_062_4561, w_062_4562, w_062_4563, w_062_4565, w_062_4566, w_062_4567, w_062_4572, w_062_4573, w_062_4577, w_062_4581, w_062_4590, w_062_4594, w_062_4601, w_062_4602, w_062_4606, w_062_4612, w_062_4614, w_062_4615, w_062_4617, w_062_4618, w_062_4619, w_062_4621, w_062_4623, w_062_4626, w_062_4627, w_062_4628, w_062_4629, w_062_4631, w_062_4633, w_062_4634, w_062_4636, w_062_4637, w_062_4640, w_062_4641, w_062_4642, w_062_4645, w_062_4647, w_062_4649, w_062_4650, w_062_4652, w_062_4655, w_062_4658, w_062_4661, w_062_4662, w_062_4663, w_062_4664, w_062_4679, w_062_4681, w_062_4683, w_062_4685, w_062_4704, w_062_4711, w_062_4712, w_062_4715, w_062_4718, w_062_4719, w_062_4720, w_062_4723, w_062_4727, w_062_4729, w_062_4739, w_062_4743, w_062_4744, w_062_4749, w_062_4751, w_062_4754, w_062_4755, w_062_4757, w_062_4758, w_062_4760, w_062_4761, w_062_4766, w_062_4769, w_062_4770, w_062_4773, w_062_4777, w_062_4779, w_062_4782, w_062_4784, w_062_4785, w_062_4790, w_062_4791, w_062_4792, w_062_4794, w_062_4795, w_062_4798, w_062_4800, w_062_4801, w_062_4805, w_062_4809, w_062_4810, w_062_4812, w_062_4813, w_062_4814, w_062_4817, w_062_4818, w_062_4819, w_062_4830, w_062_4831, w_062_4832, w_062_4833, w_062_4834, w_062_4838, w_062_4840, w_062_4842, w_062_4845, w_062_4846, w_062_4848, w_062_4849, w_062_4850, w_062_4857, w_062_4858, w_062_4859, w_062_4862, w_062_4863, w_062_4870, w_062_4871, w_062_4873, w_062_4874, w_062_4877, w_062_4879, w_062_4882, w_062_4886, w_062_4890, w_062_4892, w_062_4894, w_062_4895, w_062_4899, w_062_4900, w_062_4903, w_062_4908, w_062_4910, w_062_4914, w_062_4916, w_062_4917, w_062_4919, w_062_4921, w_062_4922, w_062_4925, w_062_4926, w_062_4939, w_062_4945, w_062_4950, w_062_4953, w_062_4954, w_062_4959, w_062_4965, w_062_4967, w_062_4971, w_062_4975, w_062_4979, w_062_4985, w_062_4986, w_062_4990, w_062_4992, w_062_4993, w_062_4994, w_062_4996, w_062_4998, w_062_5000, w_062_5002, w_062_5004, w_062_5006, w_062_5007, w_062_5010, w_062_5011, w_062_5013, w_062_5018, w_062_5021, w_062_5022, w_062_5025, w_062_5026, w_062_5027, w_062_5028, w_062_5029, w_062_5030, w_062_5034, w_062_5035, w_062_5038, w_062_5040, w_062_5043, w_062_5050, w_062_5051, w_062_5052, w_062_5055, w_062_5056, w_062_5057, w_062_5065, w_062_5066, w_062_5067, w_062_5068, w_062_5072, w_062_5074, w_062_5076, w_062_5086, w_062_5088, w_062_5089, w_062_5092, w_062_5095, w_062_5099, w_062_5100, w_062_5103, w_062_5107, w_062_5109, w_062_5110, w_062_5112, w_062_5117, w_062_5121, w_062_5124, w_062_5127, w_062_5133, w_062_5139, w_062_5141, w_062_5143, w_062_5145, w_062_5148, w_062_5149, w_062_5150, w_062_5151, w_062_5156, w_062_5159, w_062_5160, w_062_5162, w_062_5165, w_062_5166, w_062_5173, w_062_5174, w_062_5177, w_062_5179, w_062_5180, w_062_5183, w_062_5186, w_062_5188, w_062_5191, w_062_5192, w_062_5196, w_062_5200, w_062_5202, w_062_5205, w_062_5206, w_062_5207, w_062_5211, w_062_5212, w_062_5213, w_062_5214, w_062_5220, w_062_5223, w_062_5225, w_062_5227, w_062_5235, w_062_5236, w_062_5239, w_062_5244, w_062_5250, w_062_5251, w_062_5260, w_062_5263, w_062_5264, w_062_5267, w_062_5268, w_062_5272, w_062_5273, w_062_5274, w_062_5275, w_062_5276, w_062_5279, w_062_5280, w_062_5281, w_062_5287, w_062_5289, w_062_5290, w_062_5291, w_062_5293, w_062_5294, w_062_5295, w_062_5297, w_062_5313, w_062_5315, w_062_5318, w_062_5319, w_062_5323, w_062_5326, w_062_5327, w_062_5328, w_062_5336, w_062_5337, w_062_5339, w_062_5340, w_062_5341, w_062_5346, w_062_5347, w_062_5349, w_062_5354, w_062_5358, w_062_5360, w_062_5361, w_062_5362, w_062_5365, w_062_5367, w_062_5371, w_062_5376, w_062_5377, w_062_5378, w_062_5381, w_062_5383, w_062_5384, w_062_5387, w_062_5395, w_062_5400, w_062_5404, w_062_5407, w_062_5410, w_062_5411, w_062_5412, w_062_5414, w_062_5416, w_062_5417, w_062_5421, w_062_5423, w_062_5424, w_062_5426, w_062_5428, w_062_5431, w_062_5434, w_062_5439, w_062_5441, w_062_5445, w_062_5446, w_062_5447, w_062_5451, w_062_5453, w_062_5456, w_062_5461, w_062_5462, w_062_5463, w_062_5470, w_062_5473, w_062_5476, w_062_5477, w_062_5478, w_062_5481, w_062_5484, w_062_5485, w_062_5486, w_062_5488, w_062_5489, w_062_5490, w_062_5492, w_062_5493, w_062_5494, w_062_5495, w_062_5499, w_062_5500, w_062_5508, w_062_5514, w_062_5517, w_062_5518, w_062_5519, w_062_5526, w_062_5527, w_062_5529, w_062_5535, w_062_5537, w_062_5538, w_062_5540, w_062_5549, w_062_5550, w_062_5559, w_062_5560, w_062_5566, w_062_5570, w_062_5578, w_062_5579, w_062_5581, w_062_5583, w_062_5584, w_062_5586, w_062_5587, w_062_5589, w_062_5594, w_062_5597, w_062_5606, w_062_5609, w_062_5612, w_062_5618, w_062_5619, w_062_5621, w_062_5622, w_062_5626, w_062_5628, w_062_5631, w_062_5635, w_062_5639, w_062_5643, w_062_5644, w_062_5645, w_062_5646, w_062_5647, w_062_5653, w_062_5654, w_062_5658, w_062_5663, w_062_5667, w_062_5674, w_062_5675, w_062_5678, w_062_5679, w_062_5680, w_062_5682, w_062_5687, w_062_5690, w_062_5691, w_062_5698, w_062_5699, w_062_5700, w_062_5701, w_062_5703, w_062_5714, w_062_5716, w_062_5718, w_062_5722, w_062_5724, w_062_5734, w_062_5736, w_062_5737, w_062_5743, w_062_5744, w_062_5748, w_062_5750, w_062_5755, w_062_5756, w_062_5764, w_062_5767, w_062_5769, w_062_5771, w_062_5774, w_062_5775, w_062_5783, w_062_5786, w_062_5787, w_062_5789, w_062_5790, w_062_5794, w_062_5795, w_062_5797, w_062_5802, w_062_5803, w_062_5804, w_062_5805, w_062_5808, w_062_5815, w_062_5821, w_062_5822, w_062_5828, w_062_5829, w_062_5835, w_062_5837, w_062_5838, w_062_5845, w_062_5847, w_062_5848, w_062_5850, w_062_5852, w_062_5853, w_062_5855, w_062_5857, w_062_5859, w_062_5860, w_062_5861, w_062_5862, w_062_5864, w_062_5865, w_062_5868, w_062_5870, w_062_5872, w_062_5873, w_062_5875, w_062_5878, w_062_5881, w_062_5885, w_062_5891, w_062_5893, w_062_5894, w_062_5895, w_062_5896, w_062_5900, w_062_5902, w_062_5904, w_062_5905, w_062_5912, w_062_5918, w_062_5924, w_062_5927, w_062_5928, w_062_5929, w_062_5930, w_062_5931, w_062_5934, w_062_5941, w_062_5948, w_062_5951, w_062_5953, w_062_5954, w_062_5955, w_062_5958, w_062_5959, w_062_5963, w_062_5964, w_062_5965, w_062_5968, w_062_5972, w_062_5974, w_062_5980, w_062_5985, w_062_5989, w_062_5990, w_062_5991, w_062_5992, w_062_5993, w_062_5994, w_062_5995, w_062_5999, w_062_6001, w_062_6004, w_062_6007, w_062_6012, w_062_6014, w_062_6016, w_062_6019, w_062_6020, w_062_6021, w_062_6024, w_062_6026, w_062_6027, w_062_6028, w_062_6030, w_062_6034, w_062_6038, w_062_6040, w_062_6048, w_062_6050, w_062_6055, w_062_6057, w_062_6060, w_062_6062, w_062_6063, w_062_6065, w_062_6066, w_062_6067, w_062_6070, w_062_6072, w_062_6074, w_062_6076, w_062_6083, w_062_6088, w_062_6090, w_062_6091, w_062_6093, w_062_6096, w_062_6099, w_062_6102, w_062_6103, w_062_6109, w_062_6110, w_062_6111, w_062_6112, w_062_6114, w_062_6117, w_062_6120, w_062_6124, w_062_6126, w_062_6134, w_062_6136, w_062_6141, w_062_6145, w_062_6147, w_062_6149, w_062_6150, w_062_6153, w_062_6154, w_062_6156, w_062_6157, w_062_6158, w_062_6160, w_062_6163, w_062_6166, w_062_6168, w_062_6174, w_062_6175, w_062_6179, w_062_6180, w_062_6181, w_062_6188, w_062_6191, w_062_6194, w_062_6197, w_062_6201, w_062_6206, w_062_6209, w_062_6214, w_062_6221, w_062_6224, w_062_6225, w_062_6229, w_062_6230, w_062_6232, w_062_6234, w_062_6235, w_062_6237, w_062_6238, w_062_6243, w_062_6244, w_062_6250, w_062_6251, w_062_6253, w_062_6254, w_062_6255, w_062_6256, w_062_6261, w_062_6262, w_062_6270, w_062_6272, w_062_6273, w_062_6285, w_062_6287, w_062_6288, w_062_6289, w_062_6290, w_062_6293, w_062_6295, w_062_6297, w_062_6300, w_062_6303, w_062_6313, w_062_6317, w_062_6318, w_062_6319, w_062_6320, w_062_6324, w_062_6326, w_062_6329, w_062_6330, w_062_6331, w_062_6338, w_062_6340, w_062_6342, w_062_6344, w_062_6346, w_062_6353, w_062_6358, w_062_6359, w_062_6361, w_062_6363, w_062_6366, w_062_6368, w_062_6370, w_062_6374, w_062_6380, w_062_6385, w_062_6398, w_062_6400, w_062_6407, w_062_6408, w_062_6410, w_062_6412, w_062_6415, w_062_6416, w_062_6418, w_062_6419, w_062_6423, w_062_6428, w_062_6430, w_062_6431, w_062_6435, w_062_6436, w_062_6438, w_062_6442, w_062_6447, w_062_6449, w_062_6451, w_062_6454, w_062_6455, w_062_6458, w_062_6459, w_062_6464, w_062_6465, w_062_6466, w_062_6469, w_062_6471, w_062_6473, w_062_6476, w_062_6478, w_062_6485, w_062_6490, w_062_6491, w_062_6492, w_062_6496, w_062_6497, w_062_6500, w_062_6507, w_062_6509, w_062_6510, w_062_6512, w_062_6518, w_062_6520, w_062_6521, w_062_6529, w_062_6530, w_062_6531, w_062_6532, w_062_6534, w_062_6536, w_062_6540, w_062_6544, w_062_6548, w_062_6549, w_062_6550, w_062_6551, w_062_6552, w_062_6561, w_062_6564, w_062_6568, w_062_6569, w_062_6570, w_062_6571, w_062_6572, w_062_6573, w_062_6574, w_062_6580, w_062_6582, w_062_6585, w_062_6588, w_062_6589, w_062_6593, w_062_6595, w_062_6596, w_062_6597, w_062_6600, w_062_6613, w_062_6615, w_062_6616, w_062_6617, w_062_6623, w_062_6630, w_062_6631, w_062_6632, w_062_6633, w_062_6641, w_062_6642, w_062_6643, w_062_6645, w_062_6652, w_062_6655, w_062_6658, w_062_6659, w_062_6660, w_062_6666, w_062_6667, w_062_6671, w_062_6674, w_062_6677, w_062_6681, w_062_6692, w_062_6697, w_062_6698, w_062_6705, w_062_6710, w_062_6711, w_062_6712, w_062_6714, w_062_6715, w_062_6717, w_062_6720, w_062_6723, w_062_6724, w_062_6731, w_062_6734, w_062_6735, w_062_6738, w_062_6739, w_062_6741, w_062_6745, w_062_6746, w_062_6748, w_062_6750, w_062_6756, w_062_6758, w_062_6760, w_062_6763, w_062_6768, w_062_6772, w_062_6773, w_062_6775, w_062_6778, w_062_6780, w_062_6782, w_062_6783, w_062_6784, w_062_6788, w_062_6789, w_062_6791, w_062_6792, w_062_6794, w_062_6796, w_062_6797, w_062_6800, w_062_6806, w_062_6809, w_062_6814, w_062_6819, w_062_6822, w_062_6824, w_062_6827, w_062_6830, w_062_6832, w_062_6841, w_062_6842, w_062_6849, w_062_6852, w_062_6853, w_062_6856, w_062_6860, w_062_6866, w_062_6869, w_062_6871, w_062_6876, w_062_6883, w_062_6884, w_062_6885, w_062_6888, w_062_6889, w_062_6893, w_062_6894, w_062_6896, w_062_6899, w_062_6901, w_062_6905, w_062_6906, w_062_6909, w_062_6910, w_062_6911, w_062_6912, w_062_6913, w_062_6918, w_062_6922, w_062_6923, w_062_6924, w_062_6926, w_062_6927, w_062_6932, w_062_6934, w_062_6941, w_062_6943, w_062_6944, w_062_6956, w_062_6957, w_062_6963, w_062_6967, w_062_6973, w_062_6975, w_062_6978, w_062_6979, w_062_6982, w_062_6985, w_062_6986, w_062_6989, w_062_6990, w_062_6992, w_062_6996, w_062_7003, w_062_7010, w_062_7011, w_062_7014, w_062_7018, w_062_7019, w_062_7020, w_062_7021, w_062_7025, w_062_7027, w_062_7030, w_062_7031, w_062_7034, w_062_7035, w_062_7037, w_062_7038, w_062_7039, w_062_7040, w_062_7043, w_062_7045, w_062_7046, w_062_7047, w_062_7048, w_062_7049, w_062_7050, w_062_7052, w_062_7057, w_062_7060, w_062_7061, w_062_7066, w_062_7069, w_062_7075, w_062_7078, w_062_7083, w_062_7085, w_062_7086, w_062_7089, w_062_7093, w_062_7096, w_062_7097, w_062_7099, w_062_7104, w_062_7107, w_062_7109, w_062_7110, w_062_7116, w_062_7121, w_062_7123, w_062_7126, w_062_7136, w_062_7140, w_062_7142, w_062_7145, w_062_7147, w_062_7148, w_062_7149, w_062_7154, w_062_7156, w_062_7158, w_062_7159, w_062_7162, w_062_7163, w_062_7164, w_062_7178, w_062_7183, w_062_7184, w_062_7185, w_062_7186, w_062_7190, w_062_7192, w_062_7195, w_062_7197, w_062_7199, w_062_7201, w_062_7205, w_062_7210, w_062_7214, w_062_7216, w_062_7217, w_062_7232, w_062_7233, w_062_7235, w_062_7236, w_062_7241, w_062_7243, w_062_7244, w_062_7245, w_062_7249, w_062_7252, w_062_7255, w_062_7260, w_062_7266, w_062_7267, w_062_7273, w_062_7277, w_062_7278, w_062_7279, w_062_7281, w_062_7283, w_062_7286, w_062_7288, w_062_7291, w_062_7296, w_062_7301, w_062_7303, w_062_7305, w_062_7307, w_062_7308, w_062_7311, w_062_7315, w_062_7316, w_062_7317, w_062_7319, w_062_7323, w_062_7330, w_062_7332, w_062_7335, w_062_7336, w_062_7337, w_062_7338, w_062_7342, w_062_7343, w_062_7344;
  wire w_063_000, w_063_002, w_063_003, w_063_004, w_063_006, w_063_007, w_063_008, w_063_009, w_063_010, w_063_011, w_063_013, w_063_014, w_063_015, w_063_016, w_063_017, w_063_018, w_063_019, w_063_022, w_063_023, w_063_025, w_063_026, w_063_027, w_063_028, w_063_029, w_063_030, w_063_032, w_063_033, w_063_034, w_063_036, w_063_037, w_063_039, w_063_040, w_063_041, w_063_044, w_063_046, w_063_047, w_063_048, w_063_049, w_063_050, w_063_051, w_063_052, w_063_053, w_063_054, w_063_055, w_063_056, w_063_057, w_063_060, w_063_061, w_063_062, w_063_065, w_063_066, w_063_068, w_063_069, w_063_070, w_063_073, w_063_074, w_063_076, w_063_079, w_063_080, w_063_081, w_063_082, w_063_083, w_063_084, w_063_085, w_063_087, w_063_088, w_063_090, w_063_091, w_063_094, w_063_096, w_063_098, w_063_099, w_063_101, w_063_102, w_063_103, w_063_104, w_063_105, w_063_106, w_063_108, w_063_109, w_063_110, w_063_111, w_063_112, w_063_113, w_063_114, w_063_115, w_063_116, w_063_117, w_063_118, w_063_120, w_063_121, w_063_123, w_063_124, w_063_125, w_063_126, w_063_127, w_063_129, w_063_131, w_063_132, w_063_135, w_063_136, w_063_139, w_063_140, w_063_144, w_063_145, w_063_147, w_063_148, w_063_149, w_063_150, w_063_151, w_063_152, w_063_153, w_063_155, w_063_156, w_063_159, w_063_160, w_063_161, w_063_162, w_063_165, w_063_166, w_063_167, w_063_170, w_063_171, w_063_173, w_063_174, w_063_175, w_063_176, w_063_178, w_063_180, w_063_181, w_063_182, w_063_183, w_063_185, w_063_186, w_063_188, w_063_189, w_063_194, w_063_196, w_063_197, w_063_199, w_063_202, w_063_203, w_063_204, w_063_205, w_063_207, w_063_208, w_063_209, w_063_210, w_063_211, w_063_215, w_063_216, w_063_217, w_063_220, w_063_222, w_063_223, w_063_225, w_063_227, w_063_229, w_063_230, w_063_232, w_063_234, w_063_237, w_063_239, w_063_240, w_063_241, w_063_242, w_063_245, w_063_246, w_063_247, w_063_248, w_063_250, w_063_255, w_063_256, w_063_257, w_063_260, w_063_261, w_063_264, w_063_265, w_063_266, w_063_269, w_063_273, w_063_275, w_063_277, w_063_279, w_063_283, w_063_286, w_063_287, w_063_289, w_063_292, w_063_294, w_063_295, w_063_297, w_063_299, w_063_300, w_063_302, w_063_305, w_063_306, w_063_309, w_063_311, w_063_313, w_063_314, w_063_315, w_063_316, w_063_317, w_063_318, w_063_320, w_063_321, w_063_325, w_063_326, w_063_328, w_063_329, w_063_330, w_063_331, w_063_333, w_063_334, w_063_339, w_063_340, w_063_341, w_063_347, w_063_352, w_063_354, w_063_356, w_063_358, w_063_360, w_063_362, w_063_363, w_063_365, w_063_366, w_063_369, w_063_371, w_063_372, w_063_373, w_063_374, w_063_377, w_063_379, w_063_380, w_063_381, w_063_382, w_063_384, w_063_386, w_063_389, w_063_390, w_063_391, w_063_392, w_063_395, w_063_397, w_063_398, w_063_399, w_063_401, w_063_402, w_063_407, w_063_408, w_063_409, w_063_410, w_063_411, w_063_414, w_063_417, w_063_418, w_063_420, w_063_422, w_063_425, w_063_427, w_063_430, w_063_431, w_063_432, w_063_433, w_063_439, w_063_440, w_063_443, w_063_444, w_063_445, w_063_446, w_063_447, w_063_448, w_063_449, w_063_450, w_063_451, w_063_456, w_063_457, w_063_458, w_063_461, w_063_462, w_063_463, w_063_465, w_063_467, w_063_470, w_063_471, w_063_472, w_063_474, w_063_475, w_063_477, w_063_478, w_063_479, w_063_480, w_063_481, w_063_482, w_063_483, w_063_485, w_063_486, w_063_488, w_063_489, w_063_490, w_063_491, w_063_493, w_063_494, w_063_495, w_063_496, w_063_498, w_063_500, w_063_501, w_063_504, w_063_506, w_063_512, w_063_515, w_063_516, w_063_518, w_063_520, w_063_521, w_063_524, w_063_525, w_063_526, w_063_527, w_063_530, w_063_533, w_063_534, w_063_535, w_063_536, w_063_537, w_063_538, w_063_539, w_063_540, w_063_542, w_063_543, w_063_547, w_063_549, w_063_550, w_063_551, w_063_553, w_063_555, w_063_557, w_063_558, w_063_559, w_063_560, w_063_562, w_063_567, w_063_568, w_063_569, w_063_570, w_063_571, w_063_573, w_063_574, w_063_577, w_063_578, w_063_579, w_063_581, w_063_584, w_063_585, w_063_586, w_063_588, w_063_592, w_063_593, w_063_596, w_063_597, w_063_598, w_063_600, w_063_602, w_063_603, w_063_606, w_063_608, w_063_610, w_063_611, w_063_615, w_063_620, w_063_624, w_063_626, w_063_627, w_063_629, w_063_630, w_063_633, w_063_634, w_063_635, w_063_641, w_063_642, w_063_643, w_063_644, w_063_646, w_063_647, w_063_648, w_063_650, w_063_656, w_063_657, w_063_660, w_063_661, w_063_663, w_063_666, w_063_670, w_063_675, w_063_677, w_063_678, w_063_679, w_063_683, w_063_686, w_063_687, w_063_689, w_063_691, w_063_692, w_063_693, w_063_694, w_063_695, w_063_697, w_063_698, w_063_699, w_063_703, w_063_704, w_063_707, w_063_709, w_063_710, w_063_711, w_063_712, w_063_714, w_063_715, w_063_716, w_063_718, w_063_719, w_063_720, w_063_721, w_063_722, w_063_723, w_063_727, w_063_728, w_063_729, w_063_730, w_063_732, w_063_733, w_063_735, w_063_738, w_063_739, w_063_740, w_063_741, w_063_742, w_063_745, w_063_747, w_063_750, w_063_753, w_063_756, w_063_757, w_063_759, w_063_763, w_063_765, w_063_766, w_063_767, w_063_768, w_063_769, w_063_771, w_063_773, w_063_774, w_063_775, w_063_777, w_063_781, w_063_782, w_063_785, w_063_787, w_063_788, w_063_795, w_063_797, w_063_799, w_063_801, w_063_803, w_063_806, w_063_809, w_063_810, w_063_811, w_063_812, w_063_814, w_063_815, w_063_816, w_063_817, w_063_818, w_063_823, w_063_824, w_063_825, w_063_830, w_063_831, w_063_832, w_063_833, w_063_837, w_063_838, w_063_839, w_063_840, w_063_841, w_063_843, w_063_846, w_063_847, w_063_848, w_063_852, w_063_853, w_063_854, w_063_855, w_063_858, w_063_859, w_063_862, w_063_863, w_063_865, w_063_866, w_063_867, w_063_869, w_063_872, w_063_873, w_063_874, w_063_875, w_063_878, w_063_879, w_063_882, w_063_883, w_063_886, w_063_887, w_063_892, w_063_893, w_063_894, w_063_896, w_063_897, w_063_898, w_063_899, w_063_900, w_063_903, w_063_904, w_063_907, w_063_910, w_063_911, w_063_915, w_063_916, w_063_919, w_063_920, w_063_923, w_063_924, w_063_925, w_063_926, w_063_928, w_063_929, w_063_930, w_063_932, w_063_934, w_063_935, w_063_936, w_063_937, w_063_939, w_063_940, w_063_941, w_063_942, w_063_943, w_063_945, w_063_947, w_063_948, w_063_949, w_063_953, w_063_956, w_063_957, w_063_958, w_063_961, w_063_962, w_063_963, w_063_964, w_063_966, w_063_968, w_063_970, w_063_971, w_063_972, w_063_974, w_063_977, w_063_978, w_063_980, w_063_982, w_063_983, w_063_984, w_063_987, w_063_989, w_063_993, w_063_998, w_063_1000, w_063_1003, w_063_1004, w_063_1005, w_063_1007, w_063_1008, w_063_1009, w_063_1011, w_063_1014, w_063_1015, w_063_1016, w_063_1017, w_063_1018, w_063_1022, w_063_1023, w_063_1026, w_063_1027, w_063_1028, w_063_1029, w_063_1031, w_063_1032, w_063_1033, w_063_1034, w_063_1035, w_063_1038, w_063_1040, w_063_1041, w_063_1042, w_063_1045, w_063_1046, w_063_1049, w_063_1050, w_063_1051, w_063_1053, w_063_1055, w_063_1056, w_063_1062, w_063_1067, w_063_1068, w_063_1070, w_063_1073, w_063_1074, w_063_1075, w_063_1076, w_063_1077, w_063_1078, w_063_1079, w_063_1081, w_063_1084, w_063_1085, w_063_1086, w_063_1087, w_063_1093, w_063_1094, w_063_1097, w_063_1098, w_063_1100, w_063_1101, w_063_1102, w_063_1103, w_063_1104, w_063_1105, w_063_1108, w_063_1109, w_063_1110, w_063_1111, w_063_1113, w_063_1114, w_063_1115, w_063_1119, w_063_1121, w_063_1122, w_063_1125, w_063_1127, w_063_1128, w_063_1129, w_063_1131, w_063_1134, w_063_1136, w_063_1137, w_063_1139, w_063_1141, w_063_1142, w_063_1143, w_063_1144, w_063_1146, w_063_1147, w_063_1149, w_063_1150, w_063_1151, w_063_1153, w_063_1156, w_063_1157, w_063_1159, w_063_1162, w_063_1165, w_063_1172, w_063_1174, w_063_1176, w_063_1178, w_063_1179, w_063_1180, w_063_1182, w_063_1183, w_063_1185, w_063_1186, w_063_1187, w_063_1188, w_063_1190, w_063_1191, w_063_1192, w_063_1193, w_063_1195, w_063_1196, w_063_1197, w_063_1198, w_063_1201, w_063_1203, w_063_1204, w_063_1205, w_063_1207, w_063_1208, w_063_1210, w_063_1211, w_063_1212, w_063_1215, w_063_1220, w_063_1222, w_063_1225, w_063_1227, w_063_1229, w_063_1230, w_063_1232, w_063_1234, w_063_1236, w_063_1239, w_063_1242, w_063_1243, w_063_1245, w_063_1246, w_063_1247, w_063_1248, w_063_1249, w_063_1250, w_063_1254, w_063_1257, w_063_1259, w_063_1260, w_063_1261, w_063_1263, w_063_1264, w_063_1265, w_063_1266, w_063_1267, w_063_1268, w_063_1271, w_063_1273, w_063_1276, w_063_1279, w_063_1281, w_063_1285, w_063_1286, w_063_1287, w_063_1288, w_063_1293, w_063_1295, w_063_1296, w_063_1297, w_063_1298, w_063_1300, w_063_1305, w_063_1306, w_063_1308, w_063_1311, w_063_1312, w_063_1314, w_063_1315, w_063_1316, w_063_1317, w_063_1322, w_063_1323, w_063_1325, w_063_1328, w_063_1329, w_063_1330, w_063_1332, w_063_1333, w_063_1334, w_063_1335, w_063_1336, w_063_1338, w_063_1341, w_063_1342, w_063_1343, w_063_1344, w_063_1346, w_063_1347, w_063_1348, w_063_1350, w_063_1353, w_063_1354, w_063_1355, w_063_1358, w_063_1361, w_063_1362, w_063_1365, w_063_1366, w_063_1367, w_063_1368, w_063_1369, w_063_1370, w_063_1373, w_063_1375, w_063_1377, w_063_1379, w_063_1380, w_063_1382, w_063_1383, w_063_1384, w_063_1387, w_063_1388, w_063_1390, w_063_1393, w_063_1395, w_063_1396, w_063_1398, w_063_1399, w_063_1400, w_063_1401, w_063_1405, w_063_1406, w_063_1407, w_063_1411, w_063_1412, w_063_1413, w_063_1415, w_063_1416, w_063_1417, w_063_1418, w_063_1419, w_063_1421, w_063_1422, w_063_1423, w_063_1424, w_063_1426, w_063_1428, w_063_1429, w_063_1430, w_063_1431, w_063_1432, w_063_1436, w_063_1439, w_063_1441, w_063_1443, w_063_1446, w_063_1447, w_063_1449, w_063_1450, w_063_1451, w_063_1452, w_063_1454, w_063_1456, w_063_1458, w_063_1460, w_063_1461, w_063_1463, w_063_1464, w_063_1466, w_063_1467, w_063_1468, w_063_1469, w_063_1471, w_063_1474, w_063_1475, w_063_1476, w_063_1478, w_063_1480, w_063_1481, w_063_1483, w_063_1485, w_063_1486, w_063_1487, w_063_1493, w_063_1494, w_063_1495, w_063_1496, w_063_1498, w_063_1499, w_063_1500, w_063_1501, w_063_1502, w_063_1505, w_063_1507, w_063_1508, w_063_1509, w_063_1511, w_063_1512, w_063_1513, w_063_1514, w_063_1515, w_063_1516, w_063_1518, w_063_1519, w_063_1524, w_063_1526, w_063_1528, w_063_1531, w_063_1540, w_063_1541, w_063_1542, w_063_1544, w_063_1546, w_063_1547, w_063_1550, w_063_1551, w_063_1552, w_063_1553, w_063_1554, w_063_1556, w_063_1557, w_063_1558, w_063_1560, w_063_1563, w_063_1565, w_063_1567, w_063_1569, w_063_1571, w_063_1574, w_063_1577, w_063_1578, w_063_1580, w_063_1581, w_063_1582, w_063_1583, w_063_1585, w_063_1588, w_063_1589, w_063_1590, w_063_1591, w_063_1592, w_063_1595, w_063_1598, w_063_1599, w_063_1602, w_063_1603, w_063_1605, w_063_1608, w_063_1611, w_063_1612, w_063_1614, w_063_1616, w_063_1618, w_063_1619, w_063_1620, w_063_1622, w_063_1623, w_063_1624, w_063_1625, w_063_1627, w_063_1628, w_063_1633, w_063_1637, w_063_1638, w_063_1640, w_063_1644, w_063_1645, w_063_1646, w_063_1652, w_063_1655, w_063_1656, w_063_1657, w_063_1658, w_063_1659, w_063_1660, w_063_1661, w_063_1662, w_063_1671, w_063_1673, w_063_1679, w_063_1681, w_063_1682, w_063_1685, w_063_1686, w_063_1687, w_063_1690, w_063_1693, w_063_1694, w_063_1695, w_063_1697, w_063_1698, w_063_1699, w_063_1702, w_063_1705, w_063_1706, w_063_1707, w_063_1709, w_063_1710, w_063_1712, w_063_1713, w_063_1718, w_063_1719, w_063_1722, w_063_1723, w_063_1726, w_063_1729, w_063_1730, w_063_1731, w_063_1733, w_063_1735, w_063_1736, w_063_1737, w_063_1738, w_063_1740, w_063_1741, w_063_1743, w_063_1744, w_063_1746, w_063_1747, w_063_1748, w_063_1749, w_063_1750, w_063_1751, w_063_1752, w_063_1754, w_063_1755, w_063_1756, w_063_1757, w_063_1758, w_063_1761, w_063_1762, w_063_1763, w_063_1764, w_063_1765, w_063_1766, w_063_1767, w_063_1770, w_063_1775, w_063_1776, w_063_1777, w_063_1778, w_063_1782, w_063_1783, w_063_1784, w_063_1785, w_063_1786, w_063_1787, w_063_1790, w_063_1791, w_063_1792, w_063_1793, w_063_1795, w_063_1796, w_063_1797, w_063_1801, w_063_1802, w_063_1803, w_063_1804, w_063_1806, w_063_1807, w_063_1810, w_063_1812, w_063_1815, w_063_1817, w_063_1818, w_063_1819, w_063_1822, w_063_1823, w_063_1825, w_063_1826, w_063_1828, w_063_1831, w_063_1832, w_063_1834, w_063_1836, w_063_1838, w_063_1839, w_063_1841, w_063_1842, w_063_1845, w_063_1846, w_063_1849, w_063_1850, w_063_1851, w_063_1853, w_063_1854, w_063_1856, w_063_1857, w_063_1859, w_063_1863, w_063_1864, w_063_1865, w_063_1867, w_063_1869, w_063_1870, w_063_1875, w_063_1878, w_063_1880, w_063_1886, w_063_1887, w_063_1890, w_063_1892, w_063_1893, w_063_1894, w_063_1896, w_063_1897, w_063_1899, w_063_1900, w_063_1903, w_063_1904, w_063_1906, w_063_1908, w_063_1909, w_063_1911, w_063_1913, w_063_1915, w_063_1916, w_063_1917, w_063_1918, w_063_1919, w_063_1921, w_063_1922, w_063_1923, w_063_1925, w_063_1928, w_063_1929, w_063_1930, w_063_1931, w_063_1932, w_063_1933, w_063_1935, w_063_1936, w_063_1937, w_063_1939, w_063_1941, w_063_1942, w_063_1944, w_063_1945, w_063_1946, w_063_1947, w_063_1951, w_063_1952, w_063_1954, w_063_1956, w_063_1958, w_063_1959, w_063_1961, w_063_1962, w_063_1966, w_063_1967, w_063_1968, w_063_1969, w_063_1972, w_063_1976, w_063_1979, w_063_1980, w_063_1981, w_063_1983, w_063_1985, w_063_1987, w_063_1988, w_063_1989, w_063_1991, w_063_1992, w_063_1996, w_063_1998, w_063_1999, w_063_2001, w_063_2005, w_063_2007, w_063_2008, w_063_2010, w_063_2011, w_063_2012, w_063_2013, w_063_2014, w_063_2015, w_063_2018, w_063_2020, w_063_2021, w_063_2023, w_063_2026, w_063_2028, w_063_2030, w_063_2033, w_063_2036, w_063_2037, w_063_2038, w_063_2039, w_063_2040, w_063_2041, w_063_2043, w_063_2044, w_063_2046, w_063_2047, w_063_2050, w_063_2052, w_063_2060, w_063_2061, w_063_2062, w_063_2063, w_063_2065, w_063_2066, w_063_2068, w_063_2069, w_063_2072, w_063_2073, w_063_2075, w_063_2079, w_063_2080, w_063_2083, w_063_2085, w_063_2086, w_063_2088, w_063_2089, w_063_2091, w_063_2092, w_063_2093, w_063_2094, w_063_2095, w_063_2096, w_063_2097, w_063_2098, w_063_2099, w_063_2101, w_063_2103, w_063_2104, w_063_2106, w_063_2107, w_063_2111, w_063_2112, w_063_2113, w_063_2114, w_063_2115, w_063_2116, w_063_2118, w_063_2119, w_063_2121, w_063_2122, w_063_2125, w_063_2127, w_063_2128, w_063_2130, w_063_2134, w_063_2136, w_063_2137, w_063_2142, w_063_2143, w_063_2144, w_063_2145, w_063_2146, w_063_2147, w_063_2148, w_063_2151, w_063_2153, w_063_2155, w_063_2157, w_063_2158, w_063_2161, w_063_2163, w_063_2165, w_063_2168, w_063_2169, w_063_2171, w_063_2173, w_063_2180, w_063_2181, w_063_2182, w_063_2183, w_063_2184, w_063_2185, w_063_2186, w_063_2189, w_063_2190, w_063_2192, w_063_2193, w_063_2194, w_063_2196, w_063_2197, w_063_2198, w_063_2199, w_063_2200, w_063_2202, w_063_2203, w_063_2204, w_063_2205, w_063_2206, w_063_2209, w_063_2211, w_063_2212, w_063_2213, w_063_2214, w_063_2216, w_063_2221, w_063_2222, w_063_2223, w_063_2224, w_063_2225, w_063_2227, w_063_2228, w_063_2231, w_063_2232, w_063_2233, w_063_2234, w_063_2238, w_063_2241, w_063_2242, w_063_2244, w_063_2246, w_063_2248, w_063_2249, w_063_2250, w_063_2252, w_063_2254, w_063_2255, w_063_2257, w_063_2258, w_063_2259, w_063_2260, w_063_2262, w_063_2263, w_063_2264, w_063_2265, w_063_2266, w_063_2267, w_063_2270, w_063_2271, w_063_2272, w_063_2273, w_063_2275, w_063_2276, w_063_2277, w_063_2280, w_063_2282, w_063_2284, w_063_2285, w_063_2288, w_063_2290, w_063_2293, w_063_2294, w_063_2296, w_063_2297, w_063_2298, w_063_2299, w_063_2300, w_063_2301, w_063_2302, w_063_2303, w_063_2304, w_063_2307, w_063_2308, w_063_2310, w_063_2312, w_063_2315, w_063_2316, w_063_2318, w_063_2319, w_063_2321, w_063_2324, w_063_2325, w_063_2326, w_063_2327, w_063_2329, w_063_2333, w_063_2337, w_063_2338, w_063_2340, w_063_2342, w_063_2343, w_063_2344, w_063_2345, w_063_2346, w_063_2348, w_063_2350, w_063_2351, w_063_2353, w_063_2354, w_063_2355, w_063_2357, w_063_2359, w_063_2361, w_063_2366, w_063_2367, w_063_2371, w_063_2373, w_063_2374, w_063_2375, w_063_2376, w_063_2377, w_063_2378, w_063_2379, w_063_2380, w_063_2381, w_063_2382, w_063_2385, w_063_2386, w_063_2388, w_063_2390, w_063_2391, w_063_2393, w_063_2394, w_063_2398, w_063_2402, w_063_2403, w_063_2405, w_063_2406, w_063_2407, w_063_2408, w_063_2409, w_063_2411, w_063_2413, w_063_2414, w_063_2418, w_063_2421, w_063_2422, w_063_2427, w_063_2428, w_063_2429, w_063_2433, w_063_2434, w_063_2435, w_063_2436, w_063_2437, w_063_2438, w_063_2439, w_063_2441, w_063_2442, w_063_2443, w_063_2445, w_063_2446, w_063_2447, w_063_2448, w_063_2449, w_063_2451, w_063_2452, w_063_2453, w_063_2455, w_063_2456, w_063_2457, w_063_2458, w_063_2459, w_063_2461, w_063_2463, w_063_2464, w_063_2465, w_063_2467, w_063_2468, w_063_2469, w_063_2470, w_063_2472, w_063_2474, w_063_2475, w_063_2476, w_063_2477, w_063_2478, w_063_2479, w_063_2480, w_063_2482, w_063_2483, w_063_2485, w_063_2486, w_063_2487, w_063_2488, w_063_2492, w_063_2495, w_063_2497, w_063_2498, w_063_2499, w_063_2500, w_063_2501, w_063_2502, w_063_2505, w_063_2506, w_063_2510, w_063_2511, w_063_2512, w_063_2513, w_063_2514, w_063_2515, w_063_2516, w_063_2518, w_063_2520, w_063_2521, w_063_2524, w_063_2525, w_063_2527, w_063_2531, w_063_2532, w_063_2534, w_063_2535, w_063_2536, w_063_2537, w_063_2542, w_063_2544, w_063_2546, w_063_2547, w_063_2551, w_063_2553, w_063_2554, w_063_2555, w_063_2556, w_063_2559, w_063_2560, w_063_2561, w_063_2562, w_063_2564, w_063_2565, w_063_2567, w_063_2569, w_063_2571, w_063_2572, w_063_2576, w_063_2581, w_063_2582, w_063_2583, w_063_2585, w_063_2587, w_063_2588, w_063_2589, w_063_2590, w_063_2592, w_063_2594, w_063_2597, w_063_2598, w_063_2599, w_063_2600, w_063_2602, w_063_2603, w_063_2604, w_063_2607, w_063_2608, w_063_2609, w_063_2612, w_063_2613, w_063_2615, w_063_2618, w_063_2619, w_063_2620, w_063_2622, w_063_2623, w_063_2625, w_063_2627, w_063_2628, w_063_2630, w_063_2631, w_063_2633, w_063_2634, w_063_2635, w_063_2638, w_063_2640, w_063_2644, w_063_2645, w_063_2646, w_063_2648, w_063_2651, w_063_2653, w_063_2656, w_063_2658, w_063_2660, w_063_2661, w_063_2662, w_063_2663, w_063_2665, w_063_2666, w_063_2667, w_063_2669, w_063_2670, w_063_2671, w_063_2673, w_063_2674, w_063_2676, w_063_2677, w_063_2679, w_063_2680, w_063_2682, w_063_2683, w_063_2684, w_063_2685, w_063_2686, w_063_2689, w_063_2690, w_063_2692, w_063_2693, w_063_2694, w_063_2695, w_063_2700, w_063_2702, w_063_2705, w_063_2706, w_063_2707, w_063_2710, w_063_2711, w_063_2712, w_063_2714, w_063_2715, w_063_2720, w_063_2721, w_063_2722, w_063_2724, w_063_2726, w_063_2727, w_063_2729, w_063_2730, w_063_2732, w_063_2734, w_063_2735, w_063_2736, w_063_2740, w_063_2741, w_063_2742, w_063_2745, w_063_2747, w_063_2751, w_063_2754, w_063_2756, w_063_2757, w_063_2758, w_063_2761, w_063_2763, w_063_2766, w_063_2767, w_063_2768, w_063_2769, w_063_2771, w_063_2772, w_063_2774, w_063_2775, w_063_2776, w_063_2777, w_063_2778, w_063_2779, w_063_2780, w_063_2784, w_063_2786, w_063_2787, w_063_2788, w_063_2789, w_063_2790, w_063_2793, w_063_2794, w_063_2795, w_063_2796, w_063_2797, w_063_2799, w_063_2801, w_063_2802, w_063_2803, w_063_2805, w_063_2809, w_063_2810, w_063_2811, w_063_2813, w_063_2816, w_063_2817, w_063_2819, w_063_2820, w_063_2821, w_063_2822, w_063_2825, w_063_2826, w_063_2828, w_063_2830, w_063_2831, w_063_2832, w_063_2837, w_063_2839, w_063_2840, w_063_2843, w_063_2844, w_063_2845, w_063_2846, w_063_2847, w_063_2849, w_063_2850, w_063_2851, w_063_2855, w_063_2858, w_063_2860, w_063_2861, w_063_2863, w_063_2864, w_063_2865, w_063_2866, w_063_2870, w_063_2873, w_063_2875, w_063_2876, w_063_2879, w_063_2882, w_063_2883, w_063_2887, w_063_2888, w_063_2893, w_063_2894, w_063_2895, w_063_2896, w_063_2897, w_063_2898, w_063_2899, w_063_2900, w_063_2901, w_063_2902, w_063_2903, w_063_2904, w_063_2907, w_063_2908, w_063_2909, w_063_2910, w_063_2913, w_063_2915, w_063_2917, w_063_2919, w_063_2921, w_063_2922, w_063_2924, w_063_2926, w_063_2928, w_063_2932, w_063_2933, w_063_2934, w_063_2935, w_063_2938, w_063_2939, w_063_2940, w_063_2942, w_063_2943, w_063_2944, w_063_2945, w_063_2946, w_063_2947, w_063_2948, w_063_2949, w_063_2951, w_063_2953, w_063_2954, w_063_2963, w_063_2964, w_063_2966, w_063_2967, w_063_2969, w_063_2970, w_063_2971, w_063_2972, w_063_2974, w_063_2975, w_063_2977, w_063_2978, w_063_2979, w_063_2980, w_063_2981, w_063_2982, w_063_2983, w_063_2985, w_063_2986, w_063_2987, w_063_2989, w_063_2990, w_063_2993, w_063_2996, w_063_2998, w_063_3000, w_063_3002, w_063_3003, w_063_3004, w_063_3005, w_063_3007, w_063_3013, w_063_3015, w_063_3017, w_063_3019, w_063_3021, w_063_3022, w_063_3024, w_063_3025, w_063_3026, w_063_3028, w_063_3029, w_063_3030, w_063_3032, w_063_3034, w_063_3035, w_063_3038, w_063_3039, w_063_3040, w_063_3045, w_063_3048, w_063_3051, w_063_3055, w_063_3056, w_063_3058, w_063_3060, w_063_3061, w_063_3062, w_063_3065, w_063_3066, w_063_3068, w_063_3071, w_063_3072, w_063_3073, w_063_3076, w_063_3078, w_063_3080, w_063_3082, w_063_3087, w_063_3088, w_063_3092, w_063_3094, w_063_3097, w_063_3099, w_063_3101, w_063_3105, w_063_3108, w_063_3109, w_063_3110, w_063_3113, w_063_3114, w_063_3115, w_063_3119, w_063_3120, w_063_3121, w_063_3122, w_063_3124, w_063_3126, w_063_3128, w_063_3129, w_063_3131, w_063_3132, w_063_3136, w_063_3137, w_063_3139, w_063_3144, w_063_3145, w_063_3147, w_063_3149, w_063_3150, w_063_3152, w_063_3153, w_063_3154, w_063_3155, w_063_3157, w_063_3158, w_063_3160, w_063_3161, w_063_3162, w_063_3164, w_063_3165, w_063_3166, w_063_3167, w_063_3170, w_063_3171, w_063_3172, w_063_3174, w_063_3175, w_063_3176, w_063_3178, w_063_3179, w_063_3181, w_063_3182, w_063_3183, w_063_3184, w_063_3187, w_063_3188, w_063_3189, w_063_3192, w_063_3193, w_063_3196, w_063_3198, w_063_3199, w_063_3201, w_063_3202, w_063_3203, w_063_3206, w_063_3208, w_063_3211, w_063_3214, w_063_3218, w_063_3219, w_063_3221, w_063_3222, w_063_3223, w_063_3224, w_063_3226, w_063_3227, w_063_3230, w_063_3231, w_063_3232, w_063_3233, w_063_3234, w_063_3236, w_063_3237, w_063_3238, w_063_3239, w_063_3240, w_063_3244, w_063_3246, w_063_3248, w_063_3249, w_063_3250, w_063_3251, w_063_3254, w_063_3255, w_063_3256, w_063_3257, w_063_3258, w_063_3259, w_063_3263, w_063_3264, w_063_3265, w_063_3269, w_063_3270, w_063_3271, w_063_3273, w_063_3274, w_063_3276, w_063_3277, w_063_3278, w_063_3281, w_063_3284, w_063_3289, w_063_3291, w_063_3295, w_063_3296, w_063_3298, w_063_3303, w_063_3304, w_063_3306, w_063_3308, w_063_3309, w_063_3312, w_063_3313, w_063_3315, w_063_3317, w_063_3319, w_063_3320, w_063_3321, w_063_3323, w_063_3324, w_063_3325, w_063_3326, w_063_3327, w_063_3328, w_063_3329, w_063_3330, w_063_3332, w_063_3333, w_063_3334, w_063_3335, w_063_3337, w_063_3338, w_063_3339, w_063_3340, w_063_3342, w_063_3343, w_063_3344, w_063_3346, w_063_3347, w_063_3349, w_063_3350, w_063_3351, w_063_3352, w_063_3356, w_063_3357, w_063_3358, w_063_3359, w_063_3361, w_063_3362, w_063_3364, w_063_3365, w_063_3366, w_063_3367, w_063_3368, w_063_3370, w_063_3376, w_063_3377, w_063_3380, w_063_3381, w_063_3382, w_063_3385, w_063_3387, w_063_3389, w_063_3390, w_063_3391, w_063_3392, w_063_3393, w_063_3394, w_063_3397, w_063_3398, w_063_3400, w_063_3404, w_063_3405, w_063_3407, w_063_3408, w_063_3410, w_063_3412, w_063_3413, w_063_3414, w_063_3417, w_063_3418, w_063_3419, w_063_3421, w_063_3424, w_063_3425, w_063_3429, w_063_3431, w_063_3432, w_063_3433, w_063_3434, w_063_3439, w_063_3442, w_063_3443, w_063_3445, w_063_3446, w_063_3450, w_063_3451, w_063_3452, w_063_3453, w_063_3458, w_063_3459, w_063_3460, w_063_3462, w_063_3463, w_063_3464, w_063_3465, w_063_3466, w_063_3467, w_063_3469, w_063_3470, w_063_3471, w_063_3476, w_063_3477, w_063_3478, w_063_3479, w_063_3480, w_063_3481, w_063_3482, w_063_3483, w_063_3486, w_063_3487, w_063_3490, w_063_3492, w_063_3494, w_063_3495, w_063_3496, w_063_3497, w_063_3499, w_063_3500, w_063_3501, w_063_3502, w_063_3503, w_063_3504, w_063_3505, w_063_3506, w_063_3512, w_063_3514, w_063_3517, w_063_3518, w_063_3519, w_063_3520, w_063_3521, w_063_3522, w_063_3525, w_063_3526, w_063_3528, w_063_3529, w_063_3530, w_063_3532, w_063_3533, w_063_3534, w_063_3537, w_063_3539, w_063_3542, w_063_3544, w_063_3548, w_063_3550, w_063_3551, w_063_3554, w_063_3556, w_063_3557, w_063_3558, w_063_3559, w_063_3560, w_063_3561, w_063_3565, w_063_3569, w_063_3570, w_063_3572, w_063_3573, w_063_3574, w_063_3575, w_063_3576, w_063_3577, w_063_3579, w_063_3581, w_063_3583, w_063_3584, w_063_3589, w_063_3590, w_063_3591, w_063_3595, w_063_3596, w_063_3598, w_063_3601, w_063_3605, w_063_3608, w_063_3609, w_063_3612, w_063_3614, w_063_3615, w_063_3618, w_063_3619, w_063_3623, w_063_3624, w_063_3625, w_063_3626, w_063_3627, w_063_3628, w_063_3631, w_063_3632, w_063_3636, w_063_3638, w_063_3641, w_063_3642, w_063_3643, w_063_3645, w_063_3647, w_063_3648, w_063_3651, w_063_3653, w_063_3654, w_063_3655, w_063_3656, w_063_3657, w_063_3660, w_063_3662, w_063_3664, w_063_3665, w_063_3667, w_063_3668, w_063_3669, w_063_3670, w_063_3675, w_063_3677, w_063_3680, w_063_3683, w_063_3684, w_063_3685, w_063_3686, w_063_3688, w_063_3689, w_063_3690, w_063_3691, w_063_3696, w_063_3697, w_063_3698, w_063_3705, w_063_3706, w_063_3707, w_063_3711, w_063_3712, w_063_3713, w_063_3716, w_063_3717, w_063_3719, w_063_3720, w_063_3724, w_063_3725, w_063_3727, w_063_3728, w_063_3729, w_063_3730, w_063_3732, w_063_3740, w_063_3741, w_063_3742, w_063_3743, w_063_3744, w_063_3746, w_063_3748, w_063_3750, w_063_3751, w_063_3753, w_063_3754, w_063_3755, w_063_3757, w_063_3760, w_063_3763, w_063_3767, w_063_3770, w_063_3772, w_063_3773, w_063_3778, w_063_3785, w_063_3788, w_063_3790, w_063_3791, w_063_3792, w_063_3793, w_063_3794, w_063_3795, w_063_3796, w_063_3797, w_063_3799, w_063_3801, w_063_3802, w_063_3806, w_063_3809, w_063_3810, w_063_3814, w_063_3815, w_063_3816, w_063_3817, w_063_3819, w_063_3820, w_063_3821, w_063_3822, w_063_3824, w_063_3826, w_063_3829, w_063_3830, w_063_3831, w_063_3832, w_063_3834, w_063_3835, w_063_3837, w_063_3838, w_063_3839, w_063_3842, w_063_3843, w_063_3845, w_063_3848, w_063_3850, w_063_3851, w_063_3856, w_063_3857, w_063_3858, w_063_3860, w_063_3861, w_063_3862, w_063_3863, w_063_3864, w_063_3868, w_063_3871, w_063_3872, w_063_3873, w_063_3876, w_063_3877, w_063_3880, w_063_3881, w_063_3884, w_063_3885, w_063_3889, w_063_3891, w_063_3893, w_063_3898, w_063_3899, w_063_3900, w_063_3901, w_063_3903, w_063_3906, w_063_3907, w_063_3909, w_063_3911, w_063_3912, w_063_3913, w_063_3914, w_063_3915, w_063_3917, w_063_3918, w_063_3919, w_063_3921, w_063_3923, w_063_3925, w_063_3928, w_063_3930, w_063_3934, w_063_3935, w_063_3936, w_063_3938, w_063_3939, w_063_3941, w_063_3942, w_063_3944, w_063_3945, w_063_3950, w_063_3952, w_063_3954, w_063_3956, w_063_3958, w_063_3959, w_063_3960, w_063_3964, w_063_3965, w_063_3967, w_063_3968, w_063_3970, w_063_3971, w_063_3972, w_063_3975, w_063_3978, w_063_3981, w_063_3982, w_063_3984, w_063_3985, w_063_3986, w_063_3988, w_063_3990, w_063_3993, w_063_3997, w_063_4001, w_063_4003, w_063_4004, w_063_4005, w_063_4007, w_063_4009, w_063_4010, w_063_4012, w_063_4013, w_063_4014, w_063_4015, w_063_4017, w_063_4018, w_063_4019, w_063_4020, w_063_4022, w_063_4023, w_063_4024, w_063_4025, w_063_4026, w_063_4027, w_063_4028, w_063_4030, w_063_4032, w_063_4036, w_063_4037, w_063_4039, w_063_4041, w_063_4042, w_063_4043, w_063_4044, w_063_4045, w_063_4048, w_063_4049, w_063_4051, w_063_4052, w_063_4053, w_063_4054, w_063_4055, w_063_4058, w_063_4059, w_063_4060, w_063_4061, w_063_4067, w_063_4068, w_063_4071, w_063_4072, w_063_4073, w_063_4077, w_063_4078, w_063_4080, w_063_4084, w_063_4085, w_063_4086, w_063_4087, w_063_4089, w_063_4090, w_063_4091, w_063_4092, w_063_4093, w_063_4097, w_063_4102, w_063_4103, w_063_4107, w_063_4108, w_063_4111, w_063_4114, w_063_4115, w_063_4116, w_063_4118, w_063_4120, w_063_4121, w_063_4122, w_063_4123, w_063_4124, w_063_4125, w_063_4126, w_063_4131, w_063_4134, w_063_4136, w_063_4137, w_063_4141, w_063_4142, w_063_4143, w_063_4145, w_063_4146, w_063_4147, w_063_4148, w_063_4149, w_063_4150, w_063_4152, w_063_4153, w_063_4154, w_063_4155, w_063_4157, w_063_4160, w_063_4161, w_063_4165, w_063_4168, w_063_4169, w_063_4170, w_063_4171, w_063_4172, w_063_4174, w_063_4175, w_063_4176, w_063_4177, w_063_4178, w_063_4179, w_063_4182, w_063_4183, w_063_4185, w_063_4186, w_063_4187, w_063_4189, w_063_4190, w_063_4191, w_063_4192, w_063_4195, w_063_4198, w_063_4200, w_063_4201, w_063_4202, w_063_4204, w_063_4205, w_063_4207, w_063_4208, w_063_4209, w_063_4210, w_063_4215, w_063_4216, w_063_4219, w_063_4220, w_063_4224, w_063_4225, w_063_4226, w_063_4227, w_063_4231, w_063_4234, w_063_4235, w_063_4236, w_063_4237, w_063_4239, w_063_4240, w_063_4242, w_063_4243, w_063_4244, w_063_4245, w_063_4247, w_063_4248, w_063_4249, w_063_4250, w_063_4252, w_063_4253, w_063_4254, w_063_4256, w_063_4259, w_063_4260, w_063_4261, w_063_4262, w_063_4263, w_063_4264, w_063_4265, w_063_4270, w_063_4271, w_063_4276, w_063_4278, w_063_4280, w_063_4281, w_063_4285, w_063_4286, w_063_4289, w_063_4291, w_063_4292, w_063_4294, w_063_4296, w_063_4297, w_063_4300, w_063_4301, w_063_4302, w_063_4303, w_063_4304, w_063_4306, w_063_4308, w_063_4309, w_063_4311, w_063_4313, w_063_4314, w_063_4316, w_063_4318, w_063_4319, w_063_4320, w_063_4322, w_063_4324, w_063_4325, w_063_4329, w_063_4331, w_063_4332, w_063_4333, w_063_4335, w_063_4336, w_063_4337, w_063_4340, w_063_4341, w_063_4342, w_063_4343, w_063_4348, w_063_4352, w_063_4355, w_063_4357, w_063_4358, w_063_4361, w_063_4362, w_063_4363, w_063_4364, w_063_4365, w_063_4366, w_063_4367, w_063_4369, w_063_4370, w_063_4371, w_063_4372, w_063_4373, w_063_4374, w_063_4377, w_063_4379, w_063_4381, w_063_4384, w_063_4385, w_063_4386, w_063_4387, w_063_4388, w_063_4392, w_063_4393, w_063_4394, w_063_4396, w_063_4397, w_063_4398, w_063_4399, w_063_4400, w_063_4404, w_063_4405, w_063_4407, w_063_4409, w_063_4411, w_063_4412, w_063_4414, w_063_4415, w_063_4417, w_063_4419, w_063_4422, w_063_4423, w_063_4424, w_063_4425, w_063_4426, w_063_4427, w_063_4428, w_063_4429, w_063_4431, w_063_4434, w_063_4436, w_063_4438, w_063_4442, w_063_4444, w_063_4445, w_063_4446, w_063_4447, w_063_4451, w_063_4454, w_063_4456, w_063_4457, w_063_4459, w_063_4460, w_063_4463, w_063_4464, w_063_4465, w_063_4466, w_063_4467, w_063_4469, w_063_4470, w_063_4471, w_063_4472, w_063_4473, w_063_4474, w_063_4475, w_063_4476, w_063_4477, w_063_4478, w_063_4481, w_063_4482, w_063_4483, w_063_4485, w_063_4486, w_063_4487, w_063_4490, w_063_4498, w_063_4499, w_063_4501, w_063_4504, w_063_4506, w_063_4507, w_063_4508, w_063_4511, w_063_4513, w_063_4514, w_063_4516, w_063_4517, w_063_4519, w_063_4520, w_063_4521, w_063_4522, w_063_4523, w_063_4524, w_063_4526, w_063_4528, w_063_4529, w_063_4531, w_063_4532, w_063_4533, w_063_4534, w_063_4537, w_063_4540, w_063_4541, w_063_4543, w_063_4544, w_063_4545, w_063_4547, w_063_4550, w_063_4551, w_063_4552, w_063_4553, w_063_4554, w_063_4555, w_063_4557, w_063_4558, w_063_4559, w_063_4561, w_063_4562, w_063_4563, w_063_4565, w_063_4568, w_063_4569, w_063_4570, w_063_4571, w_063_4573, w_063_4574, w_063_4575, w_063_4578, w_063_4579, w_063_4580, w_063_4585, w_063_4586, w_063_4587, w_063_4589, w_063_4593, w_063_4594, w_063_4595, w_063_4596, w_063_4598, w_063_4599, w_063_4600, w_063_4604, w_063_4605, w_063_4606, w_063_4609, w_063_4612, w_063_4613, w_063_4614, w_063_4616, w_063_4617, w_063_4618, w_063_4619, w_063_4620, w_063_4623, w_063_4624, w_063_4626, w_063_4627, w_063_4629, w_063_4631, w_063_4634, w_063_4635, w_063_4639, w_063_4642, w_063_4646, w_063_4647, w_063_4650, w_063_4652, w_063_4654, w_063_4655, w_063_4658, w_063_4661, w_063_4662, w_063_4663, w_063_4664, w_063_4668, w_063_4669, w_063_4672, w_063_4674, w_063_4676, w_063_4679, w_063_4681, w_063_4685, w_063_4686, w_063_4687, w_063_4688, w_063_4689, w_063_4690, w_063_4691, w_063_4692, w_063_4693, w_063_4694, w_063_4695, w_063_4701, w_063_4702, w_063_4705, w_063_4709, w_063_4710, w_063_4711, w_063_4712, w_063_4714, w_063_4715, w_063_4716, w_063_4717, w_063_4719, w_063_4727, w_063_4728, w_063_4730, w_063_4731, w_063_4732, w_063_4733, w_063_4734, w_063_4735, w_063_4736, w_063_4738, w_063_4739, w_063_4740, w_063_4741, w_063_4743, w_063_4744, w_063_4745, w_063_4746, w_063_4747, w_063_4749, w_063_4750, w_063_4757, w_063_4758, w_063_4759, w_063_4761, w_063_4762, w_063_4765, w_063_4766, w_063_4767, w_063_4769, w_063_4775, w_063_4776, w_063_4778, w_063_4780, w_063_4783, w_063_4786, w_063_4787, w_063_4788, w_063_4789, w_063_4792, w_063_4794, w_063_4795, w_063_4797, w_063_4799, w_063_4800, w_063_4802, w_063_4803, w_063_4805, w_063_4806, w_063_4813, w_063_4814, w_063_4818, w_063_4819, w_063_4820, w_063_4823, w_063_4825, w_063_4826, w_063_4827, w_063_4828, w_063_4829, w_063_4834, w_063_4835, w_063_4836, w_063_4837, w_063_4840, w_063_4841, w_063_4843, w_063_4844, w_063_4847, w_063_4848, w_063_4851, w_063_4852, w_063_4853, w_063_4855, w_063_4856, w_063_4857, w_063_4858, w_063_4861, w_063_4862, w_063_4865, w_063_4866, w_063_4869, w_063_4870, w_063_4871, w_063_4872, w_063_4877, w_063_4878, w_063_4879, w_063_4881, w_063_4883, w_063_4884, w_063_4885, w_063_4887, w_063_4891, w_063_4893, w_063_4894, w_063_4895, w_063_4896, w_063_4897, w_063_4898, w_063_4900, w_063_4901;
  wire w_064_000, w_064_001, w_064_002, w_064_003, w_064_004, w_064_005, w_064_006, w_064_008, w_064_009, w_064_011, w_064_012, w_064_013, w_064_014, w_064_015, w_064_016, w_064_017, w_064_018, w_064_019, w_064_020, w_064_021, w_064_022, w_064_023, w_064_024, w_064_025, w_064_026, w_064_028, w_064_029, w_064_030, w_064_031, w_064_032, w_064_033, w_064_034, w_064_035, w_064_036, w_064_037, w_064_038, w_064_039, w_064_041, w_064_042, w_064_043, w_064_045, w_064_046, w_064_047, w_064_048, w_064_049, w_064_050, w_064_051, w_064_052, w_064_053, w_064_054, w_064_055, w_064_056, w_064_057, w_064_058, w_064_059, w_064_060, w_064_061, w_064_062, w_064_063, w_064_064, w_064_065, w_064_067, w_064_068, w_064_071, w_064_072, w_064_073, w_064_074, w_064_075, w_064_078, w_064_079, w_064_080, w_064_081, w_064_082, w_064_083, w_064_084, w_064_086, w_064_087, w_064_088, w_064_089, w_064_090, w_064_092, w_064_093, w_064_094, w_064_095, w_064_096, w_064_098, w_064_099, w_064_101, w_064_102, w_064_103, w_064_104, w_064_105, w_064_106, w_064_107, w_064_108, w_064_109, w_064_111, w_064_112, w_064_113, w_064_114, w_064_115, w_064_116, w_064_118, w_064_119, w_064_120, w_064_121, w_064_123, w_064_125, w_064_127, w_064_128, w_064_130, w_064_132, w_064_133, w_064_134, w_064_135, w_064_137, w_064_138, w_064_139, w_064_140, w_064_143, w_064_144, w_064_145, w_064_146, w_064_148, w_064_149, w_064_150, w_064_151, w_064_152, w_064_153, w_064_154, w_064_155, w_064_156, w_064_157, w_064_158, w_064_159, w_064_160, w_064_161, w_064_164, w_064_165, w_064_166, w_064_168, w_064_169, w_064_170, w_064_171, w_064_172, w_064_173, w_064_174, w_064_175, w_064_176, w_064_177, w_064_178, w_064_179, w_064_180, w_064_181, w_064_182, w_064_183, w_064_184, w_064_186, w_064_187, w_064_188, w_064_190, w_064_191, w_064_192, w_064_193, w_064_194, w_064_195, w_064_199, w_064_200, w_064_201, w_064_203, w_064_204, w_064_205, w_064_206, w_064_207, w_064_209, w_064_210, w_064_211, w_064_213, w_064_214, w_064_216, w_064_217, w_064_218, w_064_219, w_064_220, w_064_221, w_064_222, w_064_223, w_064_224, w_064_225, w_064_226, w_064_227, w_064_230, w_064_231, w_064_233, w_064_234, w_064_235, w_064_236, w_064_238, w_064_239, w_064_240, w_064_242, w_064_243, w_064_244, w_064_245, w_064_246, w_064_247, w_064_248, w_064_249, w_064_250, w_064_251, w_064_253, w_064_254, w_064_255, w_064_256, w_064_257, w_064_258, w_064_259, w_064_260, w_064_261, w_064_262, w_064_263, w_064_265, w_064_266, w_064_268, w_064_269, w_064_270, w_064_271, w_064_272, w_064_273, w_064_274, w_064_275, w_064_276, w_064_277, w_064_278, w_064_279, w_064_280, w_064_281, w_064_283, w_064_284, w_064_285, w_064_286, w_064_287, w_064_288, w_064_290, w_064_291, w_064_293, w_064_294, w_064_296, w_064_297, w_064_298, w_064_299, w_064_300, w_064_301, w_064_302, w_064_303, w_064_304, w_064_305, w_064_306, w_064_308, w_064_309, w_064_310, w_064_311, w_064_312, w_064_313, w_064_315, w_064_316, w_064_317, w_064_318, w_064_320, w_064_321, w_064_322, w_064_323, w_064_324, w_064_325, w_064_326, w_064_327, w_064_328, w_064_331, w_064_332, w_064_333, w_064_334, w_064_336, w_064_337, w_064_339, w_064_340, w_064_341, w_064_342, w_064_344, w_064_345, w_064_346, w_064_347, w_064_348, w_064_349, w_064_350, w_064_352, w_064_353, w_064_354, w_064_356, w_064_357, w_064_358, w_064_359, w_064_360, w_064_361, w_064_363, w_064_364, w_064_366, w_064_367, w_064_368, w_064_369, w_064_372, w_064_373, w_064_376, w_064_377, w_064_378, w_064_379, w_064_380, w_064_381, w_064_382, w_064_383, w_064_384, w_064_385, w_064_386, w_064_387, w_064_389, w_064_390, w_064_391, w_064_392, w_064_393, w_064_394, w_064_395, w_064_396, w_064_397, w_064_398, w_064_399, w_064_400, w_064_401, w_064_402, w_064_403, w_064_404, w_064_405, w_064_406, w_064_407, w_064_408, w_064_409, w_064_410, w_064_411, w_064_412, w_064_413, w_064_414, w_064_415, w_064_417, w_064_418, w_064_419, w_064_420, w_064_421, w_064_422, w_064_423, w_064_425, w_064_426, w_064_427, w_064_428, w_064_429, w_064_431, w_064_432, w_064_433, w_064_435, w_064_436, w_064_437, w_064_438, w_064_439, w_064_440, w_064_441, w_064_442, w_064_443, w_064_444, w_064_445, w_064_446, w_064_447, w_064_450, w_064_451, w_064_452, w_064_454, w_064_455, w_064_457, w_064_459, w_064_461, w_064_462, w_064_463, w_064_464, w_064_465, w_064_466, w_064_467, w_064_468, w_064_469, w_064_470, w_064_471, w_064_472, w_064_474, w_064_475, w_064_476, w_064_477, w_064_478, w_064_479, w_064_481, w_064_482, w_064_483, w_064_485, w_064_486, w_064_487, w_064_488, w_064_489, w_064_490, w_064_491, w_064_492, w_064_493, w_064_494, w_064_496, w_064_497, w_064_498, w_064_499, w_064_502, w_064_505, w_064_506, w_064_507, w_064_508, w_064_509, w_064_510, w_064_512, w_064_513, w_064_514, w_064_515, w_064_516, w_064_518, w_064_519, w_064_520, w_064_521, w_064_523, w_064_524, w_064_525, w_064_526, w_064_528, w_064_531, w_064_532, w_064_534, w_064_535, w_064_536, w_064_537, w_064_538, w_064_540, w_064_541, w_064_542, w_064_544, w_064_546, w_064_547, w_064_548, w_064_550, w_064_551, w_064_554, w_064_555, w_064_556, w_064_557, w_064_558, w_064_559, w_064_560, w_064_561, w_064_562, w_064_563, w_064_565, w_064_566, w_064_567, w_064_568, w_064_569, w_064_570, w_064_571, w_064_572, w_064_573, w_064_575, w_064_576, w_064_577, w_064_578, w_064_579, w_064_580, w_064_581, w_064_582, w_064_583, w_064_584, w_064_585, w_064_586, w_064_587, w_064_588, w_064_590, w_064_592, w_064_593, w_064_594, w_064_595, w_064_596, w_064_597, w_064_599, w_064_601, w_064_602, w_064_603, w_064_605, w_064_606, w_064_608, w_064_609, w_064_610, w_064_612, w_064_613, w_064_614, w_064_615, w_064_617, w_064_620, w_064_622, w_064_623, w_064_625, w_064_626, w_064_627, w_064_628, w_064_629, w_064_630, w_064_631, w_064_632, w_064_633, w_064_634, w_064_635, w_064_636, w_064_637, w_064_638, w_064_639, w_064_640, w_064_641, w_064_642, w_064_643, w_064_644, w_064_645, w_064_646, w_064_647, w_064_648, w_064_651, w_064_652, w_064_653, w_064_655, w_064_656, w_064_657, w_064_658, w_064_659, w_064_660, w_064_661, w_064_662, w_064_663, w_064_664, w_064_665, w_064_666, w_064_667, w_064_668, w_064_671, w_064_672, w_064_673, w_064_674, w_064_675, w_064_676, w_064_677, w_064_678, w_064_679, w_064_680, w_064_681, w_064_682, w_064_683, w_064_684, w_064_688, w_064_690, w_064_693, w_064_695, w_064_696, w_064_697, w_064_698, w_064_699, w_064_702, w_064_703, w_064_705, w_064_707, w_064_708, w_064_709, w_064_710, w_064_711, w_064_713, w_064_714, w_064_715, w_064_716, w_064_717, w_064_718, w_064_719, w_064_721, w_064_722, w_064_724, w_064_727, w_064_728, w_064_729, w_064_730, w_064_731, w_064_732, w_064_733, w_064_734, w_064_735, w_064_736, w_064_737, w_064_738, w_064_739, w_064_740, w_064_741, w_064_742, w_064_743, w_064_744, w_064_745, w_064_746, w_064_747, w_064_748, w_064_749, w_064_750, w_064_751, w_064_752, w_064_753, w_064_754, w_064_757, w_064_758, w_064_759, w_064_760, w_064_761, w_064_762, w_064_763, w_064_764, w_064_765, w_064_766, w_064_767, w_064_768, w_064_769, w_064_770, w_064_771, w_064_772, w_064_773, w_064_774, w_064_775, w_064_776, w_064_777, w_064_781, w_064_782, w_064_783, w_064_784, w_064_785, w_064_787, w_064_788, w_064_789, w_064_790, w_064_792, w_064_793, w_064_795, w_064_797, w_064_798, w_064_799, w_064_801, w_064_803, w_064_804, w_064_806, w_064_807, w_064_808, w_064_809, w_064_810, w_064_811, w_064_812, w_064_813, w_064_814, w_064_815, w_064_818, w_064_820, w_064_821, w_064_822, w_064_823, w_064_824, w_064_826, w_064_827, w_064_828, w_064_829, w_064_830, w_064_831, w_064_832, w_064_833, w_064_834, w_064_835, w_064_836, w_064_838, w_064_840, w_064_842, w_064_843, w_064_844, w_064_845, w_064_846, w_064_847, w_064_848, w_064_849, w_064_850, w_064_851, w_064_852, w_064_853, w_064_854, w_064_855, w_064_856, w_064_857, w_064_858, w_064_859, w_064_860, w_064_861, w_064_862, w_064_863, w_064_864, w_064_865, w_064_866, w_064_867, w_064_868, w_064_870, w_064_871, w_064_872, w_064_873, w_064_874, w_064_875, w_064_877, w_064_878, w_064_879, w_064_880, w_064_881, w_064_882, w_064_884, w_064_885, w_064_886, w_064_887, w_064_888, w_064_889, w_064_890, w_064_891, w_064_892, w_064_893, w_064_894, w_064_895, w_064_896, w_064_897, w_064_899, w_064_902, w_064_903, w_064_904, w_064_905, w_064_907, w_064_908, w_064_909, w_064_910, w_064_911, w_064_913, w_064_914, w_064_916, w_064_917, w_064_918, w_064_920, w_064_922, w_064_924, w_064_926, w_064_927, w_064_928, w_064_929, w_064_930, w_064_931, w_064_932, w_064_934, w_064_936, w_064_937, w_064_938, w_064_939, w_064_940, w_064_941, w_064_942, w_064_944, w_064_946, w_064_948, w_064_949, w_064_950, w_064_952, w_064_953, w_064_954, w_064_955, w_064_957, w_064_958, w_064_959, w_064_961, w_064_962, w_064_963, w_064_964, w_064_965, w_064_966, w_064_968, w_064_970, w_064_971, w_064_974, w_064_975, w_064_976, w_064_977, w_064_978, w_064_979, w_064_980, w_064_981, w_064_982, w_064_984, w_064_985, w_064_986, w_064_987, w_064_988, w_064_989, w_064_990, w_064_992, w_064_995, w_064_996, w_064_997, w_064_998, w_064_999, w_064_1000, w_064_1003, w_064_1006, w_064_1007, w_064_1008, w_064_1009, w_064_1010, w_064_1011, w_064_1013, w_064_1014, w_064_1016, w_064_1017, w_064_1018, w_064_1019, w_064_1020, w_064_1021, w_064_1022, w_064_1023, w_064_1024, w_064_1025, w_064_1026, w_064_1027, w_064_1028, w_064_1031, w_064_1032, w_064_1033, w_064_1034, w_064_1035, w_064_1036, w_064_1037, w_064_1038, w_064_1039, w_064_1041, w_064_1042, w_064_1043, w_064_1044, w_064_1045, w_064_1047, w_064_1048, w_064_1049, w_064_1050, w_064_1051, w_064_1052, w_064_1053, w_064_1055, w_064_1056, w_064_1057, w_064_1058, w_064_1059, w_064_1060, w_064_1061, w_064_1062, w_064_1063, w_064_1067, w_064_1068, w_064_1069, w_064_1070, w_064_1071, w_064_1072, w_064_1074, w_064_1076, w_064_1077, w_064_1078, w_064_1079, w_064_1080, w_064_1081, w_064_1083, w_064_1085, w_064_1086, w_064_1088, w_064_1089, w_064_1090, w_064_1093, w_064_1094, w_064_1095, w_064_1096, w_064_1097, w_064_1099, w_064_1100, w_064_1101, w_064_1102, w_064_1104, w_064_1106, w_064_1108, w_064_1109, w_064_1110, w_064_1112, w_064_1113, w_064_1115, w_064_1117, w_064_1118, w_064_1119, w_064_1120, w_064_1121, w_064_1122, w_064_1123, w_064_1124, w_064_1125, w_064_1127, w_064_1128, w_064_1129, w_064_1131, w_064_1132, w_064_1133, w_064_1135, w_064_1136, w_064_1137, w_064_1138, w_064_1139, w_064_1140, w_064_1142, w_064_1143, w_064_1145, w_064_1146, w_064_1147, w_064_1148, w_064_1149, w_064_1150, w_064_1151, w_064_1153, w_064_1154, w_064_1155, w_064_1156, w_064_1158, w_064_1160, w_064_1161, w_064_1162, w_064_1163, w_064_1164, w_064_1166, w_064_1167, w_064_1168, w_064_1169, w_064_1171, w_064_1174, w_064_1176, w_064_1177, w_064_1178, w_064_1179, w_064_1180, w_064_1182, w_064_1184, w_064_1185, w_064_1186, w_064_1187, w_064_1188, w_064_1189, w_064_1190, w_064_1191, w_064_1193, w_064_1194, w_064_1195, w_064_1196, w_064_1197, w_064_1198, w_064_1199, w_064_1200, w_064_1202, w_064_1203, w_064_1204, w_064_1205, w_064_1207, w_064_1208, w_064_1209, w_064_1211, w_064_1212, w_064_1215, w_064_1216, w_064_1217, w_064_1218, w_064_1219, w_064_1220, w_064_1221, w_064_1223, w_064_1224, w_064_1225, w_064_1227, w_064_1228, w_064_1229, w_064_1231, w_064_1233, w_064_1234, w_064_1235, w_064_1236, w_064_1237, w_064_1238, w_064_1241, w_064_1243, w_064_1244, w_064_1245, w_064_1251, w_064_1252, w_064_1254, w_064_1255, w_064_1256, w_064_1257, w_064_1258, w_064_1261, w_064_1262, w_064_1263, w_064_1264, w_064_1265, w_064_1266, w_064_1267, w_064_1268, w_064_1269, w_064_1270, w_064_1271, w_064_1272, w_064_1273, w_064_1274, w_064_1275, w_064_1276, w_064_1277, w_064_1279, w_064_1280, w_064_1281, w_064_1282, w_064_1283, w_064_1285, w_064_1287, w_064_1288, w_064_1289, w_064_1290, w_064_1291, w_064_1292, w_064_1293, w_064_1295, w_064_1297, w_064_1298, w_064_1299, w_064_1300, w_064_1301, w_064_1303, w_064_1304, w_064_1305, w_064_1306, w_064_1307, w_064_1308, w_064_1309, w_064_1310, w_064_1311, w_064_1314, w_064_1315, w_064_1316, w_064_1317, w_064_1319, w_064_1320, w_064_1321, w_064_1322, w_064_1323, w_064_1326, w_064_1327, w_064_1328, w_064_1329, w_064_1330, w_064_1332, w_064_1334, w_064_1335, w_064_1336, w_064_1337, w_064_1339, w_064_1340, w_064_1341, w_064_1342, w_064_1345, w_064_1346, w_064_1347, w_064_1349, w_064_1350, w_064_1351, w_064_1352, w_064_1353, w_064_1354, w_064_1356, w_064_1357, w_064_1359, w_064_1360, w_064_1362, w_064_1364, w_064_1365, w_064_1367, w_064_1369, w_064_1370, w_064_1371, w_064_1372, w_064_1374, w_064_1379, w_064_1380, w_064_1381, w_064_1384, w_064_1385, w_064_1386, w_064_1387, w_064_1388, w_064_1390, w_064_1391, w_064_1392, w_064_1393, w_064_1396, w_064_1397, w_064_1398, w_064_1400, w_064_1401, w_064_1402, w_064_1403, w_064_1404, w_064_1405, w_064_1408, w_064_1410, w_064_1412, w_064_1414, w_064_1415, w_064_1416, w_064_1417, w_064_1418, w_064_1419, w_064_1420, w_064_1426, w_064_1427, w_064_1428, w_064_1431, w_064_1432, w_064_1434, w_064_1435, w_064_1437, w_064_1439, w_064_1440, w_064_1441, w_064_1442, w_064_1443, w_064_1444, w_064_1445, w_064_1446, w_064_1447, w_064_1448, w_064_1449, w_064_1450, w_064_1451, w_064_1452, w_064_1453, w_064_1454, w_064_1456, w_064_1458, w_064_1459, w_064_1461, w_064_1462, w_064_1464, w_064_1468, w_064_1469, w_064_1470, w_064_1471, w_064_1472, w_064_1473, w_064_1474, w_064_1475, w_064_1477, w_064_1479, w_064_1480, w_064_1481, w_064_1483, w_064_1484, w_064_1485, w_064_1486, w_064_1487, w_064_1490, w_064_1491, w_064_1492, w_064_1493, w_064_1494, w_064_1495, w_064_1496, w_064_1497, w_064_1499, w_064_1501, w_064_1503, w_064_1504, w_064_1505, w_064_1506, w_064_1507, w_064_1508, w_064_1509, w_064_1510, w_064_1512, w_064_1513, w_064_1514, w_064_1515, w_064_1516, w_064_1517, w_064_1518, w_064_1519, w_064_1521, w_064_1522, w_064_1524, w_064_1525, w_064_1526, w_064_1528, w_064_1529, w_064_1530, w_064_1531, w_064_1533, w_064_1534, w_064_1535, w_064_1537, w_064_1538, w_064_1539, w_064_1540, w_064_1541, w_064_1542, w_064_1543, w_064_1544, w_064_1545, w_064_1546, w_064_1548, w_064_1549, w_064_1550, w_064_1551, w_064_1553, w_064_1554, w_064_1555, w_064_1556, w_064_1557, w_064_1558, w_064_1561, w_064_1562, w_064_1564, w_064_1565, w_064_1566, w_064_1567, w_064_1568, w_064_1570, w_064_1571, w_064_1572, w_064_1573, w_064_1576, w_064_1578, w_064_1580, w_064_1581, w_064_1582, w_064_1583, w_064_1584, w_064_1585, w_064_1587, w_064_1589, w_064_1592, w_064_1593, w_064_1594, w_064_1595, w_064_1596, w_064_1597, w_064_1598, w_064_1599, w_064_1600, w_064_1601, w_064_1602, w_064_1603, w_064_1604, w_064_1606, w_064_1607, w_064_1608, w_064_1609, w_064_1610, w_064_1611, w_064_1612, w_064_1613, w_064_1614, w_064_1615, w_064_1616, w_064_1617, w_064_1618, w_064_1620, w_064_1622, w_064_1623, w_064_1625, w_064_1626, w_064_1628, w_064_1629, w_064_1630, w_064_1632, w_064_1635, w_064_1636, w_064_1637, w_064_1638, w_064_1639, w_064_1641, w_064_1642, w_064_1644, w_064_1646, w_064_1647, w_064_1648, w_064_1649, w_064_1653, w_064_1654, w_064_1655, w_064_1656, w_064_1657, w_064_1658, w_064_1659, w_064_1660, w_064_1661, w_064_1662, w_064_1663, w_064_1664, w_064_1665, w_064_1666, w_064_1667, w_064_1668, w_064_1670, w_064_1671, w_064_1674, w_064_1677, w_064_1680, w_064_1681, w_064_1682, w_064_1683, w_064_1684, w_064_1685, w_064_1686, w_064_1688, w_064_1690, w_064_1691, w_064_1692, w_064_1694, w_064_1695, w_064_1697, w_064_1698, w_064_1700, w_064_1701, w_064_1703, w_064_1706, w_064_1709, w_064_1710, w_064_1711, w_064_1712, w_064_1713, w_064_1716, w_064_1717, w_064_1718, w_064_1719, w_064_1721, w_064_1722, w_064_1723, w_064_1724, w_064_1725, w_064_1727, w_064_1728, w_064_1729, w_064_1730, w_064_1731, w_064_1732, w_064_1733, w_064_1734, w_064_1736, w_064_1737, w_064_1739, w_064_1740, w_064_1741, w_064_1743, w_064_1746, w_064_1747, w_064_1748, w_064_1749, w_064_1755, w_064_1756, w_064_1757, w_064_1758, w_064_1760, w_064_1762, w_064_1765, w_064_1767, w_064_1768, w_064_1769, w_064_1770, w_064_1771, w_064_1772, w_064_1773, w_064_1774, w_064_1775, w_064_1776, w_064_1777, w_064_1779, w_064_1780, w_064_1781, w_064_1782, w_064_1783, w_064_1784, w_064_1785, w_064_1788, w_064_1789, w_064_1790, w_064_1791, w_064_1792, w_064_1793, w_064_1794, w_064_1795, w_064_1796, w_064_1797, w_064_1798, w_064_1799, w_064_1800, w_064_1801, w_064_1802, w_064_1803, w_064_1804, w_064_1808, w_064_1810, w_064_1811, w_064_1812, w_064_1814, w_064_1816, w_064_1817, w_064_1818, w_064_1820, w_064_1821, w_064_1822, w_064_1823, w_064_1824, w_064_1825, w_064_1826, w_064_1827, w_064_1828, w_064_1830, w_064_1831, w_064_1832, w_064_1834, w_064_1835, w_064_1836, w_064_1837, w_064_1838, w_064_1839, w_064_1841, w_064_1842, w_064_1843, w_064_1844, w_064_1845, w_064_1849, w_064_1850, w_064_1851, w_064_1852, w_064_1853, w_064_1855, w_064_1856, w_064_1857, w_064_1858, w_064_1859, w_064_1860, w_064_1862, w_064_1863, w_064_1864, w_064_1865, w_064_1866, w_064_1867, w_064_1868, w_064_1869, w_064_1870, w_064_1871, w_064_1872, w_064_1875, w_064_1876, w_064_1879, w_064_1881, w_064_1882, w_064_1883, w_064_1884, w_064_1885, w_064_1886, w_064_1887, w_064_1889, w_064_1890, w_064_1891, w_064_1892, w_064_1894, w_064_1896, w_064_1897, w_064_1898, w_064_1900, w_064_1901, w_064_1902, w_064_1904, w_064_1905, w_064_1906, w_064_1907, w_064_1909, w_064_1910, w_064_1912, w_064_1914, w_064_1915, w_064_1916, w_064_1918, w_064_1919, w_064_1920, w_064_1921, w_064_1922, w_064_1923, w_064_1925, w_064_1926, w_064_1928, w_064_1929, w_064_1931, w_064_1932, w_064_1933, w_064_1934, w_064_1937, w_064_1939, w_064_1940, w_064_1941, w_064_1942, w_064_1943, w_064_1944, w_064_1946, w_064_1947, w_064_1948, w_064_1949, w_064_1951, w_064_1952, w_064_1954, w_064_1955, w_064_1956, w_064_1957, w_064_1960, w_064_1961, w_064_1962, w_064_1963, w_064_1964, w_064_1965, w_064_1966, w_064_1967, w_064_1968, w_064_1969, w_064_1971, w_064_1972, w_064_1973, w_064_1974, w_064_1975, w_064_1976, w_064_1978, w_064_1980, w_064_1981, w_064_1982, w_064_1983, w_064_1984, w_064_1985, w_064_1986, w_064_1987, w_064_1988, w_064_1989, w_064_1990, w_064_1991, w_064_1992, w_064_1993, w_064_1994, w_064_1995, w_064_1996, w_064_1997, w_064_1998, w_064_1999, w_064_2001, w_064_2002, w_064_2003, w_064_2006, w_064_2007, w_064_2008, w_064_2009, w_064_2011, w_064_2012, w_064_2013, w_064_2015, w_064_2016, w_064_2017, w_064_2018, w_064_2019, w_064_2020, w_064_2021, w_064_2022, w_064_2023, w_064_2024, w_064_2026, w_064_2027, w_064_2028, w_064_2030, w_064_2031, w_064_2032, w_064_2034, w_064_2036, w_064_2037, w_064_2038, w_064_2039, w_064_2041, w_064_2042, w_064_2043, w_064_2048, w_064_2049, w_064_2050, w_064_2051, w_064_2052, w_064_2053, w_064_2055, w_064_2057, w_064_2058, w_064_2059, w_064_2060, w_064_2061, w_064_2062, w_064_2064, w_064_2066, w_064_2067, w_064_2069, w_064_2070, w_064_2071, w_064_2073, w_064_2074, w_064_2075, w_064_2077, w_064_2078, w_064_2079, w_064_2081, w_064_2086, w_064_2087, w_064_2088, w_064_2091, w_064_2092, w_064_2094, w_064_2096, w_064_2098, w_064_2099, w_064_2102, w_064_2103, w_064_2104, w_064_2105, w_064_2106, w_064_2108, w_064_2109, w_064_2111, w_064_2112, w_064_2113, w_064_2114, w_064_2115, w_064_2116, w_064_2119, w_064_2121, w_064_2122, w_064_2125, w_064_2126, w_064_2127, w_064_2128, w_064_2129, w_064_2130, w_064_2132, w_064_2133, w_064_2134, w_064_2135, w_064_2136, w_064_2137, w_064_2140, w_064_2141, w_064_2143, w_064_2144, w_064_2145, w_064_2146, w_064_2147, w_064_2148, w_064_2149, w_064_2150, w_064_2151, w_064_2152, w_064_2153, w_064_2156, w_064_2157, w_064_2158, w_064_2159, w_064_2160, w_064_2161, w_064_2162, w_064_2163, w_064_2165, w_064_2166, w_064_2168, w_064_2169, w_064_2170, w_064_2171, w_064_2174, w_064_2175, w_064_2176, w_064_2177, w_064_2178, w_064_2179, w_064_2181, w_064_2182, w_064_2185, w_064_2187, w_064_2188, w_064_2189, w_064_2190, w_064_2192, w_064_2193, w_064_2194, w_064_2196, w_064_2197, w_064_2198, w_064_2199, w_064_2200, w_064_2202, w_064_2203, w_064_2204, w_064_2207, w_064_2208, w_064_2210, w_064_2211, w_064_2212, w_064_2213, w_064_2215, w_064_2216, w_064_2217, w_064_2218, w_064_2220, w_064_2221, w_064_2224, w_064_2226, w_064_2227, w_064_2228, w_064_2229, w_064_2232, w_064_2233, w_064_2234, w_064_2235, w_064_2236, w_064_2237, w_064_2239, w_064_2240, w_064_2242, w_064_2244, w_064_2246, w_064_2247, w_064_2248, w_064_2249, w_064_2251, w_064_2253, w_064_2254, w_064_2255, w_064_2256, w_064_2257, w_064_2258, w_064_2259, w_064_2260, w_064_2261, w_064_2262, w_064_2264, w_064_2265, w_064_2266, w_064_2267, w_064_2268, w_064_2270, w_064_2271, w_064_2272, w_064_2273, w_064_2274, w_064_2275, w_064_2276, w_064_2277, w_064_2280, w_064_2281, w_064_2282, w_064_2284, w_064_2285, w_064_2286, w_064_2287, w_064_2288, w_064_2289, w_064_2292, w_064_2293, w_064_2294, w_064_2297, w_064_2299, w_064_2300, w_064_2302, w_064_2303, w_064_2304, w_064_2305, w_064_2306, w_064_2307, w_064_2308, w_064_2309, w_064_2310, w_064_2313, w_064_2314, w_064_2316, w_064_2317, w_064_2319, w_064_2320, w_064_2321, w_064_2325, w_064_2326, w_064_2327, w_064_2328, w_064_2329, w_064_2331, w_064_2332, w_064_2333, w_064_2334, w_064_2335, w_064_2336, w_064_2337, w_064_2340, w_064_2341, w_064_2343, w_064_2344, w_064_2345, w_064_2346, w_064_2348, w_064_2349, w_064_2351, w_064_2352, w_064_2353, w_064_2354, w_064_2355, w_064_2356, w_064_2358, w_064_2359, w_064_2361, w_064_2362, w_064_2363, w_064_2366, w_064_2369, w_064_2370, w_064_2371, w_064_2372, w_064_2375, w_064_2377, w_064_2378, w_064_2380, w_064_2381, w_064_2382, w_064_2383, w_064_2384, w_064_2385, w_064_2386, w_064_2388, w_064_2390, w_064_2391, w_064_2394, w_064_2395, w_064_2396, w_064_2398, w_064_2399, w_064_2400, w_064_2401, w_064_2402, w_064_2403, w_064_2404, w_064_2405, w_064_2406, w_064_2407, w_064_2408, w_064_2409, w_064_2413, w_064_2414, w_064_2415, w_064_2418, w_064_2419, w_064_2421, w_064_2423, w_064_2425, w_064_2426, w_064_2427, w_064_2428, w_064_2429, w_064_2430, w_064_2431, w_064_2432, w_064_2433, w_064_2434, w_064_2435, w_064_2438, w_064_2440, w_064_2441, w_064_2443, w_064_2444, w_064_2445, w_064_2448, w_064_2450, w_064_2452, w_064_2453, w_064_2454, w_064_2456, w_064_2457, w_064_2459, w_064_2460, w_064_2461, w_064_2462, w_064_2463, w_064_2465, w_064_2466, w_064_2467, w_064_2469, w_064_2470, w_064_2471, w_064_2472, w_064_2474, w_064_2475, w_064_2476, w_064_2478, w_064_2479, w_064_2480, w_064_2481, w_064_2482, w_064_2483, w_064_2485, w_064_2488, w_064_2489, w_064_2491, w_064_2492, w_064_2493, w_064_2494, w_064_2495, w_064_2497, w_064_2499, w_064_2500, w_064_2501, w_064_2502, w_064_2503, w_064_2505, w_064_2507, w_064_2508, w_064_2509, w_064_2510, w_064_2511, w_064_2512, w_064_2513, w_064_2515, w_064_2517, w_064_2518, w_064_2519, w_064_2520, w_064_2521, w_064_2522, w_064_2524, w_064_2525, w_064_2526, w_064_2527, w_064_2528, w_064_2529, w_064_2530, w_064_2532, w_064_2533, w_064_2534, w_064_2537, w_064_2539, w_064_2541, w_064_2542, w_064_2543, w_064_2544, w_064_2546, w_064_2548, w_064_2549, w_064_2550, w_064_2552, w_064_2554, w_064_2555, w_064_2556, w_064_2557, w_064_2561, w_064_2563, w_064_2564, w_064_2565, w_064_2566, w_064_2567, w_064_2568, w_064_2570, w_064_2571, w_064_2573, w_064_2574, w_064_2576, w_064_2577, w_064_2578, w_064_2579, w_064_2580, w_064_2581, w_064_2582, w_064_2583, w_064_2584, w_064_2585, w_064_2587, w_064_2591, w_064_2595, w_064_2596, w_064_2598, w_064_2599, w_064_2601, w_064_2602, w_064_2603, w_064_2605, w_064_2606, w_064_2607, w_064_2609, w_064_2610, w_064_2611, w_064_2612, w_064_2613, w_064_2614, w_064_2615, w_064_2616, w_064_2619, w_064_2621, w_064_2622, w_064_2623, w_064_2624, w_064_2625, w_064_2627, w_064_2628, w_064_2629, w_064_2630, w_064_2631, w_064_2632, w_064_2633, w_064_2634, w_064_2636, w_064_2637, w_064_2639, w_064_2640, w_064_2641, w_064_2642, w_064_2643, w_064_2645, w_064_2647, w_064_2648, w_064_2649, w_064_2650, w_064_2652, w_064_2654, w_064_2655, w_064_2657, w_064_2659, w_064_2660, w_064_2661, w_064_2662, w_064_2663, w_064_2664, w_064_2666, w_064_2667, w_064_2668, w_064_2669, w_064_2670, w_064_2671, w_064_2673, w_064_2674, w_064_2675, w_064_2676, w_064_2677, w_064_2678, w_064_2679, w_064_2680, w_064_2681, w_064_2682, w_064_2683, w_064_2685, w_064_2686, w_064_2688, w_064_2690, w_064_2691, w_064_2692, w_064_2693, w_064_2695, w_064_2696, w_064_2697, w_064_2698, w_064_2699, w_064_2700, w_064_2701, w_064_2702, w_064_2703, w_064_2704, w_064_2705, w_064_2707, w_064_2708, w_064_2709, w_064_2710, w_064_2711, w_064_2712, w_064_2713, w_064_2717, w_064_2718, w_064_2719, w_064_2720, w_064_2721, w_064_2722, w_064_2723, w_064_2724, w_064_2725, w_064_2727, w_064_2731, w_064_2732, w_064_2733, w_064_2734, w_064_2735, w_064_2736, w_064_2737, w_064_2739, w_064_2740, w_064_2742, w_064_2746, w_064_2747, w_064_2748, w_064_2749, w_064_2750, w_064_2751, w_064_2752, w_064_2753, w_064_2754, w_064_2757, w_064_2758, w_064_2759, w_064_2760, w_064_2763, w_064_2764, w_064_2765, w_064_2766, w_064_2769, w_064_2770, w_064_2771, w_064_2773, w_064_2774, w_064_2775, w_064_2776, w_064_2779, w_064_2780, w_064_2781, w_064_2783, w_064_2785, w_064_2786, w_064_2788, w_064_2789, w_064_2794, w_064_2795, w_064_2796, w_064_2798, w_064_2799, w_064_2800, w_064_2801, w_064_2802, w_064_2803, w_064_2804, w_064_2805, w_064_2806, w_064_2808, w_064_2809, w_064_2810, w_064_2813, w_064_2814, w_064_2815, w_064_2816, w_064_2817, w_064_2818, w_064_2820, w_064_2822, w_064_2824, w_064_2827, w_064_2828, w_064_2829, w_064_2832, w_064_2833, w_064_2836, w_064_2839, w_064_2840, w_064_2841, w_064_2842, w_064_2843, w_064_2844, w_064_2845, w_064_2847, w_064_2848, w_064_2849, w_064_2850, w_064_2853, w_064_2855, w_064_2857, w_064_2859, w_064_2860, w_064_2864, w_064_2866, w_064_2867, w_064_2868, w_064_2869, w_064_2870, w_064_2871, w_064_2872, w_064_2873, w_064_2875, w_064_2876, w_064_2877, w_064_2880, w_064_2882, w_064_2883, w_064_2884, w_064_2885, w_064_2886, w_064_2888, w_064_2889, w_064_2890, w_064_2891, w_064_2892, w_064_2893, w_064_2894, w_064_2895, w_064_2896, w_064_2897, w_064_2898, w_064_2899, w_064_2902, w_064_2904, w_064_2905, w_064_2906, w_064_2907, w_064_2909, w_064_2910, w_064_2911, w_064_2912, w_064_2913, w_064_2914, w_064_2915, w_064_2916, w_064_2917, w_064_2921, w_064_2923, w_064_2925, w_064_2926, w_064_2927, w_064_2930, w_064_2932, w_064_2935, w_064_2936, w_064_2937, w_064_2939, w_064_2942, w_064_2943, w_064_2944, w_064_2945;
  wire w_065_000, w_065_001, w_065_002, w_065_003, w_065_004, w_065_005, w_065_006, w_065_007, w_065_008, w_065_010, w_065_012, w_065_013, w_065_014, w_065_015, w_065_018, w_065_019, w_065_021, w_065_022, w_065_023, w_065_025, w_065_026, w_065_027, w_065_028, w_065_029, w_065_030, w_065_031, w_065_032, w_065_033, w_065_034, w_065_035, w_065_036, w_065_037, w_065_040, w_065_046, w_065_047, w_065_050, w_065_053, w_065_054, w_065_055, w_065_057, w_065_061, w_065_063, w_065_064, w_065_066, w_065_067, w_065_069, w_065_070, w_065_071, w_065_073, w_065_074, w_065_075, w_065_076, w_065_077, w_065_079, w_065_082, w_065_086, w_065_088, w_065_089, w_065_090, w_065_093, w_065_094, w_065_095, w_065_097, w_065_098, w_065_100, w_065_101, w_065_102, w_065_107, w_065_109, w_065_110, w_065_111, w_065_112, w_065_117, w_065_121, w_065_122, w_065_123, w_065_124, w_065_125, w_065_126, w_065_127, w_065_129, w_065_130, w_065_131, w_065_132, w_065_135, w_065_136, w_065_137, w_065_138, w_065_139, w_065_140, w_065_142, w_065_143, w_065_144, w_065_145, w_065_148, w_065_150, w_065_151, w_065_153, w_065_154, w_065_155, w_065_156, w_065_159, w_065_161, w_065_162, w_065_163, w_065_167, w_065_168, w_065_169, w_065_170, w_065_172, w_065_174, w_065_175, w_065_177, w_065_178, w_065_179, w_065_181, w_065_182, w_065_183, w_065_184, w_065_186, w_065_189, w_065_190, w_065_191, w_065_192, w_065_194, w_065_195, w_065_197, w_065_201, w_065_203, w_065_204, w_065_205, w_065_207, w_065_208, w_065_209, w_065_210, w_065_211, w_065_213, w_065_215, w_065_216, w_065_218, w_065_219, w_065_221, w_065_224, w_065_225, w_065_226, w_065_227, w_065_228, w_065_233, w_065_234, w_065_236, w_065_241, w_065_243, w_065_249, w_065_251, w_065_254, w_065_257, w_065_259, w_065_260, w_065_261, w_065_262, w_065_263, w_065_264, w_065_265, w_065_268, w_065_269, w_065_274, w_065_276, w_065_277, w_065_279, w_065_280, w_065_281, w_065_283, w_065_284, w_065_285, w_065_286, w_065_288, w_065_290, w_065_291, w_065_292, w_065_294, w_065_298, w_065_299, w_065_300, w_065_301, w_065_302, w_065_303, w_065_305, w_065_311, w_065_313, w_065_314, w_065_315, w_065_318, w_065_319, w_065_320, w_065_321, w_065_322, w_065_323, w_065_330, w_065_334, w_065_336, w_065_337, w_065_339, w_065_342, w_065_343, w_065_345, w_065_346, w_065_348, w_065_349, w_065_350, w_065_356, w_065_359, w_065_362, w_065_363, w_065_364, w_065_365, w_065_367, w_065_368, w_065_369, w_065_370, w_065_372, w_065_374, w_065_375, w_065_376, w_065_377, w_065_378, w_065_380, w_065_381, w_065_382, w_065_383, w_065_384, w_065_386, w_065_388, w_065_390, w_065_391, w_065_392, w_065_398, w_065_399, w_065_400, w_065_401, w_065_402, w_065_404, w_065_405, w_065_406, w_065_408, w_065_409, w_065_410, w_065_411, w_065_414, w_065_415, w_065_417, w_065_419, w_065_420, w_065_421, w_065_426, w_065_427, w_065_431, w_065_433, w_065_434, w_065_435, w_065_438, w_065_439, w_065_440, w_065_441, w_065_445, w_065_446, w_065_447, w_065_448, w_065_449, w_065_450, w_065_451, w_065_452, w_065_453, w_065_454, w_065_455, w_065_456, w_065_457, w_065_459, w_065_460, w_065_465, w_065_467, w_065_468, w_065_469, w_065_470, w_065_472, w_065_475, w_065_479, w_065_481, w_065_482, w_065_484, w_065_488, w_065_489, w_065_492, w_065_493, w_065_495, w_065_498, w_065_502, w_065_504, w_065_505, w_065_506, w_065_507, w_065_509, w_065_510, w_065_511, w_065_513, w_065_515, w_065_516, w_065_517, w_065_520, w_065_521, w_065_522, w_065_523, w_065_524, w_065_525, w_065_527, w_065_528, w_065_529, w_065_530, w_065_531, w_065_532, w_065_534, w_065_537, w_065_539, w_065_540, w_065_541, w_065_542, w_065_543, w_065_544, w_065_545, w_065_546, w_065_548, w_065_551, w_065_552, w_065_553, w_065_554, w_065_555, w_065_556, w_065_557, w_065_558, w_065_560, w_065_561, w_065_565, w_065_566, w_065_567, w_065_571, w_065_572, w_065_573, w_065_575, w_065_577, w_065_579, w_065_581, w_065_583, w_065_587, w_065_588, w_065_590, w_065_591, w_065_592, w_065_598, w_065_600, w_065_601, w_065_604, w_065_605, w_065_606, w_065_608, w_065_612, w_065_613, w_065_615, w_065_616, w_065_617, w_065_618, w_065_620, w_065_621, w_065_622, w_065_625, w_065_627, w_065_629, w_065_630, w_065_631, w_065_633, w_065_636, w_065_637, w_065_639, w_065_640, w_065_642, w_065_643, w_065_644, w_065_646, w_065_647, w_065_649, w_065_652, w_065_656, w_065_657, w_065_658, w_065_660, w_065_663, w_065_667, w_065_669, w_065_674, w_065_676, w_065_678, w_065_679, w_065_680, w_065_681, w_065_683, w_065_684, w_065_687, w_065_688, w_065_691, w_065_692, w_065_693, w_065_695, w_065_698, w_065_699, w_065_700, w_065_701, w_065_702, w_065_703, w_065_705, w_065_707, w_065_710, w_065_711, w_065_712, w_065_713, w_065_714, w_065_715, w_065_717, w_065_719, w_065_720, w_065_722, w_065_725, w_065_726, w_065_727, w_065_728, w_065_731, w_065_732, w_065_733, w_065_734, w_065_735, w_065_736, w_065_738, w_065_739, w_065_740, w_065_741, w_065_743, w_065_744, w_065_748, w_065_749, w_065_751, w_065_752, w_065_753, w_065_754, w_065_756, w_065_757, w_065_759, w_065_760, w_065_763, w_065_765, w_065_766, w_065_767, w_065_768, w_065_769, w_065_770, w_065_775, w_065_778, w_065_780, w_065_782, w_065_786, w_065_787, w_065_789, w_065_791, w_065_793, w_065_795, w_065_796, w_065_797, w_065_798, w_065_799, w_065_801, w_065_802, w_065_803, w_065_809, w_065_811, w_065_813, w_065_817, w_065_819, w_065_823, w_065_824, w_065_825, w_065_827, w_065_828, w_065_829, w_065_832, w_065_837, w_065_838, w_065_840, w_065_842, w_065_846, w_065_848, w_065_850, w_065_852, w_065_854, w_065_855, w_065_856, w_065_857, w_065_858, w_065_860, w_065_862, w_065_864, w_065_866, w_065_867, w_065_870, w_065_875, w_065_876, w_065_877, w_065_878, w_065_879, w_065_880, w_065_883, w_065_884, w_065_886, w_065_887, w_065_889, w_065_893, w_065_894, w_065_896, w_065_898, w_065_899, w_065_900, w_065_901, w_065_903, w_065_904, w_065_905, w_065_907, w_065_911, w_065_912, w_065_916, w_065_917, w_065_922, w_065_925, w_065_926, w_065_927, w_065_928, w_065_932, w_065_935, w_065_936, w_065_941, w_065_943, w_065_949, w_065_950, w_065_952, w_065_955, w_065_958, w_065_959, w_065_960, w_065_962, w_065_963, w_065_964, w_065_965, w_065_966, w_065_968, w_065_970, w_065_971, w_065_972, w_065_974, w_065_975, w_065_976, w_065_978, w_065_984, w_065_988, w_065_989, w_065_990, w_065_992, w_065_997, w_065_998, w_065_999, w_065_1001, w_065_1004, w_065_1006, w_065_1007, w_065_1010, w_065_1011, w_065_1012, w_065_1013, w_065_1015, w_065_1016, w_065_1017, w_065_1018, w_065_1020, w_065_1021, w_065_1023, w_065_1024, w_065_1026, w_065_1029, w_065_1030, w_065_1032, w_065_1033, w_065_1036, w_065_1037, w_065_1038, w_065_1039, w_065_1040, w_065_1043, w_065_1044, w_065_1046, w_065_1047, w_065_1049, w_065_1050, w_065_1051, w_065_1052, w_065_1053, w_065_1055, w_065_1057, w_065_1059, w_065_1060, w_065_1061, w_065_1062, w_065_1063, w_065_1064, w_065_1066, w_065_1068, w_065_1069, w_065_1070, w_065_1071, w_065_1073, w_065_1074, w_065_1075, w_065_1076, w_065_1077, w_065_1078, w_065_1079, w_065_1081, w_065_1083, w_065_1085, w_065_1090, w_065_1093, w_065_1099, w_065_1100, w_065_1102, w_065_1103, w_065_1104, w_065_1114, w_065_1115, w_065_1117, w_065_1119, w_065_1120, w_065_1121, w_065_1122, w_065_1127, w_065_1129, w_065_1132, w_065_1136, w_065_1137, w_065_1139, w_065_1140, w_065_1141, w_065_1144, w_065_1145, w_065_1146, w_065_1147, w_065_1151, w_065_1153, w_065_1154, w_065_1155, w_065_1157, w_065_1158, w_065_1160, w_065_1161, w_065_1162, w_065_1163, w_065_1168, w_065_1170, w_065_1174, w_065_1175, w_065_1176, w_065_1177, w_065_1181, w_065_1182, w_065_1184, w_065_1186, w_065_1187, w_065_1188, w_065_1193, w_065_1201, w_065_1202, w_065_1203, w_065_1204, w_065_1205, w_065_1206, w_065_1208, w_065_1210, w_065_1212, w_065_1217, w_065_1218, w_065_1220, w_065_1222, w_065_1224, w_065_1226, w_065_1227, w_065_1228, w_065_1229, w_065_1230, w_065_1232, w_065_1233, w_065_1234, w_065_1235, w_065_1236, w_065_1237, w_065_1238, w_065_1239, w_065_1240, w_065_1241, w_065_1242, w_065_1243, w_065_1246, w_065_1247, w_065_1248, w_065_1249, w_065_1250, w_065_1252, w_065_1253, w_065_1254, w_065_1255, w_065_1256, w_065_1257, w_065_1258, w_065_1260, w_065_1261, w_065_1262, w_065_1263, w_065_1265, w_065_1266, w_065_1267, w_065_1268, w_065_1270, w_065_1271, w_065_1272, w_065_1275, w_065_1278, w_065_1280, w_065_1284, w_065_1285, w_065_1286, w_065_1288, w_065_1291, w_065_1292, w_065_1293, w_065_1294, w_065_1296, w_065_1297, w_065_1298, w_065_1301, w_065_1305, w_065_1306, w_065_1307, w_065_1309, w_065_1315, w_065_1319, w_065_1327, w_065_1329, w_065_1330, w_065_1331, w_065_1333, w_065_1334, w_065_1335, w_065_1336, w_065_1341, w_065_1343, w_065_1344, w_065_1345, w_065_1346, w_065_1347, w_065_1348, w_065_1349, w_065_1351, w_065_1354, w_065_1355, w_065_1356, w_065_1357, w_065_1358, w_065_1359, w_065_1362, w_065_1364, w_065_1365, w_065_1366, w_065_1367, w_065_1369, w_065_1371, w_065_1374, w_065_1376, w_065_1377, w_065_1378, w_065_1380, w_065_1382, w_065_1383, w_065_1385, w_065_1387, w_065_1388, w_065_1389, w_065_1390, w_065_1391, w_065_1392, w_065_1396, w_065_1398, w_065_1401, w_065_1402, w_065_1407, w_065_1409, w_065_1411, w_065_1412, w_065_1413, w_065_1414, w_065_1416, w_065_1418, w_065_1419, w_065_1420, w_065_1422, w_065_1424, w_065_1427, w_065_1430, w_065_1433, w_065_1435, w_065_1436, w_065_1439, w_065_1440, w_065_1443, w_065_1445, w_065_1446, w_065_1449, w_065_1453, w_065_1456, w_065_1459, w_065_1461, w_065_1462, w_065_1464, w_065_1465, w_065_1470, w_065_1472, w_065_1473, w_065_1476, w_065_1483, w_065_1484, w_065_1485, w_065_1487, w_065_1488, w_065_1491, w_065_1492, w_065_1495, w_065_1496, w_065_1497, w_065_1498, w_065_1499, w_065_1500, w_065_1501, w_065_1502, w_065_1503, w_065_1504, w_065_1505, w_065_1506, w_065_1507, w_065_1510, w_065_1512, w_065_1513, w_065_1516, w_065_1518, w_065_1519, w_065_1521, w_065_1522, w_065_1524, w_065_1525, w_065_1529, w_065_1534, w_065_1536, w_065_1537, w_065_1538, w_065_1541, w_065_1542, w_065_1544, w_065_1547, w_065_1549, w_065_1553, w_065_1554, w_065_1555, w_065_1556, w_065_1558, w_065_1560, w_065_1562, w_065_1563, w_065_1564, w_065_1568, w_065_1569, w_065_1570, w_065_1571, w_065_1573, w_065_1574, w_065_1575, w_065_1576, w_065_1577, w_065_1578, w_065_1579, w_065_1580, w_065_1581, w_065_1582, w_065_1584, w_065_1586, w_065_1587, w_065_1589, w_065_1591, w_065_1592, w_065_1594, w_065_1595, w_065_1596, w_065_1600, w_065_1602, w_065_1605, w_065_1606, w_065_1609, w_065_1610, w_065_1611, w_065_1612, w_065_1619, w_065_1620, w_065_1621, w_065_1622, w_065_1623, w_065_1624, w_065_1626, w_065_1627, w_065_1628, w_065_1629, w_065_1630, w_065_1632, w_065_1633, w_065_1635, w_065_1637, w_065_1638, w_065_1643, w_065_1648, w_065_1649, w_065_1650, w_065_1651, w_065_1652, w_065_1653, w_065_1654, w_065_1656, w_065_1657, w_065_1659, w_065_1660, w_065_1661, w_065_1662, w_065_1663, w_065_1665, w_065_1669, w_065_1670, w_065_1675, w_065_1677, w_065_1678, w_065_1679, w_065_1680, w_065_1682, w_065_1684, w_065_1685, w_065_1686, w_065_1687, w_065_1688, w_065_1691, w_065_1692, w_065_1693, w_065_1694, w_065_1695, w_065_1696, w_065_1697, w_065_1698, w_065_1700, w_065_1705, w_065_1707, w_065_1708, w_065_1710, w_065_1711, w_065_1712, w_065_1715, w_065_1716, w_065_1717, w_065_1718, w_065_1719, w_065_1722, w_065_1724, w_065_1731, w_065_1734, w_065_1736, w_065_1738, w_065_1740, w_065_1741, w_065_1742, w_065_1743, w_065_1744, w_065_1746, w_065_1750, w_065_1754, w_065_1755, w_065_1758, w_065_1759, w_065_1760, w_065_1761, w_065_1762, w_065_1764, w_065_1767, w_065_1768, w_065_1769, w_065_1770, w_065_1773, w_065_1774, w_065_1775, w_065_1776, w_065_1778, w_065_1781, w_065_1782, w_065_1784, w_065_1785, w_065_1789, w_065_1790, w_065_1792, w_065_1793, w_065_1798, w_065_1799, w_065_1800, w_065_1801, w_065_1803, w_065_1807, w_065_1808, w_065_1809, w_065_1811, w_065_1814, w_065_1819, w_065_1823, w_065_1824, w_065_1827, w_065_1828, w_065_1829, w_065_1831, w_065_1833, w_065_1834, w_065_1835, w_065_1837, w_065_1839, w_065_1840, w_065_1841, w_065_1842, w_065_1844, w_065_1845, w_065_1846, w_065_1848, w_065_1851, w_065_1852, w_065_1854, w_065_1857, w_065_1864, w_065_1865, w_065_1867, w_065_1869, w_065_1871, w_065_1873, w_065_1874, w_065_1875, w_065_1877, w_065_1878, w_065_1880, w_065_1881, w_065_1882, w_065_1884, w_065_1885, w_065_1887, w_065_1890, w_065_1891, w_065_1894, w_065_1896, w_065_1897, w_065_1900, w_065_1906, w_065_1907, w_065_1909, w_065_1912, w_065_1913, w_065_1914, w_065_1915, w_065_1918, w_065_1920, w_065_1921, w_065_1923, w_065_1925, w_065_1929, w_065_1930, w_065_1932, w_065_1937, w_065_1938, w_065_1939, w_065_1940, w_065_1941, w_065_1943, w_065_1945, w_065_1946, w_065_1948, w_065_1952, w_065_1953, w_065_1954, w_065_1955, w_065_1956, w_065_1957, w_065_1959, w_065_1960, w_065_1961, w_065_1968, w_065_1969, w_065_1970, w_065_1975, w_065_1978, w_065_1980, w_065_1981, w_065_1983, w_065_1987, w_065_1988, w_065_1990, w_065_1993, w_065_1994, w_065_1995, w_065_1996, w_065_1997, w_065_1998, w_065_2000, w_065_2003, w_065_2004, w_065_2005, w_065_2006, w_065_2007, w_065_2013, w_065_2014, w_065_2016, w_065_2018, w_065_2019, w_065_2020, w_065_2021, w_065_2022, w_065_2024, w_065_2026, w_065_2027, w_065_2030, w_065_2031, w_065_2033, w_065_2034, w_065_2035, w_065_2036, w_065_2038, w_065_2041, w_065_2042, w_065_2043, w_065_2044, w_065_2045, w_065_2046, w_065_2047, w_065_2048, w_065_2051, w_065_2053, w_065_2054, w_065_2055, w_065_2057, w_065_2059, w_065_2062, w_065_2064, w_065_2065, w_065_2068, w_065_2069, w_065_2072, w_065_2073, w_065_2075, w_065_2076, w_065_2077, w_065_2079, w_065_2080, w_065_2083, w_065_2085, w_065_2086, w_065_2087, w_065_2088, w_065_2089, w_065_2090, w_065_2091, w_065_2092, w_065_2095, w_065_2096, w_065_2098, w_065_2100, w_065_2102, w_065_2104, w_065_2105, w_065_2106, w_065_2110, w_065_2111, w_065_2112, w_065_2114, w_065_2115, w_065_2116, w_065_2118, w_065_2119, w_065_2120, w_065_2126, w_065_2129, w_065_2130, w_065_2132, w_065_2133, w_065_2136, w_065_2137, w_065_2138, w_065_2139, w_065_2140, w_065_2141, w_065_2143, w_065_2147, w_065_2149, w_065_2150, w_065_2151, w_065_2153, w_065_2155, w_065_2156, w_065_2157, w_065_2158, w_065_2160, w_065_2161, w_065_2162, w_065_2163, w_065_2164, w_065_2165, w_065_2166, w_065_2168, w_065_2169, w_065_2172, w_065_2173, w_065_2174, w_065_2176, w_065_2178, w_065_2179, w_065_2181, w_065_2185, w_065_2187, w_065_2188, w_065_2189, w_065_2191, w_065_2192, w_065_2194, w_065_2196, w_065_2197, w_065_2201, w_065_2204, w_065_2206, w_065_2213, w_065_2214, w_065_2215, w_065_2216, w_065_2217, w_065_2218, w_065_2219, w_065_2220, w_065_2221, w_065_2223, w_065_2224, w_065_2226, w_065_2227, w_065_2228, w_065_2229, w_065_2231, w_065_2237, w_065_2240, w_065_2241, w_065_2244, w_065_2246, w_065_2248, w_065_2252, w_065_2256, w_065_2259, w_065_2262, w_065_2263, w_065_2268, w_065_2269, w_065_2270, w_065_2274, w_065_2275, w_065_2276, w_065_2277, w_065_2278, w_065_2279, w_065_2281, w_065_2282, w_065_2285, w_065_2286, w_065_2288, w_065_2289, w_065_2290, w_065_2292, w_065_2293, w_065_2295, w_065_2296, w_065_2300, w_065_2301, w_065_2302, w_065_2309, w_065_2310, w_065_2311, w_065_2313, w_065_2314, w_065_2316, w_065_2317, w_065_2318, w_065_2320, w_065_2321, w_065_2322, w_065_2323, w_065_2325, w_065_2326, w_065_2329, w_065_2330, w_065_2333, w_065_2335, w_065_2337, w_065_2338, w_065_2339, w_065_2342, w_065_2344, w_065_2345, w_065_2347, w_065_2348, w_065_2349, w_065_2350, w_065_2351, w_065_2352, w_065_2354, w_065_2356, w_065_2358, w_065_2359, w_065_2360, w_065_2361, w_065_2363, w_065_2364, w_065_2365, w_065_2367, w_065_2368, w_065_2371, w_065_2372, w_065_2373, w_065_2374, w_065_2375, w_065_2376, w_065_2377, w_065_2380, w_065_2381, w_065_2382, w_065_2385, w_065_2387, w_065_2389, w_065_2390, w_065_2393, w_065_2395, w_065_2396, w_065_2398, w_065_2399, w_065_2403, w_065_2405, w_065_2408, w_065_2410, w_065_2411, w_065_2412, w_065_2415, w_065_2417, w_065_2418, w_065_2419, w_065_2420, w_065_2421, w_065_2423, w_065_2426, w_065_2431, w_065_2432, w_065_2433, w_065_2435, w_065_2436, w_065_2437, w_065_2439, w_065_2440, w_065_2443, w_065_2444, w_065_2445, w_065_2447, w_065_2450, w_065_2451, w_065_2452, w_065_2453, w_065_2454, w_065_2455, w_065_2456, w_065_2457, w_065_2458, w_065_2464, w_065_2465, w_065_2467, w_065_2468, w_065_2469, w_065_2470, w_065_2471, w_065_2474, w_065_2476, w_065_2478, w_065_2479, w_065_2480, w_065_2483, w_065_2484, w_065_2485, w_065_2488, w_065_2489, w_065_2490, w_065_2493, w_065_2494, w_065_2495, w_065_2496, w_065_2501, w_065_2502, w_065_2504, w_065_2505, w_065_2506, w_065_2508, w_065_2509, w_065_2510, w_065_2512, w_065_2514, w_065_2515, w_065_2518, w_065_2519, w_065_2520, w_065_2523, w_065_2524, w_065_2525, w_065_2526, w_065_2527, w_065_2529, w_065_2531, w_065_2532, w_065_2533, w_065_2534, w_065_2538, w_065_2539, w_065_2540, w_065_2542, w_065_2545, w_065_2546, w_065_2547, w_065_2548, w_065_2549, w_065_2550, w_065_2551, w_065_2552, w_065_2553, w_065_2555, w_065_2556, w_065_2557, w_065_2560, w_065_2563, w_065_2569, w_065_2570, w_065_2571, w_065_2572, w_065_2579, w_065_2580, w_065_2581, w_065_2584, w_065_2585, w_065_2588, w_065_2590, w_065_2594, w_065_2597, w_065_2598, w_065_2600, w_065_2601, w_065_2603, w_065_2604, w_065_2606, w_065_2607, w_065_2608, w_065_2610, w_065_2612, w_065_2613, w_065_2614, w_065_2615, w_065_2617, w_065_2619, w_065_2620, w_065_2621, w_065_2622, w_065_2625, w_065_2628, w_065_2630, w_065_2635, w_065_2637, w_065_2639, w_065_2640, w_065_2641, w_065_2643, w_065_2646, w_065_2647, w_065_2649, w_065_2650, w_065_2651, w_065_2653, w_065_2654, w_065_2655, w_065_2656, w_065_2658, w_065_2662, w_065_2663, w_065_2666, w_065_2667, w_065_2668, w_065_2669, w_065_2671, w_065_2673, w_065_2677, w_065_2678, w_065_2679, w_065_2680, w_065_2683, w_065_2684, w_065_2687, w_065_2689, w_065_2690, w_065_2693, w_065_2694, w_065_2695, w_065_2696, w_065_2700, w_065_2703, w_065_2706, w_065_2709, w_065_2711, w_065_2712, w_065_2715, w_065_2716, w_065_2718, w_065_2719, w_065_2720, w_065_2721, w_065_2722, w_065_2724, w_065_2727, w_065_2728, w_065_2729, w_065_2730, w_065_2733, w_065_2740, w_065_2742, w_065_2746, w_065_2748, w_065_2749, w_065_2750, w_065_2753, w_065_2754, w_065_2755, w_065_2757, w_065_2760, w_065_2765, w_065_2768, w_065_2771, w_065_2773, w_065_2775, w_065_2777, w_065_2779, w_065_2780, w_065_2781, w_065_2782, w_065_2785, w_065_2788, w_065_2789, w_065_2791, w_065_2792, w_065_2793, w_065_2794, w_065_2795, w_065_2796, w_065_2797, w_065_2798, w_065_2800, w_065_2802, w_065_2803, w_065_2804, w_065_2805, w_065_2807, w_065_2810, w_065_2811, w_065_2813, w_065_2816, w_065_2817, w_065_2819, w_065_2820, w_065_2821, w_065_2822, w_065_2825, w_065_2827, w_065_2829, w_065_2831, w_065_2833, w_065_2834, w_065_2836, w_065_2837, w_065_2838, w_065_2839, w_065_2841, w_065_2846, w_065_2847, w_065_2848, w_065_2849, w_065_2852, w_065_2853, w_065_2854, w_065_2856, w_065_2857, w_065_2858, w_065_2859, w_065_2861, w_065_2862, w_065_2864, w_065_2865, w_065_2867, w_065_2868, w_065_2872, w_065_2873, w_065_2878, w_065_2879, w_065_2880, w_065_2881, w_065_2883, w_065_2885, w_065_2886, w_065_2887, w_065_2888, w_065_2891, w_065_2892, w_065_2894, w_065_2896, w_065_2897, w_065_2898, w_065_2901, w_065_2903, w_065_2904, w_065_2905, w_065_2907, w_065_2909, w_065_2910, w_065_2912, w_065_2913, w_065_2916, w_065_2917, w_065_2919, w_065_2920, w_065_2921, w_065_2924, w_065_2925, w_065_2929, w_065_2933, w_065_2935, w_065_2937, w_065_2938, w_065_2940, w_065_2942, w_065_2944, w_065_2945, w_065_2946, w_065_2949, w_065_2950, w_065_2951, w_065_2953, w_065_2954, w_065_2956, w_065_2957, w_065_2958, w_065_2960, w_065_2961, w_065_2962, w_065_2966, w_065_2967, w_065_2970, w_065_2973, w_065_2974, w_065_2975, w_065_2976, w_065_2978, w_065_2980, w_065_2981, w_065_2984, w_065_2985, w_065_2986, w_065_2992, w_065_2993, w_065_2994, w_065_2995, w_065_2998, w_065_2999, w_065_3005, w_065_3006, w_065_3007, w_065_3008, w_065_3009, w_065_3010, w_065_3012, w_065_3014, w_065_3015, w_065_3016, w_065_3018, w_065_3022, w_065_3023, w_065_3025, w_065_3027, w_065_3029, w_065_3030, w_065_3031, w_065_3034, w_065_3035, w_065_3036, w_065_3038, w_065_3039, w_065_3040, w_065_3043, w_065_3044, w_065_3046, w_065_3048, w_065_3049, w_065_3051, w_065_3052, w_065_3053, w_065_3054, w_065_3055, w_065_3056, w_065_3057, w_065_3059, w_065_3060, w_065_3062, w_065_3068, w_065_3069, w_065_3070, w_065_3072, w_065_3073, w_065_3074, w_065_3075, w_065_3077, w_065_3078, w_065_3080, w_065_3081, w_065_3083, w_065_3086, w_065_3089, w_065_3092, w_065_3095, w_065_3098, w_065_3101, w_065_3104, w_065_3105, w_065_3107, w_065_3109, w_065_3110, w_065_3111, w_065_3113, w_065_3116, w_065_3118, w_065_3119, w_065_3120, w_065_3121, w_065_3122, w_065_3124, w_065_3126, w_065_3127, w_065_3128, w_065_3129, w_065_3132, w_065_3133, w_065_3134, w_065_3135, w_065_3136, w_065_3137, w_065_3139, w_065_3140, w_065_3141, w_065_3142, w_065_3143, w_065_3144, w_065_3145, w_065_3146, w_065_3147, w_065_3150, w_065_3153, w_065_3155, w_065_3157, w_065_3158, w_065_3159, w_065_3162, w_065_3164, w_065_3166, w_065_3167, w_065_3171, w_065_3172, w_065_3174, w_065_3176, w_065_3177, w_065_3178, w_065_3180, w_065_3182, w_065_3185, w_065_3186, w_065_3188, w_065_3189, w_065_3190, w_065_3193, w_065_3196, w_065_3200, w_065_3201, w_065_3204, w_065_3208, w_065_3209, w_065_3210, w_065_3211, w_065_3213, w_065_3216, w_065_3219, w_065_3221, w_065_3222, w_065_3223, w_065_3224, w_065_3227, w_065_3228, w_065_3229, w_065_3233, w_065_3234, w_065_3237, w_065_3238, w_065_3240, w_065_3243, w_065_3244, w_065_3245, w_065_3246, w_065_3247, w_065_3248, w_065_3249, w_065_3250, w_065_3251, w_065_3256, w_065_3257, w_065_3261, w_065_3263, w_065_3264, w_065_3265, w_065_3266, w_065_3269, w_065_3270, w_065_3271, w_065_3272, w_065_3274, w_065_3275, w_065_3278, w_065_3279, w_065_3282, w_065_3283, w_065_3287, w_065_3290, w_065_3291, w_065_3292, w_065_3295, w_065_3296, w_065_3297, w_065_3298, w_065_3299, w_065_3300, w_065_3301, w_065_3304, w_065_3305, w_065_3306, w_065_3308, w_065_3309, w_065_3310, w_065_3311, w_065_3312, w_065_3318, w_065_3319, w_065_3326, w_065_3328, w_065_3330, w_065_3331, w_065_3333, w_065_3334, w_065_3343, w_065_3346, w_065_3348, w_065_3351, w_065_3352, w_065_3353, w_065_3354, w_065_3356, w_065_3358, w_065_3360, w_065_3361, w_065_3362, w_065_3363, w_065_3365, w_065_3366, w_065_3373, w_065_3374, w_065_3375, w_065_3376, w_065_3377, w_065_3381, w_065_3382, w_065_3383, w_065_3384, w_065_3385, w_065_3386, w_065_3388, w_065_3390, w_065_3392, w_065_3394, w_065_3395, w_065_3396, w_065_3398, w_065_3399, w_065_3400, w_065_3402, w_065_3404, w_065_3405, w_065_3406, w_065_3407, w_065_3410, w_065_3414, w_065_3415, w_065_3417, w_065_3418, w_065_3420, w_065_3424, w_065_3426, w_065_3428, w_065_3429, w_065_3430, w_065_3432, w_065_3434, w_065_3435, w_065_3439, w_065_3440, w_065_3442, w_065_3443, w_065_3444, w_065_3445, w_065_3447, w_065_3448, w_065_3449, w_065_3452, w_065_3454, w_065_3457, w_065_3459, w_065_3463, w_065_3464, w_065_3465, w_065_3467, w_065_3468, w_065_3469, w_065_3470, w_065_3471, w_065_3472, w_065_3473, w_065_3474, w_065_3476, w_065_3478, w_065_3479, w_065_3481, w_065_3482, w_065_3483, w_065_3484, w_065_3485, w_065_3486, w_065_3487, w_065_3489, w_065_3490, w_065_3491, w_065_3492, w_065_3496, w_065_3497, w_065_3499, w_065_3505, w_065_3507, w_065_3508, w_065_3509, w_065_3510, w_065_3512, w_065_3516, w_065_3519, w_065_3527, w_065_3530, w_065_3531, w_065_3533, w_065_3535, w_065_3539, w_065_3541, w_065_3545, w_065_3548, w_065_3551, w_065_3553, w_065_3558, w_065_3559, w_065_3564, w_065_3578, w_065_3584, w_065_3585, w_065_3589, w_065_3594, w_065_3601, w_065_3603, w_065_3604, w_065_3606, w_065_3608, w_065_3609, w_065_3614, w_065_3616, w_065_3617, w_065_3625, w_065_3627, w_065_3628, w_065_3630, w_065_3633, w_065_3636, w_065_3638, w_065_3639, w_065_3642, w_065_3643, w_065_3644, w_065_3645, w_065_3646, w_065_3650, w_065_3652, w_065_3655, w_065_3657, w_065_3658, w_065_3666, w_065_3669, w_065_3676, w_065_3677, w_065_3679, w_065_3680, w_065_3681, w_065_3682, w_065_3686, w_065_3689, w_065_3691, w_065_3693, w_065_3694, w_065_3695, w_065_3696, w_065_3697, w_065_3698, w_065_3699, w_065_3700, w_065_3701, w_065_3706, w_065_3707, w_065_3708, w_065_3709, w_065_3712, w_065_3713, w_065_3723, w_065_3724, w_065_3726, w_065_3727, w_065_3729, w_065_3730, w_065_3731, w_065_3732, w_065_3737, w_065_3738, w_065_3739, w_065_3742, w_065_3743, w_065_3748, w_065_3749, w_065_3751, w_065_3755, w_065_3759, w_065_3762, w_065_3764, w_065_3765, w_065_3766, w_065_3769, w_065_3770, w_065_3775, w_065_3777, w_065_3780, w_065_3781, w_065_3788, w_065_3791, w_065_3793, w_065_3794, w_065_3796, w_065_3799, w_065_3800, w_065_3801, w_065_3806, w_065_3808, w_065_3809, w_065_3812, w_065_3819, w_065_3822, w_065_3833, w_065_3835, w_065_3836, w_065_3841, w_065_3844, w_065_3850, w_065_3853, w_065_3856, w_065_3860, w_065_3863, w_065_3867, w_065_3870, w_065_3878, w_065_3879, w_065_3880, w_065_3886, w_065_3888, w_065_3889, w_065_3891, w_065_3893, w_065_3894, w_065_3898, w_065_3902, w_065_3907, w_065_3912, w_065_3918, w_065_3919, w_065_3921, w_065_3923, w_065_3926, w_065_3927, w_065_3931, w_065_3933, w_065_3934, w_065_3935, w_065_3940, w_065_3941, w_065_3947, w_065_3948, w_065_3949, w_065_3950, w_065_3954, w_065_3959, w_065_3960, w_065_3963, w_065_3964, w_065_3965, w_065_3967, w_065_3971, w_065_3977, w_065_3978, w_065_3983, w_065_3985, w_065_3987, w_065_3990, w_065_3992, w_065_3993, w_065_3995, w_065_3999, w_065_4001, w_065_4015, w_065_4016, w_065_4017, w_065_4019, w_065_4021, w_065_4028, w_065_4031, w_065_4032, w_065_4034, w_065_4035, w_065_4037, w_065_4044, w_065_4046, w_065_4054, w_065_4055, w_065_4056, w_065_4061, w_065_4062, w_065_4068, w_065_4069, w_065_4072, w_065_4076, w_065_4078, w_065_4079, w_065_4081, w_065_4083, w_065_4085, w_065_4086, w_065_4087, w_065_4090, w_065_4093, w_065_4097, w_065_4100, w_065_4102, w_065_4106, w_065_4108, w_065_4111, w_065_4112, w_065_4113, w_065_4115, w_065_4116, w_065_4118, w_065_4130, w_065_4131, w_065_4133, w_065_4139, w_065_4140, w_065_4146, w_065_4148, w_065_4152, w_065_4155, w_065_4159, w_065_4160, w_065_4162, w_065_4172, w_065_4173, w_065_4177, w_065_4178, w_065_4179, w_065_4181, w_065_4184, w_065_4202, w_065_4204, w_065_4205, w_065_4207, w_065_4214, w_065_4216, w_065_4218, w_065_4224, w_065_4229, w_065_4231, w_065_4232, w_065_4233, w_065_4234, w_065_4249, w_065_4252, w_065_4257, w_065_4259, w_065_4267, w_065_4269, w_065_4271, w_065_4272, w_065_4275, w_065_4276, w_065_4277, w_065_4279, w_065_4282, w_065_4283, w_065_4287, w_065_4293, w_065_4294, w_065_4296, w_065_4297, w_065_4298, w_065_4301, w_065_4304, w_065_4305, w_065_4308, w_065_4309, w_065_4314, w_065_4315, w_065_4320, w_065_4326, w_065_4327, w_065_4329, w_065_4334, w_065_4337, w_065_4340, w_065_4342, w_065_4344, w_065_4347, w_065_4350, w_065_4353, w_065_4354, w_065_4358, w_065_4359, w_065_4362, w_065_4363, w_065_4368, w_065_4369, w_065_4370, w_065_4378, w_065_4379, w_065_4399, w_065_4402, w_065_4403, w_065_4405, w_065_4406, w_065_4408, w_065_4409, w_065_4410, w_065_4411, w_065_4412, w_065_4413, w_065_4416, w_065_4419, w_065_4420, w_065_4423, w_065_4425, w_065_4435, w_065_4437, w_065_4438, w_065_4450, w_065_4451, w_065_4456, w_065_4458, w_065_4461, w_065_4463, w_065_4466, w_065_4471, w_065_4472, w_065_4473, w_065_4474, w_065_4480, w_065_4487, w_065_4488, w_065_4489, w_065_4500, w_065_4502, w_065_4509, w_065_4514, w_065_4517, w_065_4518, w_065_4521, w_065_4522, w_065_4523, w_065_4526, w_065_4536, w_065_4537, w_065_4539, w_065_4540, w_065_4542, w_065_4550, w_065_4558, w_065_4560, w_065_4562, w_065_4565, w_065_4567, w_065_4569, w_065_4571, w_065_4573, w_065_4574, w_065_4576, w_065_4580, w_065_4584, w_065_4585, w_065_4587, w_065_4595, w_065_4596, w_065_4598, w_065_4602, w_065_4604, w_065_4605, w_065_4611, w_065_4612, w_065_4614, w_065_4616, w_065_4618, w_065_4619, w_065_4620, w_065_4623, w_065_4624, w_065_4625, w_065_4626, w_065_4627, w_065_4628, w_065_4633, w_065_4635, w_065_4636, w_065_4638, w_065_4643, w_065_4644, w_065_4648, w_065_4649, w_065_4650, w_065_4654, w_065_4664, w_065_4665, w_065_4668, w_065_4669, w_065_4674, w_065_4675, w_065_4683, w_065_4687, w_065_4691, w_065_4696, w_065_4697, w_065_4698, w_065_4701, w_065_4702, w_065_4704, w_065_4705, w_065_4707, w_065_4715, w_065_4716, w_065_4717, w_065_4718, w_065_4719, w_065_4725, w_065_4726, w_065_4730, w_065_4733, w_065_4734, w_065_4736, w_065_4739, w_065_4741, w_065_4742, w_065_4746, w_065_4747, w_065_4751, w_065_4752, w_065_4754, w_065_4761, w_065_4763, w_065_4764, w_065_4767, w_065_4768, w_065_4777, w_065_4778, w_065_4779, w_065_4785, w_065_4793, w_065_4795, w_065_4799, w_065_4803, w_065_4811, w_065_4817, w_065_4818, w_065_4819, w_065_4820, w_065_4838, w_065_4839, w_065_4843, w_065_4845, w_065_4846, w_065_4847, w_065_4849, w_065_4851, w_065_4853, w_065_4859, w_065_4862, w_065_4863, w_065_4865, w_065_4866, w_065_4868, w_065_4869, w_065_4873, w_065_4874, w_065_4875, w_065_4880, w_065_4882, w_065_4883, w_065_4885, w_065_4886, w_065_4891, w_065_4900, w_065_4905, w_065_4910, w_065_4912, w_065_4922, w_065_4923, w_065_4935, w_065_4940, w_065_4941, w_065_4942, w_065_4943, w_065_4944, w_065_4946, w_065_4951, w_065_4952, w_065_4953, w_065_4955, w_065_4959, w_065_4967, w_065_4968, w_065_4969, w_065_4972, w_065_4974, w_065_4975, w_065_4982, w_065_4984, w_065_4985, w_065_4987, w_065_4988, w_065_4991, w_065_4992, w_065_4995, w_065_4996, w_065_5000, w_065_5002, w_065_5003, w_065_5008, w_065_5013, w_065_5015, w_065_5019, w_065_5020, w_065_5021, w_065_5028, w_065_5031, w_065_5034, w_065_5035, w_065_5037, w_065_5038, w_065_5041, w_065_5042, w_065_5050, w_065_5055, w_065_5057, w_065_5063, w_065_5064, w_065_5067, w_065_5069, w_065_5097, w_065_5101, w_065_5102, w_065_5107, w_065_5112, w_065_5117, w_065_5119, w_065_5120, w_065_5121, w_065_5124, w_065_5128, w_065_5134, w_065_5136, w_065_5137, w_065_5138, w_065_5140, w_065_5145, w_065_5147, w_065_5148, w_065_5149, w_065_5151, w_065_5153, w_065_5158, w_065_5163, w_065_5167, w_065_5169, w_065_5172, w_065_5174, w_065_5175, w_065_5182, w_065_5183, w_065_5186, w_065_5189, w_065_5191, w_065_5192, w_065_5193, w_065_5194, w_065_5204, w_065_5208, w_065_5209, w_065_5210, w_065_5211, w_065_5213, w_065_5215, w_065_5221, w_065_5222, w_065_5223, w_065_5225, w_065_5234, w_065_5235, w_065_5240, w_065_5241, w_065_5242, w_065_5243, w_065_5246, w_065_5249, w_065_5254, w_065_5256, w_065_5257, w_065_5262, w_065_5265, w_065_5270, w_065_5272, w_065_5274, w_065_5276, w_065_5281, w_065_5282, w_065_5283, w_065_5292, w_065_5297, w_065_5299, w_065_5305, w_065_5308, w_065_5309, w_065_5310, w_065_5311, w_065_5316, w_065_5317, w_065_5319, w_065_5320, w_065_5321, w_065_5324, w_065_5332, w_065_5333, w_065_5337, w_065_5338, w_065_5339, w_065_5342, w_065_5344, w_065_5346, w_065_5351, w_065_5358, w_065_5361, w_065_5362, w_065_5365, w_065_5368, w_065_5370, w_065_5372, w_065_5377, w_065_5378, w_065_5379, w_065_5380, w_065_5383, w_065_5385, w_065_5386, w_065_5387, w_065_5388, w_065_5389, w_065_5397, w_065_5398, w_065_5399, w_065_5400, w_065_5401, w_065_5405, w_065_5407, w_065_5412, w_065_5413, w_065_5419, w_065_5421, w_065_5423, w_065_5429, w_065_5434, w_065_5436, w_065_5438, w_065_5439, w_065_5443, w_065_5445, w_065_5448, w_065_5451, w_065_5454, w_065_5459, w_065_5461, w_065_5462, w_065_5465, w_065_5466, w_065_5467, w_065_5470, w_065_5472, w_065_5476, w_065_5478, w_065_5479, w_065_5480, w_065_5486, w_065_5489, w_065_5490, w_065_5493, w_065_5496, w_065_5498, w_065_5500, w_065_5502, w_065_5508, w_065_5510, w_065_5515, w_065_5517, w_065_5519, w_065_5520, w_065_5522, w_065_5526, w_065_5534, w_065_5535, w_065_5539, w_065_5540, w_065_5542, w_065_5544, w_065_5546, w_065_5548, w_065_5549, w_065_5554, w_065_5557, w_065_5559, w_065_5565, w_065_5573, w_065_5574, w_065_5575, w_065_5576, w_065_5578, w_065_5584, w_065_5589, w_065_5594, w_065_5595, w_065_5598, w_065_5599, w_065_5600, w_065_5602, w_065_5607, w_065_5609, w_065_5611, w_065_5613, w_065_5614, w_065_5616, w_065_5618, w_065_5619, w_065_5622, w_065_5623, w_065_5625, w_065_5628, w_065_5629, w_065_5635, w_065_5636, w_065_5638, w_065_5640, w_065_5642, w_065_5644, w_065_5648, w_065_5650, w_065_5656, w_065_5665, w_065_5669, w_065_5673, w_065_5677, w_065_5679, w_065_5680, w_065_5686, w_065_5689, w_065_5690, w_065_5691, w_065_5692, w_065_5696, w_065_5697, w_065_5699, w_065_5700, w_065_5703, w_065_5708, w_065_5714, w_065_5718, w_065_5726, w_065_5736, w_065_5737, w_065_5741, w_065_5742, w_065_5743, w_065_5744, w_065_5745, w_065_5747, w_065_5750, w_065_5751, w_065_5758, w_065_5760, w_065_5761, w_065_5762, w_065_5764, w_065_5768, w_065_5778, w_065_5779, w_065_5783, w_065_5785, w_065_5790, w_065_5792, w_065_5796, w_065_5798, w_065_5803, w_065_5805, w_065_5808, w_065_5809, w_065_5810, w_065_5814, w_065_5820, w_065_5822, w_065_5824, w_065_5828, w_065_5832, w_065_5834, w_065_5836, w_065_5837, w_065_5839, w_065_5841, w_065_5845, w_065_5846, w_065_5850, w_065_5855, w_065_5857, w_065_5860, w_065_5871, w_065_5879, w_065_5882, w_065_5883, w_065_5893, w_065_5895, w_065_5896, w_065_5897, w_065_5898, w_065_5903, w_065_5904, w_065_5906, w_065_5910, w_065_5923, w_065_5926, w_065_5927, w_065_5934, w_065_5936, w_065_5938, w_065_5944, w_065_5947, w_065_5950, w_065_5952, w_065_5953, w_065_5956, w_065_5957, w_065_5960, w_065_5962, w_065_5964, w_065_5966, w_065_5975, w_065_5976, w_065_5978, w_065_5982, w_065_5994, w_065_5995, w_065_5999, w_065_6000, w_065_6002, w_065_6005, w_065_6006, w_065_6007, w_065_6013, w_065_6016, w_065_6018, w_065_6019, w_065_6022, w_065_6023, w_065_6024, w_065_6027, w_065_6030, w_065_6033, w_065_6034, w_065_6035, w_065_6036, w_065_6040, w_065_6044, w_065_6047, w_065_6049, w_065_6051, w_065_6052, w_065_6057, w_065_6061, w_065_6063, w_065_6070, w_065_6073, w_065_6077, w_065_6085, w_065_6087, w_065_6088, w_065_6089, w_065_6097, w_065_6099, w_065_6105, w_065_6111, w_065_6112, w_065_6115, w_065_6121, w_065_6123, w_065_6131, w_065_6133, w_065_6134, w_065_6135, w_065_6136, w_065_6142, w_065_6145, w_065_6151, w_065_6157, w_065_6160, w_065_6165, w_065_6166, w_065_6169, w_065_6172, w_065_6177, w_065_6178, w_065_6182, w_065_6183, w_065_6184, w_065_6185, w_065_6187, w_065_6188, w_065_6190, w_065_6191, w_065_6197, w_065_6198, w_065_6200, w_065_6207, w_065_6209, w_065_6210, w_065_6211, w_065_6212, w_065_6219, w_065_6221, w_065_6224, w_065_6225, w_065_6229, w_065_6230, w_065_6234, w_065_6240, w_065_6241, w_065_6243, w_065_6247, w_065_6253, w_065_6256, w_065_6259, w_065_6260, w_065_6268, w_065_6274, w_065_6275, w_065_6278, w_065_6283, w_065_6286, w_065_6288, w_065_6293, w_065_6303, w_065_6314, w_065_6317, w_065_6318, w_065_6319, w_065_6320, w_065_6325, w_065_6329, w_065_6331, w_065_6333, w_065_6335, w_065_6341, w_065_6346, w_065_6353, w_065_6358, w_065_6359, w_065_6363, w_065_6365, w_065_6368, w_065_6370, w_065_6383, w_065_6385, w_065_6389, w_065_6390, w_065_6391, w_065_6396, w_065_6399, w_065_6400, w_065_6403, w_065_6405, w_065_6407, w_065_6408, w_065_6409, w_065_6410, w_065_6414, w_065_6415, w_065_6420, w_065_6422, w_065_6430, w_065_6433, w_065_6436, w_065_6445, w_065_6447, w_065_6452, w_065_6455, w_065_6457, w_065_6462, w_065_6466, w_065_6467, w_065_6468, w_065_6469, w_065_6473, w_065_6475, w_065_6478, w_065_6485, w_065_6486;
  wire w_066_000, w_066_002, w_066_005, w_066_006, w_066_007, w_066_010, w_066_011, w_066_012, w_066_013, w_066_014, w_066_015, w_066_016, w_066_018, w_066_019, w_066_020, w_066_021, w_066_022, w_066_024, w_066_027, w_066_028, w_066_029, w_066_031, w_066_032, w_066_035, w_066_036, w_066_037, w_066_038, w_066_039, w_066_042, w_066_044, w_066_045, w_066_046, w_066_047, w_066_051, w_066_052, w_066_053, w_066_054, w_066_055, w_066_056, w_066_057, w_066_058, w_066_059, w_066_061, w_066_062, w_066_063, w_066_065, w_066_067, w_066_069, w_066_071, w_066_072, w_066_073, w_066_075, w_066_076, w_066_077, w_066_078, w_066_081, w_066_082, w_066_083, w_066_085, w_066_086, w_066_088, w_066_090, w_066_091, w_066_093, w_066_094, w_066_095, w_066_097, w_066_098, w_066_099, w_066_100, w_066_101, w_066_103, w_066_104, w_066_105, w_066_106, w_066_107, w_066_108, w_066_109, w_066_110, w_066_111, w_066_113, w_066_114, w_066_117, w_066_118, w_066_119, w_066_120, w_066_123, w_066_124, w_066_126, w_066_127, w_066_128, w_066_129, w_066_130, w_066_131, w_066_133, w_066_134, w_066_135, w_066_137, w_066_138, w_066_139, w_066_140, w_066_143, w_066_145, w_066_146, w_066_147, w_066_148, w_066_149, w_066_150, w_066_151, w_066_152, w_066_155, w_066_156, w_066_157, w_066_158, w_066_160, w_066_161, w_066_162, w_066_163, w_066_164, w_066_165, w_066_166, w_066_167, w_066_168, w_066_170, w_066_171, w_066_172, w_066_173, w_066_176, w_066_177, w_066_178, w_066_179, w_066_181, w_066_183, w_066_184, w_066_185, w_066_186, w_066_187, w_066_191, w_066_193, w_066_195, w_066_197, w_066_198, w_066_199, w_066_200, w_066_202, w_066_203, w_066_204, w_066_205, w_066_207, w_066_208, w_066_210, w_066_212, w_066_216, w_066_217, w_066_218, w_066_219, w_066_221, w_066_222, w_066_223, w_066_224, w_066_225, w_066_226, w_066_227, w_066_228, w_066_229, w_066_231, w_066_233, w_066_235, w_066_236, w_066_237, w_066_238, w_066_240, w_066_241, w_066_243, w_066_244, w_066_245, w_066_248, w_066_249, w_066_250, w_066_251, w_066_252, w_066_253, w_066_254, w_066_256, w_066_258, w_066_259, w_066_260, w_066_261, w_066_262, w_066_263, w_066_265, w_066_266, w_066_267, w_066_269, w_066_273, w_066_274, w_066_275, w_066_276, w_066_278, w_066_279, w_066_280, w_066_281, w_066_282, w_066_283, w_066_284, w_066_285, w_066_286, w_066_287, w_066_288, w_066_289, w_066_291, w_066_292, w_066_293, w_066_296, w_066_298, w_066_299, w_066_300, w_066_301, w_066_302, w_066_303, w_066_304, w_066_308, w_066_314, w_066_315, w_066_318, w_066_322, w_066_323, w_066_324, w_066_325, w_066_326, w_066_327, w_066_329, w_066_330, w_066_331, w_066_333, w_066_334, w_066_335, w_066_336, w_066_338, w_066_339, w_066_340, w_066_344, w_066_345, w_066_347, w_066_348, w_066_349, w_066_350, w_066_353, w_066_354, w_066_355, w_066_356, w_066_357, w_066_358, w_066_359, w_066_360, w_066_361, w_066_365, w_066_366, w_066_369, w_066_370, w_066_373, w_066_374, w_066_375, w_066_376, w_066_377, w_066_378, w_066_379, w_066_380, w_066_381, w_066_383, w_066_384, w_066_386, w_066_391, w_066_395, w_066_396, w_066_397, w_066_398, w_066_399, w_066_400, w_066_402, w_066_403, w_066_406, w_066_407, w_066_408, w_066_409, w_066_411, w_066_412, w_066_413, w_066_417, w_066_418, w_066_421, w_066_422, w_066_423, w_066_425, w_066_426, w_066_427, w_066_428, w_066_430, w_066_432, w_066_433, w_066_434, w_066_436, w_066_437, w_066_439, w_066_440, w_066_441, w_066_443, w_066_444, w_066_445, w_066_446, w_066_447, w_066_448, w_066_450, w_066_453, w_066_455, w_066_456, w_066_457, w_066_459, w_066_460, w_066_462, w_066_464, w_066_465, w_066_466, w_066_467, w_066_469, w_066_470, w_066_471, w_066_472, w_066_473, w_066_474, w_066_475, w_066_477, w_066_478, w_066_479, w_066_480, w_066_481, w_066_482, w_066_483, w_066_484, w_066_487, w_066_490, w_066_491, w_066_492, w_066_493, w_066_495, w_066_496, w_066_498, w_066_499, w_066_500, w_066_502, w_066_504, w_066_505, w_066_506, w_066_507, w_066_508, w_066_509, w_066_511, w_066_512, w_066_513, w_066_514, w_066_515, w_066_516, w_066_517, w_066_518, w_066_519, w_066_520, w_066_521, w_066_523, w_066_524, w_066_525, w_066_526, w_066_527, w_066_529, w_066_531, w_066_532, w_066_538, w_066_539, w_066_540, w_066_541, w_066_543, w_066_545, w_066_547, w_066_548, w_066_549, w_066_550, w_066_553, w_066_556, w_066_557, w_066_563, w_066_565, w_066_566, w_066_569, w_066_571, w_066_572, w_066_573, w_066_574, w_066_575, w_066_576, w_066_577, w_066_578, w_066_579, w_066_580, w_066_581, w_066_582, w_066_583, w_066_584, w_066_585, w_066_586, w_066_587, w_066_589, w_066_590, w_066_591, w_066_593, w_066_594, w_066_595, w_066_596, w_066_597, w_066_598, w_066_601, w_066_602, w_066_603, w_066_604, w_066_605, w_066_606, w_066_607, w_066_608, w_066_609, w_066_610, w_066_612, w_066_615, w_066_616, w_066_618, w_066_619, w_066_620, w_066_621, w_066_622, w_066_623, w_066_625, w_066_627, w_066_628, w_066_629, w_066_630, w_066_632, w_066_633, w_066_634, w_066_635, w_066_637, w_066_638, w_066_639, w_066_640, w_066_641, w_066_642, w_066_643, w_066_646, w_066_647, w_066_648, w_066_650, w_066_651, w_066_652, w_066_653, w_066_655, w_066_656, w_066_657, w_066_658, w_066_659, w_066_661, w_066_663, w_066_664, w_066_665, w_066_667, w_066_668, w_066_669, w_066_670, w_066_671, w_066_672, w_066_673, w_066_674, w_066_675, w_066_678, w_066_679, w_066_680, w_066_685, w_066_686, w_066_687, w_066_688, w_066_690, w_066_691, w_066_692, w_066_694, w_066_695, w_066_697, w_066_698, w_066_703, w_066_706, w_066_707, w_066_708, w_066_709, w_066_710, w_066_712, w_066_713, w_066_714, w_066_715, w_066_716, w_066_717, w_066_719, w_066_726, w_066_727, w_066_728, w_066_729, w_066_730, w_066_731, w_066_733, w_066_734, w_066_736, w_066_738, w_066_739, w_066_740, w_066_741, w_066_743, w_066_744, w_066_745, w_066_748, w_066_750, w_066_751, w_066_752, w_066_753, w_066_754, w_066_755, w_066_756, w_066_757, w_066_758, w_066_760, w_066_762, w_066_763, w_066_764, w_066_765, w_066_767, w_066_768, w_066_771, w_066_772, w_066_773, w_066_774, w_066_775, w_066_777, w_066_778, w_066_779, w_066_780, w_066_781, w_066_783, w_066_784, w_066_785, w_066_786, w_066_788, w_066_789, w_066_790, w_066_791, w_066_792, w_066_793, w_066_795, w_066_797, w_066_800, w_066_801, w_066_802, w_066_803, w_066_805, w_066_806, w_066_809, w_066_810, w_066_812, w_066_815, w_066_816, w_066_817, w_066_818, w_066_820, w_066_821, w_066_822, w_066_823, w_066_825, w_066_826, w_066_827, w_066_828, w_066_830, w_066_831, w_066_833, w_066_834, w_066_835, w_066_836, w_066_837, w_066_838, w_066_840, w_066_841, w_066_842, w_066_844, w_066_846, w_066_847, w_066_848, w_066_849, w_066_851, w_066_853, w_066_858, w_066_859, w_066_860, w_066_862, w_066_863, w_066_864, w_066_866, w_066_867, w_066_869, w_066_870, w_066_871, w_066_872, w_066_874, w_066_875, w_066_879, w_066_880, w_066_882, w_066_884, w_066_885, w_066_889, w_066_890, w_066_891, w_066_893, w_066_895, w_066_897, w_066_899, w_066_901, w_066_902, w_066_905, w_066_907, w_066_908, w_066_909, w_066_911, w_066_914, w_066_915, w_066_916, w_066_918, w_066_919, w_066_920, w_066_922, w_066_923, w_066_925, w_066_926, w_066_927, w_066_928, w_066_929, w_066_930, w_066_932, w_066_933, w_066_934, w_066_935, w_066_937, w_066_938, w_066_939, w_066_940, w_066_943, w_066_944, w_066_946, w_066_947, w_066_949, w_066_951, w_066_953, w_066_954, w_066_957, w_066_959, w_066_960, w_066_961, w_066_962, w_066_963, w_066_964, w_066_965, w_066_966, w_066_968, w_066_969, w_066_970, w_066_971, w_066_972, w_066_973, w_066_974, w_066_976, w_066_977, w_066_978, w_066_980, w_066_981, w_066_983, w_066_984, w_066_985, w_066_986, w_066_990, w_066_993, w_066_994, w_066_995, w_066_996, w_066_997, w_066_998, w_066_999, w_066_1001, w_066_1002, w_066_1003, w_066_1004, w_066_1005, w_066_1006, w_066_1007, w_066_1008, w_066_1009, w_066_1010, w_066_1012, w_066_1013, w_066_1014, w_066_1015, w_066_1016, w_066_1018, w_066_1020, w_066_1021, w_066_1023, w_066_1024, w_066_1025, w_066_1027, w_066_1028, w_066_1029, w_066_1030, w_066_1035, w_066_1036, w_066_1037, w_066_1038, w_066_1039, w_066_1041, w_066_1045, w_066_1046, w_066_1048, w_066_1049, w_066_1050, w_066_1051, w_066_1052, w_066_1054, w_066_1055, w_066_1056, w_066_1057, w_066_1060, w_066_1061, w_066_1063, w_066_1064, w_066_1065, w_066_1070, w_066_1073, w_066_1074, w_066_1076, w_066_1077, w_066_1078, w_066_1079, w_066_1080, w_066_1081, w_066_1082, w_066_1083, w_066_1085, w_066_1087, w_066_1088, w_066_1089, w_066_1090, w_066_1093, w_066_1094, w_066_1095, w_066_1096, w_066_1097, w_066_1099, w_066_1102, w_066_1104, w_066_1105, w_066_1106, w_066_1107, w_066_1109, w_066_1110, w_066_1111, w_066_1112, w_066_1115, w_066_1116, w_066_1117, w_066_1118, w_066_1119, w_066_1121, w_066_1122, w_066_1128, w_066_1129, w_066_1131, w_066_1132, w_066_1133, w_066_1134, w_066_1138, w_066_1139, w_066_1140, w_066_1141, w_066_1142, w_066_1143, w_066_1144, w_066_1145, w_066_1146, w_066_1148, w_066_1149, w_066_1150, w_066_1151, w_066_1152, w_066_1153, w_066_1154, w_066_1155, w_066_1156, w_066_1157, w_066_1158, w_066_1159, w_066_1161, w_066_1163, w_066_1165, w_066_1166, w_066_1168, w_066_1169, w_066_1170, w_066_1171, w_066_1172, w_066_1173, w_066_1174, w_066_1175, w_066_1176, w_066_1177, w_066_1178, w_066_1180, w_066_1181, w_066_1182, w_066_1183, w_066_1184, w_066_1185, w_066_1187, w_066_1188, w_066_1189, w_066_1191, w_066_1192, w_066_1193, w_066_1194, w_066_1197, w_066_1200, w_066_1203, w_066_1206, w_066_1207, w_066_1208, w_066_1209, w_066_1213, w_066_1214, w_066_1215, w_066_1216, w_066_1218, w_066_1219, w_066_1221, w_066_1223, w_066_1225, w_066_1226, w_066_1227, w_066_1228, w_066_1230, w_066_1231, w_066_1232, w_066_1233, w_066_1235, w_066_1239, w_066_1240, w_066_1241, w_066_1242, w_066_1243, w_066_1245, w_066_1249, w_066_1251, w_066_1253, w_066_1254, w_066_1256, w_066_1257, w_066_1259, w_066_1260, w_066_1261, w_066_1264, w_066_1265, w_066_1267, w_066_1268, w_066_1272, w_066_1276, w_066_1279, w_066_1282, w_066_1284, w_066_1286, w_066_1287, w_066_1288, w_066_1289, w_066_1291, w_066_1293, w_066_1294, w_066_1295, w_066_1297, w_066_1298, w_066_1299, w_066_1300, w_066_1302, w_066_1303, w_066_1304, w_066_1307, w_066_1308, w_066_1309, w_066_1311, w_066_1312, w_066_1313, w_066_1314, w_066_1316, w_066_1317, w_066_1319, w_066_1321, w_066_1324, w_066_1325, w_066_1326, w_066_1327, w_066_1328, w_066_1330, w_066_1332, w_066_1333, w_066_1335, w_066_1336, w_066_1341, w_066_1342, w_066_1345, w_066_1347, w_066_1348, w_066_1349, w_066_1350, w_066_1351, w_066_1353, w_066_1354, w_066_1357, w_066_1358, w_066_1360, w_066_1362, w_066_1364, w_066_1365, w_066_1369, w_066_1370, w_066_1371, w_066_1372, w_066_1373, w_066_1374, w_066_1377, w_066_1379, w_066_1381, w_066_1382, w_066_1385, w_066_1386, w_066_1390, w_066_1391, w_066_1393, w_066_1394, w_066_1398, w_066_1400, w_066_1402, w_066_1407, w_066_1408, w_066_1411, w_066_1412, w_066_1415, w_066_1417, w_066_1418, w_066_1420, w_066_1422, w_066_1423, w_066_1427, w_066_1429, w_066_1431, w_066_1432, w_066_1433, w_066_1434, w_066_1435, w_066_1437, w_066_1438, w_066_1439, w_066_1443, w_066_1444, w_066_1449, w_066_1451, w_066_1455, w_066_1456, w_066_1457, w_066_1460, w_066_1465, w_066_1468, w_066_1470, w_066_1474, w_066_1475, w_066_1476, w_066_1478, w_066_1479, w_066_1480, w_066_1482, w_066_1483, w_066_1484, w_066_1487, w_066_1488, w_066_1489, w_066_1492, w_066_1493, w_066_1495, w_066_1496, w_066_1497, w_066_1498, w_066_1500, w_066_1501, w_066_1504, w_066_1505, w_066_1506, w_066_1507, w_066_1508, w_066_1510, w_066_1511, w_066_1517, w_066_1518, w_066_1519, w_066_1520, w_066_1524, w_066_1525, w_066_1527, w_066_1528, w_066_1529, w_066_1531, w_066_1532, w_066_1534, w_066_1536, w_066_1538, w_066_1539, w_066_1540, w_066_1542, w_066_1543, w_066_1544, w_066_1545, w_066_1547, w_066_1548, w_066_1549, w_066_1552, w_066_1555, w_066_1556, w_066_1558, w_066_1559, w_066_1560, w_066_1561, w_066_1567, w_066_1570, w_066_1571, w_066_1573, w_066_1576, w_066_1578, w_066_1579, w_066_1580, w_066_1582, w_066_1583, w_066_1589, w_066_1592, w_066_1593, w_066_1594, w_066_1595, w_066_1596, w_066_1597, w_066_1598, w_066_1600, w_066_1601, w_066_1602, w_066_1603, w_066_1604, w_066_1605, w_066_1609, w_066_1611, w_066_1612, w_066_1616, w_066_1618, w_066_1619, w_066_1620, w_066_1625, w_066_1626, w_066_1627, w_066_1630, w_066_1632, w_066_1633, w_066_1635, w_066_1636, w_066_1637, w_066_1638, w_066_1639, w_066_1640, w_066_1645, w_066_1646, w_066_1647, w_066_1648, w_066_1649, w_066_1651, w_066_1653, w_066_1655, w_066_1657, w_066_1659, w_066_1661, w_066_1664, w_066_1667, w_066_1670, w_066_1673, w_066_1674, w_066_1679, w_066_1684, w_066_1685, w_066_1690, w_066_1692, w_066_1695, w_066_1696, w_066_1701, w_066_1706, w_066_1709, w_066_1710, w_066_1712, w_066_1716, w_066_1717, w_066_1720, w_066_1722, w_066_1723, w_066_1724, w_066_1725, w_066_1726, w_066_1728, w_066_1730, w_066_1731, w_066_1732, w_066_1733, w_066_1734, w_066_1735, w_066_1736, w_066_1738, w_066_1740, w_066_1742, w_066_1743, w_066_1744, w_066_1748, w_066_1750, w_066_1753, w_066_1754, w_066_1756, w_066_1759, w_066_1761, w_066_1762, w_066_1763, w_066_1764, w_066_1765, w_066_1767, w_066_1768, w_066_1772, w_066_1775, w_066_1778, w_066_1779, w_066_1780, w_066_1781, w_066_1782, w_066_1783, w_066_1786, w_066_1788, w_066_1789, w_066_1791, w_066_1792, w_066_1795, w_066_1797, w_066_1798, w_066_1799, w_066_1800, w_066_1801, w_066_1803, w_066_1806, w_066_1807, w_066_1811, w_066_1813, w_066_1814, w_066_1815, w_066_1816, w_066_1819, w_066_1828, w_066_1829, w_066_1835, w_066_1836, w_066_1837, w_066_1838, w_066_1841, w_066_1842, w_066_1843, w_066_1845, w_066_1848, w_066_1849, w_066_1850, w_066_1851, w_066_1852, w_066_1853, w_066_1855, w_066_1856, w_066_1857, w_066_1858, w_066_1859, w_066_1860, w_066_1861, w_066_1864, w_066_1865, w_066_1866, w_066_1867, w_066_1870, w_066_1871, w_066_1872, w_066_1873, w_066_1876, w_066_1880, w_066_1882, w_066_1885, w_066_1886, w_066_1887, w_066_1888, w_066_1890, w_066_1891, w_066_1892, w_066_1893, w_066_1894, w_066_1898, w_066_1899, w_066_1900, w_066_1901, w_066_1902, w_066_1904, w_066_1905, w_066_1909, w_066_1910, w_066_1912, w_066_1913, w_066_1914, w_066_1920, w_066_1924, w_066_1925, w_066_1928, w_066_1931, w_066_1934, w_066_1935, w_066_1940, w_066_1941, w_066_1943, w_066_1945, w_066_1949, w_066_1950, w_066_1951, w_066_1952, w_066_1953, w_066_1954, w_066_1955, w_066_1956, w_066_1957, w_066_1958, w_066_1959, w_066_1960, w_066_1961, w_066_1962, w_066_1963, w_066_1965, w_066_1967, w_066_1969, w_066_1972, w_066_1975, w_066_1976, w_066_1977, w_066_1978, w_066_1981, w_066_1983, w_066_1984, w_066_1985, w_066_1986, w_066_1987, w_066_1989, w_066_1990, w_066_1992, w_066_1993, w_066_1996, w_066_2002, w_066_2003, w_066_2005, w_066_2006, w_066_2009, w_066_2011, w_066_2012, w_066_2015, w_066_2017, w_066_2021, w_066_2023, w_066_2026, w_066_2028, w_066_2032, w_066_2037, w_066_2038, w_066_2039, w_066_2042, w_066_2044, w_066_2047, w_066_2050, w_066_2051, w_066_2052, w_066_2057, w_066_2060, w_066_2062, w_066_2065, w_066_2066, w_066_2067, w_066_2070, w_066_2073, w_066_2074, w_066_2075, w_066_2077, w_066_2078, w_066_2079, w_066_2081, w_066_2082, w_066_2084, w_066_2086, w_066_2087, w_066_2089, w_066_2090, w_066_2091, w_066_2092, w_066_2097, w_066_2099, w_066_2100, w_066_2101, w_066_2106, w_066_2107, w_066_2109, w_066_2110, w_066_2112, w_066_2113, w_066_2114, w_066_2115, w_066_2116, w_066_2117, w_066_2119, w_066_2120, w_066_2121, w_066_2122, w_066_2123, w_066_2125, w_066_2127, w_066_2128, w_066_2129, w_066_2130, w_066_2133, w_066_2135, w_066_2136, w_066_2138, w_066_2139, w_066_2141, w_066_2142, w_066_2143, w_066_2147, w_066_2148, w_066_2149, w_066_2152, w_066_2153, w_066_2154, w_066_2155, w_066_2156, w_066_2157, w_066_2159, w_066_2161, w_066_2162, w_066_2164, w_066_2166, w_066_2167, w_066_2168, w_066_2171, w_066_2172, w_066_2173, w_066_2178, w_066_2180, w_066_2182, w_066_2184, w_066_2185, w_066_2186, w_066_2187, w_066_2188, w_066_2189, w_066_2190, w_066_2191, w_066_2192, w_066_2195, w_066_2196, w_066_2197, w_066_2200, w_066_2201, w_066_2203, w_066_2206, w_066_2207, w_066_2211, w_066_2212, w_066_2213, w_066_2214, w_066_2216, w_066_2219, w_066_2220, w_066_2221, w_066_2222, w_066_2223, w_066_2224, w_066_2226, w_066_2229, w_066_2231, w_066_2233, w_066_2234, w_066_2235, w_066_2236, w_066_2238, w_066_2239, w_066_2241, w_066_2242, w_066_2243, w_066_2245, w_066_2246, w_066_2247, w_066_2249, w_066_2251, w_066_2255, w_066_2260, w_066_2261, w_066_2263, w_066_2264, w_066_2265, w_066_2266, w_066_2267, w_066_2268, w_066_2270, w_066_2271, w_066_2272, w_066_2273, w_066_2276, w_066_2283, w_066_2284, w_066_2286, w_066_2289, w_066_2292, w_066_2295, w_066_2297, w_066_2298, w_066_2299, w_066_2301, w_066_2305, w_066_2308, w_066_2309, w_066_2310, w_066_2311, w_066_2313, w_066_2315, w_066_2316, w_066_2318, w_066_2319, w_066_2320, w_066_2321, w_066_2325, w_066_2327, w_066_2329, w_066_2330, w_066_2331, w_066_2334, w_066_2335, w_066_2336, w_066_2338, w_066_2339, w_066_2340, w_066_2342, w_066_2343, w_066_2346, w_066_2350, w_066_2351, w_066_2352, w_066_2353, w_066_2356, w_066_2358, w_066_2359, w_066_2360, w_066_2361, w_066_2362, w_066_2364, w_066_2365, w_066_2367, w_066_2369, w_066_2370, w_066_2371, w_066_2372, w_066_2375, w_066_2376, w_066_2377, w_066_2378, w_066_2381, w_066_2384, w_066_2389, w_066_2390, w_066_2391, w_066_2392, w_066_2393, w_066_2395, w_066_2397, w_066_2399, w_066_2400, w_066_2403, w_066_2404, w_066_2405, w_066_2407, w_066_2408, w_066_2411, w_066_2412, w_066_2413, w_066_2414, w_066_2421, w_066_2422, w_066_2423, w_066_2425, w_066_2426, w_066_2427, w_066_2432, w_066_2436, w_066_2437, w_066_2438, w_066_2440, w_066_2442, w_066_2444, w_066_2446, w_066_2447, w_066_2450, w_066_2454, w_066_2456, w_066_2458, w_066_2460, w_066_2461, w_066_2462, w_066_2464, w_066_2467, w_066_2468, w_066_2469, w_066_2471, w_066_2472, w_066_2474, w_066_2475, w_066_2478, w_066_2479, w_066_2480, w_066_2485, w_066_2486, w_066_2487, w_066_2488, w_066_2489, w_066_2490, w_066_2492, w_066_2495, w_066_2496, w_066_2497, w_066_2498, w_066_2499, w_066_2500, w_066_2502, w_066_2506, w_066_2508, w_066_2509, w_066_2513, w_066_2515, w_066_2518, w_066_2521, w_066_2522, w_066_2523, w_066_2524, w_066_2525, w_066_2526, w_066_2527, w_066_2530, w_066_2532, w_066_2537, w_066_2541, w_066_2543, w_066_2546, w_066_2549, w_066_2550, w_066_2552, w_066_2554, w_066_2555, w_066_2557, w_066_2558, w_066_2559, w_066_2560, w_066_2561, w_066_2562, w_066_2564, w_066_2565, w_066_2566, w_066_2567, w_066_2569, w_066_2571, w_066_2572, w_066_2573, w_066_2574, w_066_2575, w_066_2576, w_066_2577, w_066_2580, w_066_2583, w_066_2584, w_066_2585, w_066_2586, w_066_2589, w_066_2590, w_066_2591, w_066_2592, w_066_2593, w_066_2594, w_066_2595, w_066_2597, w_066_2598, w_066_2599, w_066_2600, w_066_2602, w_066_2603, w_066_2605, w_066_2606, w_066_2607, w_066_2609, w_066_2611, w_066_2613, w_066_2614, w_066_2615, w_066_2616, w_066_2620, w_066_2621, w_066_2622, w_066_2625, w_066_2626, w_066_2627, w_066_2629, w_066_2630, w_066_2633, w_066_2636, w_066_2637, w_066_2639, w_066_2642, w_066_2643, w_066_2645, w_066_2648, w_066_2649, w_066_2650, w_066_2655, w_066_2656, w_066_2657, w_066_2660, w_066_2661, w_066_2662, w_066_2663, w_066_2666, w_066_2667, w_066_2668, w_066_2679, w_066_2681, w_066_2682, w_066_2683, w_066_2685, w_066_2686, w_066_2687, w_066_2688, w_066_2689, w_066_2695, w_066_2696, w_066_2697, w_066_2699, w_066_2702, w_066_2703, w_066_2705, w_066_2706, w_066_2707, w_066_2709, w_066_2710, w_066_2716, w_066_2718, w_066_2719, w_066_2721, w_066_2724, w_066_2725, w_066_2726, w_066_2727, w_066_2730, w_066_2731, w_066_2732, w_066_2735, w_066_2740, w_066_2741, w_066_2744, w_066_2748, w_066_2749, w_066_2750, w_066_2751, w_066_2753, w_066_2754, w_066_2759, w_066_2760, w_066_2762, w_066_2763, w_066_2765, w_066_2766, w_066_2770, w_066_2772, w_066_2773, w_066_2774, w_066_2777, w_066_2778, w_066_2780, w_066_2783, w_066_2784, w_066_2785, w_066_2786, w_066_2788, w_066_2792, w_066_2794, w_066_2795, w_066_2797, w_066_2799, w_066_2800, w_066_2801, w_066_2802, w_066_2803, w_066_2805, w_066_2806, w_066_2807, w_066_2808, w_066_2809, w_066_2810, w_066_2811, w_066_2813, w_066_2816, w_066_2818, w_066_2819, w_066_2820, w_066_2823, w_066_2824, w_066_2829, w_066_2830, w_066_2831, w_066_2834, w_066_2835, w_066_2836, w_066_2838, w_066_2839, w_066_2843, w_066_2846, w_066_2847, w_066_2850, w_066_2852, w_066_2854, w_066_2855, w_066_2858, w_066_2859, w_066_2860, w_066_2861, w_066_2862, w_066_2865, w_066_2866, w_066_2867, w_066_2868, w_066_2870, w_066_2871, w_066_2873, w_066_2878, w_066_2880, w_066_2881, w_066_2883, w_066_2884, w_066_2886, w_066_2890, w_066_2891, w_066_2894, w_066_2895, w_066_2900, w_066_2901, w_066_2902, w_066_2903, w_066_2904, w_066_2907, w_066_2908, w_066_2913, w_066_2914, w_066_2915, w_066_2916, w_066_2917, w_066_2918, w_066_2919, w_066_2920, w_066_2921, w_066_2922, w_066_2923, w_066_2924, w_066_2926, w_066_2928, w_066_2930, w_066_2932, w_066_2936, w_066_2937, w_066_2939, w_066_2941, w_066_2943, w_066_2944, w_066_2946, w_066_2947, w_066_2948, w_066_2949, w_066_2950, w_066_2951, w_066_2952, w_066_2953, w_066_2954, w_066_2955, w_066_2957, w_066_2958, w_066_2959, w_066_2960, w_066_2962, w_066_2964, w_066_2965, w_066_2966, w_066_2967, w_066_2974, w_066_2977, w_066_2978, w_066_2980, w_066_2982, w_066_2983, w_066_2985, w_066_2987, w_066_2988, w_066_2989, w_066_2990, w_066_2991, w_066_2993, w_066_2994, w_066_2996, w_066_2998, w_066_3003, w_066_3004, w_066_3006, w_066_3007, w_066_3008, w_066_3009, w_066_3010, w_066_3012, w_066_3013, w_066_3014, w_066_3017, w_066_3020, w_066_3022, w_066_3028, w_066_3031, w_066_3032, w_066_3033, w_066_3035, w_066_3037, w_066_3038, w_066_3039, w_066_3040, w_066_3041, w_066_3044, w_066_3046, w_066_3048, w_066_3049, w_066_3051, w_066_3053, w_066_3054, w_066_3055, w_066_3056, w_066_3058, w_066_3059, w_066_3060, w_066_3068, w_066_3069, w_066_3070, w_066_3072, w_066_3073, w_066_3074, w_066_3078, w_066_3079, w_066_3082, w_066_3083, w_066_3084, w_066_3086, w_066_3089, w_066_3090, w_066_3093, w_066_3094, w_066_3097, w_066_3098, w_066_3100, w_066_3101, w_066_3102, w_066_3104, w_066_3105, w_066_3107, w_066_3108, w_066_3110, w_066_3112, w_066_3117, w_066_3118, w_066_3119, w_066_3120, w_066_3122, w_066_3123, w_066_3124, w_066_3125, w_066_3127, w_066_3128, w_066_3130, w_066_3131, w_066_3132, w_066_3133, w_066_3134, w_066_3136, w_066_3138, w_066_3139, w_066_3141, w_066_3142, w_066_3144, w_066_3147, w_066_3149, w_066_3150, w_066_3151, w_066_3152, w_066_3155, w_066_3157, w_066_3160, w_066_3161, w_066_3162, w_066_3163, w_066_3164, w_066_3166, w_066_3167, w_066_3172, w_066_3173, w_066_3176, w_066_3178, w_066_3179, w_066_3180, w_066_3181, w_066_3185, w_066_3187, w_066_3189, w_066_3190, w_066_3191, w_066_3192, w_066_3193, w_066_3194, w_066_3196, w_066_3197, w_066_3200, w_066_3201, w_066_3202, w_066_3204, w_066_3207, w_066_3208, w_066_3212, w_066_3214, w_066_3216, w_066_3218, w_066_3219, w_066_3220, w_066_3224, w_066_3225, w_066_3227, w_066_3228, w_066_3229, w_066_3230, w_066_3231, w_066_3235, w_066_3237, w_066_3238, w_066_3239, w_066_3244, w_066_3247, w_066_3248, w_066_3249, w_066_3251, w_066_3252, w_066_3253, w_066_3254, w_066_3255, w_066_3256, w_066_3262, w_066_3263, w_066_3264, w_066_3265, w_066_3268, w_066_3270, w_066_3274, w_066_3275, w_066_3277, w_066_3278, w_066_3281, w_066_3283, w_066_3287, w_066_3288, w_066_3289, w_066_3290, w_066_3292, w_066_3294, w_066_3295, w_066_3296, w_066_3300, w_066_3301, w_066_3307, w_066_3310, w_066_3311, w_066_3312, w_066_3313, w_066_3314, w_066_3316, w_066_3317, w_066_3323, w_066_3327, w_066_3329, w_066_3331, w_066_3332, w_066_3333, w_066_3336, w_066_3337, w_066_3338, w_066_3339, w_066_3340, w_066_3341, w_066_3343, w_066_3348, w_066_3349, w_066_3350, w_066_3351, w_066_3352, w_066_3354, w_066_3356, w_066_3357, w_066_3360, w_066_3363, w_066_3364, w_066_3368, w_066_3369, w_066_3372, w_066_3373, w_066_3376, w_066_3377, w_066_3379, w_066_3380, w_066_3381, w_066_3382, w_066_3383, w_066_3384, w_066_3385, w_066_3386, w_066_3387, w_066_3391, w_066_3392, w_066_3395, w_066_3399, w_066_3400, w_066_3401, w_066_3402, w_066_3404, w_066_3405, w_066_3406, w_066_3407, w_066_3408, w_066_3410, w_066_3411, w_066_3412, w_066_3418, w_066_3419, w_066_3421, w_066_3422, w_066_3423, w_066_3425, w_066_3426, w_066_3428, w_066_3431, w_066_3432, w_066_3433, w_066_3436, w_066_3437, w_066_3438, w_066_3440, w_066_3441, w_066_3443, w_066_3445, w_066_3446, w_066_3449, w_066_3451, w_066_3453, w_066_3454, w_066_3455, w_066_3457, w_066_3458, w_066_3461, w_066_3463, w_066_3466, w_066_3467, w_066_3468, w_066_3474, w_066_3477, w_066_3479, w_066_3481, w_066_3482, w_066_3485, w_066_3486, w_066_3487, w_066_3490, w_066_3491, w_066_3492, w_066_3494, w_066_3496, w_066_3497, w_066_3499, w_066_3502, w_066_3505, w_066_3507, w_066_3508, w_066_3509, w_066_3510, w_066_3511, w_066_3512, w_066_3513, w_066_3514, w_066_3518, w_066_3519, w_066_3520, w_066_3521, w_066_3522, w_066_3523, w_066_3525, w_066_3526, w_066_3529, w_066_3532, w_066_3534, w_066_3535, w_066_3536, w_066_3538, w_066_3539, w_066_3542, w_066_3543, w_066_3549, w_066_3552, w_066_3554, w_066_3555, w_066_3557, w_066_3558, w_066_3559, w_066_3560, w_066_3561, w_066_3562, w_066_3563, w_066_3566, w_066_3567, w_066_3568, w_066_3570, w_066_3572, w_066_3573, w_066_3575, w_066_3576, w_066_3577, w_066_3578, w_066_3579, w_066_3580, w_066_3581, w_066_3582, w_066_3583, w_066_3584, w_066_3585, w_066_3588, w_066_3590, w_066_3592, w_066_3593, w_066_3594, w_066_3596, w_066_3600, w_066_3601, w_066_3602, w_066_3604, w_066_3605, w_066_3606, w_066_3607, w_066_3609, w_066_3611, w_066_3613, w_066_3614, w_066_3615, w_066_3618, w_066_3620, w_066_3622, w_066_3626, w_066_3628, w_066_3631, w_066_3633, w_066_3634, w_066_3637, w_066_3638, w_066_3640, w_066_3641, w_066_3642, w_066_3643, w_066_3644, w_066_3648, w_066_3649, w_066_3650, w_066_3651, w_066_3653, w_066_3654, w_066_3655, w_066_3656, w_066_3659, w_066_3667, w_066_3669, w_066_3670, w_066_3672, w_066_3673, w_066_3678, w_066_3680, w_066_3681, w_066_3682, w_066_3689, w_066_3690, w_066_3695, w_066_3698, w_066_3700, w_066_3701, w_066_3703, w_066_3704, w_066_3706, w_066_3708, w_066_3709, w_066_3711, w_066_3712, w_066_3713, w_066_3714, w_066_3717, w_066_3719, w_066_3722, w_066_3723, w_066_3724, w_066_3726, w_066_3728, w_066_3730, w_066_3732, w_066_3734, w_066_3735, w_066_3737, w_066_3738, w_066_3739, w_066_3740, w_066_3742, w_066_3744, w_066_3746, w_066_3747, w_066_3751, w_066_3753, w_066_3754, w_066_3757, w_066_3758, w_066_3759, w_066_3760, w_066_3761, w_066_3763, w_066_3764, w_066_3765, w_066_3766, w_066_3767, w_066_3768, w_066_3769, w_066_3771, w_066_3776, w_066_3779, w_066_3782, w_066_3786, w_066_3787, w_066_3788, w_066_3789, w_066_3791, w_066_3792, w_066_3793, w_066_3794, w_066_3795, w_066_3798, w_066_3803, w_066_3807, w_066_3808, w_066_3809, w_066_3811, w_066_3812, w_066_3814, w_066_3817, w_066_3818, w_066_3820, w_066_3821, w_066_3823, w_066_3827, w_066_3828, w_066_3830, w_066_3831, w_066_3832, w_066_3833, w_066_3834, w_066_3836, w_066_3837, w_066_3838, w_066_3842, w_066_3846, w_066_3847, w_066_3848, w_066_3849, w_066_3850, w_066_3851, w_066_3852, w_066_3856, w_066_3857, w_066_3858, w_066_3859, w_066_3860, w_066_3862, w_066_3864, w_066_3865, w_066_3869, w_066_3870, w_066_3873, w_066_3874, w_066_3875, w_066_3877, w_066_3880, w_066_3884, w_066_3888, w_066_3889, w_066_3891, w_066_3892, w_066_3893, w_066_3895, w_066_3896, w_066_3899, w_066_3900, w_066_3904, w_066_3905, w_066_3906, w_066_3907, w_066_3911, w_066_3913, w_066_3914, w_066_3915, w_066_3916, w_066_3918, w_066_3922, w_066_3923, w_066_3924, w_066_3925, w_066_3927, w_066_3929, w_066_3932, w_066_3933, w_066_3935, w_066_3938, w_066_3940, w_066_3943, w_066_3944, w_066_3949, w_066_3953, w_066_3955, w_066_3956, w_066_3958, w_066_3961, w_066_3962, w_066_3963, w_066_3966, w_066_3969, w_066_3970, w_066_3971, w_066_3973, w_066_3975, w_066_3976, w_066_3977, w_066_3981, w_066_3982, w_066_3984, w_066_3988, w_066_3990, w_066_3991, w_066_3993, w_066_3994, w_066_3996, w_066_4001, w_066_4007, w_066_4010, w_066_4011, w_066_4012, w_066_4019, w_066_4020, w_066_4024, w_066_4025, w_066_4026, w_066_4028, w_066_4032, w_066_4033, w_066_4036, w_066_4037, w_066_4043, w_066_4044, w_066_4046, w_066_4047, w_066_4049, w_066_4050, w_066_4051, w_066_4053, w_066_4054, w_066_4055, w_066_4056, w_066_4057, w_066_4058, w_066_4059, w_066_4061, w_066_4063, w_066_4064, w_066_4067, w_066_4070, w_066_4072, w_066_4073, w_066_4074, w_066_4075, w_066_4077, w_066_4081, w_066_4082, w_066_4084, w_066_4087, w_066_4088, w_066_4091, w_066_4092, w_066_4093, w_066_4095, w_066_4096, w_066_4098, w_066_4099, w_066_4103, w_066_4105, w_066_4107, w_066_4109, w_066_4111, w_066_4112, w_066_4116, w_066_4117, w_066_4118, w_066_4120, w_066_4122, w_066_4123, w_066_4124, w_066_4125, w_066_4126, w_066_4127, w_066_4129, w_066_4130, w_066_4132, w_066_4135, w_066_4136, w_066_4139, w_066_4140, w_066_4141, w_066_4142, w_066_4145, w_066_4146, w_066_4147, w_066_4148, w_066_4149, w_066_4151, w_066_4152, w_066_4153, w_066_4155, w_066_4156, w_066_4157, w_066_4159, w_066_4161, w_066_4163, w_066_4164, w_066_4165, w_066_4168, w_066_4170, w_066_4171, w_066_4172, w_066_4175, w_066_4176, w_066_4178, w_066_4181, w_066_4185, w_066_4186, w_066_4188, w_066_4191, w_066_4195, w_066_4196, w_066_4198, w_066_4201, w_066_4202, w_066_4205, w_066_4207, w_066_4209, w_066_4210, w_066_4212, w_066_4213, w_066_4214, w_066_4215, w_066_4216, w_066_4217, w_066_4218, w_066_4219, w_066_4220, w_066_4221, w_066_4224, w_066_4225, w_066_4230, w_066_4232, w_066_4233, w_066_4240, w_066_4241, w_066_4243, w_066_4244, w_066_4247, w_066_4250, w_066_4252, w_066_4253, w_066_4258, w_066_4259, w_066_4260, w_066_4261, w_066_4265, w_066_4268, w_066_4270, w_066_4272, w_066_4275, w_066_4276, w_066_4280, w_066_4283, w_066_4285, w_066_4286, w_066_4288, w_066_4289, w_066_4291, w_066_4292, w_066_4295, w_066_4297, w_066_4298, w_066_4303, w_066_4304, w_066_4305, w_066_4306, w_066_4309, w_066_4310, w_066_4311, w_066_4313, w_066_4314, w_066_4318, w_066_4319, w_066_4321, w_066_4323, w_066_4324, w_066_4325, w_066_4326, w_066_4327, w_066_4330, w_066_4331, w_066_4332, w_066_4336, w_066_4337, w_066_4338, w_066_4339, w_066_4340, w_066_4342, w_066_4343, w_066_4344, w_066_4348, w_066_4350, w_066_4353, w_066_4354, w_066_4358, w_066_4359, w_066_4360, w_066_4361, w_066_4364, w_066_4365, w_066_4366, w_066_4369;
  wire w_067_000, w_067_001, w_067_002, w_067_003, w_067_004, w_067_005, w_067_006, w_067_007, w_067_008, w_067_009, w_067_010, w_067_011, w_067_012, w_067_016, w_067_017, w_067_019, w_067_021, w_067_022, w_067_023, w_067_024, w_067_025, w_067_026, w_067_027, w_067_028, w_067_029, w_067_031, w_067_032, w_067_034, w_067_035, w_067_036, w_067_038, w_067_040, w_067_041, w_067_043, w_067_044, w_067_045, w_067_049, w_067_050, w_067_051, w_067_052, w_067_054, w_067_055, w_067_057, w_067_058, w_067_059, w_067_061, w_067_062, w_067_063, w_067_064, w_067_065, w_067_066, w_067_070, w_067_071, w_067_072, w_067_074, w_067_075, w_067_076, w_067_077, w_067_080, w_067_081, w_067_082, w_067_083, w_067_084, w_067_085, w_067_088, w_067_091, w_067_092, w_067_093, w_067_095, w_067_096, w_067_098, w_067_099, w_067_100, w_067_101, w_067_102, w_067_103, w_067_105, w_067_106, w_067_107, w_067_108, w_067_110, w_067_111, w_067_112, w_067_113, w_067_114, w_067_115, w_067_116, w_067_117, w_067_119, w_067_120, w_067_121, w_067_123, w_067_124, w_067_125, w_067_126, w_067_127, w_067_128, w_067_129, w_067_130, w_067_132, w_067_133, w_067_134, w_067_135, w_067_136, w_067_138, w_067_139, w_067_140, w_067_141, w_067_142, w_067_143, w_067_144, w_067_145, w_067_146, w_067_147, w_067_149, w_067_150, w_067_151, w_067_152, w_067_154, w_067_155, w_067_156, w_067_157, w_067_158, w_067_159, w_067_161, w_067_164, w_067_165, w_067_166, w_067_168, w_067_169, w_067_170, w_067_171, w_067_173, w_067_174, w_067_176, w_067_177, w_067_179, w_067_182, w_067_184, w_067_185, w_067_187, w_067_188, w_067_189, w_067_190, w_067_191, w_067_192, w_067_196, w_067_197, w_067_198, w_067_199, w_067_200, w_067_201, w_067_202, w_067_203, w_067_204, w_067_205, w_067_206, w_067_207, w_067_208, w_067_209, w_067_211, w_067_212, w_067_213, w_067_214, w_067_215, w_067_216, w_067_217, w_067_218, w_067_219, w_067_220, w_067_221, w_067_222, w_067_223, w_067_224, w_067_225, w_067_226, w_067_227, w_067_228, w_067_229, w_067_230, w_067_231, w_067_232, w_067_233, w_067_236, w_067_237, w_067_239, w_067_240, w_067_243, w_067_245, w_067_247, w_067_248, w_067_249, w_067_250, w_067_251, w_067_252, w_067_253, w_067_254, w_067_256, w_067_257, w_067_258, w_067_259, w_067_260, w_067_261, w_067_262, w_067_263, w_067_264, w_067_265, w_067_266, w_067_267, w_067_268, w_067_269, w_067_272, w_067_273, w_067_275, w_067_278, w_067_279, w_067_280, w_067_281, w_067_282, w_067_284, w_067_285, w_067_286, w_067_287, w_067_289, w_067_291, w_067_292, w_067_293, w_067_294, w_067_296, w_067_297, w_067_298, w_067_300, w_067_303, w_067_305, w_067_306, w_067_307, w_067_309, w_067_310, w_067_311, w_067_312, w_067_315, w_067_316, w_067_318, w_067_319, w_067_320, w_067_321, w_067_323, w_067_324, w_067_325, w_067_326, w_067_327, w_067_328, w_067_329, w_067_330, w_067_331, w_067_334, w_067_336, w_067_337, w_067_338, w_067_340, w_067_341, w_067_343, w_067_344, w_067_345, w_067_346, w_067_347, w_067_348, w_067_349, w_067_350, w_067_351, w_067_352, w_067_353, w_067_354, w_067_355, w_067_356, w_067_357, w_067_360, w_067_361, w_067_363, w_067_364, w_067_366, w_067_367, w_067_368, w_067_369, w_067_370, w_067_371, w_067_372, w_067_373, w_067_375, w_067_376, w_067_377, w_067_378, w_067_379, w_067_380, w_067_381, w_067_382, w_067_383, w_067_384, w_067_385, w_067_386, w_067_388, w_067_389, w_067_390, w_067_391, w_067_393, w_067_394, w_067_395, w_067_396, w_067_397, w_067_398, w_067_399, w_067_401, w_067_403, w_067_404, w_067_405, w_067_406, w_067_407, w_067_410, w_067_414, w_067_415, w_067_416, w_067_418, w_067_419, w_067_420, w_067_421, w_067_422, w_067_423, w_067_424, w_067_425, w_067_426, w_067_428, w_067_429, w_067_430, w_067_431, w_067_432, w_067_433, w_067_434, w_067_435, w_067_436, w_067_437, w_067_439, w_067_440, w_067_441, w_067_442, w_067_443, w_067_444, w_067_445, w_067_446, w_067_447, w_067_448, w_067_449, w_067_450, w_067_451, w_067_452, w_067_453, w_067_455, w_067_456, w_067_457, w_067_459, w_067_460, w_067_461, w_067_462, w_067_463, w_067_464, w_067_466, w_067_467, w_067_468, w_067_469, w_067_471, w_067_472, w_067_473, w_067_474, w_067_476, w_067_477, w_067_478, w_067_479, w_067_480, w_067_481, w_067_482, w_067_483, w_067_484, w_067_487, w_067_488, w_067_489, w_067_490, w_067_491, w_067_494, w_067_495, w_067_496, w_067_497, w_067_498, w_067_500, w_067_501, w_067_502, w_067_504, w_067_508, w_067_509, w_067_510, w_067_511, w_067_512, w_067_514, w_067_515, w_067_516, w_067_517, w_067_518, w_067_521, w_067_522, w_067_523, w_067_524, w_067_525, w_067_526, w_067_527, w_067_528, w_067_529, w_067_530, w_067_531, w_067_532, w_067_534, w_067_535, w_067_536, w_067_537, w_067_538, w_067_539, w_067_540, w_067_541, w_067_542, w_067_543, w_067_545, w_067_546, w_067_547, w_067_548, w_067_549, w_067_550, w_067_552, w_067_553, w_067_554, w_067_555, w_067_556, w_067_557, w_067_558, w_067_559, w_067_560, w_067_561, w_067_562, w_067_563, w_067_564, w_067_568, w_067_569, w_067_570, w_067_571, w_067_572, w_067_573, w_067_575, w_067_576, w_067_577, w_067_579, w_067_580, w_067_581, w_067_583, w_067_584, w_067_586, w_067_587, w_067_588, w_067_589, w_067_590, w_067_592, w_067_593, w_067_594, w_067_595, w_067_596, w_067_598, w_067_599, w_067_600, w_067_601, w_067_602, w_067_604, w_067_605, w_067_607, w_067_608, w_067_609, w_067_611, w_067_612, w_067_613, w_067_614, w_067_615, w_067_616, w_067_617, w_067_619, w_067_621, w_067_622, w_067_623, w_067_624, w_067_625, w_067_626, w_067_627, w_067_628, w_067_629, w_067_630, w_067_631, w_067_632, w_067_633, w_067_634, w_067_637, w_067_639, w_067_640, w_067_641, w_067_643, w_067_644, w_067_645, w_067_646, w_067_648, w_067_649, w_067_650, w_067_652, w_067_653, w_067_655, w_067_657, w_067_658, w_067_659, w_067_660, w_067_661, w_067_662, w_067_664, w_067_666, w_067_667, w_067_668, w_067_669, w_067_670, w_067_671, w_067_673, w_067_675, w_067_676, w_067_677, w_067_678, w_067_679, w_067_681, w_067_682, w_067_683, w_067_684, w_067_685, w_067_686, w_067_689, w_067_691, w_067_694, w_067_696, w_067_698, w_067_699, w_067_700, w_067_701, w_067_702, w_067_703, w_067_704, w_067_705, w_067_706, w_067_707, w_067_708, w_067_709, w_067_710, w_067_712, w_067_713, w_067_714, w_067_715, w_067_716, w_067_717, w_067_718, w_067_719, w_067_720, w_067_721, w_067_722, w_067_724, w_067_725, w_067_726, w_067_727, w_067_728, w_067_729, w_067_732, w_067_733, w_067_737, w_067_739, w_067_740, w_067_741, w_067_742, w_067_743, w_067_744, w_067_745, w_067_746, w_067_748, w_067_752, w_067_753, w_067_755, w_067_756, w_067_757, w_067_758, w_067_759, w_067_760, w_067_763, w_067_764, w_067_765, w_067_766, w_067_767, w_067_770, w_067_771, w_067_773, w_067_775, w_067_776, w_067_777, w_067_779, w_067_780, w_067_782, w_067_783, w_067_784, w_067_786, w_067_787, w_067_788, w_067_789, w_067_790, w_067_791, w_067_792, w_067_793, w_067_794, w_067_795, w_067_797, w_067_798, w_067_799, w_067_800, w_067_802, w_067_803, w_067_804, w_067_805, w_067_806, w_067_807, w_067_808, w_067_809, w_067_810, w_067_811, w_067_812, w_067_813, w_067_814, w_067_815, w_067_817, w_067_818, w_067_819, w_067_821, w_067_823, w_067_824, w_067_825, w_067_826, w_067_828, w_067_829, w_067_830, w_067_831, w_067_832, w_067_834, w_067_835, w_067_836, w_067_837, w_067_838, w_067_840, w_067_841, w_067_843, w_067_844, w_067_845, w_067_846, w_067_847, w_067_849, w_067_851, w_067_852, w_067_854, w_067_855, w_067_856, w_067_857, w_067_858, w_067_861, w_067_862, w_067_863, w_067_864, w_067_865, w_067_867, w_067_868, w_067_869, w_067_870, w_067_871, w_067_872, w_067_873, w_067_874, w_067_875, w_067_876, w_067_877, w_067_878, w_067_879, w_067_880, w_067_881, w_067_882, w_067_883, w_067_885, w_067_887, w_067_888, w_067_889, w_067_892, w_067_893, w_067_894, w_067_895, w_067_897, w_067_899, w_067_900, w_067_901, w_067_902, w_067_904, w_067_905, w_067_906, w_067_907, w_067_908, w_067_910, w_067_913, w_067_914, w_067_915, w_067_916, w_067_917, w_067_919, w_067_920, w_067_921, w_067_922, w_067_923, w_067_924, w_067_925, w_067_927, w_067_928, w_067_929, w_067_931, w_067_932, w_067_933, w_067_934, w_067_935, w_067_936, w_067_937, w_067_940, w_067_941, w_067_942, w_067_943, w_067_944, w_067_945, w_067_946, w_067_947, w_067_948, w_067_949, w_067_950, w_067_951, w_067_952, w_067_953, w_067_955, w_067_956, w_067_957, w_067_958, w_067_959, w_067_960, w_067_961, w_067_963, w_067_965, w_067_967, w_067_968, w_067_969, w_067_974, w_067_975, w_067_976, w_067_977, w_067_979, w_067_982, w_067_983, w_067_984, w_067_985, w_067_986, w_067_987, w_067_989, w_067_990, w_067_991, w_067_992, w_067_993, w_067_994, w_067_995, w_067_996, w_067_997, w_067_998, w_067_999, w_067_1000, w_067_1001, w_067_1002, w_067_1003, w_067_1004, w_067_1005, w_067_1006, w_067_1007, w_067_1009, w_067_1010, w_067_1011, w_067_1012, w_067_1013, w_067_1014, w_067_1015, w_067_1016, w_067_1017, w_067_1019, w_067_1021, w_067_1022, w_067_1023, w_067_1025, w_067_1026, w_067_1027, w_067_1029, w_067_1030, w_067_1031, w_067_1032, w_067_1033, w_067_1034, w_067_1036, w_067_1039, w_067_1042, w_067_1043, w_067_1045, w_067_1046, w_067_1047, w_067_1049, w_067_1050, w_067_1052, w_067_1053, w_067_1054, w_067_1055, w_067_1056, w_067_1057, w_067_1058, w_067_1059, w_067_1060, w_067_1061, w_067_1063, w_067_1064, w_067_1066, w_067_1067, w_067_1068, w_067_1070, w_067_1071, w_067_1072, w_067_1073, w_067_1074, w_067_1075, w_067_1077, w_067_1079, w_067_1080, w_067_1082, w_067_1083, w_067_1084, w_067_1085, w_067_1086, w_067_1087, w_067_1088, w_067_1089, w_067_1090, w_067_1091, w_067_1092, w_067_1093, w_067_1094, w_067_1095, w_067_1096, w_067_1097, w_067_1098, w_067_1102, w_067_1103, w_067_1104, w_067_1106, w_067_1107, w_067_1110, w_067_1111, w_067_1112, w_067_1113, w_067_1114, w_067_1115, w_067_1116, w_067_1118, w_067_1119, w_067_1121, w_067_1122, w_067_1123, w_067_1124, w_067_1126, w_067_1127, w_067_1128, w_067_1129, w_067_1132, w_067_1134, w_067_1135, w_067_1136, w_067_1137, w_067_1138, w_067_1139, w_067_1140, w_067_1141, w_067_1142, w_067_1143, w_067_1147, w_067_1150, w_067_1151, w_067_1152, w_067_1154, w_067_1156, w_067_1158, w_067_1159, w_067_1161, w_067_1162, w_067_1165, w_067_1166, w_067_1167, w_067_1168, w_067_1169, w_067_1174, w_067_1175, w_067_1176, w_067_1177, w_067_1178, w_067_1179, w_067_1181, w_067_1182, w_067_1183, w_067_1184, w_067_1185, w_067_1186, w_067_1187, w_067_1188, w_067_1189, w_067_1191, w_067_1192, w_067_1194, w_067_1195, w_067_1196, w_067_1197, w_067_1199, w_067_1201, w_067_1202, w_067_1203, w_067_1205, w_067_1207, w_067_1208, w_067_1209, w_067_1210, w_067_1212, w_067_1214, w_067_1215, w_067_1216, w_067_1217, w_067_1218, w_067_1219, w_067_1220, w_067_1223, w_067_1224, w_067_1225, w_067_1226, w_067_1227, w_067_1228, w_067_1229, w_067_1230, w_067_1231, w_067_1232, w_067_1233, w_067_1235, w_067_1236, w_067_1237, w_067_1239, w_067_1240, w_067_1241, w_067_1242, w_067_1243, w_067_1244, w_067_1245, w_067_1246, w_067_1247, w_067_1248, w_067_1250, w_067_1251, w_067_1252, w_067_1253, w_067_1255, w_067_1257, w_067_1258, w_067_1259, w_067_1260, w_067_1262, w_067_1263, w_067_1264, w_067_1267, w_067_1268, w_067_1269, w_067_1270, w_067_1271, w_067_1272, w_067_1274, w_067_1277, w_067_1278, w_067_1281, w_067_1283, w_067_1284, w_067_1285, w_067_1286, w_067_1289, w_067_1290, w_067_1292, w_067_1293, w_067_1294, w_067_1295, w_067_1296, w_067_1298, w_067_1299, w_067_1300, w_067_1301, w_067_1302, w_067_1304, w_067_1305, w_067_1307, w_067_1310, w_067_1311, w_067_1313, w_067_1314, w_067_1315, w_067_1320, w_067_1321, w_067_1322, w_067_1323, w_067_1324, w_067_1325, w_067_1326, w_067_1327, w_067_1328, w_067_1329, w_067_1331, w_067_1332, w_067_1333, w_067_1334, w_067_1335, w_067_1336, w_067_1337, w_067_1338, w_067_1339, w_067_1341, w_067_1342, w_067_1346, w_067_1349, w_067_1350, w_067_1352, w_067_1353, w_067_1354, w_067_1355, w_067_1359, w_067_1360, w_067_1361, w_067_1362, w_067_1365, w_067_1367, w_067_1368, w_067_1369, w_067_1373, w_067_1374, w_067_1375, w_067_1377, w_067_1378, w_067_1379, w_067_1380, w_067_1381, w_067_1382, w_067_1383, w_067_1384, w_067_1387, w_067_1388, w_067_1389, w_067_1390, w_067_1391, w_067_1392, w_067_1393, w_067_1394, w_067_1395, w_067_1396, w_067_1397, w_067_1399, w_067_1401, w_067_1402, w_067_1403, w_067_1404, w_067_1405, w_067_1406, w_067_1407, w_067_1409, w_067_1410, w_067_1413, w_067_1414, w_067_1416, w_067_1417, w_067_1418, w_067_1422, w_067_1423, w_067_1424, w_067_1425, w_067_1426, w_067_1427, w_067_1428, w_067_1429, w_067_1431, w_067_1432, w_067_1435, w_067_1436, w_067_1437, w_067_1438, w_067_1439, w_067_1440, w_067_1441, w_067_1442, w_067_1443, w_067_1445, w_067_1451, w_067_1454, w_067_1455, w_067_1458, w_067_1459, w_067_1460, w_067_1461, w_067_1462, w_067_1464, w_067_1465, w_067_1466, w_067_1467, w_067_1471, w_067_1473, w_067_1474, w_067_1477, w_067_1478, w_067_1479, w_067_1480, w_067_1481, w_067_1482, w_067_1486, w_067_1487, w_067_1488, w_067_1490, w_067_1491, w_067_1492, w_067_1493, w_067_1494, w_067_1495, w_067_1496, w_067_1497, w_067_1498, w_067_1499, w_067_1500, w_067_1502, w_067_1503, w_067_1504, w_067_1505, w_067_1506, w_067_1507, w_067_1508, w_067_1510, w_067_1512, w_067_1513, w_067_1514, w_067_1515, w_067_1516, w_067_1518, w_067_1519, w_067_1520, w_067_1521, w_067_1522, w_067_1525, w_067_1526, w_067_1529, w_067_1530, w_067_1531, w_067_1532, w_067_1533, w_067_1535, w_067_1536, w_067_1539, w_067_1540, w_067_1541, w_067_1543, w_067_1544, w_067_1545, w_067_1546, w_067_1547, w_067_1548, w_067_1549, w_067_1550, w_067_1551, w_067_1552, w_067_1554, w_067_1556, w_067_1558, w_067_1559, w_067_1560, w_067_1561, w_067_1562, w_067_1563, w_067_1566, w_067_1568, w_067_1570, w_067_1571, w_067_1575, w_067_1576, w_067_1577, w_067_1578, w_067_1579, w_067_1580, w_067_1582, w_067_1583, w_067_1584, w_067_1585, w_067_1586, w_067_1587, w_067_1588, w_067_1589, w_067_1590, w_067_1591, w_067_1592, w_067_1593, w_067_1594, w_067_1596, w_067_1598, w_067_1599, w_067_1600, w_067_1602, w_067_1603, w_067_1604, w_067_1605, w_067_1607, w_067_1608, w_067_1609, w_067_1611, w_067_1612, w_067_1614, w_067_1615, w_067_1616, w_067_1617, w_067_1618, w_067_1619, w_067_1621, w_067_1622, w_067_1623, w_067_1624, w_067_1625, w_067_1626, w_067_1627, w_067_1630, w_067_1631, w_067_1632, w_067_1633, w_067_1634, w_067_1635, w_067_1636, w_067_1637, w_067_1638, w_067_1639, w_067_1640, w_067_1641, w_067_1642, w_067_1643, w_067_1646, w_067_1647, w_067_1648, w_067_1650, w_067_1651, w_067_1656, w_067_1658, w_067_1659, w_067_1660, w_067_1661, w_067_1662, w_067_1664, w_067_1665, w_067_1666, w_067_1667, w_067_1668, w_067_1669, w_067_1670, w_067_1671, w_067_1673, w_067_1675, w_067_1676, w_067_1677, w_067_1678, w_067_1680, w_067_1681, w_067_1683, w_067_1684, w_067_1685, w_067_1687, w_067_1688, w_067_1689, w_067_1690, w_067_1693, w_067_1695, w_067_1696, w_067_1697, w_067_1700, w_067_1701, w_067_1702, w_067_1703, w_067_1704, w_067_1705, w_067_1707, w_067_1708, w_067_1709, w_067_1710, w_067_1711, w_067_1713, w_067_1714, w_067_1715, w_067_1716, w_067_1717, w_067_1719, w_067_1720, w_067_1721, w_067_1723, w_067_1724, w_067_1727, w_067_1728, w_067_1729, w_067_1731, w_067_1732, w_067_1734, w_067_1736, w_067_1737, w_067_1738, w_067_1739, w_067_1740, w_067_1742, w_067_1743, w_067_1744, w_067_1746, w_067_1747, w_067_1748, w_067_1751, w_067_1752, w_067_1753, w_067_1754, w_067_1755, w_067_1758, w_067_1759, w_067_1762, w_067_1763, w_067_1764, w_067_1766, w_067_1767, w_067_1768, w_067_1771, w_067_1772, w_067_1773, w_067_1774, w_067_1775, w_067_1777, w_067_1778, w_067_1779, w_067_1781, w_067_1783, w_067_1785, w_067_1786, w_067_1787, w_067_1788, w_067_1789, w_067_1790, w_067_1791, w_067_1792, w_067_1794, w_067_1796, w_067_1797, w_067_1798, w_067_1799, w_067_1800, w_067_1801, w_067_1802, w_067_1803, w_067_1804, w_067_1805, w_067_1806, w_067_1808, w_067_1809, w_067_1810, w_067_1813, w_067_1815, w_067_1817, w_067_1818, w_067_1819, w_067_1820, w_067_1821, w_067_1823, w_067_1827, w_067_1828, w_067_1829, w_067_1830, w_067_1831, w_067_1833, w_067_1834, w_067_1837, w_067_1838, w_067_1840, w_067_1841, w_067_1843, w_067_1844, w_067_1845, w_067_1847, w_067_1848, w_067_1849, w_067_1851, w_067_1854, w_067_1855, w_067_1856, w_067_1858, w_067_1861, w_067_1864, w_067_1866, w_067_1867, w_067_1868, w_067_1869, w_067_1870, w_067_1872, w_067_1877, w_067_1880, w_067_1881, w_067_1882, w_067_1885, w_067_1886, w_067_1887, w_067_1888, w_067_1890, w_067_1891, w_067_1892, w_067_1893, w_067_1894, w_067_1895, w_067_1896, w_067_1898, w_067_1899, w_067_1900, w_067_1901, w_067_1902, w_067_1903, w_067_1906, w_067_1907, w_067_1908, w_067_1909, w_067_1910, w_067_1911, w_067_1913, w_067_1914, w_067_1915, w_067_1917, w_067_1920, w_067_1923, w_067_1925, w_067_1926, w_067_1927, w_067_1928, w_067_1929, w_067_1930, w_067_1932, w_067_1933, w_067_1935, w_067_1936, w_067_1938, w_067_1939, w_067_1940, w_067_1941, w_067_1943, w_067_1944, w_067_1945, w_067_1946, w_067_1947, w_067_1949, w_067_1950, w_067_1951, w_067_1953, w_067_1955, w_067_1956, w_067_1957, w_067_1958, w_067_1959, w_067_1960, w_067_1962, w_067_1963, w_067_1966, w_067_1967, w_067_1968, w_067_1969, w_067_1970, w_067_1972, w_067_1973, w_067_1974, w_067_1975, w_067_1976, w_067_1978, w_067_1981, w_067_1982, w_067_1983, w_067_1984, w_067_1985, w_067_1986, w_067_1989, w_067_1991, w_067_1992, w_067_1994, w_067_1997, w_067_1998, w_067_2000, w_067_2001, w_067_2002, w_067_2003, w_067_2005, w_067_2006, w_067_2007, w_067_2008, w_067_2010, w_067_2011, w_067_2012, w_067_2013, w_067_2014, w_067_2017, w_067_2018, w_067_2019, w_067_2021, w_067_2022, w_067_2023, w_067_2027, w_067_2028, w_067_2029, w_067_2031, w_067_2033, w_067_2034, w_067_2035, w_067_2038, w_067_2039, w_067_2041, w_067_2042, w_067_2043, w_067_2044, w_067_2045, w_067_2046, w_067_2047, w_067_2048, w_067_2050, w_067_2051, w_067_2052, w_067_2054, w_067_2055, w_067_2056, w_067_2057, w_067_2059, w_067_2060, w_067_2061, w_067_2062, w_067_2064, w_067_2065, w_067_2067, w_067_2069, w_067_2071, w_067_2072, w_067_2073, w_067_2074, w_067_2077, w_067_2078, w_067_2081, w_067_2083, w_067_2085, w_067_2087, w_067_2088, w_067_2089, w_067_2090, w_067_2091, w_067_2093, w_067_2094, w_067_2095, w_067_2096, w_067_2097, w_067_2098, w_067_2099, w_067_2100, w_067_2101, w_067_2102, w_067_2104, w_067_2106, w_067_2113, w_067_2115, w_067_2118, w_067_2123, w_067_2124, w_067_2125, w_067_2126, w_067_2128, w_067_2129, w_067_2130, w_067_2133, w_067_2134, w_067_2136, w_067_2137, w_067_2138, w_067_2140, w_067_2141, w_067_2142, w_067_2143, w_067_2144, w_067_2145, w_067_2146, w_067_2148, w_067_2149, w_067_2150, w_067_2151, w_067_2152, w_067_2153, w_067_2154, w_067_2155, w_067_2156, w_067_2157, w_067_2158, w_067_2160, w_067_2161, w_067_2163, w_067_2164, w_067_2165, w_067_2166, w_067_2168, w_067_2169, w_067_2171, w_067_2172, w_067_2173, w_067_2174, w_067_2175, w_067_2177, w_067_2179, w_067_2180, w_067_2181, w_067_2182, w_067_2183, w_067_2185, w_067_2190, w_067_2191, w_067_2193, w_067_2194, w_067_2195, w_067_2196, w_067_2197, w_067_2200, w_067_2202, w_067_2203, w_067_2206, w_067_2207, w_067_2208, w_067_2209, w_067_2210, w_067_2211, w_067_2213, w_067_2214, w_067_2215, w_067_2216, w_067_2218, w_067_2219, w_067_2220, w_067_2221, w_067_2223, w_067_2224, w_067_2226, w_067_2227, w_067_2230, w_067_2231, w_067_2232, w_067_2233, w_067_2234, w_067_2236, w_067_2240, w_067_2241, w_067_2242, w_067_2243, w_067_2246, w_067_2247, w_067_2248, w_067_2249, w_067_2251, w_067_2252, w_067_2253, w_067_2255, w_067_2258, w_067_2259, w_067_2261, w_067_2262, w_067_2263, w_067_2264, w_067_2265, w_067_2266, w_067_2267, w_067_2269, w_067_2271, w_067_2273, w_067_2274, w_067_2275, w_067_2276, w_067_2277, w_067_2278, w_067_2279, w_067_2280, w_067_2281, w_067_2283, w_067_2284, w_067_2285, w_067_2287, w_067_2288, w_067_2289, w_067_2291, w_067_2292, w_067_2293, w_067_2294, w_067_2296, w_067_2298, w_067_2299, w_067_2301, w_067_2302, w_067_2303, w_067_2305, w_067_2307, w_067_2308, w_067_2309, w_067_2310, w_067_2311, w_067_2312, w_067_2313, w_067_2315, w_067_2316, w_067_2317, w_067_2318, w_067_2321, w_067_2322, w_067_2324, w_067_2325, w_067_2326, w_067_2327, w_067_2328, w_067_2329, w_067_2330, w_067_2331, w_067_2332, w_067_2333, w_067_2334, w_067_2337, w_067_2338, w_067_2339, w_067_2340, w_067_2341, w_067_2342, w_067_2343, w_067_2344, w_067_2345, w_067_2346, w_067_2347, w_067_2348, w_067_2349, w_067_2350, w_067_2354, w_067_2355, w_067_2356, w_067_2357, w_067_2358, w_067_2359, w_067_2363, w_067_2364, w_067_2365, w_067_2367, w_067_2368, w_067_2369, w_067_2371, w_067_2372, w_067_2374, w_067_2375, w_067_2376, w_067_2379, w_067_2380, w_067_2381, w_067_2383, w_067_2384, w_067_2385, w_067_2389, w_067_2392, w_067_2393, w_067_2394, w_067_2395, w_067_2396, w_067_2397, w_067_2399, w_067_2400, w_067_2403, w_067_2405, w_067_2406, w_067_2408, w_067_2410, w_067_2413, w_067_2414, w_067_2415, w_067_2416, w_067_2420, w_067_2421, w_067_2423, w_067_2424, w_067_2426, w_067_2428, w_067_2430, w_067_2432, w_067_2433, w_067_2434, w_067_2435, w_067_2436, w_067_2437, w_067_2439, w_067_2441, w_067_2445, w_067_2447, w_067_2448, w_067_2449, w_067_2451, w_067_2452, w_067_2453, w_067_2454, w_067_2455, w_067_2457, w_067_2458, w_067_2460, w_067_2461, w_067_2464, w_067_2467, w_067_2468, w_067_2469, w_067_2472, w_067_2474, w_067_2475, w_067_2477, w_067_2479, w_067_2480, w_067_2481, w_067_2482, w_067_2483, w_067_2484, w_067_2485, w_067_2486, w_067_2487, w_067_2488, w_067_2490, w_067_2491, w_067_2494, w_067_2496, w_067_2497, w_067_2498, w_067_2499, w_067_2501, w_067_2502, w_067_2504, w_067_2505, w_067_2506, w_067_2507, w_067_2508, w_067_2509, w_067_2511, w_067_2512, w_067_2513, w_067_2515, w_067_2519, w_067_2520, w_067_2522, w_067_2523, w_067_2525, w_067_2527, w_067_2528, w_067_2530, w_067_2531, w_067_2532, w_067_2533, w_067_2534, w_067_2536, w_067_2537, w_067_2539, w_067_2540, w_067_2541, w_067_2542, w_067_2543, w_067_2545, w_067_2546, w_067_2547, w_067_2548, w_067_2550, w_067_2552, w_067_2553, w_067_2555, w_067_2556, w_067_2557, w_067_2558, w_067_2559, w_067_2562, w_067_2565, w_067_2566, w_067_2568, w_067_2569, w_067_2570, w_067_2572, w_067_2573, w_067_2577, w_067_2578, w_067_2579, w_067_2580, w_067_2582, w_067_2584, w_067_2585, w_067_2586, w_067_2587, w_067_2590, w_067_2592, w_067_2593, w_067_2595, w_067_2596, w_067_2597, w_067_2599, w_067_2600, w_067_2601, w_067_2602, w_067_2604, w_067_2605, w_067_2606, w_067_2607, w_067_2608, w_067_2609, w_067_2610, w_067_2611, w_067_2612, w_067_2613, w_067_2614, w_067_2615, w_067_2616, w_067_2617, w_067_2619, w_067_2620, w_067_2622, w_067_2623, w_067_2624, w_067_2625, w_067_2628, w_067_2629, w_067_2630, w_067_2631, w_067_2632, w_067_2633, w_067_2634, w_067_2635, w_067_2636, w_067_2637, w_067_2638, w_067_2640, w_067_2641, w_067_2643, w_067_2644, w_067_2646, w_067_2647, w_067_2648, w_067_2649, w_067_2652, w_067_2654, w_067_2656, w_067_2657, w_067_2659, w_067_2660, w_067_2662, w_067_2666, w_067_2667, w_067_2668, w_067_2671, w_067_2672, w_067_2673, w_067_2674, w_067_2675, w_067_2676, w_067_2678, w_067_2680, w_067_2681, w_067_2682, w_067_2684, w_067_2685, w_067_2686, w_067_2687, w_067_2690, w_067_2694, w_067_2695, w_067_2696, w_067_2697, w_067_2699, w_067_2700, w_067_2702, w_067_2704, w_067_2705, w_067_2706, w_067_2707, w_067_2708, w_067_2709, w_067_2710, w_067_2711, w_067_2714, w_067_2715, w_067_2716, w_067_2717, w_067_2719, w_067_2720, w_067_2721, w_067_2724, w_067_2725, w_067_2726, w_067_2727, w_067_2729, w_067_2733, w_067_2735, w_067_2738, w_067_2740, w_067_2741, w_067_2742, w_067_2743, w_067_2744, w_067_2746, w_067_2747, w_067_2749, w_067_2752, w_067_2753, w_067_2754, w_067_2756, w_067_2758, w_067_2759, w_067_2760, w_067_2761, w_067_2762, w_067_2763, w_067_2764, w_067_2765, w_067_2768, w_067_2769, w_067_2770, w_067_2771, w_067_2772, w_067_2773, w_067_2774, w_067_2775, w_067_2776, w_067_2777, w_067_2778, w_067_2779, w_067_2780, w_067_2782, w_067_2783, w_067_2784, w_067_2785, w_067_2786, w_067_2787, w_067_2788, w_067_2789, w_067_2790, w_067_2791, w_067_2792, w_067_2793, w_067_2794, w_067_2795, w_067_2796, w_067_2797, w_067_2799, w_067_2801, w_067_2802, w_067_2803, w_067_2804, w_067_2805, w_067_2809, w_067_2810, w_067_2812, w_067_2813, w_067_2814, w_067_2815, w_067_2816, w_067_2817, w_067_2818, w_067_2820, w_067_2822, w_067_2823, w_067_2824, w_067_2825, w_067_2827, w_067_2828, w_067_2830, w_067_2831, w_067_2832, w_067_2833, w_067_2835, w_067_2837, w_067_2838, w_067_2839, w_067_2842, w_067_2843, w_067_2844, w_067_2846, w_067_2847, w_067_2848, w_067_2850, w_067_2851, w_067_2852, w_067_2853, w_067_2854, w_067_2856, w_067_2857, w_067_2858, w_067_2859, w_067_2861, w_067_2863, w_067_2865, w_067_2866, w_067_2867, w_067_2870, w_067_2871, w_067_2872, w_067_2873, w_067_2874, w_067_2876, w_067_2877, w_067_2879, w_067_2881, w_067_2882, w_067_2883, w_067_2884, w_067_2885, w_067_2888, w_067_2889, w_067_2890, w_067_2891, w_067_2892, w_067_2894, w_067_2895, w_067_2896;
  wire w_068_002, w_068_006, w_068_008, w_068_012, w_068_013, w_068_014, w_068_015, w_068_017, w_068_018, w_068_020, w_068_021, w_068_022, w_068_023, w_068_024, w_068_025, w_068_028, w_068_029, w_068_030, w_068_032, w_068_033, w_068_034, w_068_036, w_068_039, w_068_040, w_068_041, w_068_045, w_068_049, w_068_050, w_068_054, w_068_055, w_068_056, w_068_057, w_068_059, w_068_062, w_068_063, w_068_064, w_068_066, w_068_069, w_068_070, w_068_071, w_068_073, w_068_074, w_068_075, w_068_076, w_068_079, w_068_083, w_068_085, w_068_087, w_068_089, w_068_090, w_068_092, w_068_093, w_068_094, w_068_096, w_068_097, w_068_100, w_068_101, w_068_103, w_068_104, w_068_106, w_068_107, w_068_108, w_068_112, w_068_113, w_068_114, w_068_115, w_068_118, w_068_119, w_068_120, w_068_122, w_068_123, w_068_124, w_068_125, w_068_126, w_068_127, w_068_130, w_068_131, w_068_133, w_068_134, w_068_136, w_068_140, w_068_141, w_068_142, w_068_143, w_068_144, w_068_145, w_068_150, w_068_153, w_068_154, w_068_157, w_068_159, w_068_160, w_068_163, w_068_164, w_068_165, w_068_167, w_068_168, w_068_169, w_068_171, w_068_172, w_068_174, w_068_175, w_068_177, w_068_178, w_068_180, w_068_181, w_068_182, w_068_183, w_068_186, w_068_189, w_068_190, w_068_191, w_068_192, w_068_194, w_068_196, w_068_198, w_068_200, w_068_204, w_068_207, w_068_210, w_068_212, w_068_213, w_068_216, w_068_220, w_068_225, w_068_226, w_068_228, w_068_231, w_068_233, w_068_234, w_068_236, w_068_237, w_068_238, w_068_239, w_068_241, w_068_244, w_068_245, w_068_251, w_068_252, w_068_254, w_068_255, w_068_257, w_068_258, w_068_259, w_068_260, w_068_261, w_068_262, w_068_263, w_068_264, w_068_274, w_068_275, w_068_280, w_068_281, w_068_282, w_068_283, w_068_284, w_068_285, w_068_288, w_068_289, w_068_290, w_068_291, w_068_293, w_068_294, w_068_295, w_068_297, w_068_299, w_068_300, w_068_301, w_068_302, w_068_303, w_068_307, w_068_310, w_068_311, w_068_315, w_068_318, w_068_319, w_068_320, w_068_321, w_068_322, w_068_324, w_068_325, w_068_328, w_068_333, w_068_334, w_068_335, w_068_337, w_068_338, w_068_340, w_068_342, w_068_344, w_068_346, w_068_350, w_068_351, w_068_354, w_068_356, w_068_357, w_068_358, w_068_359, w_068_364, w_068_368, w_068_371, w_068_376, w_068_377, w_068_378, w_068_379, w_068_380, w_068_381, w_068_386, w_068_389, w_068_390, w_068_391, w_068_392, w_068_393, w_068_394, w_068_396, w_068_397, w_068_398, w_068_399, w_068_401, w_068_402, w_068_404, w_068_409, w_068_410, w_068_411, w_068_413, w_068_415, w_068_416, w_068_417, w_068_420, w_068_421, w_068_424, w_068_425, w_068_429, w_068_434, w_068_436, w_068_437, w_068_438, w_068_439, w_068_441, w_068_442, w_068_443, w_068_445, w_068_446, w_068_448, w_068_449, w_068_450, w_068_451, w_068_452, w_068_453, w_068_454, w_068_457, w_068_458, w_068_459, w_068_462, w_068_466, w_068_469, w_068_470, w_068_471, w_068_473, w_068_476, w_068_478, w_068_479, w_068_481, w_068_482, w_068_483, w_068_484, w_068_486, w_068_491, w_068_493, w_068_494, w_068_495, w_068_496, w_068_497, w_068_499, w_068_500, w_068_502, w_068_504, w_068_505, w_068_506, w_068_507, w_068_508, w_068_509, w_068_510, w_068_511, w_068_512, w_068_515, w_068_516, w_068_517, w_068_518, w_068_520, w_068_521, w_068_522, w_068_530, w_068_531, w_068_533, w_068_534, w_068_535, w_068_537, w_068_538, w_068_540, w_068_543, w_068_545, w_068_547, w_068_548, w_068_550, w_068_553, w_068_554, w_068_555, w_068_558, w_068_563, w_068_568, w_068_569, w_068_570, w_068_571, w_068_572, w_068_573, w_068_574, w_068_576, w_068_577, w_068_578, w_068_579, w_068_581, w_068_582, w_068_583, w_068_584, w_068_586, w_068_587, w_068_589, w_068_593, w_068_594, w_068_595, w_068_596, w_068_597, w_068_598, w_068_599, w_068_600, w_068_601, w_068_602, w_068_603, w_068_605, w_068_606, w_068_607, w_068_608, w_068_609, w_068_610, w_068_612, w_068_615, w_068_616, w_068_617, w_068_621, w_068_622, w_068_625, w_068_626, w_068_627, w_068_632, w_068_636, w_068_638, w_068_640, w_068_641, w_068_645, w_068_647, w_068_648, w_068_651, w_068_652, w_068_653, w_068_654, w_068_658, w_068_659, w_068_660, w_068_661, w_068_666, w_068_668, w_068_670, w_068_671, w_068_675, w_068_676, w_068_677, w_068_680, w_068_682, w_068_685, w_068_689, w_068_690, w_068_691, w_068_692, w_068_697, w_068_699, w_068_700, w_068_701, w_068_702, w_068_703, w_068_704, w_068_706, w_068_708, w_068_711, w_068_712, w_068_715, w_068_716, w_068_717, w_068_718, w_068_719, w_068_722, w_068_723, w_068_726, w_068_727, w_068_728, w_068_729, w_068_732, w_068_733, w_068_736, w_068_741, w_068_742, w_068_744, w_068_746, w_068_749, w_068_751, w_068_754, w_068_756, w_068_757, w_068_758, w_068_759, w_068_760, w_068_761, w_068_763, w_068_764, w_068_765, w_068_768, w_068_769, w_068_771, w_068_773, w_068_774, w_068_776, w_068_777, w_068_778, w_068_779, w_068_780, w_068_782, w_068_784, w_068_785, w_068_786, w_068_787, w_068_789, w_068_790, w_068_791, w_068_792, w_068_794, w_068_795, w_068_796, w_068_801, w_068_802, w_068_803, w_068_804, w_068_805, w_068_806, w_068_807, w_068_809, w_068_810, w_068_812, w_068_813, w_068_814, w_068_815, w_068_816, w_068_817, w_068_818, w_068_819, w_068_820, w_068_822, w_068_823, w_068_827, w_068_829, w_068_830, w_068_834, w_068_839, w_068_840, w_068_841, w_068_842, w_068_843, w_068_844, w_068_845, w_068_846, w_068_847, w_068_850, w_068_851, w_068_852, w_068_854, w_068_855, w_068_856, w_068_858, w_068_861, w_068_862, w_068_863, w_068_865, w_068_866, w_068_869, w_068_872, w_068_873, w_068_876, w_068_878, w_068_883, w_068_885, w_068_886, w_068_887, w_068_889, w_068_892, w_068_893, w_068_895, w_068_898, w_068_900, w_068_901, w_068_905, w_068_906, w_068_909, w_068_910, w_068_912, w_068_913, w_068_918, w_068_920, w_068_921, w_068_922, w_068_923, w_068_924, w_068_926, w_068_927, w_068_930, w_068_933, w_068_934, w_068_936, w_068_937, w_068_939, w_068_940, w_068_944, w_068_946, w_068_948, w_068_952, w_068_954, w_068_955, w_068_957, w_068_958, w_068_959, w_068_963, w_068_964, w_068_965, w_068_967, w_068_971, w_068_972, w_068_974, w_068_975, w_068_976, w_068_977, w_068_978, w_068_979, w_068_980, w_068_982, w_068_984, w_068_985, w_068_988, w_068_989, w_068_990, w_068_991, w_068_992, w_068_995, w_068_996, w_068_997, w_068_998, w_068_999, w_068_1000, w_068_1001, w_068_1002, w_068_1004, w_068_1009, w_068_1011, w_068_1012, w_068_1014, w_068_1015, w_068_1018, w_068_1019, w_068_1022, w_068_1024, w_068_1027, w_068_1030, w_068_1031, w_068_1032, w_068_1033, w_068_1034, w_068_1036, w_068_1039, w_068_1041, w_068_1042, w_068_1044, w_068_1045, w_068_1046, w_068_1048, w_068_1049, w_068_1050, w_068_1052, w_068_1053, w_068_1054, w_068_1055, w_068_1056, w_068_1058, w_068_1063, w_068_1067, w_068_1069, w_068_1070, w_068_1071, w_068_1073, w_068_1074, w_068_1076, w_068_1077, w_068_1080, w_068_1081, w_068_1082, w_068_1083, w_068_1085, w_068_1086, w_068_1091, w_068_1093, w_068_1095, w_068_1098, w_068_1099, w_068_1100, w_068_1101, w_068_1102, w_068_1103, w_068_1104, w_068_1105, w_068_1110, w_068_1111, w_068_1112, w_068_1115, w_068_1116, w_068_1117, w_068_1119, w_068_1124, w_068_1125, w_068_1127, w_068_1128, w_068_1129, w_068_1130, w_068_1131, w_068_1134, w_068_1135, w_068_1137, w_068_1138, w_068_1140, w_068_1143, w_068_1144, w_068_1145, w_068_1146, w_068_1148, w_068_1149, w_068_1150, w_068_1152, w_068_1153, w_068_1154, w_068_1155, w_068_1156, w_068_1157, w_068_1158, w_068_1160, w_068_1161, w_068_1163, w_068_1175, w_068_1176, w_068_1179, w_068_1183, w_068_1185, w_068_1187, w_068_1188, w_068_1190, w_068_1191, w_068_1193, w_068_1194, w_068_1196, w_068_1199, w_068_1201, w_068_1204, w_068_1206, w_068_1209, w_068_1210, w_068_1212, w_068_1215, w_068_1216, w_068_1218, w_068_1219, w_068_1220, w_068_1221, w_068_1222, w_068_1224, w_068_1226, w_068_1229, w_068_1230, w_068_1233, w_068_1234, w_068_1235, w_068_1239, w_068_1242, w_068_1244, w_068_1245, w_068_1247, w_068_1248, w_068_1250, w_068_1253, w_068_1254, w_068_1256, w_068_1257, w_068_1259, w_068_1260, w_068_1262, w_068_1265, w_068_1266, w_068_1267, w_068_1274, w_068_1275, w_068_1276, w_068_1277, w_068_1278, w_068_1280, w_068_1282, w_068_1285, w_068_1286, w_068_1287, w_068_1288, w_068_1289, w_068_1294, w_068_1295, w_068_1296, w_068_1298, w_068_1299, w_068_1302, w_068_1304, w_068_1305, w_068_1306, w_068_1308, w_068_1309, w_068_1312, w_068_1314, w_068_1315, w_068_1317, w_068_1321, w_068_1323, w_068_1324, w_068_1325, w_068_1327, w_068_1328, w_068_1329, w_068_1331, w_068_1332, w_068_1334, w_068_1335, w_068_1337, w_068_1339, w_068_1340, w_068_1341, w_068_1343, w_068_1348, w_068_1349, w_068_1350, w_068_1354, w_068_1355, w_068_1357, w_068_1358, w_068_1359, w_068_1360, w_068_1361, w_068_1363, w_068_1365, w_068_1368, w_068_1370, w_068_1371, w_068_1372, w_068_1373, w_068_1374, w_068_1375, w_068_1376, w_068_1377, w_068_1380, w_068_1382, w_068_1383, w_068_1387, w_068_1388, w_068_1389, w_068_1390, w_068_1391, w_068_1394, w_068_1399, w_068_1400, w_068_1401, w_068_1402, w_068_1403, w_068_1406, w_068_1407, w_068_1408, w_068_1409, w_068_1413, w_068_1415, w_068_1416, w_068_1418, w_068_1419, w_068_1420, w_068_1421, w_068_1422, w_068_1424, w_068_1425, w_068_1426, w_068_1427, w_068_1431, w_068_1433, w_068_1435, w_068_1440, w_068_1442, w_068_1444, w_068_1445, w_068_1446, w_068_1447, w_068_1448, w_068_1450, w_068_1451, w_068_1455, w_068_1456, w_068_1460, w_068_1461, w_068_1465, w_068_1466, w_068_1467, w_068_1468, w_068_1469, w_068_1470, w_068_1471, w_068_1478, w_068_1479, w_068_1480, w_068_1481, w_068_1482, w_068_1483, w_068_1485, w_068_1486, w_068_1487, w_068_1488, w_068_1490, w_068_1491, w_068_1494, w_068_1496, w_068_1497, w_068_1499, w_068_1500, w_068_1504, w_068_1507, w_068_1508, w_068_1509, w_068_1512, w_068_1513, w_068_1517, w_068_1518, w_068_1519, w_068_1520, w_068_1522, w_068_1523, w_068_1524, w_068_1526, w_068_1527, w_068_1528, w_068_1534, w_068_1536, w_068_1539, w_068_1540, w_068_1542, w_068_1543, w_068_1545, w_068_1547, w_068_1549, w_068_1550, w_068_1551, w_068_1553, w_068_1554, w_068_1560, w_068_1561, w_068_1562, w_068_1566, w_068_1567, w_068_1568, w_068_1569, w_068_1570, w_068_1571, w_068_1572, w_068_1577, w_068_1578, w_068_1579, w_068_1580, w_068_1582, w_068_1586, w_068_1588, w_068_1589, w_068_1591, w_068_1593, w_068_1594, w_068_1596, w_068_1597, w_068_1598, w_068_1599, w_068_1600, w_068_1601, w_068_1603, w_068_1605, w_068_1606, w_068_1607, w_068_1611, w_068_1612, w_068_1613, w_068_1615, w_068_1618, w_068_1620, w_068_1621, w_068_1623, w_068_1624, w_068_1625, w_068_1626, w_068_1627, w_068_1628, w_068_1629, w_068_1631, w_068_1632, w_068_1635, w_068_1636, w_068_1637, w_068_1642, w_068_1643, w_068_1644, w_068_1647, w_068_1648, w_068_1650, w_068_1652, w_068_1656, w_068_1658, w_068_1660, w_068_1661, w_068_1662, w_068_1665, w_068_1668, w_068_1670, w_068_1672, w_068_1676, w_068_1677, w_068_1680, w_068_1681, w_068_1682, w_068_1683, w_068_1684, w_068_1685, w_068_1687, w_068_1690, w_068_1691, w_068_1692, w_068_1694, w_068_1695, w_068_1696, w_068_1697, w_068_1698, w_068_1699, w_068_1700, w_068_1701, w_068_1702, w_068_1704, w_068_1705, w_068_1706, w_068_1708, w_068_1709, w_068_1710, w_068_1712, w_068_1715, w_068_1717, w_068_1722, w_068_1724, w_068_1727, w_068_1731, w_068_1732, w_068_1734, w_068_1739, w_068_1741, w_068_1743, w_068_1744, w_068_1745, w_068_1747, w_068_1749, w_068_1750, w_068_1752, w_068_1753, w_068_1755, w_068_1758, w_068_1760, w_068_1762, w_068_1765, w_068_1767, w_068_1768, w_068_1769, w_068_1770, w_068_1773, w_068_1776, w_068_1778, w_068_1779, w_068_1783, w_068_1784, w_068_1785, w_068_1786, w_068_1789, w_068_1792, w_068_1793, w_068_1794, w_068_1795, w_068_1796, w_068_1797, w_068_1798, w_068_1799, w_068_1801, w_068_1802, w_068_1805, w_068_1809, w_068_1812, w_068_1813, w_068_1815, w_068_1816, w_068_1817, w_068_1818, w_068_1820, w_068_1821, w_068_1822, w_068_1824, w_068_1826, w_068_1827, w_068_1830, w_068_1836, w_068_1838, w_068_1839, w_068_1840, w_068_1842, w_068_1847, w_068_1848, w_068_1850, w_068_1852, w_068_1853, w_068_1854, w_068_1856, w_068_1858, w_068_1860, w_068_1863, w_068_1864, w_068_1865, w_068_1868, w_068_1872, w_068_1875, w_068_1876, w_068_1877, w_068_1881, w_068_1882, w_068_1883, w_068_1884, w_068_1886, w_068_1887, w_068_1888, w_068_1889, w_068_1891, w_068_1892, w_068_1895, w_068_1899, w_068_1900, w_068_1902, w_068_1903, w_068_1904, w_068_1906, w_068_1907, w_068_1908, w_068_1909, w_068_1911, w_068_1914, w_068_1915, w_068_1917, w_068_1918, w_068_1919, w_068_1921, w_068_1922, w_068_1923, w_068_1924, w_068_1927, w_068_1928, w_068_1929, w_068_1931, w_068_1934, w_068_1935, w_068_1936, w_068_1940, w_068_1941, w_068_1942, w_068_1943, w_068_1944, w_068_1945, w_068_1946, w_068_1947, w_068_1948, w_068_1949, w_068_1951, w_068_1952, w_068_1954, w_068_1955, w_068_1956, w_068_1957, w_068_1960, w_068_1961, w_068_1963, w_068_1967, w_068_1968, w_068_1969, w_068_1975, w_068_1979, w_068_1980, w_068_1981, w_068_1982, w_068_1985, w_068_1988, w_068_1990, w_068_1991, w_068_1992, w_068_1993, w_068_1994, w_068_1996, w_068_1997, w_068_2000, w_068_2002, w_068_2005, w_068_2006, w_068_2007, w_068_2008, w_068_2009, w_068_2010, w_068_2011, w_068_2012, w_068_2013, w_068_2014, w_068_2015, w_068_2016, w_068_2022, w_068_2023, w_068_2027, w_068_2028, w_068_2029, w_068_2030, w_068_2031, w_068_2032, w_068_2033, w_068_2034, w_068_2037, w_068_2038, w_068_2041, w_068_2045, w_068_2048, w_068_2051, w_068_2053, w_068_2054, w_068_2055, w_068_2058, w_068_2059, w_068_2060, w_068_2061, w_068_2062, w_068_2066, w_068_2068, w_068_2073, w_068_2074, w_068_2075, w_068_2076, w_068_2077, w_068_2078, w_068_2080, w_068_2081, w_068_2084, w_068_2085, w_068_2086, w_068_2090, w_068_2091, w_068_2092, w_068_2095, w_068_2096, w_068_2100, w_068_2101, w_068_2102, w_068_2103, w_068_2104, w_068_2109, w_068_2110, w_068_2111, w_068_2117, w_068_2121, w_068_2122, w_068_2126, w_068_2129, w_068_2132, w_068_2133, w_068_2135, w_068_2137, w_068_2138, w_068_2139, w_068_2140, w_068_2141, w_068_2142, w_068_2143, w_068_2144, w_068_2145, w_068_2146, w_068_2147, w_068_2148, w_068_2150, w_068_2151, w_068_2153, w_068_2154, w_068_2155, w_068_2156, w_068_2158, w_068_2159, w_068_2161, w_068_2162, w_068_2163, w_068_2164, w_068_2165, w_068_2166, w_068_2169, w_068_2171, w_068_2172, w_068_2174, w_068_2175, w_068_2177, w_068_2178, w_068_2179, w_068_2180, w_068_2181, w_068_2182, w_068_2183, w_068_2185, w_068_2186, w_068_2187, w_068_2190, w_068_2192, w_068_2197, w_068_2198, w_068_2200, w_068_2201, w_068_2202, w_068_2203, w_068_2204, w_068_2205, w_068_2206, w_068_2208, w_068_2209, w_068_2210, w_068_2211, w_068_2212, w_068_2214, w_068_2215, w_068_2216, w_068_2219, w_068_2220, w_068_2225, w_068_2227, w_068_2231, w_068_2235, w_068_2236, w_068_2237, w_068_2238, w_068_2239, w_068_2241, w_068_2242, w_068_2243, w_068_2248, w_068_2249, w_068_2250, w_068_2253, w_068_2255, w_068_2256, w_068_2260, w_068_2261, w_068_2262, w_068_2264, w_068_2266, w_068_2271, w_068_2273, w_068_2275, w_068_2278, w_068_2279, w_068_2283, w_068_2284, w_068_2285, w_068_2288, w_068_2292, w_068_2293, w_068_2295, w_068_2296, w_068_2297, w_068_2298, w_068_2299, w_068_2303, w_068_2304, w_068_2305, w_068_2306, w_068_2310, w_068_2314, w_068_2315, w_068_2316, w_068_2318, w_068_2319, w_068_2321, w_068_2322, w_068_2325, w_068_2326, w_068_2327, w_068_2328, w_068_2329, w_068_2331, w_068_2332, w_068_2333, w_068_2336, w_068_2337, w_068_2339, w_068_2344, w_068_2345, w_068_2346, w_068_2349, w_068_2351, w_068_2352, w_068_2353, w_068_2356, w_068_2357, w_068_2358, w_068_2359, w_068_2360, w_068_2361, w_068_2362, w_068_2364, w_068_2365, w_068_2366, w_068_2367, w_068_2368, w_068_2370, w_068_2372, w_068_2373, w_068_2376, w_068_2377, w_068_2378, w_068_2382, w_068_2383, w_068_2384, w_068_2385, w_068_2386, w_068_2389, w_068_2390, w_068_2393, w_068_2394, w_068_2397, w_068_2398, w_068_2401, w_068_2402, w_068_2404, w_068_2407, w_068_2410, w_068_2412, w_068_2413, w_068_2414, w_068_2416, w_068_2418, w_068_2421, w_068_2422, w_068_2423, w_068_2424, w_068_2426, w_068_2427, w_068_2428, w_068_2430, w_068_2432, w_068_2435, w_068_2439, w_068_2442, w_068_2444, w_068_2446, w_068_2447, w_068_2448, w_068_2449, w_068_2450, w_068_2451, w_068_2452, w_068_2454, w_068_2456, w_068_2457, w_068_2458, w_068_2459, w_068_2460, w_068_2461, w_068_2463, w_068_2465, w_068_2466, w_068_2467, w_068_2469, w_068_2470, w_068_2472, w_068_2474, w_068_2480, w_068_2484, w_068_2486, w_068_2487, w_068_2490, w_068_2491, w_068_2493, w_068_2496, w_068_2497, w_068_2501, w_068_2502, w_068_2503, w_068_2504, w_068_2505, w_068_2507, w_068_2510, w_068_2513, w_068_2514, w_068_2515, w_068_2517, w_068_2519, w_068_2520, w_068_2521, w_068_2522, w_068_2523, w_068_2525, w_068_2531, w_068_2532, w_068_2534, w_068_2535, w_068_2537, w_068_2538, w_068_2540, w_068_2541, w_068_2542, w_068_2544, w_068_2546, w_068_2547, w_068_2550, w_068_2552, w_068_2553, w_068_2556, w_068_2557, w_068_2562, w_068_2563, w_068_2565, w_068_2566, w_068_2568, w_068_2570, w_068_2571, w_068_2572, w_068_2574, w_068_2575, w_068_2578, w_068_2579, w_068_2582, w_068_2584, w_068_2589, w_068_2590, w_068_2591, w_068_2592, w_068_2593, w_068_2595, w_068_2598, w_068_2599, w_068_2600, w_068_2601, w_068_2603, w_068_2604, w_068_2605, w_068_2606, w_068_2607, w_068_2613, w_068_2614, w_068_2615, w_068_2618, w_068_2619, w_068_2620, w_068_2621, w_068_2623, w_068_2626, w_068_2627, w_068_2628, w_068_2632, w_068_2633, w_068_2635, w_068_2636, w_068_2637, w_068_2639, w_068_2640, w_068_2643, w_068_2646, w_068_2647, w_068_2650, w_068_2653, w_068_2654, w_068_2656, w_068_2657, w_068_2658, w_068_2660, w_068_2664, w_068_2667, w_068_2670, w_068_2671, w_068_2673, w_068_2674, w_068_2676, w_068_2680, w_068_2682, w_068_2684, w_068_2685, w_068_2686, w_068_2687, w_068_2690, w_068_2691, w_068_2692, w_068_2693, w_068_2694, w_068_2697, w_068_2698, w_068_2700, w_068_2701, w_068_2703, w_068_2705, w_068_2707, w_068_2708, w_068_2710, w_068_2712, w_068_2713, w_068_2714, w_068_2715, w_068_2716, w_068_2717, w_068_2718, w_068_2719, w_068_2722, w_068_2723, w_068_2724, w_068_2725, w_068_2726, w_068_2729, w_068_2731, w_068_2737, w_068_2743, w_068_2744, w_068_2748, w_068_2750, w_068_2752, w_068_2753, w_068_2755, w_068_2756, w_068_2757, w_068_2760, w_068_2761, w_068_2762, w_068_2764, w_068_2765, w_068_2769, w_068_2770, w_068_2772, w_068_2773, w_068_2774, w_068_2775, w_068_2776, w_068_2777, w_068_2778, w_068_2780, w_068_2781, w_068_2784, w_068_2785, w_068_2788, w_068_2789, w_068_2790, w_068_2791, w_068_2793, w_068_2797, w_068_2798, w_068_2800, w_068_2803, w_068_2805, w_068_2807, w_068_2808, w_068_2809, w_068_2811, w_068_2813, w_068_2814, w_068_2815, w_068_2816, w_068_2817, w_068_2823, w_068_2825, w_068_2828, w_068_2830, w_068_2832, w_068_2833, w_068_2834, w_068_2838, w_068_2840, w_068_2841, w_068_2842, w_068_2843, w_068_2844, w_068_2846, w_068_2847, w_068_2849, w_068_2851, w_068_2853, w_068_2855, w_068_2856, w_068_2857, w_068_2858, w_068_2859, w_068_2860, w_068_2861, w_068_2863, w_068_2864, w_068_2865, w_068_2866, w_068_2867, w_068_2869, w_068_2870, w_068_2874, w_068_2876, w_068_2882, w_068_2884, w_068_2885, w_068_2888, w_068_2893, w_068_2897, w_068_2901, w_068_2903, w_068_2905, w_068_2906, w_068_2910, w_068_2911, w_068_2913, w_068_2915, w_068_2917, w_068_2919, w_068_2922, w_068_2924, w_068_2926, w_068_2927, w_068_2928, w_068_2931, w_068_2933, w_068_2934, w_068_2935, w_068_2936, w_068_2937, w_068_2938, w_068_2941, w_068_2942, w_068_2944, w_068_2945, w_068_2949, w_068_2953, w_068_2954, w_068_2955, w_068_2956, w_068_2958, w_068_2959, w_068_2962, w_068_2963, w_068_2964, w_068_2965, w_068_2966, w_068_2967, w_068_2968, w_068_2970, w_068_2972, w_068_2975, w_068_2977, w_068_2978, w_068_2979, w_068_2982, w_068_2984, w_068_2987, w_068_2989, w_068_2990, w_068_2992, w_068_2993, w_068_2994, w_068_2995, w_068_2996, w_068_2997, w_068_2999, w_068_3000, w_068_3001, w_068_3002, w_068_3003, w_068_3006, w_068_3007, w_068_3010, w_068_3011, w_068_3013, w_068_3015, w_068_3016, w_068_3018, w_068_3019, w_068_3023, w_068_3025, w_068_3027, w_068_3028, w_068_3029, w_068_3030, w_068_3031, w_068_3032, w_068_3033, w_068_3035, w_068_3036, w_068_3039, w_068_3040, w_068_3043, w_068_3044, w_068_3047, w_068_3050, w_068_3051, w_068_3053, w_068_3056, w_068_3058, w_068_3059, w_068_3065, w_068_3066, w_068_3067, w_068_3069, w_068_3071, w_068_3072, w_068_3073, w_068_3075, w_068_3076, w_068_3077, w_068_3078, w_068_3080, w_068_3082, w_068_3083, w_068_3084, w_068_3085, w_068_3086, w_068_3087, w_068_3088, w_068_3090, w_068_3091, w_068_3092, w_068_3093, w_068_3095, w_068_3096, w_068_3099, w_068_3100, w_068_3101, w_068_3103, w_068_3104, w_068_3106, w_068_3107, w_068_3109, w_068_3111, w_068_3112, w_068_3113, w_068_3114, w_068_3119, w_068_3120, w_068_3121, w_068_3122, w_068_3125, w_068_3126, w_068_3128, w_068_3129, w_068_3130, w_068_3132, w_068_3133, w_068_3134, w_068_3135, w_068_3136, w_068_3141, w_068_3143, w_068_3144, w_068_3145, w_068_3146, w_068_3148, w_068_3149, w_068_3150, w_068_3151, w_068_3153, w_068_3155, w_068_3156, w_068_3161, w_068_3162, w_068_3164, w_068_3165, w_068_3167, w_068_3169, w_068_3173, w_068_3174, w_068_3177, w_068_3178, w_068_3180, w_068_3181, w_068_3182, w_068_3184, w_068_3185, w_068_3188, w_068_3191, w_068_3192, w_068_3193, w_068_3194, w_068_3195, w_068_3199, w_068_3201, w_068_3202, w_068_3203, w_068_3204, w_068_3205, w_068_3206, w_068_3207, w_068_3208, w_068_3210, w_068_3213, w_068_3214, w_068_3215, w_068_3216, w_068_3217, w_068_3218, w_068_3226, w_068_3227, w_068_3229, w_068_3231, w_068_3232, w_068_3233, w_068_3234, w_068_3235, w_068_3236, w_068_3237, w_068_3238, w_068_3241, w_068_3243, w_068_3244, w_068_3247, w_068_3248, w_068_3253, w_068_3255, w_068_3259, w_068_3260, w_068_3264, w_068_3268, w_068_3270, w_068_3271, w_068_3275, w_068_3276, w_068_3278, w_068_3279, w_068_3280, w_068_3281, w_068_3282, w_068_3285, w_068_3286, w_068_3287, w_068_3288, w_068_3291, w_068_3294, w_068_3295, w_068_3298, w_068_3302, w_068_3307, w_068_3309, w_068_3310, w_068_3312, w_068_3317, w_068_3318, w_068_3319, w_068_3320, w_068_3321, w_068_3323, w_068_3325, w_068_3327, w_068_3329, w_068_3332, w_068_3335, w_068_3336, w_068_3337, w_068_3338, w_068_3339, w_068_3340, w_068_3342, w_068_3343, w_068_3344, w_068_3346, w_068_3349, w_068_3350, w_068_3352, w_068_3353, w_068_3354, w_068_3360, w_068_3362, w_068_3370, w_068_3371, w_068_3372, w_068_3377, w_068_3379, w_068_3380, w_068_3381, w_068_3383, w_068_3386, w_068_3388, w_068_3393, w_068_3396, w_068_3400, w_068_3402, w_068_3404, w_068_3406, w_068_3407, w_068_3410, w_068_3411, w_068_3412, w_068_3414, w_068_3415, w_068_3420, w_068_3421, w_068_3422, w_068_3423, w_068_3424, w_068_3425, w_068_3428, w_068_3430, w_068_3431, w_068_3433, w_068_3437, w_068_3439, w_068_3440, w_068_3441, w_068_3442, w_068_3444, w_068_3448, w_068_3450, w_068_3451, w_068_3452, w_068_3453, w_068_3455, w_068_3456, w_068_3457, w_068_3458, w_068_3461, w_068_3464, w_068_3465, w_068_3466, w_068_3468, w_068_3469, w_068_3471, w_068_3472, w_068_3474, w_068_3475, w_068_3477, w_068_3478, w_068_3479, w_068_3480, w_068_3482, w_068_3486, w_068_3489, w_068_3490, w_068_3491, w_068_3493, w_068_3494, w_068_3495, w_068_3496, w_068_3497, w_068_3501, w_068_3503, w_068_3504, w_068_3505, w_068_3506, w_068_3511, w_068_3518, w_068_3524, w_068_3525, w_068_3527, w_068_3528, w_068_3529, w_068_3533, w_068_3535, w_068_3537, w_068_3539, w_068_3540, w_068_3541, w_068_3542, w_068_3543, w_068_3546, w_068_3547, w_068_3550, w_068_3553, w_068_3554, w_068_3555, w_068_3562, w_068_3563, w_068_3565, w_068_3567, w_068_3568, w_068_3569, w_068_3571, w_068_3572, w_068_3576, w_068_3577, w_068_3578, w_068_3579, w_068_3582, w_068_3583, w_068_3587, w_068_3592, w_068_3594, w_068_3601, w_068_3602, w_068_3603, w_068_3606, w_068_3607, w_068_3608, w_068_3609, w_068_3610, w_068_3613, w_068_3614, w_068_3615, w_068_3616, w_068_3618, w_068_3621, w_068_3622, w_068_3624, w_068_3627, w_068_3628, w_068_3630, w_068_3631, w_068_3632, w_068_3633, w_068_3635, w_068_3636, w_068_3639, w_068_3641, w_068_3643, w_068_3646, w_068_3647, w_068_3649, w_068_3651, w_068_3652, w_068_3653, w_068_3657, w_068_3658, w_068_3659, w_068_3661, w_068_3662, w_068_3663, w_068_3668, w_068_3671, w_068_3672, w_068_3673, w_068_3674, w_068_3676, w_068_3677, w_068_3679, w_068_3682, w_068_3685, w_068_3686, w_068_3687, w_068_3689, w_068_3690, w_068_3692, w_068_3695, w_068_3699, w_068_3700, w_068_3702, w_068_3705, w_068_3707, w_068_3708, w_068_3710, w_068_3711, w_068_3712, w_068_3714, w_068_3716, w_068_3717, w_068_3719, w_068_3721, w_068_3722, w_068_3730, w_068_3731, w_068_3734, w_068_3739, w_068_3740, w_068_3741, w_068_3743, w_068_3744, w_068_3747, w_068_3748, w_068_3749, w_068_3753, w_068_3755, w_068_3757, w_068_3758, w_068_3759, w_068_3760, w_068_3764, w_068_3765, w_068_3766, w_068_3767, w_068_3774, w_068_3775, w_068_3776, w_068_3779, w_068_3780, w_068_3782, w_068_3784, w_068_3785, w_068_3786, w_068_3789, w_068_3790, w_068_3791, w_068_3792, w_068_3794, w_068_3797, w_068_3800, w_068_3802, w_068_3803, w_068_3804, w_068_3805, w_068_3806, w_068_3810, w_068_3812, w_068_3815, w_068_3816, w_068_3817, w_068_3818, w_068_3826, w_068_3827, w_068_3828, w_068_3832, w_068_3833, w_068_3835, w_068_3836, w_068_3837, w_068_3838, w_068_3839, w_068_3841, w_068_3843, w_068_3844, w_068_3847, w_068_3849, w_068_3851, w_068_3852, w_068_3853, w_068_3855, w_068_3858, w_068_3859, w_068_3860, w_068_3864, w_068_3865, w_068_3868, w_068_3869, w_068_3870, w_068_3871, w_068_3872, w_068_3874, w_068_3875, w_068_3877, w_068_3879, w_068_3882, w_068_3883, w_068_3887, w_068_3889, w_068_3890, w_068_3891, w_068_3894, w_068_3896, w_068_3898, w_068_3899, w_068_3900, w_068_3901, w_068_3905, w_068_3907, w_068_3908, w_068_3911, w_068_3913, w_068_3916, w_068_3917, w_068_3922, w_068_3923, w_068_3927, w_068_3931, w_068_3933, w_068_3934, w_068_3936, w_068_3938, w_068_3939, w_068_3940, w_068_3941, w_068_3942, w_068_3943, w_068_3945, w_068_3946, w_068_3948, w_068_3949, w_068_3951, w_068_3952, w_068_3954, w_068_3955, w_068_3956, w_068_3957, w_068_3959, w_068_3961, w_068_3962, w_068_3963, w_068_3965, w_068_3966, w_068_3967, w_068_3969, w_068_3970, w_068_3971, w_068_3972, w_068_3973, w_068_3974, w_068_3975, w_068_3978, w_068_3979, w_068_3981, w_068_3982, w_068_3983, w_068_3984, w_068_3990, w_068_3992, w_068_3993, w_068_3995, w_068_3996, w_068_3997, w_068_4000, w_068_4002, w_068_4004, w_068_4005, w_068_4007, w_068_4008, w_068_4010, w_068_4011, w_068_4018, w_068_4023, w_068_4024, w_068_4025, w_068_4026, w_068_4028, w_068_4031, w_068_4035, w_068_4036, w_068_4037, w_068_4040, w_068_4042, w_068_4044, w_068_4045, w_068_4046, w_068_4047, w_068_4049, w_068_4050, w_068_4051, w_068_4053, w_068_4055, w_068_4060, w_068_4063, w_068_4064, w_068_4065, w_068_4066, w_068_4067, w_068_4068, w_068_4070, w_068_4071, w_068_4074, w_068_4076, w_068_4078, w_068_4079, w_068_4081, w_068_4082, w_068_4083, w_068_4084, w_068_4085, w_068_4088, w_068_4090, w_068_4093, w_068_4094, w_068_4095, w_068_4098, w_068_4099, w_068_4103, w_068_4106, w_068_4109, w_068_4112, w_068_4113, w_068_4115, w_068_4118, w_068_4121, w_068_4122, w_068_4123, w_068_4126, w_068_4129, w_068_4130, w_068_4133, w_068_4134, w_068_4135, w_068_4136, w_068_4137, w_068_4140, w_068_4141, w_068_4143, w_068_4145, w_068_4146, w_068_4147, w_068_4149, w_068_4150, w_068_4153, w_068_4155, w_068_4156, w_068_4160, w_068_4161, w_068_4162, w_068_4163, w_068_4164, w_068_4166, w_068_4172, w_068_4178, w_068_4180, w_068_4185, w_068_4187, w_068_4188, w_068_4189, w_068_4190, w_068_4191, w_068_4192, w_068_4195, w_068_4197, w_068_4200, w_068_4201, w_068_4203, w_068_4205, w_068_4206, w_068_4209, w_068_4210, w_068_4215, w_068_4216, w_068_4219, w_068_4220, w_068_4223, w_068_4224, w_068_4225, w_068_4226, w_068_4227, w_068_4229, w_068_4230, w_068_4232, w_068_4237, w_068_4240, w_068_4242, w_068_4243, w_068_4244, w_068_4245, w_068_4246, w_068_4247, w_068_4248, w_068_4251, w_068_4256, w_068_4260, w_068_4263, w_068_4264, w_068_4265, w_068_4266, w_068_4270, w_068_4272, w_068_4273, w_068_4274, w_068_4276, w_068_4277, w_068_4279, w_068_4280, w_068_4281, w_068_4287, w_068_4289, w_068_4290, w_068_4294, w_068_4295, w_068_4297, w_068_4299, w_068_4301, w_068_4302, w_068_4303, w_068_4305, w_068_4306, w_068_4308, w_068_4310, w_068_4311, w_068_4312, w_068_4313, w_068_4314, w_068_4315, w_068_4317, w_068_4319, w_068_4320, w_068_4324, w_068_4327, w_068_4332, w_068_4333, w_068_4338, w_068_4340, w_068_4341, w_068_4342, w_068_4343, w_068_4344, w_068_4345, w_068_4346, w_068_4348, w_068_4349, w_068_4351, w_068_4352, w_068_4353, w_068_4355, w_068_4356, w_068_4357, w_068_4359, w_068_4362, w_068_4364, w_068_4365, w_068_4367, w_068_4368, w_068_4369, w_068_4370, w_068_4373, w_068_4375, w_068_4376, w_068_4377, w_068_4379, w_068_4380, w_068_4381, w_068_4382, w_068_4383, w_068_4386, w_068_4387, w_068_4388, w_068_4389, w_068_4391, w_068_4392, w_068_4393, w_068_4394, w_068_4395, w_068_4396, w_068_4397, w_068_4398, w_068_4399, w_068_4400, w_068_4402, w_068_4403, w_068_4404, w_068_4408, w_068_4409, w_068_4410, w_068_4412, w_068_4413, w_068_4414, w_068_4415, w_068_4416, w_068_4418, w_068_4419, w_068_4420, w_068_4422, w_068_4423, w_068_4426, w_068_4428, w_068_4431, w_068_4432, w_068_4433, w_068_4437, w_068_4438, w_068_4440, w_068_4441, w_068_4442, w_068_4444, w_068_4445, w_068_4446, w_068_4448, w_068_4449, w_068_4450, w_068_4451, w_068_4452, w_068_4457, w_068_4462, w_068_4463, w_068_4464, w_068_4466, w_068_4472, w_068_4475, w_068_4476, w_068_4477, w_068_4480, w_068_4482, w_068_4485, w_068_4486, w_068_4489, w_068_4491, w_068_4492, w_068_4496, w_068_4497, w_068_4500, w_068_4503, w_068_4504, w_068_4507, w_068_4508, w_068_4510, w_068_4511, w_068_4512, w_068_4514, w_068_4515, w_068_4516, w_068_4517, w_068_4522, w_068_4523, w_068_4524, w_068_4526, w_068_4530, w_068_4531, w_068_4533, w_068_4534, w_068_4536, w_068_4537, w_068_4540, w_068_4542, w_068_4543, w_068_4544, w_068_4550, w_068_4551, w_068_4555, w_068_4556, w_068_4557, w_068_4558, w_068_4559, w_068_4561, w_068_4562, w_068_4564, w_068_4565, w_068_4566, w_068_4567, w_068_4569, w_068_4570, w_068_4571, w_068_4572, w_068_4573, w_068_4574, w_068_4575, w_068_4576, w_068_4577, w_068_4578, w_068_4582, w_068_4583, w_068_4587, w_068_4591, w_068_4592, w_068_4593, w_068_4594, w_068_4595, w_068_4596, w_068_4597, w_068_4598, w_068_4601, w_068_4602, w_068_4603, w_068_4611, w_068_4612, w_068_4613, w_068_4616, w_068_4620, w_068_4622, w_068_4624, w_068_4625, w_068_4626, w_068_4627, w_068_4629, w_068_4634, w_068_4635, w_068_4636, w_068_4637, w_068_4640, w_068_4642, w_068_4645, w_068_4646, w_068_4648, w_068_4650, w_068_4651, w_068_4652, w_068_4653, w_068_4654, w_068_4655, w_068_4656, w_068_4658, w_068_4663, w_068_4666, w_068_4668, w_068_4669, w_068_4671, w_068_4672, w_068_4673, w_068_4675, w_068_4676, w_068_4678, w_068_4679, w_068_4682, w_068_4683, w_068_4684, w_068_4688, w_068_4692, w_068_4693, w_068_4694, w_068_4696, w_068_4700, w_068_4702, w_068_4703, w_068_4704, w_068_4705, w_068_4707, w_068_4709, w_068_4710, w_068_4711, w_068_4717, w_068_4718, w_068_4719, w_068_4721, w_068_4724, w_068_4726, w_068_4729, w_068_4731, w_068_4733, w_068_4734, w_068_4740, w_068_4743, w_068_4745, w_068_4749, w_068_4750, w_068_4751, w_068_4753, w_068_4754, w_068_4755, w_068_4756, w_068_4759, w_068_4760, w_068_4767, w_068_4769, w_068_4773, w_068_4779, w_068_4787, w_068_4791, w_068_4794, w_068_4801, w_068_4802, w_068_4804, w_068_4806, w_068_4808, w_068_4809, w_068_4810, w_068_4811, w_068_4817, w_068_4820, w_068_4825, w_068_4828, w_068_4829, w_068_4830, w_068_4831, w_068_4833, w_068_4835, w_068_4838, w_068_4839, w_068_4844, w_068_4846, w_068_4847, w_068_4848, w_068_4850, w_068_4855, w_068_4860, w_068_4861, w_068_4862, w_068_4863, w_068_4864, w_068_4865, w_068_4870, w_068_4871, w_068_4875, w_068_4876, w_068_4877, w_068_4888, w_068_4889, w_068_4890, w_068_4892, w_068_4898, w_068_4899, w_068_4905, w_068_4916, w_068_4919, w_068_4923, w_068_4925, w_068_4927, w_068_4929, w_068_4930, w_068_4931, w_068_4936, w_068_4937, w_068_4942, w_068_4943, w_068_4952, w_068_4955, w_068_4957, w_068_4961, w_068_4963, w_068_4965, w_068_4966, w_068_4968, w_068_4970, w_068_4973, w_068_4975, w_068_4981, w_068_4982, w_068_5001, w_068_5003, w_068_5007, w_068_5009, w_068_5010, w_068_5013, w_068_5014, w_068_5018, w_068_5019, w_068_5021, w_068_5024, w_068_5034, w_068_5044, w_068_5045, w_068_5047, w_068_5048, w_068_5052, w_068_5053, w_068_5054, w_068_5059, w_068_5060, w_068_5061, w_068_5062, w_068_5065, w_068_5067, w_068_5068, w_068_5071, w_068_5072, w_068_5077, w_068_5078, w_068_5081, w_068_5082, w_068_5083, w_068_5084, w_068_5085, w_068_5088, w_068_5093, w_068_5094, w_068_5100, w_068_5104, w_068_5108, w_068_5115, w_068_5116, w_068_5118, w_068_5122, w_068_5124, w_068_5125, w_068_5129, w_068_5130, w_068_5132, w_068_5135, w_068_5137, w_068_5138, w_068_5150, w_068_5158, w_068_5166, w_068_5171, w_068_5177, w_068_5180, w_068_5181, w_068_5184, w_068_5185, w_068_5191, w_068_5196, w_068_5202, w_068_5203, w_068_5205, w_068_5206, w_068_5207, w_068_5210, w_068_5213, w_068_5214, w_068_5218, w_068_5220, w_068_5228, w_068_5231, w_068_5232, w_068_5237, w_068_5241, w_068_5253, w_068_5254, w_068_5255, w_068_5256, w_068_5264, w_068_5273, w_068_5276, w_068_5278, w_068_5282, w_068_5283, w_068_5284, w_068_5285, w_068_5289, w_068_5290, w_068_5298, w_068_5307, w_068_5310, w_068_5311;
  wire w_069_002, w_069_004, w_069_005, w_069_006, w_069_009, w_069_011, w_069_012, w_069_016, w_069_017, w_069_018, w_069_020, w_069_021, w_069_022, w_069_025, w_069_029, w_069_030, w_069_034, w_069_036, w_069_037, w_069_039, w_069_040, w_069_041, w_069_043, w_069_044, w_069_045, w_069_046, w_069_047, w_069_048, w_069_049, w_069_051, w_069_052, w_069_053, w_069_056, w_069_057, w_069_059, w_069_064, w_069_067, w_069_069, w_069_072, w_069_074, w_069_075, w_069_078, w_069_079, w_069_080, w_069_082, w_069_084, w_069_088, w_069_089, w_069_090, w_069_093, w_069_096, w_069_097, w_069_098, w_069_100, w_069_101, w_069_102, w_069_104, w_069_106, w_069_108, w_069_109, w_069_110, w_069_113, w_069_114, w_069_115, w_069_116, w_069_118, w_069_121, w_069_122, w_069_123, w_069_124, w_069_125, w_069_126, w_069_131, w_069_133, w_069_136, w_069_137, w_069_138, w_069_139, w_069_140, w_069_143, w_069_144, w_069_148, w_069_150, w_069_152, w_069_154, w_069_157, w_069_160, w_069_161, w_069_162, w_069_163, w_069_168, w_069_169, w_069_170, w_069_172, w_069_173, w_069_174, w_069_175, w_069_176, w_069_178, w_069_180, w_069_182, w_069_183, w_069_184, w_069_188, w_069_191, w_069_194, w_069_200, w_069_201, w_069_202, w_069_203, w_069_205, w_069_206, w_069_207, w_069_208, w_069_209, w_069_210, w_069_213, w_069_214, w_069_216, w_069_217, w_069_220, w_069_222, w_069_228, w_069_229, w_069_230, w_069_231, w_069_233, w_069_236, w_069_237, w_069_238, w_069_239, w_069_241, w_069_245, w_069_246, w_069_247, w_069_250, w_069_251, w_069_252, w_069_253, w_069_255, w_069_258, w_069_259, w_069_261, w_069_262, w_069_264, w_069_266, w_069_268, w_069_270, w_069_271, w_069_272, w_069_273, w_069_275, w_069_277, w_069_280, w_069_281, w_069_282, w_069_283, w_069_284, w_069_285, w_069_287, w_069_288, w_069_290, w_069_291, w_069_292, w_069_294, w_069_296, w_069_297, w_069_298, w_069_300, w_069_303, w_069_304, w_069_305, w_069_308, w_069_310, w_069_311, w_069_312, w_069_315, w_069_319, w_069_320, w_069_321, w_069_322, w_069_325, w_069_326, w_069_327, w_069_329, w_069_332, w_069_334, w_069_338, w_069_341, w_069_342, w_069_343, w_069_344, w_069_346, w_069_347, w_069_348, w_069_351, w_069_352, w_069_355, w_069_356, w_069_357, w_069_359, w_069_360, w_069_361, w_069_362, w_069_363, w_069_364, w_069_365, w_069_366, w_069_367, w_069_368, w_069_370, w_069_371, w_069_372, w_069_373, w_069_377, w_069_379, w_069_380, w_069_381, w_069_386, w_069_389, w_069_390, w_069_391, w_069_394, w_069_396, w_069_400, w_069_401, w_069_403, w_069_405, w_069_408, w_069_409, w_069_411, w_069_412, w_069_413, w_069_416, w_069_417, w_069_418, w_069_420, w_069_421, w_069_422, w_069_423, w_069_425, w_069_426, w_069_427, w_069_428, w_069_431, w_069_434, w_069_439, w_069_441, w_069_445, w_069_446, w_069_447, w_069_448, w_069_449, w_069_450, w_069_460, w_069_461, w_069_463, w_069_465, w_069_466, w_069_467, w_069_474, w_069_480, w_069_481, w_069_482, w_069_484, w_069_485, w_069_488, w_069_489, w_069_493, w_069_494, w_069_497, w_069_499, w_069_500, w_069_501, w_069_502, w_069_507, w_069_511, w_069_512, w_069_514, w_069_516, w_069_520, w_069_522, w_069_523, w_069_526, w_069_527, w_069_529, w_069_531, w_069_532, w_069_533, w_069_536, w_069_540, w_069_545, w_069_546, w_069_547, w_069_549, w_069_550, w_069_552, w_069_554, w_069_556, w_069_557, w_069_558, w_069_559, w_069_560, w_069_563, w_069_564, w_069_566, w_069_567, w_069_569, w_069_571, w_069_574, w_069_575, w_069_576, w_069_577, w_069_578, w_069_579, w_069_581, w_069_582, w_069_583, w_069_586, w_069_587, w_069_592, w_069_594, w_069_597, w_069_598, w_069_599, w_069_600, w_069_602, w_069_603, w_069_605, w_069_606, w_069_608, w_069_609, w_069_611, w_069_612, w_069_613, w_069_614, w_069_615, w_069_620, w_069_621, w_069_622, w_069_624, w_069_626, w_069_627, w_069_628, w_069_631, w_069_632, w_069_637, w_069_638, w_069_639, w_069_640, w_069_643, w_069_649, w_069_650, w_069_651, w_069_652, w_069_653, w_069_654, w_069_655, w_069_657, w_069_658, w_069_659, w_069_660, w_069_662, w_069_663, w_069_665, w_069_666, w_069_669, w_069_670, w_069_671, w_069_672, w_069_673, w_069_675, w_069_676, w_069_677, w_069_682, w_069_685, w_069_687, w_069_688, w_069_689, w_069_691, w_069_693, w_069_694, w_069_695, w_069_696, w_069_699, w_069_700, w_069_701, w_069_703, w_069_704, w_069_705, w_069_706, w_069_710, w_069_712, w_069_713, w_069_714, w_069_715, w_069_728, w_069_730, w_069_731, w_069_738, w_069_739, w_069_742, w_069_743, w_069_745, w_069_746, w_069_748, w_069_749, w_069_752, w_069_753, w_069_758, w_069_763, w_069_764, w_069_766, w_069_771, w_069_772, w_069_775, w_069_776, w_069_778, w_069_781, w_069_782, w_069_784, w_069_786, w_069_787, w_069_789, w_069_792, w_069_795, w_069_796, w_069_798, w_069_800, w_069_801, w_069_804, w_069_807, w_069_810, w_069_811, w_069_814, w_069_818, w_069_819, w_069_822, w_069_823, w_069_824, w_069_825, w_069_826, w_069_828, w_069_830, w_069_834, w_069_835, w_069_836, w_069_837, w_069_839, w_069_840, w_069_841, w_069_842, w_069_843, w_069_845, w_069_847, w_069_848, w_069_850, w_069_851, w_069_852, w_069_853, w_069_854, w_069_855, w_069_857, w_069_860, w_069_861, w_069_862, w_069_864, w_069_865, w_069_866, w_069_868, w_069_870, w_069_871, w_069_874, w_069_875, w_069_878, w_069_883, w_069_884, w_069_887, w_069_888, w_069_889, w_069_890, w_069_891, w_069_896, w_069_897, w_069_898, w_069_899, w_069_900, w_069_904, w_069_905, w_069_906, w_069_909, w_069_913, w_069_914, w_069_920, w_069_923, w_069_924, w_069_926, w_069_929, w_069_930, w_069_931, w_069_933, w_069_934, w_069_935, w_069_938, w_069_939, w_069_940, w_069_942, w_069_943, w_069_948, w_069_951, w_069_952, w_069_953, w_069_955, w_069_956, w_069_957, w_069_958, w_069_959, w_069_960, w_069_961, w_069_962, w_069_963, w_069_965, w_069_967, w_069_970, w_069_971, w_069_973, w_069_976, w_069_977, w_069_981, w_069_985, w_069_987, w_069_988, w_069_989, w_069_991, w_069_993, w_069_995, w_069_996, w_069_997, w_069_998, w_069_1000, w_069_1002, w_069_1004, w_069_1005, w_069_1008, w_069_1009, w_069_1010, w_069_1012, w_069_1013, w_069_1014, w_069_1015, w_069_1016, w_069_1018, w_069_1019, w_069_1022, w_069_1023, w_069_1025, w_069_1028, w_069_1029, w_069_1030, w_069_1034, w_069_1038, w_069_1039, w_069_1042, w_069_1045, w_069_1047, w_069_1048, w_069_1049, w_069_1050, w_069_1052, w_069_1053, w_069_1055, w_069_1059, w_069_1060, w_069_1061, w_069_1063, w_069_1065, w_069_1072, w_069_1073, w_069_1075, w_069_1076, w_069_1077, w_069_1078, w_069_1079, w_069_1080, w_069_1085, w_069_1086, w_069_1087, w_069_1088, w_069_1090, w_069_1091, w_069_1092, w_069_1093, w_069_1094, w_069_1095, w_069_1096, w_069_1098, w_069_1099, w_069_1100, w_069_1102, w_069_1103, w_069_1106, w_069_1107, w_069_1108, w_069_1111, w_069_1113, w_069_1114, w_069_1115, w_069_1116, w_069_1117, w_069_1118, w_069_1119, w_069_1120, w_069_1122, w_069_1123, w_069_1124, w_069_1125, w_069_1127, w_069_1128, w_069_1130, w_069_1134, w_069_1135, w_069_1139, w_069_1140, w_069_1143, w_069_1145, w_069_1146, w_069_1149, w_069_1152, w_069_1153, w_069_1154, w_069_1157, w_069_1161, w_069_1163, w_069_1164, w_069_1166, w_069_1167, w_069_1168, w_069_1170, w_069_1171, w_069_1172, w_069_1173, w_069_1175, w_069_1176, w_069_1177, w_069_1178, w_069_1180, w_069_1181, w_069_1183, w_069_1186, w_069_1189, w_069_1190, w_069_1192, w_069_1193, w_069_1197, w_069_1198, w_069_1200, w_069_1203, w_069_1204, w_069_1205, w_069_1206, w_069_1207, w_069_1208, w_069_1209, w_069_1212, w_069_1214, w_069_1216, w_069_1217, w_069_1219, w_069_1220, w_069_1221, w_069_1222, w_069_1224, w_069_1226, w_069_1227, w_069_1229, w_069_1230, w_069_1232, w_069_1233, w_069_1236, w_069_1237, w_069_1238, w_069_1240, w_069_1241, w_069_1244, w_069_1246, w_069_1248, w_069_1253, w_069_1255, w_069_1256, w_069_1258, w_069_1260, w_069_1261, w_069_1263, w_069_1266, w_069_1268, w_069_1270, w_069_1274, w_069_1276, w_069_1278, w_069_1280, w_069_1281, w_069_1282, w_069_1285, w_069_1289, w_069_1290, w_069_1291, w_069_1293, w_069_1295, w_069_1297, w_069_1298, w_069_1300, w_069_1303, w_069_1304, w_069_1308, w_069_1309, w_069_1310, w_069_1311, w_069_1312, w_069_1313, w_069_1315, w_069_1316, w_069_1317, w_069_1318, w_069_1319, w_069_1320, w_069_1322, w_069_1324, w_069_1326, w_069_1329, w_069_1331, w_069_1332, w_069_1333, w_069_1334, w_069_1335, w_069_1337, w_069_1338, w_069_1340, w_069_1343, w_069_1344, w_069_1347, w_069_1349, w_069_1350, w_069_1351, w_069_1352, w_069_1355, w_069_1356, w_069_1357, w_069_1358, w_069_1359, w_069_1360, w_069_1361, w_069_1363, w_069_1364, w_069_1365, w_069_1370, w_069_1371, w_069_1373, w_069_1375, w_069_1376, w_069_1378, w_069_1379, w_069_1380, w_069_1382, w_069_1383, w_069_1387, w_069_1389, w_069_1391, w_069_1392, w_069_1394, w_069_1397, w_069_1398, w_069_1400, w_069_1402, w_069_1403, w_069_1405, w_069_1406, w_069_1408, w_069_1410, w_069_1411, w_069_1412, w_069_1414, w_069_1417, w_069_1419, w_069_1421, w_069_1422, w_069_1423, w_069_1431, w_069_1434, w_069_1435, w_069_1436, w_069_1437, w_069_1438, w_069_1439, w_069_1441, w_069_1442, w_069_1444, w_069_1445, w_069_1447, w_069_1448, w_069_1449, w_069_1450, w_069_1451, w_069_1456, w_069_1457, w_069_1460, w_069_1464, w_069_1471, w_069_1473, w_069_1476, w_069_1477, w_069_1479, w_069_1480, w_069_1481, w_069_1482, w_069_1483, w_069_1485, w_069_1488, w_069_1491, w_069_1493, w_069_1494, w_069_1495, w_069_1498, w_069_1499, w_069_1500, w_069_1501, w_069_1502, w_069_1503, w_069_1505, w_069_1507, w_069_1508, w_069_1513, w_069_1514, w_069_1517, w_069_1519, w_069_1524, w_069_1527, w_069_1529, w_069_1531, w_069_1532, w_069_1533, w_069_1536, w_069_1537, w_069_1538, w_069_1540, w_069_1542, w_069_1543, w_069_1544, w_069_1545, w_069_1546, w_069_1548, w_069_1549, w_069_1552, w_069_1559, w_069_1561, w_069_1563, w_069_1565, w_069_1568, w_069_1569, w_069_1570, w_069_1573, w_069_1574, w_069_1575, w_069_1576, w_069_1577, w_069_1578, w_069_1579, w_069_1580, w_069_1582, w_069_1583, w_069_1584, w_069_1585, w_069_1586, w_069_1587, w_069_1589, w_069_1590, w_069_1593, w_069_1596, w_069_1600, w_069_1608, w_069_1612, w_069_1613, w_069_1615, w_069_1618, w_069_1619, w_069_1622, w_069_1623, w_069_1626, w_069_1627, w_069_1628, w_069_1629, w_069_1630, w_069_1631, w_069_1633, w_069_1637, w_069_1638, w_069_1641, w_069_1642, w_069_1643, w_069_1644, w_069_1645, w_069_1647, w_069_1648, w_069_1650, w_069_1652, w_069_1655, w_069_1660, w_069_1661, w_069_1662, w_069_1664, w_069_1665, w_069_1666, w_069_1667, w_069_1668, w_069_1669, w_069_1673, w_069_1674, w_069_1675, w_069_1678, w_069_1679, w_069_1681, w_069_1684, w_069_1686, w_069_1689, w_069_1691, w_069_1693, w_069_1694, w_069_1699, w_069_1701, w_069_1702, w_069_1703, w_069_1704, w_069_1705, w_069_1706, w_069_1707, w_069_1708, w_069_1709, w_069_1711, w_069_1712, w_069_1714, w_069_1716, w_069_1719, w_069_1720, w_069_1721, w_069_1722, w_069_1724, w_069_1725, w_069_1728, w_069_1729, w_069_1730, w_069_1731, w_069_1733, w_069_1734, w_069_1735, w_069_1740, w_069_1741, w_069_1742, w_069_1745, w_069_1746, w_069_1749, w_069_1752, w_069_1753, w_069_1754, w_069_1755, w_069_1756, w_069_1757, w_069_1758, w_069_1759, w_069_1760, w_069_1761, w_069_1762, w_069_1763, w_069_1766, w_069_1768, w_069_1771, w_069_1775, w_069_1776, w_069_1777, w_069_1781, w_069_1783, w_069_1786, w_069_1787, w_069_1791, w_069_1793, w_069_1794, w_069_1797, w_069_1799, w_069_1801, w_069_1811, w_069_1813, w_069_1814, w_069_1817, w_069_1819, w_069_1820, w_069_1821, w_069_1823, w_069_1825, w_069_1826, w_069_1827, w_069_1829, w_069_1830, w_069_1832, w_069_1837, w_069_1838, w_069_1841, w_069_1845, w_069_1846, w_069_1848, w_069_1849, w_069_1852, w_069_1854, w_069_1857, w_069_1858, w_069_1859, w_069_1860, w_069_1862, w_069_1863, w_069_1864, w_069_1865, w_069_1866, w_069_1867, w_069_1868, w_069_1869, w_069_1870, w_069_1871, w_069_1874, w_069_1875, w_069_1876, w_069_1878, w_069_1880, w_069_1882, w_069_1884, w_069_1887, w_069_1889, w_069_1892, w_069_1893, w_069_1894, w_069_1895, w_069_1898, w_069_1899, w_069_1902, w_069_1904, w_069_1905, w_069_1907, w_069_1908, w_069_1910, w_069_1912, w_069_1913, w_069_1915, w_069_1918, w_069_1920, w_069_1922, w_069_1924, w_069_1925, w_069_1926, w_069_1927, w_069_1928, w_069_1929, w_069_1931, w_069_1932, w_069_1933, w_069_1934, w_069_1937, w_069_1938, w_069_1942, w_069_1946, w_069_1947, w_069_1948, w_069_1950, w_069_1951, w_069_1953, w_069_1954, w_069_1955, w_069_1958, w_069_1959, w_069_1960, w_069_1962, w_069_1965, w_069_1968, w_069_1969, w_069_1970, w_069_1971, w_069_1972, w_069_1977, w_069_1978, w_069_1983, w_069_1987, w_069_1992, w_069_1993, w_069_1994, w_069_1997, w_069_1998, w_069_2001, w_069_2002, w_069_2003, w_069_2006, w_069_2008, w_069_2010, w_069_2014, w_069_2015, w_069_2016, w_069_2019, w_069_2020, w_069_2021, w_069_2022, w_069_2023, w_069_2024, w_069_2026, w_069_2027, w_069_2028, w_069_2031, w_069_2032, w_069_2033, w_069_2034, w_069_2037, w_069_2039, w_069_2040, w_069_2041, w_069_2042, w_069_2044, w_069_2045, w_069_2047, w_069_2050, w_069_2051, w_069_2052, w_069_2055, w_069_2059, w_069_2060, w_069_2061, w_069_2062, w_069_2063, w_069_2064, w_069_2065, w_069_2066, w_069_2067, w_069_2068, w_069_2069, w_069_2070, w_069_2076, w_069_2077, w_069_2079, w_069_2080, w_069_2081, w_069_2082, w_069_2086, w_069_2090, w_069_2091, w_069_2092, w_069_2093, w_069_2094, w_069_2096, w_069_2097, w_069_2098, w_069_2099, w_069_2100, w_069_2102, w_069_2103, w_069_2108, w_069_2113, w_069_2114, w_069_2115, w_069_2116, w_069_2121, w_069_2122, w_069_2124, w_069_2125, w_069_2127, w_069_2131, w_069_2132, w_069_2133, w_069_2137, w_069_2139, w_069_2140, w_069_2141, w_069_2143, w_069_2144, w_069_2145, w_069_2147, w_069_2148, w_069_2150, w_069_2157, w_069_2158, w_069_2160, w_069_2163, w_069_2164, w_069_2165, w_069_2167, w_069_2169, w_069_2170, w_069_2175, w_069_2176, w_069_2177, w_069_2179, w_069_2185, w_069_2190, w_069_2191, w_069_2192, w_069_2193, w_069_2194, w_069_2195, w_069_2197, w_069_2198, w_069_2199, w_069_2200, w_069_2201, w_069_2202, w_069_2203, w_069_2205, w_069_2206, w_069_2208, w_069_2209, w_069_2212, w_069_2213, w_069_2214, w_069_2215, w_069_2217, w_069_2218, w_069_2220, w_069_2222, w_069_2230, w_069_2231, w_069_2234, w_069_2236, w_069_2238, w_069_2239, w_069_2240, w_069_2242, w_069_2243, w_069_2244, w_069_2246, w_069_2247, w_069_2248, w_069_2250, w_069_2251, w_069_2253, w_069_2255, w_069_2256, w_069_2257, w_069_2258, w_069_2260, w_069_2261, w_069_2262, w_069_2265, w_069_2271, w_069_2272, w_069_2273, w_069_2275, w_069_2276, w_069_2277, w_069_2281, w_069_2282, w_069_2284, w_069_2286, w_069_2291, w_069_2292, w_069_2293, w_069_2295, w_069_2296, w_069_2297, w_069_2301, w_069_2302, w_069_2305, w_069_2307, w_069_2308, w_069_2309, w_069_2311, w_069_2312, w_069_2317, w_069_2318, w_069_2319, w_069_2320, w_069_2322, w_069_2327, w_069_2328, w_069_2329, w_069_2330, w_069_2331, w_069_2332, w_069_2333, w_069_2337, w_069_2338, w_069_2339, w_069_2340, w_069_2341, w_069_2344, w_069_2348, w_069_2349, w_069_2350, w_069_2351, w_069_2355, w_069_2357, w_069_2358, w_069_2363, w_069_2364, w_069_2366, w_069_2367, w_069_2372, w_069_2373, w_069_2374, w_069_2378, w_069_2379, w_069_2380, w_069_2383, w_069_2385, w_069_2388, w_069_2390, w_069_2391, w_069_2392, w_069_2393, w_069_2394, w_069_2396, w_069_2398, w_069_2400, w_069_2401, w_069_2402, w_069_2404, w_069_2406, w_069_2408, w_069_2409, w_069_2411, w_069_2412, w_069_2419, w_069_2421, w_069_2423, w_069_2424, w_069_2425, w_069_2429, w_069_2437, w_069_2440, w_069_2443, w_069_2444, w_069_2445, w_069_2446, w_069_2447, w_069_2450, w_069_2451, w_069_2452, w_069_2453, w_069_2454, w_069_2455, w_069_2456, w_069_2457, w_069_2459, w_069_2460, w_069_2461, w_069_2462, w_069_2464, w_069_2465, w_069_2470, w_069_2472, w_069_2474, w_069_2477, w_069_2481, w_069_2482, w_069_2483, w_069_2485, w_069_2486, w_069_2487, w_069_2491, w_069_2496, w_069_2499, w_069_2501, w_069_2506, w_069_2509, w_069_2510, w_069_2514, w_069_2515, w_069_2519, w_069_2520, w_069_2523, w_069_2524, w_069_2525, w_069_2526, w_069_2527, w_069_2536, w_069_2542, w_069_2547, w_069_2549, w_069_2550, w_069_2551, w_069_2552, w_069_2553, w_069_2554, w_069_2555, w_069_2557, w_069_2559, w_069_2560, w_069_2564, w_069_2565, w_069_2567, w_069_2568, w_069_2570, w_069_2571, w_069_2572, w_069_2573, w_069_2574, w_069_2576, w_069_2579, w_069_2580, w_069_2581, w_069_2583, w_069_2584, w_069_2585, w_069_2592, w_069_2593, w_069_2595, w_069_2598, w_069_2600, w_069_2602, w_069_2605, w_069_2606, w_069_2607, w_069_2608, w_069_2609, w_069_2610, w_069_2612, w_069_2614, w_069_2615, w_069_2618, w_069_2620, w_069_2621, w_069_2622, w_069_2625, w_069_2626, w_069_2627, w_069_2629, w_069_2632, w_069_2633, w_069_2637, w_069_2638, w_069_2639, w_069_2643, w_069_2647, w_069_2648, w_069_2649, w_069_2651, w_069_2654, w_069_2655, w_069_2657, w_069_2659, w_069_2660, w_069_2661, w_069_2662, w_069_2663, w_069_2665, w_069_2668, w_069_2669, w_069_2670, w_069_2671, w_069_2672, w_069_2674, w_069_2675, w_069_2676, w_069_2677, w_069_2678, w_069_2679, w_069_2681, w_069_2682, w_069_2683, w_069_2687, w_069_2688, w_069_2689, w_069_2692, w_069_2694, w_069_2695, w_069_2696, w_069_2699, w_069_2700, w_069_2701, w_069_2702, w_069_2703, w_069_2704, w_069_2708, w_069_2712, w_069_2717, w_069_2719, w_069_2720, w_069_2722, w_069_2726, w_069_2727, w_069_2728, w_069_2730, w_069_2732, w_069_2733, w_069_2734, w_069_2735, w_069_2736, w_069_2737, w_069_2743, w_069_2745, w_069_2748, w_069_2751, w_069_2752, w_069_2753, w_069_2754, w_069_2756, w_069_2757, w_069_2758, w_069_2761, w_069_2763, w_069_2764, w_069_2766, w_069_2767, w_069_2768, w_069_2770, w_069_2772, w_069_2774, w_069_2776, w_069_2778, w_069_2779, w_069_2784, w_069_2788, w_069_2789, w_069_2795, w_069_2801, w_069_2802, w_069_2803, w_069_2804, w_069_2805, w_069_2808, w_069_2810, w_069_2813, w_069_2817, w_069_2819, w_069_2820, w_069_2821, w_069_2822, w_069_2824, w_069_2826, w_069_2827, w_069_2828, w_069_2829, w_069_2830, w_069_2835, w_069_2837, w_069_2838, w_069_2841, w_069_2842, w_069_2845, w_069_2846, w_069_2849, w_069_2850, w_069_2851, w_069_2853, w_069_2854, w_069_2858, w_069_2863, w_069_2865, w_069_2867, w_069_2869, w_069_2871, w_069_2873, w_069_2875, w_069_2876, w_069_2877, w_069_2880, w_069_2885, w_069_2887, w_069_2890, w_069_2896, w_069_2897, w_069_2898, w_069_2900, w_069_2901, w_069_2902, w_069_2903, w_069_2904, w_069_2905, w_069_2906, w_069_2907, w_069_2908, w_069_2910, w_069_2912, w_069_2920, w_069_2921, w_069_2925, w_069_2927, w_069_2931, w_069_2933, w_069_2934, w_069_2935, w_069_2936, w_069_2937, w_069_2942, w_069_2946, w_069_2947, w_069_2948, w_069_2949, w_069_2952, w_069_2954, w_069_2955, w_069_2956, w_069_2958, w_069_2967, w_069_2968, w_069_2969, w_069_2971, w_069_2975, w_069_2976, w_069_2977, w_069_2978, w_069_2979, w_069_2980, w_069_2982, w_069_2984, w_069_2987, w_069_2988, w_069_2989, w_069_2992, w_069_2994, w_069_2995, w_069_2998, w_069_2999, w_069_3001, w_069_3002, w_069_3003, w_069_3005, w_069_3006, w_069_3008, w_069_3009, w_069_3010, w_069_3013, w_069_3014, w_069_3015, w_069_3018, w_069_3021, w_069_3024, w_069_3027, w_069_3028, w_069_3029, w_069_3030, w_069_3031, w_069_3032, w_069_3034, w_069_3036, w_069_3037, w_069_3039, w_069_3041, w_069_3045, w_069_3047, w_069_3048, w_069_3053, w_069_3054, w_069_3057, w_069_3058, w_069_3059, w_069_3061, w_069_3062, w_069_3063, w_069_3064, w_069_3066, w_069_3069, w_069_3071, w_069_3074, w_069_3075, w_069_3076, w_069_3077, w_069_3078, w_069_3080, w_069_3082, w_069_3083, w_069_3084, w_069_3086, w_069_3087, w_069_3089, w_069_3090, w_069_3091, w_069_3094, w_069_3096, w_069_3097, w_069_3098, w_069_3099, w_069_3102, w_069_3103, w_069_3106, w_069_3108, w_069_3110, w_069_3111, w_069_3112, w_069_3114, w_069_3115, w_069_3116, w_069_3118, w_069_3119, w_069_3120, w_069_3121, w_069_3122, w_069_3123, w_069_3125, w_069_3126, w_069_3127, w_069_3128, w_069_3129, w_069_3130, w_069_3132, w_069_3136, w_069_3137, w_069_3138, w_069_3144, w_069_3146, w_069_3147, w_069_3150, w_069_3151, w_069_3155, w_069_3156, w_069_3159, w_069_3160, w_069_3162, w_069_3169, w_069_3173, w_069_3176, w_069_3177, w_069_3179, w_069_3180, w_069_3181, w_069_3182, w_069_3184, w_069_3185, w_069_3186, w_069_3188, w_069_3189, w_069_3190, w_069_3193, w_069_3194, w_069_3196, w_069_3197, w_069_3198, w_069_3199, w_069_3203, w_069_3204, w_069_3205, w_069_3207, w_069_3208, w_069_3209, w_069_3211, w_069_3212, w_069_3213, w_069_3214, w_069_3216, w_069_3217, w_069_3224, w_069_3226, w_069_3230, w_069_3231, w_069_3232, w_069_3235, w_069_3236, w_069_3237, w_069_3239, w_069_3241, w_069_3242, w_069_3243, w_069_3245, w_069_3247, w_069_3248, w_069_3250, w_069_3254, w_069_3258, w_069_3261, w_069_3262, w_069_3263, w_069_3266, w_069_3267, w_069_3269, w_069_3270, w_069_3272, w_069_3273, w_069_3274, w_069_3275, w_069_3277, w_069_3281, w_069_3283, w_069_3284, w_069_3285, w_069_3287, w_069_3288, w_069_3291, w_069_3292, w_069_3293, w_069_3297, w_069_3298, w_069_3299, w_069_3300, w_069_3303, w_069_3305, w_069_3306, w_069_3308, w_069_3309, w_069_3311, w_069_3313, w_069_3314, w_069_3316, w_069_3321, w_069_3324, w_069_3325, w_069_3327, w_069_3329, w_069_3332, w_069_3335, w_069_3337, w_069_3339, w_069_3341, w_069_3342, w_069_3343, w_069_3345, w_069_3347, w_069_3350, w_069_3354, w_069_3355, w_069_3357, w_069_3362, w_069_3366, w_069_3368, w_069_3369, w_069_3370, w_069_3371, w_069_3372, w_069_3373, w_069_3374, w_069_3375, w_069_3376, w_069_3377, w_069_3380, w_069_3381, w_069_3385, w_069_3386, w_069_3387, w_069_3388, w_069_3391, w_069_3392, w_069_3395, w_069_3397, w_069_3398, w_069_3399, w_069_3400, w_069_3402, w_069_3404, w_069_3405, w_069_3406, w_069_3407, w_069_3409, w_069_3410, w_069_3412, w_069_3414, w_069_3417, w_069_3419, w_069_3420, w_069_3422, w_069_3424, w_069_3425, w_069_3426, w_069_3427, w_069_3428, w_069_3429, w_069_3434, w_069_3435, w_069_3436, w_069_3437, w_069_3438, w_069_3439, w_069_3441, w_069_3442, w_069_3443, w_069_3445, w_069_3446, w_069_3447, w_069_3449, w_069_3453, w_069_3456, w_069_3458, w_069_3461, w_069_3462, w_069_3464, w_069_3466, w_069_3467, w_069_3468, w_069_3470, w_069_3471, w_069_3474, w_069_3477, w_069_3478, w_069_3479, w_069_3485, w_069_3486, w_069_3489, w_069_3491, w_069_3492, w_069_3496, w_069_3497, w_069_3498, w_069_3499, w_069_3500, w_069_3501, w_069_3502, w_069_3504, w_069_3505, w_069_3507, w_069_3509, w_069_3510, w_069_3514, w_069_3516, w_069_3518, w_069_3519, w_069_3520, w_069_3521, w_069_3522, w_069_3524, w_069_3526, w_069_3528, w_069_3529, w_069_3533, w_069_3534, w_069_3538, w_069_3539, w_069_3540, w_069_3542, w_069_3543, w_069_3545, w_069_3546, w_069_3548, w_069_3549, w_069_3550, w_069_3551, w_069_3554, w_069_3556, w_069_3558, w_069_3559, w_069_3561, w_069_3563, w_069_3564, w_069_3569, w_069_3573, w_069_3576, w_069_3578, w_069_3579, w_069_3582, w_069_3583, w_069_3585, w_069_3586, w_069_3587, w_069_3588, w_069_3589, w_069_3590, w_069_3592, w_069_3597, w_069_3598, w_069_3601, w_069_3602, w_069_3603, w_069_3604, w_069_3605, w_069_3606, w_069_3608, w_069_3612, w_069_3613, w_069_3614, w_069_3616, w_069_3617, w_069_3618, w_069_3619, w_069_3624, w_069_3625, w_069_3626, w_069_3628, w_069_3629, w_069_3631, w_069_3633, w_069_3634, w_069_3638, w_069_3639, w_069_3641, w_069_3645, w_069_3647, w_069_3648, w_069_3650, w_069_3652, w_069_3653, w_069_3655, w_069_3657, w_069_3660, w_069_3662, w_069_3663, w_069_3664, w_069_3665, w_069_3666, w_069_3667, w_069_3671, w_069_3673, w_069_3676, w_069_3677, w_069_3678, w_069_3680, w_069_3682, w_069_3683, w_069_3684, w_069_3687, w_069_3691, w_069_3692, w_069_3694, w_069_3696, w_069_3697, w_069_3698, w_069_3700, w_069_3703, w_069_3704, w_069_3707, w_069_3709, w_069_3711, w_069_3712, w_069_3715, w_069_3718, w_069_3722, w_069_3723, w_069_3725, w_069_3726, w_069_3727, w_069_3730, w_069_3733, w_069_3734, w_069_3737, w_069_3738, w_069_3740, w_069_3743, w_069_3745, w_069_3748, w_069_3749, w_069_3750, w_069_3752, w_069_3753, w_069_3755, w_069_3756, w_069_3757, w_069_3759, w_069_3762, w_069_3764, w_069_3765, w_069_3767, w_069_3768, w_069_3770, w_069_3771, w_069_3776, w_069_3780, w_069_3784, w_069_3786, w_069_3787, w_069_3789, w_069_3790, w_069_3793, w_069_3794, w_069_3797, w_069_3798, w_069_3800, w_069_3801, w_069_3804, w_069_3805, w_069_3807, w_069_3809, w_069_3811, w_069_3813, w_069_3816, w_069_3824, w_069_3826, w_069_3830, w_069_3832, w_069_3834, w_069_3835, w_069_3838, w_069_3840, w_069_3841, w_069_3851, w_069_3853, w_069_3856, w_069_3857, w_069_3860, w_069_3863, w_069_3866, w_069_3871, w_069_3877, w_069_3884, w_069_3885, w_069_3886, w_069_3888, w_069_3889, w_069_3890, w_069_3894, w_069_3896, w_069_3897, w_069_3898, w_069_3900, w_069_3902, w_069_3906, w_069_3907, w_069_3908, w_069_3910, w_069_3911, w_069_3912, w_069_3913, w_069_3915, w_069_3917, w_069_3920, w_069_3924, w_069_3927, w_069_3929, w_069_3936, w_069_3944, w_069_3947, w_069_3948, w_069_3954, w_069_3955, w_069_3960, w_069_3964, w_069_3965, w_069_3966, w_069_3967, w_069_3970, w_069_3971, w_069_3978, w_069_3981, w_069_3982, w_069_3984, w_069_3986, w_069_3987, w_069_3990, w_069_3991, w_069_3994, w_069_3995, w_069_3996, w_069_3998, w_069_4000, w_069_4003, w_069_4004, w_069_4005, w_069_4013, w_069_4015, w_069_4020, w_069_4021, w_069_4024, w_069_4027, w_069_4031, w_069_4037, w_069_4038, w_069_4042, w_069_4051, w_069_4062, w_069_4064, w_069_4065, w_069_4067, w_069_4069, w_069_4070, w_069_4072, w_069_4078, w_069_4081, w_069_4082, w_069_4088, w_069_4093, w_069_4096, w_069_4100, w_069_4102, w_069_4111, w_069_4113, w_069_4116, w_069_4118, w_069_4127, w_069_4128, w_069_4129, w_069_4132, w_069_4134, w_069_4136, w_069_4137, w_069_4143, w_069_4144, w_069_4146, w_069_4149, w_069_4152, w_069_4155, w_069_4159, w_069_4161, w_069_4162, w_069_4165, w_069_4168, w_069_4170, w_069_4171, w_069_4172, w_069_4173, w_069_4176, w_069_4180, w_069_4184, w_069_4187, w_069_4189, w_069_4190, w_069_4192, w_069_4207, w_069_4210, w_069_4214, w_069_4220, w_069_4221, w_069_4223, w_069_4224, w_069_4225, w_069_4228, w_069_4238, w_069_4240, w_069_4242, w_069_4244, w_069_4249, w_069_4250, w_069_4252, w_069_4253, w_069_4254, w_069_4255, w_069_4256, w_069_4257, w_069_4260, w_069_4268, w_069_4271, w_069_4273, w_069_4275, w_069_4277, w_069_4281, w_069_4283, w_069_4291, w_069_4292, w_069_4297, w_069_4302, w_069_4310, w_069_4311, w_069_4315, w_069_4318, w_069_4320, w_069_4324, w_069_4326, w_069_4336, w_069_4341, w_069_4342, w_069_4344, w_069_4346, w_069_4349, w_069_4352, w_069_4362, w_069_4371, w_069_4372, w_069_4376, w_069_4377, w_069_4380, w_069_4385, w_069_4388, w_069_4389, w_069_4390, w_069_4391, w_069_4393, w_069_4394, w_069_4405, w_069_4407, w_069_4408, w_069_4410, w_069_4411, w_069_4414, w_069_4415, w_069_4416, w_069_4418, w_069_4422, w_069_4425, w_069_4428, w_069_4434, w_069_4435, w_069_4444, w_069_4449, w_069_4450, w_069_4452, w_069_4460, w_069_4461, w_069_4463, w_069_4467, w_069_4468, w_069_4472, w_069_4473, w_069_4476, w_069_4477, w_069_4478, w_069_4479, w_069_4481, w_069_4482, w_069_4483, w_069_4485, w_069_4490, w_069_4491, w_069_4492, w_069_4493, w_069_4497, w_069_4504, w_069_4506, w_069_4507, w_069_4508, w_069_4512, w_069_4513, w_069_4514, w_069_4516, w_069_4531, w_069_4540, w_069_4542, w_069_4543, w_069_4544, w_069_4545, w_069_4550, w_069_4551, w_069_4552, w_069_4553, w_069_4554, w_069_4555, w_069_4559, w_069_4563, w_069_4565, w_069_4566, w_069_4567, w_069_4571, w_069_4573, w_069_4575, w_069_4576, w_069_4579, w_069_4580, w_069_4591, w_069_4595, w_069_4599, w_069_4602, w_069_4609, w_069_4611, w_069_4613, w_069_4616, w_069_4617, w_069_4618, w_069_4619, w_069_4620, w_069_4623, w_069_4626, w_069_4629, w_069_4639, w_069_4640, w_069_4641, w_069_4642, w_069_4645, w_069_4647, w_069_4649, w_069_4654, w_069_4655, w_069_4658, w_069_4660, w_069_4662, w_069_4664, w_069_4668, w_069_4671, w_069_4675, w_069_4681, w_069_4683, w_069_4684, w_069_4686, w_069_4689, w_069_4690, w_069_4691, w_069_4692, w_069_4693, w_069_4694, w_069_4699, w_069_4700, w_069_4704, w_069_4705, w_069_4706, w_069_4707, w_069_4710, w_069_4713, w_069_4714, w_069_4717, w_069_4721, w_069_4723, w_069_4724, w_069_4725, w_069_4728, w_069_4729, w_069_4734, w_069_4737, w_069_4744, w_069_4752, w_069_4754, w_069_4760, w_069_4761, w_069_4763, w_069_4765, w_069_4778, w_069_4781, w_069_4782, w_069_4783, w_069_4787, w_069_4793, w_069_4796, w_069_4802, w_069_4808, w_069_4809, w_069_4811, w_069_4812, w_069_4813, w_069_4815, w_069_4816, w_069_4822, w_069_4823, w_069_4825, w_069_4826, w_069_4829, w_069_4831, w_069_4840, w_069_4847, w_069_4848, w_069_4849, w_069_4851, w_069_4852, w_069_4854, w_069_4857, w_069_4860, w_069_4862, w_069_4867, w_069_4871, w_069_4873, w_069_4877, w_069_4883, w_069_4892, w_069_4893, w_069_4894, w_069_4896, w_069_4902, w_069_4903, w_069_4907, w_069_4921, w_069_4924, w_069_4928, w_069_4929, w_069_4930, w_069_4933, w_069_4937, w_069_4941, w_069_4946, w_069_4947, w_069_4948, w_069_4950, w_069_4952, w_069_4956, w_069_4963, w_069_4967, w_069_4970, w_069_4971, w_069_4973, w_069_4974, w_069_4978, w_069_4979, w_069_4985, w_069_4988, w_069_4989, w_069_4990, w_069_4991, w_069_4993, w_069_4996, w_069_4998, w_069_5002, w_069_5004, w_069_5005, w_069_5017, w_069_5026, w_069_5027, w_069_5028, w_069_5034, w_069_5037, w_069_5042, w_069_5044, w_069_5046, w_069_5047, w_069_5048, w_069_5052, w_069_5053, w_069_5058, w_069_5067, w_069_5073, w_069_5078, w_069_5085, w_069_5089, w_069_5091, w_069_5094, w_069_5095, w_069_5097, w_069_5103, w_069_5113, w_069_5117, w_069_5123, w_069_5127, w_069_5129, w_069_5130, w_069_5132, w_069_5133, w_069_5134, w_069_5137, w_069_5140, w_069_5144, w_069_5145, w_069_5146, w_069_5148, w_069_5150, w_069_5153, w_069_5154, w_069_5156, w_069_5161, w_069_5164, w_069_5166, w_069_5173, w_069_5174, w_069_5178, w_069_5184, w_069_5186, w_069_5194, w_069_5195, w_069_5200, w_069_5201, w_069_5209, w_069_5210, w_069_5228, w_069_5230, w_069_5235, w_069_5237, w_069_5243, w_069_5245, w_069_5250, w_069_5251, w_069_5254, w_069_5255, w_069_5258, w_069_5259, w_069_5260, w_069_5262, w_069_5264, w_069_5266, w_069_5272, w_069_5274, w_069_5278, w_069_5281, w_069_5283, w_069_5289, w_069_5290, w_069_5295, w_069_5298, w_069_5301, w_069_5304, w_069_5312, w_069_5318, w_069_5321, w_069_5323, w_069_5325, w_069_5330, w_069_5337, w_069_5338, w_069_5346, w_069_5351, w_069_5353, w_069_5358, w_069_5360, w_069_5372, w_069_5375, w_069_5377, w_069_5378, w_069_5379, w_069_5386, w_069_5388, w_069_5390, w_069_5392, w_069_5393, w_069_5394, w_069_5401, w_069_5406, w_069_5412, w_069_5413, w_069_5419, w_069_5420, w_069_5421, w_069_5427, w_069_5429, w_069_5438, w_069_5447, w_069_5449, w_069_5450, w_069_5451, w_069_5456, w_069_5458, w_069_5460, w_069_5461, w_069_5462, w_069_5471, w_069_5477, w_069_5479, w_069_5481, w_069_5484, w_069_5485, w_069_5486, w_069_5488, w_069_5492, w_069_5494, w_069_5496, w_069_5497, w_069_5498, w_069_5501, w_069_5502, w_069_5504, w_069_5506, w_069_5507, w_069_5510, w_069_5516, w_069_5517, w_069_5522, w_069_5525, w_069_5526, w_069_5529, w_069_5532, w_069_5534, w_069_5535, w_069_5536, w_069_5537, w_069_5538, w_069_5545, w_069_5546, w_069_5553, w_069_5555, w_069_5562, w_069_5566, w_069_5569, w_069_5570, w_069_5573, w_069_5576, w_069_5577, w_069_5579, w_069_5581, w_069_5583, w_069_5587, w_069_5592, w_069_5594, w_069_5599, w_069_5603, w_069_5606, w_069_5607, w_069_5615, w_069_5617, w_069_5619, w_069_5624, w_069_5625, w_069_5631, w_069_5632, w_069_5636, w_069_5639, w_069_5640, w_069_5643, w_069_5645, w_069_5649, w_069_5651, w_069_5654, w_069_5660, w_069_5661, w_069_5664, w_069_5668, w_069_5669, w_069_5671, w_069_5679, w_069_5682, w_069_5684, w_069_5693, w_069_5694, w_069_5697, w_069_5702, w_069_5705, w_069_5707, w_069_5709, w_069_5712, w_069_5713, w_069_5722, w_069_5725, w_069_5728, w_069_5729, w_069_5741, w_069_5746, w_069_5749, w_069_5751, w_069_5755, w_069_5756, w_069_5759, w_069_5764, w_069_5765, w_069_5768, w_069_5769, w_069_5770, w_069_5771, w_069_5772, w_069_5773, w_069_5776, w_069_5777, w_069_5782, w_069_5783, w_069_5792, w_069_5793, w_069_5795, w_069_5806, w_069_5809, w_069_5815, w_069_5816, w_069_5817, w_069_5820, w_069_5825, w_069_5838, w_069_5844, w_069_5850, w_069_5852, w_069_5859, w_069_5864, w_069_5874, w_069_5878, w_069_5881, w_069_5882, w_069_5883, w_069_5884, w_069_5885, w_069_5891, w_069_5893, w_069_5894, w_069_5896, w_069_5897, w_069_5898, w_069_5899, w_069_5901, w_069_5902, w_069_5904, w_069_5910, w_069_5920, w_069_5924, w_069_5926, w_069_5931, w_069_5933, w_069_5939, w_069_5940, w_069_5945, w_069_5949, w_069_5951, w_069_5952, w_069_5953, w_069_5956, w_069_5961, w_069_5962, w_069_5964, w_069_5965, w_069_5970, w_069_5971, w_069_5973, w_069_5984, w_069_5987, w_069_5990, w_069_5995, w_069_6001, w_069_6002, w_069_6003, w_069_6004, w_069_6008, w_069_6010, w_069_6011, w_069_6016, w_069_6017, w_069_6022, w_069_6024, w_069_6025, w_069_6027, w_069_6028, w_069_6029, w_069_6031, w_069_6032, w_069_6034, w_069_6037, w_069_6043, w_069_6044, w_069_6051, w_069_6052, w_069_6054, w_069_6059, w_069_6063, w_069_6066, w_069_6068, w_069_6070, w_069_6075, w_069_6079, w_069_6082, w_069_6083, w_069_6086, w_069_6087, w_069_6091, w_069_6093, w_069_6097, w_069_6101, w_069_6102, w_069_6105, w_069_6107, w_069_6108, w_069_6109, w_069_6113, w_069_6116, w_069_6120, w_069_6123, w_069_6127, w_069_6131, w_069_6132, w_069_6133, w_069_6135, w_069_6138, w_069_6142, w_069_6147, w_069_6153, w_069_6159, w_069_6162, w_069_6166, w_069_6168, w_069_6169, w_069_6170, w_069_6171, w_069_6179, w_069_6181, w_069_6184, w_069_6189, w_069_6192;
  wire w_070_000, w_070_002, w_070_004, w_070_005, w_070_007, w_070_010, w_070_011, w_070_012, w_070_013, w_070_015, w_070_020, w_070_023, w_070_024, w_070_025, w_070_028, w_070_030, w_070_031, w_070_033, w_070_034, w_070_035, w_070_036, w_070_038, w_070_040, w_070_042, w_070_044, w_070_047, w_070_049, w_070_051, w_070_052, w_070_054, w_070_061, w_070_062, w_070_064, w_070_065, w_070_066, w_070_068, w_070_069, w_070_070, w_070_073, w_070_078, w_070_079, w_070_081, w_070_083, w_070_084, w_070_086, w_070_090, w_070_091, w_070_092, w_070_093, w_070_096, w_070_097, w_070_098, w_070_099, w_070_100, w_070_101, w_070_106, w_070_107, w_070_109, w_070_111, w_070_117, w_070_120, w_070_122, w_070_125, w_070_126, w_070_127, w_070_129, w_070_131, w_070_137, w_070_138, w_070_139, w_070_140, w_070_142, w_070_148, w_070_149, w_070_151, w_070_152, w_070_153, w_070_155, w_070_156, w_070_157, w_070_158, w_070_159, w_070_161, w_070_164, w_070_166, w_070_168, w_070_169, w_070_170, w_070_171, w_070_172, w_070_173, w_070_176, w_070_180, w_070_181, w_070_185, w_070_186, w_070_187, w_070_188, w_070_191, w_070_193, w_070_194, w_070_195, w_070_196, w_070_197, w_070_198, w_070_199, w_070_200, w_070_204, w_070_205, w_070_206, w_070_207, w_070_209, w_070_211, w_070_213, w_070_214, w_070_215, w_070_218, w_070_219, w_070_221, w_070_222, w_070_224, w_070_225, w_070_229, w_070_230, w_070_233, w_070_234, w_070_236, w_070_237, w_070_239, w_070_241, w_070_242, w_070_243, w_070_244, w_070_247, w_070_250, w_070_251, w_070_252, w_070_253, w_070_254, w_070_255, w_070_256, w_070_257, w_070_258, w_070_259, w_070_260, w_070_261, w_070_263, w_070_265, w_070_268, w_070_271, w_070_272, w_070_273, w_070_274, w_070_275, w_070_277, w_070_280, w_070_281, w_070_290, w_070_293, w_070_297, w_070_298, w_070_300, w_070_302, w_070_305, w_070_306, w_070_309, w_070_310, w_070_311, w_070_312, w_070_316, w_070_317, w_070_319, w_070_321, w_070_323, w_070_325, w_070_329, w_070_331, w_070_332, w_070_334, w_070_335, w_070_338, w_070_339, w_070_342, w_070_344, w_070_347, w_070_350, w_070_353, w_070_358, w_070_359, w_070_361, w_070_364, w_070_365, w_070_367, w_070_371, w_070_372, w_070_373, w_070_375, w_070_379, w_070_380, w_070_381, w_070_383, w_070_384, w_070_386, w_070_387, w_070_388, w_070_390, w_070_392, w_070_394, w_070_397, w_070_399, w_070_406, w_070_408, w_070_410, w_070_411, w_070_412, w_070_413, w_070_415, w_070_416, w_070_418, w_070_419, w_070_421, w_070_423, w_070_427, w_070_428, w_070_429, w_070_430, w_070_432, w_070_433, w_070_434, w_070_437, w_070_439, w_070_440, w_070_442, w_070_443, w_070_444, w_070_445, w_070_447, w_070_448, w_070_454, w_070_459, w_070_461, w_070_462, w_070_463, w_070_464, w_070_465, w_070_468, w_070_469, w_070_470, w_070_471, w_070_472, w_070_473, w_070_474, w_070_477, w_070_478, w_070_480, w_070_482, w_070_485, w_070_491, w_070_493, w_070_495, w_070_496, w_070_497, w_070_498, w_070_499, w_070_500, w_070_503, w_070_504, w_070_505, w_070_506, w_070_507, w_070_510, w_070_515, w_070_516, w_070_517, w_070_518, w_070_519, w_070_520, w_070_522, w_070_523, w_070_527, w_070_528, w_070_530, w_070_533, w_070_534, w_070_536, w_070_537, w_070_538, w_070_539, w_070_546, w_070_549, w_070_551, w_070_553, w_070_556, w_070_561, w_070_562, w_070_565, w_070_570, w_070_571, w_070_574, w_070_575, w_070_577, w_070_578, w_070_579, w_070_580, w_070_582, w_070_583, w_070_584, w_070_586, w_070_587, w_070_589, w_070_591, w_070_595, w_070_597, w_070_598, w_070_599, w_070_600, w_070_605, w_070_607, w_070_609, w_070_611, w_070_614, w_070_617, w_070_618, w_070_619, w_070_621, w_070_622, w_070_624, w_070_626, w_070_629, w_070_630, w_070_632, w_070_634, w_070_636, w_070_638, w_070_639, w_070_640, w_070_642, w_070_644, w_070_648, w_070_653, w_070_657, w_070_658, w_070_665, w_070_667, w_070_668, w_070_669, w_070_671, w_070_672, w_070_673, w_070_674, w_070_675, w_070_677, w_070_678, w_070_681, w_070_682, w_070_683, w_070_684, w_070_686, w_070_687, w_070_688, w_070_689, w_070_690, w_070_691, w_070_695, w_070_696, w_070_697, w_070_700, w_070_701, w_070_703, w_070_704, w_070_706, w_070_707, w_070_708, w_070_709, w_070_710, w_070_711, w_070_715, w_070_716, w_070_717, w_070_719, w_070_720, w_070_727, w_070_728, w_070_729, w_070_737, w_070_738, w_070_739, w_070_741, w_070_742, w_070_743, w_070_745, w_070_746, w_070_747, w_070_749, w_070_750, w_070_751, w_070_752, w_070_757, w_070_758, w_070_759, w_070_762, w_070_763, w_070_764, w_070_765, w_070_766, w_070_768, w_070_769, w_070_770, w_070_771, w_070_773, w_070_774, w_070_775, w_070_778, w_070_779, w_070_780, w_070_781, w_070_784, w_070_786, w_070_788, w_070_790, w_070_791, w_070_792, w_070_793, w_070_794, w_070_795, w_070_796, w_070_797, w_070_798, w_070_799, w_070_801, w_070_803, w_070_804, w_070_808, w_070_809, w_070_810, w_070_811, w_070_813, w_070_815, w_070_819, w_070_820, w_070_821, w_070_822, w_070_829, w_070_833, w_070_834, w_070_835, w_070_840, w_070_842, w_070_843, w_070_845, w_070_850, w_070_851, w_070_855, w_070_856, w_070_857, w_070_860, w_070_861, w_070_862, w_070_865, w_070_866, w_070_867, w_070_872, w_070_875, w_070_876, w_070_878, w_070_880, w_070_883, w_070_886, w_070_888, w_070_889, w_070_890, w_070_891, w_070_892, w_070_894, w_070_895, w_070_896, w_070_897, w_070_899, w_070_901, w_070_902, w_070_903, w_070_907, w_070_910, w_070_913, w_070_920, w_070_924, w_070_928, w_070_929, w_070_930, w_070_931, w_070_932, w_070_933, w_070_935, w_070_936, w_070_938, w_070_939, w_070_941, w_070_942, w_070_946, w_070_947, w_070_949, w_070_950, w_070_951, w_070_952, w_070_954, w_070_956, w_070_957, w_070_960, w_070_961, w_070_965, w_070_967, w_070_968, w_070_969, w_070_971, w_070_976, w_070_977, w_070_978, w_070_980, w_070_982, w_070_983, w_070_984, w_070_986, w_070_988, w_070_989, w_070_992, w_070_994, w_070_999, w_070_1000, w_070_1002, w_070_1003, w_070_1004, w_070_1007, w_070_1008, w_070_1015, w_070_1016, w_070_1017, w_070_1019, w_070_1022, w_070_1025, w_070_1029, w_070_1030, w_070_1033, w_070_1034, w_070_1035, w_070_1037, w_070_1046, w_070_1048, w_070_1049, w_070_1050, w_070_1054, w_070_1059, w_070_1060, w_070_1062, w_070_1063, w_070_1064, w_070_1066, w_070_1068, w_070_1071, w_070_1075, w_070_1076, w_070_1078, w_070_1079, w_070_1081, w_070_1082, w_070_1083, w_070_1085, w_070_1090, w_070_1091, w_070_1092, w_070_1093, w_070_1094, w_070_1095, w_070_1098, w_070_1103, w_070_1104, w_070_1105, w_070_1106, w_070_1110, w_070_1111, w_070_1112, w_070_1115, w_070_1116, w_070_1117, w_070_1118, w_070_1121, w_070_1123, w_070_1124, w_070_1126, w_070_1127, w_070_1128, w_070_1130, w_070_1131, w_070_1134, w_070_1135, w_070_1136, w_070_1138, w_070_1139, w_070_1140, w_070_1141, w_070_1144, w_070_1148, w_070_1149, w_070_1150, w_070_1151, w_070_1153, w_070_1154, w_070_1155, w_070_1157, w_070_1163, w_070_1164, w_070_1166, w_070_1167, w_070_1168, w_070_1176, w_070_1180, w_070_1181, w_070_1184, w_070_1185, w_070_1190, w_070_1191, w_070_1192, w_070_1195, w_070_1196, w_070_1200, w_070_1201, w_070_1203, w_070_1204, w_070_1208, w_070_1209, w_070_1210, w_070_1211, w_070_1212, w_070_1215, w_070_1216, w_070_1217, w_070_1219, w_070_1220, w_070_1221, w_070_1222, w_070_1224, w_070_1225, w_070_1226, w_070_1227, w_070_1228, w_070_1230, w_070_1231, w_070_1232, w_070_1233, w_070_1234, w_070_1236, w_070_1237, w_070_1240, w_070_1243, w_070_1247, w_070_1252, w_070_1253, w_070_1254, w_070_1256, w_070_1259, w_070_1264, w_070_1268, w_070_1269, w_070_1270, w_070_1271, w_070_1274, w_070_1276, w_070_1277, w_070_1280, w_070_1281, w_070_1283, w_070_1284, w_070_1285, w_070_1286, w_070_1287, w_070_1288, w_070_1291, w_070_1292, w_070_1294, w_070_1295, w_070_1297, w_070_1301, w_070_1304, w_070_1305, w_070_1306, w_070_1307, w_070_1308, w_070_1309, w_070_1311, w_070_1313, w_070_1316, w_070_1319, w_070_1322, w_070_1326, w_070_1328, w_070_1331, w_070_1333, w_070_1334, w_070_1335, w_070_1336, w_070_1337, w_070_1338, w_070_1339, w_070_1341, w_070_1342, w_070_1344, w_070_1345, w_070_1347, w_070_1348, w_070_1349, w_070_1350, w_070_1353, w_070_1356, w_070_1358, w_070_1360, w_070_1361, w_070_1363, w_070_1364, w_070_1366, w_070_1370, w_070_1371, w_070_1372, w_070_1374, w_070_1378, w_070_1379, w_070_1380, w_070_1381, w_070_1382, w_070_1384, w_070_1385, w_070_1386, w_070_1387, w_070_1388, w_070_1389, w_070_1390, w_070_1391, w_070_1393, w_070_1394, w_070_1396, w_070_1399, w_070_1400, w_070_1401, w_070_1402, w_070_1404, w_070_1405, w_070_1409, w_070_1410, w_070_1411, w_070_1413, w_070_1415, w_070_1416, w_070_1420, w_070_1423, w_070_1425, w_070_1426, w_070_1432, w_070_1433, w_070_1439, w_070_1441, w_070_1442, w_070_1443, w_070_1444, w_070_1446, w_070_1447, w_070_1448, w_070_1451, w_070_1452, w_070_1457, w_070_1460, w_070_1465, w_070_1469, w_070_1470, w_070_1471, w_070_1474, w_070_1479, w_070_1482, w_070_1483, w_070_1486, w_070_1487, w_070_1488, w_070_1489, w_070_1490, w_070_1492, w_070_1493, w_070_1494, w_070_1496, w_070_1500, w_070_1501, w_070_1502, w_070_1503, w_070_1505, w_070_1506, w_070_1510, w_070_1512, w_070_1513, w_070_1515, w_070_1516, w_070_1518, w_070_1519, w_070_1520, w_070_1521, w_070_1523, w_070_1525, w_070_1527, w_070_1528, w_070_1530, w_070_1532, w_070_1533, w_070_1535, w_070_1536, w_070_1539, w_070_1540, w_070_1541, w_070_1542, w_070_1543, w_070_1544, w_070_1546, w_070_1548, w_070_1549, w_070_1550, w_070_1553, w_070_1554, w_070_1558, w_070_1560, w_070_1561, w_070_1563, w_070_1564, w_070_1565, w_070_1567, w_070_1570, w_070_1571, w_070_1572, w_070_1574, w_070_1576, w_070_1577, w_070_1578, w_070_1580, w_070_1581, w_070_1582, w_070_1583, w_070_1584, w_070_1587, w_070_1589, w_070_1590, w_070_1593, w_070_1594, w_070_1596, w_070_1598, w_070_1599, w_070_1600, w_070_1601, w_070_1604, w_070_1606, w_070_1608, w_070_1609, w_070_1610, w_070_1611, w_070_1612, w_070_1613, w_070_1616, w_070_1617, w_070_1618, w_070_1620, w_070_1621, w_070_1622, w_070_1625, w_070_1626, w_070_1630, w_070_1632, w_070_1633, w_070_1635, w_070_1637, w_070_1638, w_070_1639, w_070_1640, w_070_1647, w_070_1649, w_070_1650, w_070_1653, w_070_1655, w_070_1656, w_070_1658, w_070_1662, w_070_1664, w_070_1665, w_070_1667, w_070_1670, w_070_1673, w_070_1674, w_070_1678, w_070_1679, w_070_1680, w_070_1681, w_070_1682, w_070_1686, w_070_1687, w_070_1689, w_070_1691, w_070_1695, w_070_1696, w_070_1699, w_070_1701, w_070_1702, w_070_1703, w_070_1704, w_070_1705, w_070_1706, w_070_1707, w_070_1709, w_070_1711, w_070_1712, w_070_1715, w_070_1716, w_070_1718, w_070_1719, w_070_1725, w_070_1727, w_070_1729, w_070_1730, w_070_1732, w_070_1733, w_070_1735, w_070_1736, w_070_1737, w_070_1738, w_070_1740, w_070_1743, w_070_1745, w_070_1748, w_070_1749, w_070_1750, w_070_1756, w_070_1758, w_070_1760, w_070_1761, w_070_1762, w_070_1763, w_070_1766, w_070_1767, w_070_1768, w_070_1769, w_070_1771, w_070_1772, w_070_1773, w_070_1774, w_070_1776, w_070_1777, w_070_1783, w_070_1784, w_070_1786, w_070_1787, w_070_1788, w_070_1790, w_070_1793, w_070_1794, w_070_1795, w_070_1798, w_070_1799, w_070_1803, w_070_1804, w_070_1805, w_070_1806, w_070_1809, w_070_1812, w_070_1813, w_070_1814, w_070_1816, w_070_1818, w_070_1819, w_070_1820, w_070_1822, w_070_1823, w_070_1826, w_070_1829, w_070_1830, w_070_1831, w_070_1834, w_070_1835, w_070_1836, w_070_1837, w_070_1839, w_070_1840, w_070_1841, w_070_1842, w_070_1843, w_070_1844, w_070_1846, w_070_1848, w_070_1850, w_070_1852, w_070_1853, w_070_1854, w_070_1856, w_070_1857, w_070_1858, w_070_1859, w_070_1863, w_070_1866, w_070_1867, w_070_1869, w_070_1870, w_070_1871, w_070_1872, w_070_1874, w_070_1876, w_070_1877, w_070_1878, w_070_1879, w_070_1881, w_070_1882, w_070_1884, w_070_1885, w_070_1888, w_070_1891, w_070_1893, w_070_1894, w_070_1895, w_070_1896, w_070_1900, w_070_1902, w_070_1903, w_070_1906, w_070_1909, w_070_1912, w_070_1915, w_070_1917, w_070_1922, w_070_1923, w_070_1924, w_070_1927, w_070_1929, w_070_1930, w_070_1932, w_070_1933, w_070_1934, w_070_1935, w_070_1936, w_070_1937, w_070_1940, w_070_1943, w_070_1946, w_070_1949, w_070_1950, w_070_1951, w_070_1953, w_070_1954, w_070_1956, w_070_1958, w_070_1959, w_070_1960, w_070_1961, w_070_1962, w_070_1963, w_070_1964, w_070_1971, w_070_1972, w_070_1973, w_070_1976, w_070_1983, w_070_1985, w_070_1986, w_070_1987, w_070_1988, w_070_1990, w_070_1991, w_070_1993, w_070_1995, w_070_1996, w_070_1997, w_070_1998, w_070_1999, w_070_2000, w_070_2001, w_070_2002, w_070_2004, w_070_2006, w_070_2009, w_070_2012, w_070_2013, w_070_2014, w_070_2015, w_070_2025, w_070_2026, w_070_2027, w_070_2028, w_070_2029, w_070_2033, w_070_2034, w_070_2036, w_070_2039, w_070_2040, w_070_2041, w_070_2042, w_070_2043, w_070_2044, w_070_2045, w_070_2052, w_070_2053, w_070_2055, w_070_2057, w_070_2064, w_070_2065, w_070_2067, w_070_2068, w_070_2070, w_070_2072, w_070_2073, w_070_2075, w_070_2078, w_070_2080, w_070_2081, w_070_2082, w_070_2083, w_070_2085, w_070_2086, w_070_2087, w_070_2090, w_070_2092, w_070_2093, w_070_2097, w_070_2098, w_070_2100, w_070_2103, w_070_2105, w_070_2106, w_070_2108, w_070_2110, w_070_2112, w_070_2115, w_070_2116, w_070_2120, w_070_2124, w_070_2126, w_070_2128, w_070_2129, w_070_2130, w_070_2133, w_070_2134, w_070_2136, w_070_2138, w_070_2142, w_070_2145, w_070_2149, w_070_2151, w_070_2152, w_070_2153, w_070_2156, w_070_2158, w_070_2159, w_070_2160, w_070_2161, w_070_2166, w_070_2168, w_070_2170, w_070_2171, w_070_2172, w_070_2174, w_070_2178, w_070_2180, w_070_2182, w_070_2183, w_070_2185, w_070_2187, w_070_2190, w_070_2191, w_070_2192, w_070_2193, w_070_2195, w_070_2197, w_070_2204, w_070_2205, w_070_2206, w_070_2209, w_070_2210, w_070_2211, w_070_2213, w_070_2215, w_070_2217, w_070_2218, w_070_2219, w_070_2224, w_070_2225, w_070_2226, w_070_2228, w_070_2231, w_070_2232, w_070_2233, w_070_2234, w_070_2238, w_070_2239, w_070_2240, w_070_2243, w_070_2246, w_070_2247, w_070_2248, w_070_2249, w_070_2250, w_070_2252, w_070_2254, w_070_2255, w_070_2259, w_070_2264, w_070_2266, w_070_2270, w_070_2276, w_070_2280, w_070_2281, w_070_2282, w_070_2283, w_070_2284, w_070_2287, w_070_2288, w_070_2298, w_070_2299, w_070_2300, w_070_2301, w_070_2305, w_070_2307, w_070_2310, w_070_2313, w_070_2316, w_070_2317, w_070_2319, w_070_2320, w_070_2321, w_070_2322, w_070_2326, w_070_2327, w_070_2329, w_070_2331, w_070_2332, w_070_2334, w_070_2336, w_070_2337, w_070_2339, w_070_2342, w_070_2343, w_070_2344, w_070_2346, w_070_2351, w_070_2353, w_070_2354, w_070_2355, w_070_2356, w_070_2358, w_070_2359, w_070_2361, w_070_2363, w_070_2364, w_070_2365, w_070_2367, w_070_2373, w_070_2375, w_070_2376, w_070_2377, w_070_2378, w_070_2380, w_070_2381, w_070_2382, w_070_2383, w_070_2387, w_070_2390, w_070_2392, w_070_2393, w_070_2395, w_070_2396, w_070_2397, w_070_2399, w_070_2402, w_070_2405, w_070_2406, w_070_2407, w_070_2410, w_070_2411, w_070_2413, w_070_2414, w_070_2415, w_070_2416, w_070_2418, w_070_2419, w_070_2422, w_070_2424, w_070_2426, w_070_2428, w_070_2429, w_070_2433, w_070_2435, w_070_2437, w_070_2439, w_070_2440, w_070_2441, w_070_2443, w_070_2446, w_070_2447, w_070_2449, w_070_2452, w_070_2454, w_070_2458, w_070_2465, w_070_2466, w_070_2468, w_070_2473, w_070_2474, w_070_2476, w_070_2477, w_070_2478, w_070_2479, w_070_2481, w_070_2482, w_070_2483, w_070_2486, w_070_2487, w_070_2488, w_070_2491, w_070_2493, w_070_2494, w_070_2497, w_070_2498, w_070_2499, w_070_2500, w_070_2503, w_070_2504, w_070_2505, w_070_2506, w_070_2508, w_070_2510, w_070_2512, w_070_2513, w_070_2515, w_070_2518, w_070_2519, w_070_2520, w_070_2521, w_070_2522, w_070_2523, w_070_2525, w_070_2526, w_070_2527, w_070_2528, w_070_2529, w_070_2530, w_070_2531, w_070_2532, w_070_2533, w_070_2536, w_070_2537, w_070_2539, w_070_2540, w_070_2541, w_070_2543, w_070_2545, w_070_2549, w_070_2552, w_070_2554, w_070_2556, w_070_2557, w_070_2561, w_070_2564, w_070_2566, w_070_2567, w_070_2568, w_070_2569, w_070_2570, w_070_2571, w_070_2572, w_070_2581, w_070_2582, w_070_2584, w_070_2586, w_070_2587, w_070_2588, w_070_2593, w_070_2595, w_070_2596, w_070_2599, w_070_2603, w_070_2605, w_070_2606, w_070_2609, w_070_2610, w_070_2611, w_070_2612, w_070_2615, w_070_2617, w_070_2621, w_070_2622, w_070_2625, w_070_2626, w_070_2627, w_070_2629, w_070_2631, w_070_2633, w_070_2634, w_070_2635, w_070_2638, w_070_2640, w_070_2642, w_070_2646, w_070_2647, w_070_2648, w_070_2649, w_070_2651, w_070_2652, w_070_2653, w_070_2654, w_070_2657, w_070_2658, w_070_2659, w_070_2665, w_070_2667, w_070_2669, w_070_2671, w_070_2673, w_070_2677, w_070_2678, w_070_2680, w_070_2681, w_070_2682, w_070_2685, w_070_2690, w_070_2695, w_070_2701, w_070_2703, w_070_2704, w_070_2706, w_070_2709, w_070_2710, w_070_2711, w_070_2713, w_070_2716, w_070_2717, w_070_2718, w_070_2719, w_070_2720, w_070_2724, w_070_2726, w_070_2727, w_070_2729, w_070_2730, w_070_2731, w_070_2734, w_070_2737, w_070_2739, w_070_2740, w_070_2746, w_070_2748, w_070_2749, w_070_2751, w_070_2753, w_070_2756, w_070_2758, w_070_2759, w_070_2762, w_070_2763, w_070_2764, w_070_2765, w_070_2767, w_070_2769, w_070_2770, w_070_2772, w_070_2774, w_070_2776, w_070_2778, w_070_2781, w_070_2782, w_070_2784, w_070_2785, w_070_2786, w_070_2788, w_070_2789, w_070_2790, w_070_2791, w_070_2792, w_070_2793, w_070_2796, w_070_2797, w_070_2798, w_070_2799, w_070_2800, w_070_2802, w_070_2803, w_070_2804, w_070_2805, w_070_2808, w_070_2811, w_070_2812, w_070_2814, w_070_2816, w_070_2817, w_070_2821, w_070_2822, w_070_2823, w_070_2825, w_070_2826, w_070_2827, w_070_2828, w_070_2829, w_070_2831, w_070_2832, w_070_2834, w_070_2835, w_070_2838, w_070_2839, w_070_2840, w_070_2841, w_070_2842, w_070_2843, w_070_2844, w_070_2845, w_070_2846, w_070_2847, w_070_2848, w_070_2852, w_070_2853, w_070_2857, w_070_2860, w_070_2861, w_070_2862, w_070_2864, w_070_2865, w_070_2866, w_070_2867, w_070_2868, w_070_2869, w_070_2874, w_070_2875, w_070_2876, w_070_2878, w_070_2879, w_070_2880, w_070_2884, w_070_2885, w_070_2892, w_070_2893, w_070_2894, w_070_2897, w_070_2899, w_070_2901, w_070_2902, w_070_2904, w_070_2906, w_070_2910, w_070_2911, w_070_2912, w_070_2913, w_070_2914, w_070_2919, w_070_2921, w_070_2923, w_070_2925, w_070_2928, w_070_2932, w_070_2935, w_070_2937, w_070_2939, w_070_2941, w_070_2942, w_070_2943, w_070_2949, w_070_2953, w_070_2956, w_070_2962, w_070_2963, w_070_2965, w_070_2967, w_070_2968, w_070_2970, w_070_2973, w_070_2977, w_070_2983, w_070_2984, w_070_2986, w_070_2988, w_070_2989, w_070_2990, w_070_2991, w_070_2995, w_070_2997, w_070_2999, w_070_3000, w_070_3001, w_070_3003, w_070_3005, w_070_3007, w_070_3011, w_070_3012, w_070_3013, w_070_3014, w_070_3016, w_070_3017, w_070_3019, w_070_3021, w_070_3027, w_070_3030, w_070_3033, w_070_3034, w_070_3036, w_070_3039, w_070_3040, w_070_3043, w_070_3045, w_070_3046, w_070_3047, w_070_3049, w_070_3051, w_070_3052, w_070_3053, w_070_3054, w_070_3057, w_070_3058, w_070_3060, w_070_3061, w_070_3069, w_070_3070, w_070_3071, w_070_3072, w_070_3073, w_070_3077, w_070_3079, w_070_3080, w_070_3085, w_070_3086, w_070_3087, w_070_3090, w_070_3092, w_070_3095, w_070_3096, w_070_3097, w_070_3100, w_070_3103, w_070_3104, w_070_3105, w_070_3108, w_070_3110, w_070_3115, w_070_3122, w_070_3129, w_070_3130, w_070_3131, w_070_3132, w_070_3134, w_070_3136, w_070_3137, w_070_3140, w_070_3142, w_070_3144, w_070_3147, w_070_3148, w_070_3149, w_070_3150, w_070_3152, w_070_3154, w_070_3155, w_070_3156, w_070_3157, w_070_3159, w_070_3161, w_070_3164, w_070_3167, w_070_3168, w_070_3169, w_070_3171, w_070_3173, w_070_3175, w_070_3182, w_070_3183, w_070_3184, w_070_3186, w_070_3187, w_070_3188, w_070_3190, w_070_3191, w_070_3192, w_070_3194, w_070_3199, w_070_3202, w_070_3204, w_070_3205, w_070_3208, w_070_3210, w_070_3211, w_070_3213, w_070_3215, w_070_3217, w_070_3219, w_070_3222, w_070_3223, w_070_3224, w_070_3225, w_070_3226, w_070_3227, w_070_3230, w_070_3233, w_070_3234, w_070_3235, w_070_3241, w_070_3243, w_070_3244, w_070_3245, w_070_3246, w_070_3247, w_070_3248, w_070_3251, w_070_3252, w_070_3254, w_070_3255, w_070_3256, w_070_3257, w_070_3259, w_070_3260, w_070_3262, w_070_3266, w_070_3268, w_070_3271, w_070_3272, w_070_3274, w_070_3275, w_070_3276, w_070_3278, w_070_3279, w_070_3281, w_070_3283, w_070_3285, w_070_3287, w_070_3291, w_070_3293, w_070_3295, w_070_3298, w_070_3300, w_070_3301, w_070_3303, w_070_3305, w_070_3308, w_070_3311, w_070_3312, w_070_3313, w_070_3314, w_070_3316, w_070_3317, w_070_3322, w_070_3323, w_070_3328, w_070_3329, w_070_3330, w_070_3333, w_070_3336, w_070_3337, w_070_3339, w_070_3342, w_070_3343, w_070_3344, w_070_3345, w_070_3349, w_070_3351, w_070_3353, w_070_3355, w_070_3358, w_070_3359, w_070_3364, w_070_3368, w_070_3369, w_070_3370, w_070_3371, w_070_3372, w_070_3373, w_070_3375, w_070_3379, w_070_3380, w_070_3385, w_070_3386, w_070_3390, w_070_3391, w_070_3392, w_070_3393, w_070_3396, w_070_3397, w_070_3402, w_070_3403, w_070_3405, w_070_3406, w_070_3407, w_070_3408, w_070_3409, w_070_3411, w_070_3412, w_070_3415, w_070_3416, w_070_3418, w_070_3419, w_070_3421, w_070_3422, w_070_3423, w_070_3425, w_070_3426, w_070_3430, w_070_3432, w_070_3433, w_070_3437, w_070_3438, w_070_3440, w_070_3441, w_070_3445, w_070_3446, w_070_3447, w_070_3450, w_070_3451, w_070_3452, w_070_3454, w_070_3456, w_070_3457, w_070_3458, w_070_3460, w_070_3462, w_070_3463, w_070_3470, w_070_3471, w_070_3475, w_070_3476, w_070_3478, w_070_3480, w_070_3485, w_070_3486, w_070_3487, w_070_3488, w_070_3493, w_070_3494, w_070_3495, w_070_3497, w_070_3498, w_070_3502, w_070_3503, w_070_3504, w_070_3505, w_070_3506, w_070_3507, w_070_3513, w_070_3515, w_070_3517, w_070_3518, w_070_3520, w_070_3521, w_070_3522, w_070_3523, w_070_3529, w_070_3531, w_070_3532, w_070_3533, w_070_3534, w_070_3535, w_070_3546, w_070_3548, w_070_3549, w_070_3550, w_070_3552, w_070_3554, w_070_3556, w_070_3557, w_070_3558, w_070_3560, w_070_3561, w_070_3562, w_070_3563, w_070_3565, w_070_3567, w_070_3568, w_070_3569, w_070_3571, w_070_3572, w_070_3573, w_070_3574, w_070_3575, w_070_3576, w_070_3579, w_070_3581, w_070_3586, w_070_3588, w_070_3591, w_070_3592, w_070_3593, w_070_3596, w_070_3597, w_070_3599, w_070_3602, w_070_3603, w_070_3604, w_070_3609, w_070_3611, w_070_3612, w_070_3614, w_070_3618, w_070_3619, w_070_3625, w_070_3628, w_070_3629, w_070_3632, w_070_3633, w_070_3635, w_070_3637, w_070_3638, w_070_3643, w_070_3644, w_070_3646, w_070_3649, w_070_3650, w_070_3651, w_070_3652, w_070_3656, w_070_3657, w_070_3658, w_070_3659, w_070_3660, w_070_3661, w_070_3663, w_070_3665, w_070_3667, w_070_3671, w_070_3672, w_070_3674, w_070_3675, w_070_3676, w_070_3677, w_070_3678, w_070_3679, w_070_3680, w_070_3681, w_070_3682, w_070_3683, w_070_3685, w_070_3690, w_070_3692, w_070_3693, w_070_3694, w_070_3696, w_070_3700, w_070_3701, w_070_3702, w_070_3704, w_070_3707, w_070_3709, w_070_3710, w_070_3712, w_070_3713, w_070_3716, w_070_3718, w_070_3721, w_070_3723, w_070_3724, w_070_3726, w_070_3727, w_070_3728, w_070_3729, w_070_3731, w_070_3732, w_070_3733, w_070_3737, w_070_3741, w_070_3742, w_070_3743, w_070_3744, w_070_3746, w_070_3749, w_070_3752, w_070_3753, w_070_3754, w_070_3756, w_070_3757, w_070_3758, w_070_3759, w_070_3761, w_070_3762, w_070_3763, w_070_3764, w_070_3765, w_070_3766, w_070_3768, w_070_3771, w_070_3773, w_070_3775, w_070_3777, w_070_3779, w_070_3780, w_070_3782, w_070_3783, w_070_3786, w_070_3787, w_070_3790, w_070_3791, w_070_3794, w_070_3797, w_070_3800, w_070_3801, w_070_3803, w_070_3804, w_070_3806, w_070_3810, w_070_3811, w_070_3812, w_070_3815, w_070_3816, w_070_3819, w_070_3820, w_070_3823, w_070_3824, w_070_3828, w_070_3830, w_070_3831, w_070_3832, w_070_3833, w_070_3834, w_070_3835, w_070_3838, w_070_3841, w_070_3844, w_070_3846, w_070_3847, w_070_3848, w_070_3850, w_070_3851, w_070_3852, w_070_3854, w_070_3855, w_070_3856, w_070_3857, w_070_3858, w_070_3859, w_070_3860, w_070_3861, w_070_3862, w_070_3863, w_070_3864, w_070_3866, w_070_3869, w_070_3873, w_070_3874, w_070_3876, w_070_3877, w_070_3879, w_070_3881, w_070_3882, w_070_3883, w_070_3885, w_070_3886, w_070_3888, w_070_3889, w_070_3890, w_070_3892, w_070_3895, w_070_3896, w_070_3897, w_070_3898, w_070_3900, w_070_3901, w_070_3902, w_070_3903, w_070_3906, w_070_3909, w_070_3911, w_070_3914, w_070_3922, w_070_3923, w_070_3925, w_070_3926, w_070_3928, w_070_3932, w_070_3937, w_070_3939, w_070_3940, w_070_3941, w_070_3943, w_070_3944, w_070_3946, w_070_3947, w_070_3949, w_070_3951, w_070_3952, w_070_3953, w_070_3956, w_070_3957, w_070_3958, w_070_3962, w_070_3963, w_070_3965, w_070_3966, w_070_3969, w_070_3972, w_070_3973, w_070_3974, w_070_3975, w_070_3976, w_070_3981, w_070_3982, w_070_3983, w_070_3985, w_070_3987, w_070_3988, w_070_3989, w_070_3993, w_070_3995, w_070_3997, w_070_3999, w_070_4000, w_070_4002, w_070_4003, w_070_4005, w_070_4007, w_070_4008, w_070_4010, w_070_4012, w_070_4014, w_070_4016, w_070_4018, w_070_4020, w_070_4024, w_070_4025, w_070_4028, w_070_4029, w_070_4032, w_070_4033, w_070_4034, w_070_4035, w_070_4036, w_070_4038, w_070_4039, w_070_4041, w_070_4042, w_070_4043, w_070_4044, w_070_4046, w_070_4048, w_070_4049, w_070_4051, w_070_4052, w_070_4053, w_070_4054, w_070_4057, w_070_4060, w_070_4062, w_070_4063, w_070_4065, w_070_4066, w_070_4068, w_070_4069, w_070_4071, w_070_4072, w_070_4075, w_070_4077, w_070_4079, w_070_4081, w_070_4086, w_070_4089, w_070_4090, w_070_4091, w_070_4092, w_070_4093, w_070_4094, w_070_4095, w_070_4096, w_070_4097, w_070_4099, w_070_4100, w_070_4105, w_070_4107, w_070_4108, w_070_4109, w_070_4113, w_070_4115, w_070_4116, w_070_4119, w_070_4126, w_070_4128, w_070_4131, w_070_4136, w_070_4137, w_070_4138, w_070_4139, w_070_4140, w_070_4141, w_070_4143, w_070_4145, w_070_4146, w_070_4147, w_070_4148, w_070_4149, w_070_4150, w_070_4151, w_070_4153, w_070_4156, w_070_4158, w_070_4160, w_070_4163, w_070_4164, w_070_4167, w_070_4168, w_070_4169, w_070_4171, w_070_4172, w_070_4174, w_070_4175, w_070_4180, w_070_4184, w_070_4186, w_070_4188, w_070_4189, w_070_4190, w_070_4192, w_070_4196, w_070_4197, w_070_4198, w_070_4199, w_070_4201, w_070_4203, w_070_4204, w_070_4205, w_070_4208, w_070_4211, w_070_4212, w_070_4213, w_070_4215, w_070_4217, w_070_4219, w_070_4220, w_070_4222, w_070_4223, w_070_4224, w_070_4225, w_070_4226, w_070_4227, w_070_4228, w_070_4229, w_070_4230, w_070_4231, w_070_4233, w_070_4234, w_070_4235, w_070_4236, w_070_4238, w_070_4239, w_070_4240, w_070_4241, w_070_4245, w_070_4246, w_070_4248, w_070_4249, w_070_4250, w_070_4251, w_070_4253, w_070_4257, w_070_4258, w_070_4259, w_070_4260, w_070_4261, w_070_4266, w_070_4267, w_070_4271, w_070_4272, w_070_4273, w_070_4275, w_070_4277, w_070_4278, w_070_4279, w_070_4283, w_070_4284, w_070_4286, w_070_4288, w_070_4293, w_070_4295, w_070_4296, w_070_4297, w_070_4298, w_070_4299, w_070_4302, w_070_4303, w_070_4305, w_070_4308, w_070_4309, w_070_4310, w_070_4311, w_070_4312, w_070_4314, w_070_4316, w_070_4317, w_070_4319, w_070_4320, w_070_4323, w_070_4325, w_070_4326, w_070_4328, w_070_4331, w_070_4336, w_070_4344, w_070_4346, w_070_4347, w_070_4360, w_070_4362, w_070_4363, w_070_4369, w_070_4374, w_070_4376, w_070_4379, w_070_4380, w_070_4381, w_070_4387, w_070_4389, w_070_4395, w_070_4399, w_070_4404, w_070_4408, w_070_4409, w_070_4410, w_070_4414, w_070_4422, w_070_4423, w_070_4426, w_070_4435, w_070_4442, w_070_4445, w_070_4447, w_070_4455, w_070_4456, w_070_4457, w_070_4461, w_070_4463, w_070_4467, w_070_4470, w_070_4471, w_070_4472, w_070_4473, w_070_4477, w_070_4478, w_070_4489, w_070_4495, w_070_4497, w_070_4504, w_070_4505, w_070_4506, w_070_4508, w_070_4519, w_070_4523, w_070_4527, w_070_4528, w_070_4533, w_070_4543, w_070_4544, w_070_4546, w_070_4553, w_070_4561, w_070_4567, w_070_4574, w_070_4578, w_070_4583, w_070_4585, w_070_4587, w_070_4590, w_070_4591, w_070_4602, w_070_4604, w_070_4605, w_070_4606, w_070_4609, w_070_4614, w_070_4618, w_070_4624, w_070_4625, w_070_4629, w_070_4635, w_070_4637, w_070_4638, w_070_4640, w_070_4647, w_070_4648, w_070_4650, w_070_4652, w_070_4654, w_070_4657, w_070_4660, w_070_4662, w_070_4663, w_070_4669, w_070_4670, w_070_4672, w_070_4676, w_070_4680, w_070_4682, w_070_4684, w_070_4688, w_070_4699, w_070_4701, w_070_4706, w_070_4707, w_070_4709, w_070_4713, w_070_4715, w_070_4717, w_070_4718, w_070_4719, w_070_4720, w_070_4721, w_070_4725, w_070_4727, w_070_4728, w_070_4729, w_070_4731, w_070_4732, w_070_4736, w_070_4737, w_070_4740, w_070_4741, w_070_4742, w_070_4749, w_070_4753, w_070_4760, w_070_4766, w_070_4767, w_070_4770, w_070_4772, w_070_4775, w_070_4777, w_070_4778, w_070_4780, w_070_4783, w_070_4784, w_070_4786, w_070_4789, w_070_4791, w_070_4793, w_070_4795, w_070_4797, w_070_4799, w_070_4803, w_070_4807, w_070_4811, w_070_4813, w_070_4816, w_070_4817, w_070_4818, w_070_4819, w_070_4821, w_070_4830, w_070_4832, w_070_4838, w_070_4841, w_070_4842, w_070_4843, w_070_4845, w_070_4847, w_070_4850, w_070_4851, w_070_4853, w_070_4855, w_070_4858, w_070_4860, w_070_4861, w_070_4863, w_070_4867, w_070_4872, w_070_4873, w_070_4875, w_070_4881, w_070_4887, w_070_4889, w_070_4890, w_070_4892, w_070_4895, w_070_4899, w_070_4906, w_070_4909, w_070_4912, w_070_4913, w_070_4915, w_070_4918, w_070_4919, w_070_4921, w_070_4923, w_070_4925, w_070_4927, w_070_4932, w_070_4933, w_070_4938, w_070_4947, w_070_4949, w_070_4958, w_070_4960, w_070_4962, w_070_4967, w_070_4971, w_070_4972, w_070_4973, w_070_4982, w_070_4983, w_070_4985, w_070_4987, w_070_4993, w_070_4995, w_070_5004, w_070_5009, w_070_5014, w_070_5019, w_070_5020, w_070_5022, w_070_5023, w_070_5024, w_070_5029, w_070_5030, w_070_5032, w_070_5034, w_070_5036, w_070_5037, w_070_5042, w_070_5045, w_070_5051, w_070_5052, w_070_5055, w_070_5059, w_070_5063, w_070_5064, w_070_5065, w_070_5069, w_070_5075, w_070_5076, w_070_5079, w_070_5080, w_070_5083, w_070_5086, w_070_5087, w_070_5088, w_070_5089, w_070_5093, w_070_5094, w_070_5109, w_070_5111, w_070_5117, w_070_5118, w_070_5121, w_070_5126, w_070_5129, w_070_5133, w_070_5137, w_070_5138, w_070_5146, w_070_5149, w_070_5150, w_070_5151, w_070_5152, w_070_5157, w_070_5158, w_070_5160, w_070_5165, w_070_5166, w_070_5170, w_070_5173, w_070_5174, w_070_5178, w_070_5179, w_070_5187, w_070_5188, w_070_5198, w_070_5200, w_070_5202, w_070_5203, w_070_5205, w_070_5207, w_070_5211, w_070_5214, w_070_5219, w_070_5221, w_070_5226, w_070_5228, w_070_5229, w_070_5230, w_070_5238, w_070_5242, w_070_5245, w_070_5248, w_070_5251, w_070_5252, w_070_5253, w_070_5263, w_070_5264, w_070_5265, w_070_5267, w_070_5269, w_070_5284, w_070_5288, w_070_5289, w_070_5290, w_070_5291, w_070_5295, w_070_5296, w_070_5298, w_070_5299, w_070_5300, w_070_5302, w_070_5305, w_070_5309, w_070_5310, w_070_5311, w_070_5312, w_070_5313, w_070_5315, w_070_5316, w_070_5317, w_070_5318, w_070_5321, w_070_5325, w_070_5328, w_070_5339, w_070_5350, w_070_5353, w_070_5355, w_070_5356, w_070_5359, w_070_5368, w_070_5370, w_070_5372, w_070_5373, w_070_5390, w_070_5395, w_070_5396, w_070_5399, w_070_5402, w_070_5413, w_070_5421, w_070_5423, w_070_5424, w_070_5426, w_070_5427, w_070_5428, w_070_5431, w_070_5435, w_070_5441, w_070_5442, w_070_5448, w_070_5449, w_070_5451, w_070_5453, w_070_5454, w_070_5456, w_070_5460, w_070_5461, w_070_5472, w_070_5473, w_070_5475, w_070_5479, w_070_5492, w_070_5493, w_070_5495, w_070_5497, w_070_5498, w_070_5501, w_070_5502, w_070_5503, w_070_5504, w_070_5506, w_070_5511, w_070_5513, w_070_5516, w_070_5520, w_070_5524, w_070_5525, w_070_5528, w_070_5530, w_070_5531, w_070_5534, w_070_5537, w_070_5538, w_070_5541, w_070_5544, w_070_5546, w_070_5553, w_070_5556, w_070_5561, w_070_5562, w_070_5563, w_070_5566, w_070_5567, w_070_5570, w_070_5572, w_070_5573, w_070_5577, w_070_5578, w_070_5580, w_070_5582, w_070_5583, w_070_5588, w_070_5594, w_070_5597, w_070_5599, w_070_5600, w_070_5601, w_070_5602, w_070_5604, w_070_5605, w_070_5609, w_070_5613, w_070_5614, w_070_5623, w_070_5624, w_070_5635, w_070_5637, w_070_5639, w_070_5645, w_070_5650, w_070_5655, w_070_5656, w_070_5657, w_070_5660;
  wire w_071_000, w_071_001, w_071_002, w_071_003, w_071_004, w_071_006, w_071_007, w_071_009, w_071_010, w_071_011, w_071_012, w_071_013, w_071_014, w_071_015, w_071_016, w_071_017, w_071_019, w_071_021, w_071_022, w_071_023, w_071_024, w_071_025, w_071_027, w_071_028, w_071_029, w_071_030, w_071_031, w_071_032, w_071_033, w_071_034, w_071_035, w_071_037, w_071_038, w_071_039, w_071_040, w_071_041, w_071_043, w_071_044, w_071_045, w_071_046, w_071_047, w_071_049, w_071_050, w_071_051, w_071_052, w_071_054, w_071_056, w_071_057, w_071_059, w_071_060, w_071_061, w_071_062, w_071_063, w_071_064, w_071_065, w_071_066, w_071_067, w_071_068, w_071_069, w_071_070, w_071_071, w_071_073, w_071_075, w_071_076, w_071_077, w_071_078, w_071_080, w_071_081, w_071_082, w_071_083, w_071_084, w_071_085, w_071_086, w_071_087, w_071_088, w_071_090, w_071_091, w_071_092, w_071_093, w_071_094, w_071_095, w_071_096, w_071_097, w_071_098, w_071_099, w_071_100, w_071_102, w_071_103, w_071_104, w_071_105, w_071_106, w_071_107, w_071_109, w_071_110, w_071_111, w_071_112, w_071_113, w_071_114, w_071_115, w_071_116, w_071_117, w_071_118, w_071_119, w_071_121, w_071_123, w_071_124, w_071_125, w_071_126, w_071_127, w_071_128, w_071_129, w_071_130, w_071_131, w_071_132, w_071_133, w_071_134, w_071_135, w_071_136, w_071_137, w_071_138, w_071_139, w_071_142, w_071_144, w_071_145, w_071_146, w_071_148, w_071_149, w_071_151, w_071_152, w_071_153, w_071_154, w_071_155, w_071_156, w_071_157, w_071_159, w_071_160, w_071_161, w_071_162, w_071_163, w_071_164, w_071_165, w_071_167, w_071_168, w_071_169, w_071_170, w_071_171, w_071_173, w_071_174, w_071_175, w_071_177, w_071_178, w_071_180, w_071_182, w_071_183, w_071_184, w_071_185, w_071_186, w_071_187, w_071_189, w_071_190, w_071_191, w_071_192, w_071_193, w_071_194, w_071_195, w_071_196, w_071_197, w_071_198, w_071_199, w_071_201, w_071_202, w_071_205, w_071_206, w_071_207, w_071_210, w_071_211, w_071_212, w_071_213, w_071_214, w_071_216, w_071_217, w_071_218, w_071_219, w_071_220, w_071_221, w_071_222, w_071_223, w_071_224, w_071_225, w_071_226, w_071_227, w_071_228, w_071_229, w_071_230, w_071_231, w_071_232, w_071_233, w_071_235, w_071_238, w_071_239, w_071_240, w_071_242, w_071_244, w_071_245, w_071_246, w_071_247, w_071_248, w_071_250, w_071_252, w_071_254, w_071_255, w_071_256, w_071_258, w_071_259, w_071_261, w_071_262, w_071_264, w_071_265, w_071_266, w_071_267, w_071_268, w_071_269, w_071_270, w_071_271, w_071_272, w_071_273, w_071_275, w_071_276, w_071_277, w_071_278, w_071_279, w_071_280, w_071_281, w_071_282, w_071_283, w_071_284, w_071_285, w_071_286, w_071_287, w_071_289, w_071_290, w_071_291, w_071_292, w_071_293, w_071_294, w_071_297, w_071_299, w_071_300, w_071_301, w_071_302, w_071_303, w_071_304, w_071_305, w_071_306, w_071_307, w_071_308, w_071_309, w_071_310, w_071_311, w_071_312, w_071_313, w_071_314, w_071_315, w_071_316, w_071_317, w_071_318, w_071_319, w_071_320, w_071_321, w_071_322, w_071_324, w_071_326, w_071_327, w_071_328, w_071_329, w_071_330, w_071_331, w_071_332, w_071_336, w_071_337, w_071_339, w_071_341, w_071_342, w_071_343, w_071_344, w_071_345, w_071_346, w_071_347, w_071_348, w_071_349, w_071_350, w_071_351, w_071_352, w_071_353, w_071_355, w_071_356, w_071_357, w_071_360, w_071_361, w_071_363, w_071_364, w_071_365, w_071_367, w_071_368, w_071_370, w_071_371, w_071_374, w_071_375, w_071_376, w_071_378, w_071_379, w_071_380, w_071_381, w_071_382, w_071_383, w_071_384, w_071_385, w_071_386, w_071_387, w_071_388, w_071_389, w_071_390, w_071_391, w_071_392, w_071_393, w_071_394, w_071_395, w_071_396, w_071_397, w_071_398, w_071_399, w_071_400, w_071_402, w_071_404, w_071_405, w_071_406, w_071_409, w_071_410, w_071_411, w_071_412, w_071_413, w_071_414, w_071_415, w_071_416, w_071_417, w_071_418, w_071_419, w_071_420, w_071_421, w_071_422, w_071_423, w_071_424, w_071_425, w_071_426, w_071_427, w_071_429, w_071_430, w_071_431, w_071_432, w_071_433, w_071_434, w_071_436, w_071_437, w_071_438, w_071_439, w_071_440, w_071_441, w_071_444, w_071_445, w_071_446, w_071_447, w_071_448, w_071_449, w_071_450, w_071_451, w_071_452, w_071_453, w_071_454, w_071_455, w_071_456, w_071_457, w_071_458, w_071_459, w_071_461, w_071_462, w_071_464, w_071_465, w_071_466, w_071_467, w_071_468, w_071_469, w_071_470, w_071_471, w_071_472, w_071_473, w_071_475, w_071_476, w_071_477, w_071_479, w_071_480, w_071_481, w_071_482, w_071_483, w_071_484, w_071_485, w_071_486, w_071_487, w_071_488, w_071_489, w_071_491, w_071_492, w_071_493, w_071_494, w_071_495, w_071_496, w_071_497, w_071_498, w_071_501, w_071_502, w_071_504, w_071_505, w_071_506, w_071_507, w_071_508, w_071_509, w_071_510, w_071_511, w_071_513, w_071_514, w_071_516, w_071_518, w_071_520, w_071_521, w_071_522, w_071_523, w_071_524, w_071_525, w_071_526, w_071_527, w_071_528, w_071_529, w_071_530, w_071_531, w_071_532, w_071_533, w_071_534, w_071_536, w_071_537, w_071_538, w_071_539, w_071_540, w_071_541, w_071_542, w_071_543, w_071_544, w_071_545, w_071_546, w_071_547, w_071_548, w_071_550, w_071_552, w_071_555, w_071_558, w_071_560, w_071_562, w_071_564, w_071_565, w_071_567, w_071_568, w_071_569, w_071_570, w_071_571, w_071_573, w_071_574, w_071_575, w_071_576, w_071_577, w_071_579, w_071_580, w_071_584, w_071_585, w_071_586, w_071_590, w_071_591, w_071_592, w_071_594, w_071_595, w_071_597, w_071_598, w_071_599, w_071_600, w_071_601, w_071_602, w_071_603, w_071_604, w_071_606, w_071_607, w_071_608, w_071_609, w_071_610, w_071_612, w_071_616, w_071_617, w_071_618, w_071_619, w_071_620, w_071_623, w_071_625, w_071_626, w_071_627, w_071_630, w_071_632, w_071_633, w_071_634, w_071_635, w_071_637, w_071_638, w_071_639, w_071_641, w_071_642, w_071_643, w_071_644, w_071_645, w_071_646, w_071_647, w_071_648, w_071_650, w_071_651, w_071_652, w_071_653, w_071_654, w_071_655, w_071_656, w_071_657, w_071_660, w_071_661, w_071_664, w_071_665, w_071_667, w_071_668, w_071_669, w_071_670, w_071_672, w_071_673, w_071_674, w_071_675, w_071_676, w_071_677, w_071_678, w_071_679, w_071_681, w_071_682, w_071_683, w_071_684, w_071_685, w_071_686, w_071_687, w_071_688, w_071_689, w_071_690, w_071_691, w_071_693, w_071_694, w_071_695, w_071_697, w_071_698, w_071_701, w_071_702, w_071_704, w_071_705, w_071_708, w_071_709, w_071_711, w_071_712, w_071_713, w_071_714, w_071_716, w_071_717, w_071_719, w_071_723, w_071_725, w_071_726, w_071_727, w_071_728, w_071_729, w_071_730, w_071_731, w_071_732, w_071_733, w_071_734, w_071_735, w_071_737, w_071_738, w_071_739, w_071_740, w_071_741, w_071_742, w_071_745, w_071_746, w_071_747, w_071_748, w_071_750, w_071_751, w_071_752, w_071_753, w_071_755, w_071_756, w_071_757, w_071_758, w_071_759, w_071_762, w_071_763, w_071_764, w_071_765, w_071_766, w_071_767, w_071_768, w_071_770, w_071_771, w_071_772, w_071_776, w_071_777, w_071_778, w_071_779, w_071_780, w_071_782, w_071_783, w_071_784, w_071_785, w_071_786, w_071_787, w_071_788, w_071_789, w_071_790, w_071_791, w_071_793, w_071_795, w_071_796, w_071_797, w_071_798, w_071_800, w_071_801, w_071_802, w_071_803, w_071_804, w_071_806, w_071_807, w_071_808, w_071_809, w_071_810, w_071_812, w_071_813, w_071_815, w_071_817, w_071_818, w_071_819, w_071_823, w_071_824, w_071_825, w_071_827, w_071_828, w_071_829, w_071_831, w_071_832, w_071_833, w_071_834, w_071_835, w_071_836, w_071_837, w_071_838, w_071_839, w_071_840, w_071_841, w_071_842, w_071_843, w_071_845, w_071_847, w_071_848, w_071_849, w_071_850, w_071_851, w_071_852, w_071_853, w_071_855, w_071_856, w_071_857, w_071_858, w_071_859, w_071_860, w_071_861, w_071_862, w_071_864, w_071_866, w_071_869, w_071_871, w_071_872, w_071_873, w_071_874, w_071_875, w_071_876, w_071_877, w_071_878, w_071_879, w_071_880, w_071_881, w_071_884, w_071_885, w_071_887, w_071_888, w_071_890, w_071_892, w_071_893, w_071_894, w_071_895, w_071_896, w_071_897, w_071_898, w_071_900, w_071_902, w_071_904, w_071_905, w_071_908, w_071_910, w_071_911, w_071_912, w_071_914, w_071_915, w_071_916, w_071_917, w_071_919, w_071_920, w_071_922, w_071_923, w_071_924, w_071_925, w_071_928, w_071_929, w_071_930, w_071_933, w_071_934, w_071_935, w_071_936, w_071_940, w_071_941, w_071_943, w_071_944, w_071_946, w_071_947, w_071_948, w_071_950, w_071_951, w_071_952, w_071_953, w_071_954, w_071_955, w_071_956, w_071_957, w_071_959, w_071_962, w_071_964, w_071_965, w_071_966, w_071_967, w_071_968, w_071_969, w_071_971, w_071_972, w_071_973, w_071_974, w_071_975, w_071_976, w_071_977, w_071_979, w_071_980, w_071_981, w_071_982, w_071_984, w_071_985, w_071_989, w_071_992, w_071_993, w_071_995, w_071_996, w_071_997, w_071_999, w_071_1000, w_071_1001, w_071_1002, w_071_1003, w_071_1005, w_071_1006, w_071_1009, w_071_1012, w_071_1014, w_071_1015, w_071_1016, w_071_1017, w_071_1018, w_071_1019, w_071_1020, w_071_1021, w_071_1022, w_071_1023, w_071_1024, w_071_1025, w_071_1027, w_071_1028, w_071_1029, w_071_1030, w_071_1031, w_071_1032, w_071_1033, w_071_1034, w_071_1035, w_071_1036, w_071_1037, w_071_1040, w_071_1041, w_071_1042, w_071_1043, w_071_1044, w_071_1045, w_071_1046, w_071_1047, w_071_1048, w_071_1050, w_071_1051, w_071_1052, w_071_1053, w_071_1054, w_071_1055, w_071_1056, w_071_1058, w_071_1059, w_071_1060, w_071_1061, w_071_1062, w_071_1064, w_071_1065, w_071_1067, w_071_1068, w_071_1069, w_071_1070, w_071_1071, w_071_1072, w_071_1073, w_071_1074, w_071_1076, w_071_1077, w_071_1078, w_071_1079, w_071_1081, w_071_1082, w_071_1083, w_071_1084, w_071_1085, w_071_1086, w_071_1087, w_071_1088, w_071_1091, w_071_1092, w_071_1093, w_071_1094, w_071_1095, w_071_1099, w_071_1100, w_071_1101, w_071_1102, w_071_1104, w_071_1105, w_071_1106, w_071_1107, w_071_1109, w_071_1110, w_071_1111, w_071_1113, w_071_1114, w_071_1115, w_071_1116, w_071_1117, w_071_1119, w_071_1121, w_071_1122, w_071_1123, w_071_1124, w_071_1125, w_071_1127, w_071_1130, w_071_1131, w_071_1133, w_071_1134, w_071_1135, w_071_1139, w_071_1142, w_071_1143, w_071_1144, w_071_1145, w_071_1146, w_071_1148, w_071_1150, w_071_1151, w_071_1152, w_071_1153, w_071_1154, w_071_1156, w_071_1157, w_071_1159, w_071_1161, w_071_1162, w_071_1163, w_071_1165, w_071_1166, w_071_1167, w_071_1168, w_071_1169, w_071_1170, w_071_1171, w_071_1175, w_071_1176, w_071_1177, w_071_1179, w_071_1180, w_071_1181, w_071_1183, w_071_1184, w_071_1185, w_071_1186, w_071_1188, w_071_1189, w_071_1191, w_071_1193, w_071_1194, w_071_1195, w_071_1196, w_071_1197, w_071_1198, w_071_1200, w_071_1203, w_071_1204, w_071_1206, w_071_1207, w_071_1208, w_071_1209, w_071_1210, w_071_1211, w_071_1213, w_071_1215, w_071_1216, w_071_1217, w_071_1218, w_071_1219, w_071_1220, w_071_1221, w_071_1222, w_071_1223, w_071_1224, w_071_1226, w_071_1227, w_071_1228, w_071_1229, w_071_1230, w_071_1231, w_071_1232, w_071_1233, w_071_1234, w_071_1237, w_071_1238, w_071_1239, w_071_1240, w_071_1241, w_071_1242, w_071_1243, w_071_1244, w_071_1245, w_071_1247, w_071_1249, w_071_1250, w_071_1251, w_071_1252, w_071_1255, w_071_1256, w_071_1257, w_071_1259, w_071_1260, w_071_1261, w_071_1266, w_071_1267, w_071_1268, w_071_1269, w_071_1270, w_071_1271, w_071_1272, w_071_1273, w_071_1274, w_071_1275, w_071_1276, w_071_1277, w_071_1279, w_071_1280, w_071_1281, w_071_1282, w_071_1283, w_071_1285, w_071_1286, w_071_1287, w_071_1288, w_071_1289, w_071_1290, w_071_1291, w_071_1292, w_071_1293, w_071_1294, w_071_1295, w_071_1297, w_071_1298, w_071_1299, w_071_1300, w_071_1301, w_071_1302, w_071_1303, w_071_1304, w_071_1306, w_071_1307, w_071_1309, w_071_1311, w_071_1312, w_071_1314, w_071_1315, w_071_1317, w_071_1318, w_071_1320, w_071_1321, w_071_1322, w_071_1323, w_071_1324, w_071_1326, w_071_1327, w_071_1330, w_071_1332, w_071_1334, w_071_1335, w_071_1337, w_071_1338, w_071_1339, w_071_1340, w_071_1341, w_071_1342, w_071_1343, w_071_1344, w_071_1345, w_071_1346, w_071_1347, w_071_1348, w_071_1349, w_071_1350, w_071_1351, w_071_1354, w_071_1355, w_071_1356, w_071_1357, w_071_1358, w_071_1359, w_071_1360, w_071_1361, w_071_1362, w_071_1363, w_071_1364, w_071_1365, w_071_1366, w_071_1367, w_071_1368, w_071_1369, w_071_1370, w_071_1371, w_071_1372, w_071_1373, w_071_1375, w_071_1377, w_071_1378, w_071_1379, w_071_1380, w_071_1381, w_071_1382, w_071_1383, w_071_1385, w_071_1387, w_071_1388, w_071_1389, w_071_1390, w_071_1391, w_071_1394, w_071_1395, w_071_1396, w_071_1397, w_071_1398, w_071_1399, w_071_1400, w_071_1401, w_071_1403, w_071_1404, w_071_1407, w_071_1408, w_071_1409, w_071_1410, w_071_1411, w_071_1413, w_071_1414, w_071_1415, w_071_1416, w_071_1417, w_071_1419, w_071_1420, w_071_1421, w_071_1422, w_071_1423, w_071_1424, w_071_1425, w_071_1428, w_071_1429, w_071_1430, w_071_1431, w_071_1432, w_071_1434, w_071_1435, w_071_1436, w_071_1437, w_071_1438, w_071_1439, w_071_1440, w_071_1441, w_071_1442, w_071_1443, w_071_1444, w_071_1446, w_071_1448, w_071_1449, w_071_1450, w_071_1452, w_071_1454, w_071_1457, w_071_1458, w_071_1459, w_071_1460, w_071_1461, w_071_1462, w_071_1463, w_071_1464, w_071_1465, w_071_1466, w_071_1469, w_071_1470, w_071_1471, w_071_1473, w_071_1474, w_071_1476, w_071_1477, w_071_1478, w_071_1479, w_071_1480, w_071_1482, w_071_1484, w_071_1485, w_071_1486, w_071_1487, w_071_1488, w_071_1489, w_071_1491, w_071_1492, w_071_1493, w_071_1494, w_071_1495, w_071_1496, w_071_1497, w_071_1498, w_071_1499, w_071_1500, w_071_1503, w_071_1505, w_071_1506, w_071_1507, w_071_1509, w_071_1511, w_071_1512, w_071_1513, w_071_1517, w_071_1518, w_071_1519, w_071_1520, w_071_1521, w_071_1522, w_071_1523, w_071_1525, w_071_1526, w_071_1527, w_071_1528, w_071_1529, w_071_1532, w_071_1534, w_071_1535, w_071_1536, w_071_1537, w_071_1540, w_071_1542, w_071_1543, w_071_1544, w_071_1545, w_071_1546, w_071_1547, w_071_1548, w_071_1550, w_071_1551, w_071_1554, w_071_1555, w_071_1556, w_071_1557, w_071_1559, w_071_1560, w_071_1561, w_071_1562, w_071_1563, w_071_1566, w_071_1567, w_071_1568, w_071_1571, w_071_1572, w_071_1573, w_071_1574, w_071_1576, w_071_1577, w_071_1578, w_071_1579, w_071_1580, w_071_1581, w_071_1582, w_071_1583, w_071_1584, w_071_1585, w_071_1588, w_071_1589, w_071_1590, w_071_1591, w_071_1593, w_071_1594, w_071_1595, w_071_1596, w_071_1597, w_071_1598, w_071_1600, w_071_1602, w_071_1603, w_071_1605, w_071_1606, w_071_1607, w_071_1609, w_071_1611, w_071_1612, w_071_1613, w_071_1615, w_071_1618, w_071_1619, w_071_1620, w_071_1622, w_071_1623, w_071_1625, w_071_1626, w_071_1627, w_071_1628, w_071_1630, w_071_1631, w_071_1632, w_071_1633, w_071_1634, w_071_1635, w_071_1636, w_071_1637, w_071_1639, w_071_1640, w_071_1643, w_071_1644, w_071_1646, w_071_1647, w_071_1649, w_071_1650, w_071_1651, w_071_1652, w_071_1654, w_071_1655, w_071_1656, w_071_1657, w_071_1658, w_071_1662, w_071_1663, w_071_1664, w_071_1665, w_071_1668, w_071_1669, w_071_1670, w_071_1671, w_071_1672, w_071_1675, w_071_1676, w_071_1677, w_071_1680, w_071_1681, w_071_1682, w_071_1683, w_071_1684, w_071_1685, w_071_1686, w_071_1688, w_071_1689, w_071_1690, w_071_1691, w_071_1692, w_071_1693, w_071_1694, w_071_1696, w_071_1697, w_071_1698, w_071_1699, w_071_1700, w_071_1701, w_071_1702, w_071_1703, w_071_1704, w_071_1706, w_071_1707, w_071_1708, w_071_1709, w_071_1710, w_071_1711, w_071_1712, w_071_1713, w_071_1715, w_071_1716, w_071_1717, w_071_1718, w_071_1719, w_071_1720, w_071_1721, w_071_1723, w_071_1725, w_071_1727, w_071_1728, w_071_1729, w_071_1730, w_071_1731, w_071_1732, w_071_1733, w_071_1734, w_071_1735, w_071_1736, w_071_1737, w_071_1739, w_071_1740, w_071_1741, w_071_1742, w_071_1743, w_071_1747, w_071_1749, w_071_1750, w_071_1751, w_071_1753, w_071_1754, w_071_1756, w_071_1757, w_071_1758, w_071_1760, w_071_1762, w_071_1763, w_071_1764, w_071_1765, w_071_1766, w_071_1767, w_071_1768, w_071_1770, w_071_1771, w_071_1772, w_071_1773, w_071_1774, w_071_1775, w_071_1776, w_071_1777, w_071_1778, w_071_1779, w_071_1781, w_071_1784, w_071_1787, w_071_1788, w_071_1790, w_071_1791, w_071_1792, w_071_1793, w_071_1795, w_071_1796, w_071_1797, w_071_1798, w_071_1799, w_071_1803, w_071_1804, w_071_1805, w_071_1806, w_071_1807, w_071_1808, w_071_1809, w_071_1810, w_071_1812, w_071_1813, w_071_1816, w_071_1818, w_071_1820, w_071_1821, w_071_1822, w_071_1823, w_071_1824, w_071_1825, w_071_1827, w_071_1831, w_071_1833, w_071_1834, w_071_1835, w_071_1838, w_071_1839, w_071_1841, w_071_1842, w_071_1843, w_071_1844, w_071_1845, w_071_1846, w_071_1847, w_071_1848, w_071_1852, w_071_1853, w_071_1854, w_071_1855, w_071_1856, w_071_1857, w_071_1858, w_071_1860, w_071_1862, w_071_1863, w_071_1864, w_071_1865, w_071_1866, w_071_1867, w_071_1868, w_071_1869, w_071_1871, w_071_1872, w_071_1873, w_071_1874, w_071_1876, w_071_1877, w_071_1878, w_071_1880, w_071_1881, w_071_1882, w_071_1884, w_071_1885, w_071_1887, w_071_1888, w_071_1889, w_071_1890, w_071_1891, w_071_1893, w_071_1894, w_071_1895, w_071_1896, w_071_1898, w_071_1899, w_071_1900, w_071_1901, w_071_1904, w_071_1905, w_071_1906, w_071_1907, w_071_1908, w_071_1909, w_071_1910, w_071_1911, w_071_1912, w_071_1913, w_071_1914, w_071_1915, w_071_1918, w_071_1919, w_071_1920, w_071_1921, w_071_1922, w_071_1923, w_071_1924, w_071_1925, w_071_1926, w_071_1927, w_071_1928, w_071_1929, w_071_1930, w_071_1932, w_071_1933, w_071_1935, w_071_1936, w_071_1937, w_071_1939, w_071_1940, w_071_1941, w_071_1942, w_071_1944, w_071_1946, w_071_1947, w_071_1948, w_071_1949, w_071_1950, w_071_1951, w_071_1952, w_071_1953, w_071_1954, w_071_1955, w_071_1956, w_071_1957, w_071_1958, w_071_1959, w_071_1960, w_071_1961, w_071_1962, w_071_1963, w_071_1965, w_071_1966, w_071_1968, w_071_1970, w_071_1971, w_071_1973, w_071_1974, w_071_1975, w_071_1976, w_071_1977, w_071_1978, w_071_1979, w_071_1980, w_071_1981, w_071_1982, w_071_1984, w_071_1985, w_071_1986, w_071_1987, w_071_1988, w_071_1989, w_071_1990, w_071_1991, w_071_1995, w_071_1996, w_071_1997, w_071_1998, w_071_1999, w_071_2001, w_071_2002, w_071_2003, w_071_2004, w_071_2005, w_071_2006, w_071_2008, w_071_2010, w_071_2011, w_071_2012, w_071_2013, w_071_2014, w_071_2015, w_071_2018, w_071_2019, w_071_2022, w_071_2023, w_071_2024, w_071_2027, w_071_2028, w_071_2029, w_071_2030, w_071_2032, w_071_2034, w_071_2035, w_071_2038, w_071_2040, w_071_2041, w_071_2042, w_071_2044, w_071_2046, w_071_2047, w_071_2048, w_071_2049, w_071_2050, w_071_2051, w_071_2055, w_071_2058, w_071_2059, w_071_2060, w_071_2062, w_071_2063, w_071_2065, w_071_2067, w_071_2068, w_071_2069, w_071_2070, w_071_2072, w_071_2073, w_071_2074, w_071_2075, w_071_2076, w_071_2078, w_071_2079, w_071_2080, w_071_2081, w_071_2085, w_071_2086, w_071_2087, w_071_2088, w_071_2089, w_071_2090, w_071_2092, w_071_2093, w_071_2094, w_071_2095, w_071_2096, w_071_2097, w_071_2098, w_071_2099, w_071_2100, w_071_2101, w_071_2103, w_071_2104, w_071_2107, w_071_2108, w_071_2109, w_071_2110, w_071_2111, w_071_2115, w_071_2116, w_071_2117, w_071_2118, w_071_2119, w_071_2122, w_071_2124, w_071_2126, w_071_2127, w_071_2128, w_071_2129, w_071_2130, w_071_2131, w_071_2133, w_071_2134, w_071_2135, w_071_2136, w_071_2137, w_071_2139, w_071_2140, w_071_2141, w_071_2143, w_071_2144, w_071_2145, w_071_2146, w_071_2147, w_071_2148, w_071_2149, w_071_2150, w_071_2152, w_071_2155, w_071_2157, w_071_2159, w_071_2160, w_071_2161, w_071_2162, w_071_2164, w_071_2165, w_071_2168, w_071_2169, w_071_2170, w_071_2171, w_071_2172, w_071_2173, w_071_2177, w_071_2178, w_071_2180, w_071_2182, w_071_2185, w_071_2186, w_071_2188, w_071_2189, w_071_2190, w_071_2191, w_071_2192, w_071_2193, w_071_2194, w_071_2195, w_071_2198, w_071_2199, w_071_2200, w_071_2201, w_071_2202, w_071_2203, w_071_2205, w_071_2206, w_071_2207, w_071_2208, w_071_2209, w_071_2210, w_071_2211, w_071_2212, w_071_2213, w_071_2214, w_071_2215, w_071_2216, w_071_2217, w_071_2218, w_071_2219, w_071_2220, w_071_2221, w_071_2222, w_071_2224, w_071_2225, w_071_2229, w_071_2230, w_071_2232, w_071_2233, w_071_2236, w_071_2237, w_071_2238, w_071_2239, w_071_2240, w_071_2243, w_071_2244, w_071_2246, w_071_2247, w_071_2248, w_071_2249, w_071_2250, w_071_2251, w_071_2253, w_071_2254, w_071_2255, w_071_2256, w_071_2257, w_071_2258, w_071_2259, w_071_2260, w_071_2261, w_071_2263, w_071_2264, w_071_2265, w_071_2266, w_071_2267, w_071_2268, w_071_2269, w_071_2270, w_071_2271, w_071_2273, w_071_2274, w_071_2275, w_071_2276, w_071_2278, w_071_2279, w_071_2280, w_071_2282, w_071_2284, w_071_2286, w_071_2288, w_071_2291, w_071_2292, w_071_2293, w_071_2294, w_071_2295, w_071_2296, w_071_2297, w_071_2298, w_071_2299, w_071_2300, w_071_2301, w_071_2303, w_071_2304, w_071_2306, w_071_2308, w_071_2310, w_071_2311, w_071_2312, w_071_2315, w_071_2316, w_071_2318, w_071_2319, w_071_2320, w_071_2321, w_071_2322, w_071_2323, w_071_2324, w_071_2325, w_071_2326, w_071_2327, w_071_2328, w_071_2329, w_071_2330, w_071_2331, w_071_2332, w_071_2333, w_071_2335, w_071_2336, w_071_2337, w_071_2338, w_071_2339, w_071_2340, w_071_2341, w_071_2342, w_071_2343, w_071_2344, w_071_2345, w_071_2346, w_071_2347, w_071_2348, w_071_2349, w_071_2350, w_071_2351, w_071_2353, w_071_2354, w_071_2355, w_071_2356, w_071_2357, w_071_2358, w_071_2359, w_071_2360, w_071_2361, w_071_2362, w_071_2363, w_071_2365, w_071_2366, w_071_2367, w_071_2369, w_071_2370, w_071_2373, w_071_2375, w_071_2376, w_071_2378, w_071_2379, w_071_2380, w_071_2381, w_071_2382, w_071_2383, w_071_2385, w_071_2386, w_071_2387;
  wire w_072_000, w_072_002, w_072_005, w_072_006, w_072_007, w_072_009, w_072_010, w_072_011, w_072_012, w_072_014, w_072_015, w_072_016, w_072_021, w_072_022, w_072_025, w_072_026, w_072_027, w_072_029, w_072_030, w_072_031, w_072_032, w_072_034, w_072_035, w_072_036, w_072_037, w_072_039, w_072_040, w_072_044, w_072_046, w_072_047, w_072_048, w_072_049, w_072_051, w_072_055, w_072_058, w_072_060, w_072_061, w_072_062, w_072_063, w_072_064, w_072_066, w_072_069, w_072_073, w_072_075, w_072_077, w_072_081, w_072_082, w_072_085, w_072_087, w_072_093, w_072_094, w_072_096, w_072_097, w_072_098, w_072_099, w_072_102, w_072_103, w_072_107, w_072_109, w_072_110, w_072_112, w_072_114, w_072_117, w_072_118, w_072_120, w_072_121, w_072_122, w_072_124, w_072_125, w_072_128, w_072_129, w_072_133, w_072_135, w_072_136, w_072_138, w_072_140, w_072_141, w_072_142, w_072_144, w_072_156, w_072_159, w_072_161, w_072_165, w_072_166, w_072_172, w_072_174, w_072_178, w_072_182, w_072_189, w_072_192, w_072_195, w_072_199, w_072_200, w_072_202, w_072_203, w_072_204, w_072_210, w_072_213, w_072_216, w_072_219, w_072_220, w_072_223, w_072_227, w_072_228, w_072_241, w_072_243, w_072_244, w_072_246, w_072_248, w_072_254, w_072_266, w_072_269, w_072_270, w_072_271, w_072_272, w_072_273, w_072_276, w_072_278, w_072_282, w_072_283, w_072_284, w_072_285, w_072_288, w_072_292, w_072_297, w_072_298, w_072_300, w_072_302, w_072_305, w_072_310, w_072_312, w_072_314, w_072_316, w_072_318, w_072_320, w_072_325, w_072_326, w_072_327, w_072_328, w_072_332, w_072_333, w_072_340, w_072_348, w_072_349, w_072_352, w_072_357, w_072_371, w_072_373, w_072_374, w_072_375, w_072_376, w_072_377, w_072_381, w_072_388, w_072_389, w_072_390, w_072_391, w_072_398, w_072_403, w_072_406, w_072_407, w_072_416, w_072_420, w_072_428, w_072_435, w_072_437, w_072_439, w_072_440, w_072_441, w_072_444, w_072_451, w_072_457, w_072_462, w_072_474, w_072_483, w_072_489, w_072_492, w_072_493, w_072_494, w_072_496, w_072_499, w_072_500, w_072_502, w_072_503, w_072_506, w_072_507, w_072_511, w_072_512, w_072_513, w_072_519, w_072_520, w_072_521, w_072_523, w_072_524, w_072_526, w_072_532, w_072_535, w_072_542, w_072_552, w_072_557, w_072_559, w_072_564, w_072_565, w_072_572, w_072_574, w_072_576, w_072_587, w_072_588, w_072_590, w_072_592, w_072_596, w_072_598, w_072_599, w_072_600, w_072_601, w_072_603, w_072_606, w_072_607, w_072_609, w_072_610, w_072_611, w_072_614, w_072_630, w_072_632, w_072_634, w_072_638, w_072_640, w_072_644, w_072_646, w_072_648, w_072_649, w_072_651, w_072_655, w_072_662, w_072_665, w_072_667, w_072_670, w_072_673, w_072_675, w_072_679, w_072_681, w_072_685, w_072_686, w_072_691, w_072_697, w_072_698, w_072_702, w_072_703, w_072_705, w_072_707, w_072_708, w_072_710, w_072_711, w_072_713, w_072_715, w_072_725, w_072_727, w_072_728, w_072_730, w_072_737, w_072_738, w_072_748, w_072_759, w_072_760, w_072_762, w_072_763, w_072_766, w_072_770, w_072_774, w_072_777, w_072_780, w_072_783, w_072_784, w_072_793, w_072_795, w_072_796, w_072_797, w_072_802, w_072_805, w_072_806, w_072_807, w_072_808, w_072_809, w_072_817, w_072_818, w_072_819, w_072_820, w_072_821, w_072_825, w_072_826, w_072_829, w_072_830, w_072_831, w_072_833, w_072_835, w_072_840, w_072_847, w_072_848, w_072_849, w_072_853, w_072_854, w_072_856, w_072_858, w_072_868, w_072_870, w_072_871, w_072_873, w_072_877, w_072_878, w_072_879, w_072_880, w_072_886, w_072_887, w_072_888, w_072_893, w_072_895, w_072_896, w_072_898, w_072_899, w_072_900, w_072_903, w_072_905, w_072_909, w_072_913, w_072_919, w_072_925, w_072_930, w_072_931, w_072_933, w_072_942, w_072_948, w_072_949, w_072_951, w_072_953, w_072_957, w_072_961, w_072_963, w_072_965, w_072_966, w_072_968, w_072_971, w_072_972, w_072_973, w_072_982, w_072_983, w_072_987, w_072_989, w_072_992, w_072_1003, w_072_1004, w_072_1006, w_072_1007, w_072_1013, w_072_1018, w_072_1019, w_072_1021, w_072_1023, w_072_1028, w_072_1030, w_072_1033, w_072_1034, w_072_1035, w_072_1036, w_072_1037, w_072_1041, w_072_1042, w_072_1044, w_072_1045, w_072_1049, w_072_1058, w_072_1059, w_072_1061, w_072_1062, w_072_1069, w_072_1071, w_072_1072, w_072_1075, w_072_1077, w_072_1078, w_072_1081, w_072_1087, w_072_1088, w_072_1097, w_072_1101, w_072_1103, w_072_1108, w_072_1115, w_072_1116, w_072_1119, w_072_1122, w_072_1123, w_072_1125, w_072_1135, w_072_1139, w_072_1140, w_072_1141, w_072_1142, w_072_1143, w_072_1144, w_072_1148, w_072_1149, w_072_1150, w_072_1151, w_072_1156, w_072_1157, w_072_1158, w_072_1159, w_072_1160, w_072_1167, w_072_1169, w_072_1172, w_072_1182, w_072_1184, w_072_1185, w_072_1186, w_072_1188, w_072_1190, w_072_1194, w_072_1195, w_072_1205, w_072_1207, w_072_1209, w_072_1212, w_072_1213, w_072_1217, w_072_1219, w_072_1220, w_072_1222, w_072_1223, w_072_1225, w_072_1226, w_072_1228, w_072_1232, w_072_1233, w_072_1234, w_072_1235, w_072_1242, w_072_1243, w_072_1249, w_072_1252, w_072_1253, w_072_1254, w_072_1265, w_072_1266, w_072_1267, w_072_1269, w_072_1270, w_072_1271, w_072_1283, w_072_1288, w_072_1292, w_072_1294, w_072_1295, w_072_1298, w_072_1300, w_072_1301, w_072_1302, w_072_1303, w_072_1304, w_072_1307, w_072_1310, w_072_1318, w_072_1322, w_072_1325, w_072_1328, w_072_1329, w_072_1330, w_072_1335, w_072_1337, w_072_1338, w_072_1344, w_072_1351, w_072_1354, w_072_1357, w_072_1360, w_072_1366, w_072_1370, w_072_1374, w_072_1378, w_072_1381, w_072_1390, w_072_1395, w_072_1400, w_072_1403, w_072_1404, w_072_1410, w_072_1411, w_072_1413, w_072_1415, w_072_1417, w_072_1418, w_072_1422, w_072_1423, w_072_1424, w_072_1426, w_072_1427, w_072_1428, w_072_1433, w_072_1443, w_072_1444, w_072_1457, w_072_1460, w_072_1469, w_072_1470, w_072_1471, w_072_1472, w_072_1478, w_072_1479, w_072_1486, w_072_1488, w_072_1492, w_072_1495, w_072_1496, w_072_1497, w_072_1498, w_072_1500, w_072_1502, w_072_1504, w_072_1508, w_072_1512, w_072_1515, w_072_1517, w_072_1518, w_072_1521, w_072_1522, w_072_1526, w_072_1542, w_072_1548, w_072_1552, w_072_1556, w_072_1562, w_072_1564, w_072_1568, w_072_1573, w_072_1575, w_072_1582, w_072_1587, w_072_1589, w_072_1591, w_072_1593, w_072_1595, w_072_1597, w_072_1599, w_072_1613, w_072_1619, w_072_1622, w_072_1623, w_072_1624, w_072_1627, w_072_1628, w_072_1630, w_072_1634, w_072_1637, w_072_1638, w_072_1641, w_072_1649, w_072_1656, w_072_1657, w_072_1658, w_072_1666, w_072_1669, w_072_1671, w_072_1674, w_072_1679, w_072_1685, w_072_1689, w_072_1690, w_072_1694, w_072_1696, w_072_1697, w_072_1699, w_072_1701, w_072_1705, w_072_1710, w_072_1711, w_072_1716, w_072_1723, w_072_1731, w_072_1733, w_072_1739, w_072_1743, w_072_1746, w_072_1749, w_072_1754, w_072_1758, w_072_1762, w_072_1767, w_072_1768, w_072_1774, w_072_1783, w_072_1788, w_072_1791, w_072_1797, w_072_1798, w_072_1799, w_072_1806, w_072_1809, w_072_1811, w_072_1812, w_072_1813, w_072_1817, w_072_1818, w_072_1819, w_072_1834, w_072_1836, w_072_1838, w_072_1840, w_072_1845, w_072_1847, w_072_1852, w_072_1853, w_072_1856, w_072_1861, w_072_1868, w_072_1870, w_072_1878, w_072_1880, w_072_1885, w_072_1888, w_072_1892, w_072_1902, w_072_1903, w_072_1904, w_072_1915, w_072_1917, w_072_1918, w_072_1919, w_072_1928, w_072_1938, w_072_1939, w_072_1945, w_072_1947, w_072_1950, w_072_1951, w_072_1954, w_072_1955, w_072_1958, w_072_1960, w_072_1961, w_072_1969, w_072_1971, w_072_1974, w_072_1976, w_072_1980, w_072_1994, w_072_2000, w_072_2003, w_072_2008, w_072_2014, w_072_2029, w_072_2038, w_072_2041, w_072_2049, w_072_2054, w_072_2056, w_072_2067, w_072_2079, w_072_2080, w_072_2095, w_072_2096, w_072_2098, w_072_2099, w_072_2100, w_072_2105, w_072_2112, w_072_2114, w_072_2115, w_072_2116, w_072_2119, w_072_2120, w_072_2126, w_072_2129, w_072_2131, w_072_2132, w_072_2137, w_072_2140, w_072_2144, w_072_2146, w_072_2148, w_072_2149, w_072_2151, w_072_2167, w_072_2170, w_072_2171, w_072_2173, w_072_2174, w_072_2175, w_072_2176, w_072_2184, w_072_2185, w_072_2192, w_072_2195, w_072_2196, w_072_2201, w_072_2204, w_072_2208, w_072_2216, w_072_2219, w_072_2220, w_072_2222, w_072_2228, w_072_2230, w_072_2235, w_072_2242, w_072_2247, w_072_2248, w_072_2251, w_072_2252, w_072_2253, w_072_2257, w_072_2261, w_072_2262, w_072_2265, w_072_2267, w_072_2274, w_072_2275, w_072_2277, w_072_2288, w_072_2290, w_072_2292, w_072_2299, w_072_2301, w_072_2305, w_072_2308, w_072_2309, w_072_2311, w_072_2318, w_072_2319, w_072_2330, w_072_2331, w_072_2334, w_072_2339, w_072_2347, w_072_2348, w_072_2349, w_072_2351, w_072_2353, w_072_2354, w_072_2356, w_072_2366, w_072_2368, w_072_2371, w_072_2372, w_072_2373, w_072_2375, w_072_2377, w_072_2380, w_072_2383, w_072_2388, w_072_2390, w_072_2394, w_072_2399, w_072_2403, w_072_2407, w_072_2409, w_072_2412, w_072_2413, w_072_2420, w_072_2421, w_072_2424, w_072_2429, w_072_2432, w_072_2434, w_072_2435, w_072_2438, w_072_2442, w_072_2443, w_072_2444, w_072_2445, w_072_2446, w_072_2448, w_072_2453, w_072_2455, w_072_2456, w_072_2467, w_072_2468, w_072_2471, w_072_2474, w_072_2475, w_072_2476, w_072_2478, w_072_2480, w_072_2482, w_072_2484, w_072_2491, w_072_2494, w_072_2495, w_072_2501, w_072_2504, w_072_2514, w_072_2515, w_072_2519, w_072_2521, w_072_2528, w_072_2529, w_072_2530, w_072_2532, w_072_2533, w_072_2537, w_072_2545, w_072_2558, w_072_2560, w_072_2564, w_072_2566, w_072_2579, w_072_2581, w_072_2582, w_072_2586, w_072_2589, w_072_2591, w_072_2594, w_072_2601, w_072_2602, w_072_2610, w_072_2617, w_072_2622, w_072_2626, w_072_2631, w_072_2634, w_072_2635, w_072_2637, w_072_2639, w_072_2640, w_072_2646, w_072_2651, w_072_2660, w_072_2661, w_072_2664, w_072_2669, w_072_2671, w_072_2672, w_072_2673, w_072_2674, w_072_2680, w_072_2682, w_072_2683, w_072_2684, w_072_2689, w_072_2692, w_072_2694, w_072_2697, w_072_2699, w_072_2701, w_072_2708, w_072_2709, w_072_2710, w_072_2711, w_072_2715, w_072_2717, w_072_2722, w_072_2725, w_072_2727, w_072_2729, w_072_2743, w_072_2749, w_072_2753, w_072_2756, w_072_2757, w_072_2758, w_072_2759, w_072_2761, w_072_2764, w_072_2766, w_072_2767, w_072_2773, w_072_2775, w_072_2782, w_072_2793, w_072_2798, w_072_2804, w_072_2813, w_072_2814, w_072_2815, w_072_2816, w_072_2817, w_072_2818, w_072_2819, w_072_2821, w_072_2824, w_072_2827, w_072_2833, w_072_2839, w_072_2851, w_072_2852, w_072_2855, w_072_2856, w_072_2861, w_072_2863, w_072_2865, w_072_2866, w_072_2872, w_072_2876, w_072_2877, w_072_2884, w_072_2886, w_072_2887, w_072_2890, w_072_2892, w_072_2895, w_072_2897, w_072_2898, w_072_2901, w_072_2907, w_072_2911, w_072_2917, w_072_2918, w_072_2920, w_072_2928, w_072_2931, w_072_2932, w_072_2939, w_072_2944, w_072_2949, w_072_2950, w_072_2954, w_072_2957, w_072_2961, w_072_2962, w_072_2968, w_072_2972, w_072_2979, w_072_2982, w_072_2984, w_072_2985, w_072_2993, w_072_2995, w_072_3000, w_072_3006, w_072_3009, w_072_3011, w_072_3013, w_072_3014, w_072_3015, w_072_3016, w_072_3017, w_072_3018, w_072_3021, w_072_3022, w_072_3024, w_072_3030, w_072_3031, w_072_3033, w_072_3034, w_072_3039, w_072_3041, w_072_3043, w_072_3045, w_072_3053, w_072_3057, w_072_3059, w_072_3061, w_072_3062, w_072_3065, w_072_3066, w_072_3067, w_072_3068, w_072_3069, w_072_3070, w_072_3072, w_072_3074, w_072_3076, w_072_3078, w_072_3079, w_072_3084, w_072_3086, w_072_3087, w_072_3088, w_072_3090, w_072_3091, w_072_3092, w_072_3093, w_072_3094, w_072_3098, w_072_3101, w_072_3105, w_072_3106, w_072_3107, w_072_3109, w_072_3110, w_072_3111, w_072_3120, w_072_3122, w_072_3127, w_072_3128, w_072_3134, w_072_3136, w_072_3137, w_072_3142, w_072_3146, w_072_3149, w_072_3151, w_072_3156, w_072_3161, w_072_3169, w_072_3171, w_072_3176, w_072_3177, w_072_3181, w_072_3184, w_072_3186, w_072_3195, w_072_3199, w_072_3201, w_072_3203, w_072_3208, w_072_3211, w_072_3214, w_072_3217, w_072_3220, w_072_3224, w_072_3234, w_072_3236, w_072_3237, w_072_3244, w_072_3246, w_072_3250, w_072_3258, w_072_3259, w_072_3261, w_072_3263, w_072_3265, w_072_3268, w_072_3273, w_072_3275, w_072_3276, w_072_3277, w_072_3278, w_072_3283, w_072_3285, w_072_3289, w_072_3293, w_072_3294, w_072_3296, w_072_3297, w_072_3303, w_072_3304, w_072_3308, w_072_3309, w_072_3310, w_072_3311, w_072_3313, w_072_3315, w_072_3316, w_072_3318, w_072_3320, w_072_3321, w_072_3322, w_072_3323, w_072_3324, w_072_3325, w_072_3326, w_072_3330, w_072_3332, w_072_3339, w_072_3344, w_072_3346, w_072_3349, w_072_3350, w_072_3352, w_072_3355, w_072_3356, w_072_3364, w_072_3369, w_072_3371, w_072_3372, w_072_3377, w_072_3381, w_072_3384, w_072_3385, w_072_3388, w_072_3394, w_072_3396, w_072_3408, w_072_3410, w_072_3414, w_072_3415, w_072_3417, w_072_3422, w_072_3424, w_072_3425, w_072_3427, w_072_3430, w_072_3431, w_072_3434, w_072_3435, w_072_3437, w_072_3440, w_072_3441, w_072_3442, w_072_3443, w_072_3445, w_072_3446, w_072_3449, w_072_3451, w_072_3453, w_072_3461, w_072_3463, w_072_3465, w_072_3468, w_072_3470, w_072_3471, w_072_3473, w_072_3476, w_072_3481, w_072_3494, w_072_3497, w_072_3498, w_072_3502, w_072_3507, w_072_3510, w_072_3523, w_072_3524, w_072_3527, w_072_3530, w_072_3534, w_072_3538, w_072_3540, w_072_3541, w_072_3543, w_072_3545, w_072_3546, w_072_3552, w_072_3562, w_072_3565, w_072_3566, w_072_3571, w_072_3573, w_072_3577, w_072_3579, w_072_3580, w_072_3583, w_072_3584, w_072_3588, w_072_3590, w_072_3592, w_072_3598, w_072_3608, w_072_3609, w_072_3610, w_072_3612, w_072_3613, w_072_3614, w_072_3618, w_072_3632, w_072_3635, w_072_3636, w_072_3637, w_072_3639, w_072_3640, w_072_3643, w_072_3646, w_072_3647, w_072_3649, w_072_3653, w_072_3654, w_072_3656, w_072_3659, w_072_3661, w_072_3662, w_072_3664, w_072_3665, w_072_3668, w_072_3673, w_072_3674, w_072_3675, w_072_3676, w_072_3679, w_072_3682, w_072_3689, w_072_3693, w_072_3695, w_072_3696, w_072_3700, w_072_3701, w_072_3702, w_072_3705, w_072_3707, w_072_3709, w_072_3711, w_072_3713, w_072_3723, w_072_3727, w_072_3728, w_072_3729, w_072_3730, w_072_3736, w_072_3737, w_072_3738, w_072_3742, w_072_3743, w_072_3745, w_072_3748, w_072_3751, w_072_3759, w_072_3761, w_072_3762, w_072_3763, w_072_3764, w_072_3765, w_072_3766, w_072_3768, w_072_3773, w_072_3774, w_072_3777, w_072_3779, w_072_3790, w_072_3791, w_072_3795, w_072_3796, w_072_3798, w_072_3803, w_072_3804, w_072_3805, w_072_3808, w_072_3812, w_072_3813, w_072_3814, w_072_3816, w_072_3817, w_072_3819, w_072_3822, w_072_3824, w_072_3830, w_072_3831, w_072_3834, w_072_3835, w_072_3836, w_072_3842, w_072_3846, w_072_3847, w_072_3856, w_072_3862, w_072_3863, w_072_3867, w_072_3874, w_072_3875, w_072_3876, w_072_3877, w_072_3878, w_072_3879, w_072_3883, w_072_3887, w_072_3901, w_072_3904, w_072_3909, w_072_3911, w_072_3914, w_072_3918, w_072_3921, w_072_3922, w_072_3924, w_072_3931, w_072_3944, w_072_3949, w_072_3950, w_072_3951, w_072_3952, w_072_3955, w_072_3959, w_072_3966, w_072_3969, w_072_3970, w_072_3973, w_072_3978, w_072_3981, w_072_3984, w_072_3994, w_072_3995, w_072_4000, w_072_4013, w_072_4014, w_072_4016, w_072_4025, w_072_4026, w_072_4027, w_072_4029, w_072_4038, w_072_4041, w_072_4042, w_072_4044, w_072_4045, w_072_4054, w_072_4059, w_072_4062, w_072_4065, w_072_4068, w_072_4069, w_072_4075, w_072_4079, w_072_4085, w_072_4089, w_072_4092, w_072_4109, w_072_4110, w_072_4112, w_072_4118, w_072_4120, w_072_4121, w_072_4123, w_072_4125, w_072_4127, w_072_4130, w_072_4137, w_072_4138, w_072_4140, w_072_4142, w_072_4144, w_072_4148, w_072_4158, w_072_4159, w_072_4162, w_072_4167, w_072_4172, w_072_4176, w_072_4180, w_072_4181, w_072_4182, w_072_4192, w_072_4196, w_072_4202, w_072_4207, w_072_4210, w_072_4222, w_072_4223, w_072_4226, w_072_4228, w_072_4243, w_072_4244, w_072_4249, w_072_4251, w_072_4255, w_072_4257, w_072_4260, w_072_4261, w_072_4267, w_072_4274, w_072_4278, w_072_4280, w_072_4281, w_072_4284, w_072_4291, w_072_4295, w_072_4300, w_072_4301, w_072_4302, w_072_4305, w_072_4306, w_072_4307, w_072_4309, w_072_4311, w_072_4314, w_072_4316, w_072_4318, w_072_4320, w_072_4323, w_072_4325, w_072_4326, w_072_4331, w_072_4332, w_072_4333, w_072_4337, w_072_4338, w_072_4345, w_072_4351, w_072_4359, w_072_4364, w_072_4367, w_072_4369, w_072_4372, w_072_4373, w_072_4376, w_072_4378, w_072_4380, w_072_4388, w_072_4389, w_072_4393, w_072_4395, w_072_4396, w_072_4397, w_072_4399, w_072_4400, w_072_4405, w_072_4412, w_072_4416, w_072_4418, w_072_4427, w_072_4428, w_072_4430, w_072_4432, w_072_4434, w_072_4436, w_072_4446, w_072_4447, w_072_4448, w_072_4451, w_072_4462, w_072_4467, w_072_4468, w_072_4472, w_072_4475, w_072_4479, w_072_4483, w_072_4484, w_072_4487, w_072_4491, w_072_4492, w_072_4494, w_072_4495, w_072_4496, w_072_4513, w_072_4517, w_072_4519, w_072_4521, w_072_4528, w_072_4530, w_072_4539, w_072_4542, w_072_4544, w_072_4545, w_072_4547, w_072_4549, w_072_4561, w_072_4564, w_072_4569, w_072_4570, w_072_4571, w_072_4574, w_072_4575, w_072_4577, w_072_4580, w_072_4582, w_072_4586, w_072_4587, w_072_4591, w_072_4592, w_072_4593, w_072_4595, w_072_4597, w_072_4599, w_072_4608, w_072_4612, w_072_4613, w_072_4614, w_072_4616, w_072_4620, w_072_4639, w_072_4641, w_072_4642, w_072_4646, w_072_4653, w_072_4655, w_072_4662, w_072_4666, w_072_4667, w_072_4669, w_072_4677, w_072_4682, w_072_4689, w_072_4692, w_072_4695, w_072_4698, w_072_4699, w_072_4703, w_072_4706, w_072_4710, w_072_4713, w_072_4715, w_072_4722, w_072_4724, w_072_4726, w_072_4729, w_072_4730, w_072_4734, w_072_4735, w_072_4736, w_072_4737, w_072_4742, w_072_4749, w_072_4751, w_072_4752, w_072_4755, w_072_4757, w_072_4758, w_072_4759, w_072_4765, w_072_4766, w_072_4769, w_072_4770, w_072_4774, w_072_4775, w_072_4779, w_072_4784, w_072_4785, w_072_4793, w_072_4795, w_072_4797, w_072_4799, w_072_4800, w_072_4801, w_072_4802, w_072_4804, w_072_4815, w_072_4817, w_072_4818, w_072_4819, w_072_4821, w_072_4822, w_072_4825, w_072_4829, w_072_4830, w_072_4833, w_072_4835, w_072_4836, w_072_4837, w_072_4840, w_072_4851, w_072_4852, w_072_4853, w_072_4856, w_072_4865, w_072_4866, w_072_4870, w_072_4871, w_072_4874, w_072_4883, w_072_4892, w_072_4895, w_072_4896, w_072_4901, w_072_4904, w_072_4905, w_072_4906, w_072_4909, w_072_4913, w_072_4928, w_072_4930, w_072_4934, w_072_4940, w_072_4944, w_072_4947, w_072_4951, w_072_4962, w_072_4963, w_072_4968, w_072_4971, w_072_4979, w_072_4985, w_072_4989, w_072_4995, w_072_4996, w_072_5005, w_072_5009, w_072_5013, w_072_5017, w_072_5019, w_072_5020, w_072_5021, w_072_5022, w_072_5024, w_072_5026, w_072_5027, w_072_5031, w_072_5034, w_072_5036, w_072_5037, w_072_5041, w_072_5043, w_072_5052, w_072_5058, w_072_5060, w_072_5066, w_072_5067, w_072_5069, w_072_5075, w_072_5077, w_072_5079, w_072_5082, w_072_5089, w_072_5092, w_072_5093, w_072_5096, w_072_5100, w_072_5101, w_072_5102, w_072_5108, w_072_5115, w_072_5119, w_072_5120, w_072_5121, w_072_5124, w_072_5126, w_072_5127, w_072_5128, w_072_5132, w_072_5136, w_072_5137, w_072_5138, w_072_5139, w_072_5150, w_072_5151, w_072_5152, w_072_5155, w_072_5157, w_072_5160, w_072_5168, w_072_5170, w_072_5171, w_072_5175, w_072_5176, w_072_5179, w_072_5182, w_072_5192, w_072_5197, w_072_5200, w_072_5201, w_072_5203, w_072_5209, w_072_5212, w_072_5215, w_072_5217, w_072_5225, w_072_5228, w_072_5235, w_072_5236, w_072_5237, w_072_5238, w_072_5239, w_072_5240, w_072_5241, w_072_5243, w_072_5244, w_072_5245, w_072_5247, w_072_5253, w_072_5256, w_072_5262, w_072_5269, w_072_5270, w_072_5274, w_072_5279, w_072_5280, w_072_5281, w_072_5285, w_072_5289, w_072_5292, w_072_5299, w_072_5304, w_072_5309, w_072_5316, w_072_5319, w_072_5327, w_072_5330, w_072_5332, w_072_5334, w_072_5335, w_072_5338, w_072_5339, w_072_5340, w_072_5343, w_072_5345, w_072_5346, w_072_5348, w_072_5349, w_072_5350, w_072_5351, w_072_5353, w_072_5360, w_072_5361, w_072_5368, w_072_5370, w_072_5375, w_072_5380, w_072_5382, w_072_5387, w_072_5388, w_072_5391, w_072_5395, w_072_5397, w_072_5402, w_072_5403, w_072_5404, w_072_5407, w_072_5411, w_072_5412, w_072_5413, w_072_5429, w_072_5432, w_072_5433, w_072_5436, w_072_5439, w_072_5442, w_072_5447, w_072_5449, w_072_5453, w_072_5454, w_072_5455, w_072_5458, w_072_5459, w_072_5460, w_072_5461, w_072_5464, w_072_5467, w_072_5470, w_072_5471, w_072_5472, w_072_5473, w_072_5474, w_072_5477, w_072_5480, w_072_5485, w_072_5487, w_072_5488, w_072_5493, w_072_5500, w_072_5501, w_072_5504, w_072_5506, w_072_5508, w_072_5509, w_072_5510, w_072_5515, w_072_5516, w_072_5519, w_072_5522, w_072_5523, w_072_5524, w_072_5530, w_072_5533, w_072_5538, w_072_5539, w_072_5542, w_072_5543, w_072_5545, w_072_5558, w_072_5563, w_072_5568, w_072_5570, w_072_5571, w_072_5574, w_072_5582, w_072_5586, w_072_5591, w_072_5592, w_072_5596, w_072_5597, w_072_5599, w_072_5600, w_072_5603, w_072_5606, w_072_5607, w_072_5608, w_072_5614, w_072_5617, w_072_5618, w_072_5623, w_072_5627, w_072_5633, w_072_5634, w_072_5637, w_072_5638, w_072_5648, w_072_5649, w_072_5650, w_072_5659, w_072_5662, w_072_5665, w_072_5671, w_072_5675, w_072_5682, w_072_5683, w_072_5686, w_072_5687, w_072_5689, w_072_5691, w_072_5692, w_072_5694, w_072_5697, w_072_5706, w_072_5709, w_072_5711, w_072_5717, w_072_5720, w_072_5725, w_072_5727, w_072_5728, w_072_5729, w_072_5735, w_072_5739, w_072_5740, w_072_5741, w_072_5744, w_072_5747, w_072_5751, w_072_5756, w_072_5760, w_072_5765, w_072_5767, w_072_5768, w_072_5770, w_072_5773, w_072_5775, w_072_5778, w_072_5783, w_072_5796, w_072_5797, w_072_5805, w_072_5807, w_072_5812, w_072_5816, w_072_5818, w_072_5819, w_072_5820, w_072_5826, w_072_5827, w_072_5830, w_072_5832, w_072_5833, w_072_5838, w_072_5843, w_072_5844, w_072_5848, w_072_5850, w_072_5855, w_072_5858, w_072_5866, w_072_5872, w_072_5879, w_072_5882, w_072_5887, w_072_5891, w_072_5900, w_072_5901, w_072_5903, w_072_5905, w_072_5906, w_072_5915, w_072_5931, w_072_5932, w_072_5933, w_072_5937, w_072_5939, w_072_5941, w_072_5943, w_072_5945, w_072_5947, w_072_5953, w_072_5959, w_072_5960, w_072_5965, w_072_5967, w_072_5970, w_072_5975, w_072_5976, w_072_5977, w_072_5978, w_072_5980, w_072_5983, w_072_5984, w_072_5988, w_072_5989, w_072_5990, w_072_5991, w_072_5996, w_072_6002, w_072_6009, w_072_6013, w_072_6014, w_072_6016, w_072_6023, w_072_6026, w_072_6029, w_072_6030, w_072_6034, w_072_6036, w_072_6037, w_072_6039, w_072_6042, w_072_6044, w_072_6050, w_072_6051, w_072_6056, w_072_6061, w_072_6065, w_072_6066, w_072_6069, w_072_6072, w_072_6074, w_072_6080, w_072_6081, w_072_6086, w_072_6088, w_072_6092, w_072_6093, w_072_6094, w_072_6099, w_072_6102, w_072_6108, w_072_6110, w_072_6111, w_072_6112, w_072_6115, w_072_6118, w_072_6122, w_072_6123, w_072_6124, w_072_6127, w_072_6133, w_072_6141, w_072_6142, w_072_6150, w_072_6154, w_072_6155, w_072_6158, w_072_6159, w_072_6164, w_072_6167, w_072_6173, w_072_6176, w_072_6177, w_072_6178, w_072_6179, w_072_6183, w_072_6185, w_072_6188, w_072_6189, w_072_6191, w_072_6205, w_072_6209, w_072_6215, w_072_6216, w_072_6218, w_072_6227, w_072_6229, w_072_6233, w_072_6235, w_072_6236, w_072_6248, w_072_6250, w_072_6264, w_072_6265, w_072_6266, w_072_6271, w_072_6278, w_072_6282, w_072_6284, w_072_6289, w_072_6290, w_072_6293, w_072_6298, w_072_6300, w_072_6302, w_072_6303, w_072_6306, w_072_6311, w_072_6321, w_072_6330, w_072_6336, w_072_6339, w_072_6340, w_072_6341, w_072_6342, w_072_6343, w_072_6345, w_072_6354, w_072_6359, w_072_6360, w_072_6363, w_072_6365, w_072_6378, w_072_6380, w_072_6381, w_072_6382, w_072_6383, w_072_6388, w_072_6393, w_072_6398, w_072_6406, w_072_6410, w_072_6411, w_072_6418, w_072_6422, w_072_6423, w_072_6424, w_072_6432, w_072_6433, w_072_6434, w_072_6446, w_072_6447, w_072_6448, w_072_6450, w_072_6452, w_072_6455, w_072_6456, w_072_6461, w_072_6462, w_072_6465, w_072_6467, w_072_6471, w_072_6473, w_072_6474, w_072_6477, w_072_6480, w_072_6483, w_072_6489, w_072_6492, w_072_6493, w_072_6500, w_072_6502, w_072_6506, w_072_6507, w_072_6513, w_072_6517, w_072_6518, w_072_6519, w_072_6520, w_072_6523, w_072_6528, w_072_6531, w_072_6534, w_072_6540, w_072_6547, w_072_6548, w_072_6554, w_072_6555, w_072_6560, w_072_6565, w_072_6566, w_072_6570, w_072_6572, w_072_6574, w_072_6576, w_072_6578, w_072_6580, w_072_6581, w_072_6583, w_072_6585, w_072_6586, w_072_6591, w_072_6596, w_072_6602, w_072_6604, w_072_6606, w_072_6607, w_072_6608, w_072_6609, w_072_6610, w_072_6614, w_072_6616, w_072_6617, w_072_6622, w_072_6628, w_072_6632, w_072_6633, w_072_6643, w_072_6649, w_072_6652, w_072_6655, w_072_6659, w_072_6662, w_072_6663, w_072_6665, w_072_6667, w_072_6669, w_072_6673, w_072_6674, w_072_6677, w_072_6680, w_072_6683, w_072_6687, w_072_6694, w_072_6695, w_072_6696, w_072_6702, w_072_6707, w_072_6713, w_072_6714, w_072_6719, w_072_6720, w_072_6721, w_072_6722, w_072_6726, w_072_6739, w_072_6741, w_072_6751, w_072_6753, w_072_6755, w_072_6759, w_072_6760, w_072_6770, w_072_6771, w_072_6775, w_072_6783, w_072_6786, w_072_6789, w_072_6792, w_072_6793, w_072_6794, w_072_6795, w_072_6805, w_072_6806, w_072_6807, w_072_6811, w_072_6812, w_072_6813, w_072_6814, w_072_6816, w_072_6817, w_072_6819, w_072_6822, w_072_6823, w_072_6826, w_072_6830, w_072_6842, w_072_6845, w_072_6846, w_072_6847, w_072_6851, w_072_6858, w_072_6859, w_072_6860, w_072_6868, w_072_6871, w_072_6879, w_072_6880, w_072_6882, w_072_6883, w_072_6886, w_072_6889, w_072_6893, w_072_6894, w_072_6895, w_072_6897, w_072_6900, w_072_6902, w_072_6903, w_072_6905, w_072_6906, w_072_6907, w_072_6908, w_072_6909, w_072_6911, w_072_6914, w_072_6917, w_072_6918, w_072_6926, w_072_6927, w_072_6933, w_072_6934, w_072_6937, w_072_6944, w_072_6945, w_072_6951, w_072_6957, w_072_6958, w_072_6959, w_072_6965, w_072_6968, w_072_6970, w_072_6971, w_072_6972, w_072_6980, w_072_6982, w_072_6984, w_072_6986, w_072_6987, w_072_6988, w_072_6990, w_072_6991, w_072_6992, w_072_7004, w_072_7008, w_072_7009, w_072_7010, w_072_7011, w_072_7015, w_072_7019, w_072_7025, w_072_7027, w_072_7029, w_072_7032, w_072_7039, w_072_7040, w_072_7042, w_072_7043, w_072_7048, w_072_7049, w_072_7056, w_072_7060, w_072_7064, w_072_7067, w_072_7069, w_072_7072, w_072_7082, w_072_7085, w_072_7088, w_072_7093, w_072_7094, w_072_7100, w_072_7106, w_072_7108, w_072_7110, w_072_7112, w_072_7113, w_072_7115, w_072_7116, w_072_7119, w_072_7120, w_072_7128, w_072_7129, w_072_7131, w_072_7132, w_072_7135, w_072_7137, w_072_7141, w_072_7142, w_072_7143, w_072_7149, w_072_7151, w_072_7157, w_072_7159, w_072_7162, w_072_7177, w_072_7179, w_072_7184, w_072_7189, w_072_7194, w_072_7198, w_072_7213, w_072_7216, w_072_7217, w_072_7219, w_072_7220, w_072_7222, w_072_7223, w_072_7224, w_072_7226, w_072_7227, w_072_7234, w_072_7235, w_072_7236, w_072_7238, w_072_7239, w_072_7241, w_072_7247, w_072_7249, w_072_7252, w_072_7257, w_072_7264, w_072_7270, w_072_7271, w_072_7273, w_072_7276, w_072_7281, w_072_7282, w_072_7283, w_072_7287, w_072_7293, w_072_7297, w_072_7299, w_072_7302, w_072_7303, w_072_7304, w_072_7309, w_072_7311, w_072_7312, w_072_7323, w_072_7324, w_072_7329, w_072_7335, w_072_7340, w_072_7342, w_072_7343, w_072_7346, w_072_7349, w_072_7354, w_072_7355, w_072_7359, w_072_7364, w_072_7369, w_072_7372, w_072_7376, w_072_7385, w_072_7386, w_072_7393, w_072_7397, w_072_7401, w_072_7402, w_072_7406, w_072_7407, w_072_7409, w_072_7410, w_072_7411, w_072_7417, w_072_7419, w_072_7420, w_072_7421, w_072_7423, w_072_7424, w_072_7427, w_072_7431, w_072_7434, w_072_7436, w_072_7440, w_072_7442, w_072_7450, w_072_7454, w_072_7460, w_072_7461, w_072_7462, w_072_7463, w_072_7464, w_072_7468, w_072_7471, w_072_7476, w_072_7480, w_072_7481, w_072_7484, w_072_7490, w_072_7491, w_072_7493, w_072_7497, w_072_7500, w_072_7513, w_072_7514, w_072_7516, w_072_7517, w_072_7518, w_072_7519, w_072_7520, w_072_7523, w_072_7532, w_072_7534, w_072_7538, w_072_7539, w_072_7540, w_072_7549, w_072_7550, w_072_7553, w_072_7554, w_072_7555, w_072_7556, w_072_7558, w_072_7559, w_072_7563, w_072_7566, w_072_7567, w_072_7569, w_072_7572, w_072_7577, w_072_7580, w_072_7584, w_072_7588, w_072_7592, w_072_7595, w_072_7599, w_072_7602, w_072_7607, w_072_7608, w_072_7611, w_072_7612, w_072_7613, w_072_7615, w_072_7617, w_072_7624, w_072_7627, w_072_7629, w_072_7630, w_072_7638, w_072_7640, w_072_7647, w_072_7656, w_072_7662, w_072_7663, w_072_7668, w_072_7669, w_072_7670, w_072_7676, w_072_7681, w_072_7690, w_072_7692, w_072_7693, w_072_7694, w_072_7696, w_072_7698, w_072_7700, w_072_7702, w_072_7709, w_072_7710, w_072_7715, w_072_7719, w_072_7723, w_072_7725, w_072_7727, w_072_7735, w_072_7737, w_072_7749, w_072_7750, w_072_7754, w_072_7755, w_072_7758, w_072_7759, w_072_7762, w_072_7766, w_072_7771, w_072_7773, w_072_7774, w_072_7777, w_072_7781, w_072_7782, w_072_7788, w_072_7790, w_072_7791, w_072_7792, w_072_7793, w_072_7795, w_072_7796, w_072_7799, w_072_7801, w_072_7804, w_072_7805, w_072_7807, w_072_7808, w_072_7810, w_072_7811, w_072_7818, w_072_7824, w_072_7828, w_072_7834, w_072_7835, w_072_7838, w_072_7839, w_072_7844, w_072_7845, w_072_7846, w_072_7848, w_072_7849, w_072_7852, w_072_7853, w_072_7854, w_072_7855, w_072_7860, w_072_7861, w_072_7865, w_072_7869, w_072_7872, w_072_7876, w_072_7877, w_072_7882, w_072_7887, w_072_7888, w_072_7890, w_072_7899, w_072_7902, w_072_7903, w_072_7906, w_072_7912, w_072_7913, w_072_7915, w_072_7925, w_072_7935, w_072_7936, w_072_7937, w_072_7941, w_072_7942, w_072_7943, w_072_7952, w_072_7954, w_072_7958, w_072_7961, w_072_7967, w_072_7970, w_072_7975, w_072_7982, w_072_7987, w_072_7990, w_072_7993, w_072_7994, w_072_7996, w_072_8002, w_072_8003, w_072_8004, w_072_8007, w_072_8008, w_072_8013, w_072_8014, w_072_8017, w_072_8020, w_072_8022, w_072_8026, w_072_8027, w_072_8028, w_072_8033, w_072_8034, w_072_8044, w_072_8047, w_072_8048, w_072_8050, w_072_8051, w_072_8058, w_072_8060, w_072_8061, w_072_8063, w_072_8065, w_072_8066, w_072_8073, w_072_8075, w_072_8076, w_072_8081, w_072_8082, w_072_8088, w_072_8093, w_072_8095, w_072_8097, w_072_8101, w_072_8106, w_072_8108, w_072_8109, w_072_8114, w_072_8118, w_072_8120, w_072_8121, w_072_8123, w_072_8124, w_072_8129, w_072_8130, w_072_8134, w_072_8142, w_072_8143, w_072_8146, w_072_8150, w_072_8153, w_072_8154, w_072_8155, w_072_8158, w_072_8165, w_072_8168, w_072_8177, w_072_8178, w_072_8187, w_072_8194, w_072_8195, w_072_8196, w_072_8197, w_072_8199, w_072_8200, w_072_8203, w_072_8205, w_072_8207, w_072_8214, w_072_8215, w_072_8217, w_072_8218, w_072_8221, w_072_8226, w_072_8235, w_072_8236, w_072_8238, w_072_8239, w_072_8241, w_072_8244, w_072_8252, w_072_8254, w_072_8260, w_072_8261, w_072_8262, w_072_8266, w_072_8267, w_072_8269, w_072_8272, w_072_8276, w_072_8277, w_072_8279, w_072_8284, w_072_8286, w_072_8287, w_072_8294, w_072_8297, w_072_8299, w_072_8302, w_072_8309, w_072_8310, w_072_8311, w_072_8312, w_072_8313, w_072_8318, w_072_8320, w_072_8322, w_072_8324, w_072_8325, w_072_8326, w_072_8332, w_072_8337, w_072_8346, w_072_8350, w_072_8358, w_072_8364, w_072_8370, w_072_8371, w_072_8377, w_072_8380, w_072_8381, w_072_8391, w_072_8395, w_072_8397, w_072_8398, w_072_8403, w_072_8415, w_072_8417, w_072_8418, w_072_8425, w_072_8427, w_072_8428, w_072_8429, w_072_8431, w_072_8433, w_072_8439, w_072_8443, w_072_8445, w_072_8450, w_072_8454, w_072_8459, w_072_8461, w_072_8463, w_072_8464, w_072_8469, w_072_8470, w_072_8473, w_072_8477, w_072_8479, w_072_8483, w_072_8485, w_072_8486, w_072_8487, w_072_8489, w_072_8490, w_072_8492, w_072_8498, w_072_8501, w_072_8504, w_072_8505, w_072_8510, w_072_8516, w_072_8517, w_072_8518, w_072_8523, w_072_8524, w_072_8526, w_072_8527, w_072_8528, w_072_8529, w_072_8530, w_072_8535, w_072_8538, w_072_8539, w_072_8548, w_072_8549, w_072_8555, w_072_8558, w_072_8559, w_072_8562, w_072_8564, w_072_8567, w_072_8576, w_072_8578, w_072_8579, w_072_8583, w_072_8584, w_072_8595, w_072_8596, w_072_8600, w_072_8603, w_072_8604, w_072_8605, w_072_8606, w_072_8607, w_072_8610, w_072_8617, w_072_8618, w_072_8622, w_072_8623, w_072_8624, w_072_8627, w_072_8632, w_072_8636, w_072_8638, w_072_8639, w_072_8641, w_072_8646, w_072_8650, w_072_8656, w_072_8658, w_072_8663, w_072_8665, w_072_8674, w_072_8675, w_072_8679, w_072_8684, w_072_8693, w_072_8695, w_072_8702, w_072_8708, w_072_8710, w_072_8711, w_072_8714, w_072_8727, w_072_8729, w_072_8730, w_072_8732, w_072_8734, w_072_8735, w_072_8736, w_072_8741, w_072_8750, w_072_8752, w_072_8755, w_072_8758, w_072_8761, w_072_8763, w_072_8766, w_072_8768, w_072_8770, w_072_8771, w_072_8773, w_072_8774, w_072_8776, w_072_8779, w_072_8780, w_072_8783, w_072_8785, w_072_8786, w_072_8794, w_072_8797, w_072_8801, w_072_8803, w_072_8804, w_072_8807, w_072_8809, w_072_8812, w_072_8816, w_072_8817, w_072_8818, w_072_8820, w_072_8822, w_072_8823, w_072_8825, w_072_8826, w_072_8836, w_072_8840, w_072_8847, w_072_8851, w_072_8852, w_072_8854, w_072_8855, w_072_8856, w_072_8859, w_072_8860, w_072_8865, w_072_8866, w_072_8867, w_072_8868, w_072_8869, w_072_8884, w_072_8886, w_072_8889, w_072_8893, w_072_8898, w_072_8902, w_072_8905, w_072_8907, w_072_8910, w_072_8919, w_072_8923, w_072_8925, w_072_8931, w_072_8934, w_072_8936, w_072_8938, w_072_8939, w_072_8942, w_072_8943, w_072_8948, w_072_8952, w_072_8955, w_072_8957, w_072_8966, w_072_8975, w_072_8976, w_072_8977, w_072_8978, w_072_8982, w_072_8985, w_072_8986, w_072_8989, w_072_8990, w_072_8995, w_072_9001, w_072_9004, w_072_9005, w_072_9008, w_072_9017, w_072_9019, w_072_9020, w_072_9023, w_072_9024, w_072_9026, w_072_9029, w_072_9035, w_072_9037, w_072_9040, w_072_9047, w_072_9048, w_072_9051, w_072_9053, w_072_9058, w_072_9060, w_072_9061, w_072_9069, w_072_9071, w_072_9073, w_072_9075, w_072_9081, w_072_9084, w_072_9086, w_072_9088, w_072_9092, w_072_9094, w_072_9097, w_072_9098, w_072_9106, w_072_9107, w_072_9109, w_072_9110, w_072_9113, w_072_9114, w_072_9118, w_072_9121, w_072_9124, w_072_9127, w_072_9131, w_072_9133, w_072_9140, w_072_9143, w_072_9145, w_072_9150, w_072_9151, w_072_9156, w_072_9163, w_072_9166, w_072_9167, w_072_9168, w_072_9171, w_072_9174, w_072_9177, w_072_9178, w_072_9182, w_072_9185, w_072_9187, w_072_9188, w_072_9189, w_072_9191, w_072_9192, w_072_9194, w_072_9202, w_072_9203, w_072_9208, w_072_9212, w_072_9217, w_072_9220, w_072_9228, w_072_9229, w_072_9230, w_072_9232, w_072_9239, w_072_9242, w_072_9247, w_072_9252, w_072_9258, w_072_9264, w_072_9267, w_072_9269, w_072_9270, w_072_9271, w_072_9274, w_072_9277, w_072_9283, w_072_9285, w_072_9289, w_072_9298, w_072_9299, w_072_9302, w_072_9303, w_072_9304, w_072_9310, w_072_9313, w_072_9316, w_072_9317, w_072_9320, w_072_9322, w_072_9323, w_072_9325, w_072_9327, w_072_9329, w_072_9333, w_072_9337, w_072_9338, w_072_9343, w_072_9345, w_072_9349, w_072_9360, w_072_9361, w_072_9367, w_072_9382, w_072_9383, w_072_9384, w_072_9391, w_072_9398, w_072_9400, w_072_9413, w_072_9416, w_072_9421, w_072_9425, w_072_9426, w_072_9429, w_072_9431, w_072_9433, w_072_9435, w_072_9436, w_072_9437, w_072_9438, w_072_9439, w_072_9444, w_072_9446, w_072_9448, w_072_9449, w_072_9457, w_072_9459, w_072_9460, w_072_9461, w_072_9465, w_072_9467, w_072_9468, w_072_9470, w_072_9471, w_072_9472, w_072_9473, w_072_9479, w_072_9481, w_072_9482, w_072_9486, w_072_9493, w_072_9501, w_072_9505, w_072_9508, w_072_9510, w_072_9512, w_072_9517, w_072_9533, w_072_9535, w_072_9536, w_072_9542, w_072_9543, w_072_9544, w_072_9548, w_072_9556, w_072_9557, w_072_9559, w_072_9569, w_072_9570, w_072_9571, w_072_9576, w_072_9577, w_072_9580, w_072_9581, w_072_9584, w_072_9586, w_072_9604, w_072_9607, w_072_9611, w_072_9615, w_072_9616, w_072_9617, w_072_9621, w_072_9622, w_072_9634, w_072_9641, w_072_9642, w_072_9643, w_072_9646, w_072_9647, w_072_9648, w_072_9651, w_072_9653, w_072_9654, w_072_9655, w_072_9658, w_072_9663, w_072_9664, w_072_9666, w_072_9671, w_072_9675, w_072_9677, w_072_9680, w_072_9684, w_072_9688, w_072_9691, w_072_9693, w_072_9697, w_072_9699, w_072_9700, w_072_9701, w_072_9702, w_072_9710, w_072_9712, w_072_9716, w_072_9719, w_072_9726, w_072_9735, w_072_9740, w_072_9743, w_072_9744, w_072_9745, w_072_9750, w_072_9752, w_072_9757, w_072_9759, w_072_9769, w_072_9772, w_072_9779, w_072_9780, w_072_9789, w_072_9794, w_072_9802, w_072_9803, w_072_9810, w_072_9811, w_072_9814, w_072_9815, w_072_9816, w_072_9819, w_072_9823;
  wire w_073_002, w_073_005, w_073_006, w_073_007, w_073_008, w_073_009, w_073_010, w_073_011, w_073_014, w_073_018, w_073_019, w_073_020, w_073_025, w_073_027, w_073_028, w_073_029, w_073_030, w_073_031, w_073_032, w_073_035, w_073_039, w_073_041, w_073_043, w_073_047, w_073_049, w_073_055, w_073_057, w_073_060, w_073_061, w_073_062, w_073_064, w_073_066, w_073_078, w_073_079, w_073_081, w_073_083, w_073_084, w_073_085, w_073_086, w_073_088, w_073_090, w_073_091, w_073_093, w_073_094, w_073_095, w_073_096, w_073_099, w_073_100, w_073_102, w_073_103, w_073_104, w_073_108, w_073_110, w_073_111, w_073_112, w_073_116, w_073_117, w_073_118, w_073_120, w_073_121, w_073_123, w_073_125, w_073_126, w_073_127, w_073_128, w_073_131, w_073_132, w_073_133, w_073_134, w_073_135, w_073_136, w_073_137, w_073_139, w_073_140, w_073_141, w_073_142, w_073_145, w_073_146, w_073_147, w_073_149, w_073_152, w_073_153, w_073_154, w_073_156, w_073_158, w_073_160, w_073_161, w_073_166, w_073_169, w_073_173, w_073_174, w_073_178, w_073_179, w_073_180, w_073_181, w_073_183, w_073_184, w_073_186, w_073_187, w_073_188, w_073_190, w_073_195, w_073_198, w_073_202, w_073_204, w_073_208, w_073_215, w_073_216, w_073_217, w_073_222, w_073_223, w_073_224, w_073_225, w_073_231, w_073_232, w_073_235, w_073_237, w_073_238, w_073_241, w_073_243, w_073_244, w_073_245, w_073_246, w_073_247, w_073_248, w_073_249, w_073_251, w_073_253, w_073_254, w_073_258, w_073_259, w_073_261, w_073_262, w_073_263, w_073_268, w_073_270, w_073_271, w_073_272, w_073_275, w_073_278, w_073_281, w_073_282, w_073_283, w_073_284, w_073_287, w_073_288, w_073_289, w_073_290, w_073_293, w_073_296, w_073_297, w_073_299, w_073_300, w_073_301, w_073_302, w_073_303, w_073_304, w_073_307, w_073_308, w_073_311, w_073_312, w_073_316, w_073_318, w_073_321, w_073_323, w_073_324, w_073_325, w_073_327, w_073_331, w_073_332, w_073_333, w_073_334, w_073_335, w_073_336, w_073_337, w_073_338, w_073_341, w_073_343, w_073_344, w_073_345, w_073_346, w_073_347, w_073_349, w_073_351, w_073_352, w_073_355, w_073_358, w_073_361, w_073_362, w_073_365, w_073_368, w_073_369, w_073_371, w_073_372, w_073_374, w_073_379, w_073_381, w_073_382, w_073_384, w_073_385, w_073_386, w_073_387, w_073_388, w_073_389, w_073_396, w_073_397, w_073_399, w_073_401, w_073_402, w_073_405, w_073_411, w_073_414, w_073_417, w_073_418, w_073_419, w_073_421, w_073_422, w_073_423, w_073_425, w_073_426, w_073_434, w_073_435, w_073_436, w_073_437, w_073_438, w_073_439, w_073_440, w_073_441, w_073_442, w_073_443, w_073_444, w_073_448, w_073_451, w_073_452, w_073_453, w_073_455, w_073_456, w_073_457, w_073_459, w_073_460, w_073_464, w_073_467, w_073_468, w_073_470, w_073_472, w_073_475, w_073_480, w_073_481, w_073_483, w_073_485, w_073_486, w_073_488, w_073_489, w_073_491, w_073_492, w_073_493, w_073_495, w_073_496, w_073_497, w_073_502, w_073_505, w_073_506, w_073_507, w_073_508, w_073_510, w_073_512, w_073_513, w_073_514, w_073_517, w_073_520, w_073_522, w_073_524, w_073_526, w_073_529, w_073_531, w_073_533, w_073_534, w_073_535, w_073_537, w_073_540, w_073_541, w_073_543, w_073_544, w_073_549, w_073_550, w_073_553, w_073_555, w_073_556, w_073_557, w_073_559, w_073_560, w_073_561, w_073_564, w_073_565, w_073_569, w_073_571, w_073_574, w_073_575, w_073_577, w_073_579, w_073_583, w_073_584, w_073_585, w_073_589, w_073_592, w_073_593, w_073_594, w_073_596, w_073_597, w_073_599, w_073_600, w_073_602, w_073_603, w_073_605, w_073_606, w_073_608, w_073_610, w_073_611, w_073_613, w_073_618, w_073_619, w_073_620, w_073_622, w_073_623, w_073_626, w_073_631, w_073_632, w_073_633, w_073_635, w_073_636, w_073_638, w_073_643, w_073_646, w_073_648, w_073_650, w_073_651, w_073_652, w_073_653, w_073_654, w_073_655, w_073_657, w_073_658, w_073_659, w_073_664, w_073_665, w_073_667, w_073_673, w_073_674, w_073_675, w_073_676, w_073_678, w_073_679, w_073_681, w_073_684, w_073_688, w_073_690, w_073_691, w_073_698, w_073_702, w_073_703, w_073_704, w_073_707, w_073_708, w_073_709, w_073_711, w_073_715, w_073_716, w_073_717, w_073_718, w_073_720, w_073_722, w_073_725, w_073_727, w_073_731, w_073_732, w_073_735, w_073_737, w_073_739, w_073_745, w_073_746, w_073_751, w_073_753, w_073_754, w_073_756, w_073_757, w_073_758, w_073_762, w_073_763, w_073_764, w_073_765, w_073_768, w_073_770, w_073_772, w_073_773, w_073_774, w_073_775, w_073_776, w_073_778, w_073_779, w_073_780, w_073_782, w_073_783, w_073_784, w_073_786, w_073_788, w_073_790, w_073_792, w_073_793, w_073_795, w_073_797, w_073_799, w_073_801, w_073_804, w_073_806, w_073_807, w_073_808, w_073_810, w_073_811, w_073_812, w_073_814, w_073_815, w_073_816, w_073_817, w_073_818, w_073_821, w_073_822, w_073_823, w_073_824, w_073_826, w_073_828, w_073_829, w_073_830, w_073_835, w_073_836, w_073_837, w_073_839, w_073_840, w_073_844, w_073_845, w_073_846, w_073_847, w_073_849, w_073_850, w_073_852, w_073_857, w_073_859, w_073_860, w_073_861, w_073_862, w_073_869, w_073_870, w_073_872, w_073_873, w_073_874, w_073_875, w_073_876, w_073_877, w_073_878, w_073_879, w_073_880, w_073_885, w_073_894, w_073_895, w_073_898, w_073_900, w_073_901, w_073_903, w_073_904, w_073_905, w_073_908, w_073_912, w_073_913, w_073_914, w_073_917, w_073_919, w_073_920, w_073_921, w_073_922, w_073_923, w_073_924, w_073_927, w_073_928, w_073_930, w_073_933, w_073_937, w_073_938, w_073_940, w_073_941, w_073_942, w_073_946, w_073_947, w_073_948, w_073_949, w_073_951, w_073_952, w_073_953, w_073_954, w_073_955, w_073_957, w_073_958, w_073_959, w_073_965, w_073_966, w_073_969, w_073_972, w_073_973, w_073_975, w_073_976, w_073_978, w_073_979, w_073_980, w_073_981, w_073_983, w_073_986, w_073_987, w_073_988, w_073_990, w_073_991, w_073_993, w_073_995, w_073_996, w_073_997, w_073_998, w_073_999, w_073_1001, w_073_1003, w_073_1004, w_073_1005, w_073_1006, w_073_1007, w_073_1009, w_073_1010, w_073_1015, w_073_1016, w_073_1018, w_073_1019, w_073_1020, w_073_1021, w_073_1022, w_073_1024, w_073_1025, w_073_1027, w_073_1028, w_073_1029, w_073_1031, w_073_1033, w_073_1037, w_073_1040, w_073_1042, w_073_1045, w_073_1048, w_073_1050, w_073_1051, w_073_1052, w_073_1053, w_073_1054, w_073_1055, w_073_1057, w_073_1058, w_073_1060, w_073_1062, w_073_1064, w_073_1068, w_073_1070, w_073_1071, w_073_1077, w_073_1079, w_073_1080, w_073_1081, w_073_1085, w_073_1086, w_073_1087, w_073_1090, w_073_1091, w_073_1093, w_073_1097, w_073_1098, w_073_1099, w_073_1100, w_073_1104, w_073_1105, w_073_1106, w_073_1107, w_073_1109, w_073_1112, w_073_1113, w_073_1114, w_073_1115, w_073_1116, w_073_1117, w_073_1118, w_073_1121, w_073_1123, w_073_1125, w_073_1128, w_073_1130, w_073_1131, w_073_1132, w_073_1145, w_073_1147, w_073_1148, w_073_1151, w_073_1152, w_073_1153, w_073_1154, w_073_1155, w_073_1156, w_073_1158, w_073_1160, w_073_1161, w_073_1163, w_073_1166, w_073_1170, w_073_1171, w_073_1172, w_073_1174, w_073_1176, w_073_1178, w_073_1179, w_073_1180, w_073_1181, w_073_1185, w_073_1188, w_073_1189, w_073_1190, w_073_1191, w_073_1193, w_073_1196, w_073_1198, w_073_1199, w_073_1200, w_073_1208, w_073_1210, w_073_1212, w_073_1213, w_073_1214, w_073_1217, w_073_1219, w_073_1222, w_073_1223, w_073_1233, w_073_1234, w_073_1236, w_073_1237, w_073_1238, w_073_1239, w_073_1241, w_073_1242, w_073_1244, w_073_1245, w_073_1247, w_073_1249, w_073_1251, w_073_1254, w_073_1255, w_073_1256, w_073_1257, w_073_1259, w_073_1260, w_073_1262, w_073_1263, w_073_1266, w_073_1268, w_073_1270, w_073_1273, w_073_1274, w_073_1275, w_073_1276, w_073_1277, w_073_1278, w_073_1279, w_073_1282, w_073_1287, w_073_1288, w_073_1290, w_073_1291, w_073_1292, w_073_1293, w_073_1294, w_073_1295, w_073_1296, w_073_1297, w_073_1298, w_073_1299, w_073_1306, w_073_1307, w_073_1309, w_073_1311, w_073_1312, w_073_1313, w_073_1315, w_073_1316, w_073_1321, w_073_1322, w_073_1323, w_073_1325, w_073_1327, w_073_1328, w_073_1330, w_073_1332, w_073_1334, w_073_1338, w_073_1339, w_073_1340, w_073_1341, w_073_1342, w_073_1343, w_073_1344, w_073_1345, w_073_1348, w_073_1350, w_073_1351, w_073_1353, w_073_1354, w_073_1355, w_073_1358, w_073_1359, w_073_1361, w_073_1362, w_073_1363, w_073_1366, w_073_1368, w_073_1371, w_073_1374, w_073_1376, w_073_1378, w_073_1379, w_073_1381, w_073_1382, w_073_1387, w_073_1388, w_073_1389, w_073_1390, w_073_1393, w_073_1394, w_073_1395, w_073_1396, w_073_1399, w_073_1400, w_073_1403, w_073_1404, w_073_1405, w_073_1406, w_073_1408, w_073_1411, w_073_1412, w_073_1414, w_073_1415, w_073_1416, w_073_1420, w_073_1422, w_073_1426, w_073_1428, w_073_1429, w_073_1430, w_073_1432, w_073_1439, w_073_1440, w_073_1441, w_073_1443, w_073_1444, w_073_1447, w_073_1448, w_073_1450, w_073_1453, w_073_1455, w_073_1458, w_073_1460, w_073_1461, w_073_1462, w_073_1466, w_073_1468, w_073_1478, w_073_1481, w_073_1484, w_073_1486, w_073_1488, w_073_1491, w_073_1492, w_073_1494, w_073_1497, w_073_1498, w_073_1499, w_073_1500, w_073_1503, w_073_1504, w_073_1505, w_073_1506, w_073_1511, w_073_1514, w_073_1515, w_073_1516, w_073_1517, w_073_1518, w_073_1523, w_073_1524, w_073_1525, w_073_1526, w_073_1528, w_073_1531, w_073_1533, w_073_1535, w_073_1537, w_073_1539, w_073_1540, w_073_1541, w_073_1554, w_073_1559, w_073_1561, w_073_1567, w_073_1568, w_073_1569, w_073_1572, w_073_1578, w_073_1579, w_073_1581, w_073_1583, w_073_1584, w_073_1586, w_073_1590, w_073_1591, w_073_1592, w_073_1594, w_073_1595, w_073_1596, w_073_1599, w_073_1600, w_073_1603, w_073_1607, w_073_1608, w_073_1610, w_073_1613, w_073_1615, w_073_1617, w_073_1619, w_073_1621, w_073_1623, w_073_1626, w_073_1628, w_073_1630, w_073_1634, w_073_1635, w_073_1636, w_073_1638, w_073_1640, w_073_1643, w_073_1645, w_073_1648, w_073_1650, w_073_1651, w_073_1652, w_073_1653, w_073_1654, w_073_1655, w_073_1656, w_073_1657, w_073_1659, w_073_1660, w_073_1664, w_073_1666, w_073_1667, w_073_1669, w_073_1670, w_073_1671, w_073_1672, w_073_1673, w_073_1674, w_073_1677, w_073_1680, w_073_1681, w_073_1682, w_073_1683, w_073_1684, w_073_1686, w_073_1687, w_073_1688, w_073_1691, w_073_1692, w_073_1693, w_073_1694, w_073_1695, w_073_1696, w_073_1698, w_073_1701, w_073_1702, w_073_1704, w_073_1706, w_073_1707, w_073_1710, w_073_1711, w_073_1712, w_073_1715, w_073_1716, w_073_1718, w_073_1720, w_073_1722, w_073_1723, w_073_1725, w_073_1726, w_073_1727, w_073_1729, w_073_1731, w_073_1734, w_073_1735, w_073_1736, w_073_1737, w_073_1738, w_073_1740, w_073_1741, w_073_1742, w_073_1743, w_073_1744, w_073_1746, w_073_1747, w_073_1749, w_073_1751, w_073_1752, w_073_1754, w_073_1755, w_073_1758, w_073_1760, w_073_1761, w_073_1765, w_073_1766, w_073_1768, w_073_1769, w_073_1770, w_073_1771, w_073_1776, w_073_1777, w_073_1780, w_073_1782, w_073_1786, w_073_1787, w_073_1788, w_073_1791, w_073_1795, w_073_1797, w_073_1799, w_073_1805, w_073_1806, w_073_1807, w_073_1809, w_073_1810, w_073_1815, w_073_1817, w_073_1819, w_073_1820, w_073_1821, w_073_1822, w_073_1823, w_073_1824, w_073_1825, w_073_1827, w_073_1829, w_073_1830, w_073_1831, w_073_1832, w_073_1833, w_073_1835, w_073_1839, w_073_1842, w_073_1846, w_073_1847, w_073_1848, w_073_1850, w_073_1851, w_073_1852, w_073_1854, w_073_1855, w_073_1858, w_073_1862, w_073_1866, w_073_1869, w_073_1870, w_073_1871, w_073_1874, w_073_1876, w_073_1877, w_073_1879, w_073_1881, w_073_1884, w_073_1885, w_073_1886, w_073_1887, w_073_1888, w_073_1889, w_073_1891, w_073_1893, w_073_1897, w_073_1899, w_073_1900, w_073_1901, w_073_1902, w_073_1903, w_073_1904, w_073_1905, w_073_1906, w_073_1907, w_073_1909, w_073_1910, w_073_1911, w_073_1912, w_073_1914, w_073_1915, w_073_1916, w_073_1917, w_073_1918, w_073_1920, w_073_1921, w_073_1922, w_073_1923, w_073_1924, w_073_1926, w_073_1927, w_073_1929, w_073_1931, w_073_1940, w_073_1944, w_073_1945, w_073_1946, w_073_1955, w_073_1956, w_073_1958, w_073_1960, w_073_1961, w_073_1963, w_073_1965, w_073_1966, w_073_1968, w_073_1971, w_073_1972, w_073_1974, w_073_1977, w_073_1978, w_073_1981, w_073_1983, w_073_1985, w_073_1986, w_073_1987, w_073_1989, w_073_1990, w_073_1991, w_073_1993, w_073_1995, w_073_1996, w_073_1997, w_073_1999, w_073_2000, w_073_2004, w_073_2005, w_073_2007, w_073_2008, w_073_2010, w_073_2011, w_073_2012, w_073_2016, w_073_2017, w_073_2018, w_073_2019, w_073_2022, w_073_2023, w_073_2026, w_073_2027, w_073_2029, w_073_2031, w_073_2032, w_073_2033, w_073_2035, w_073_2037, w_073_2038, w_073_2039, w_073_2043, w_073_2044, w_073_2045, w_073_2046, w_073_2047, w_073_2048, w_073_2050, w_073_2051, w_073_2052, w_073_2053, w_073_2055, w_073_2057, w_073_2058, w_073_2059, w_073_2061, w_073_2064, w_073_2065, w_073_2066, w_073_2067, w_073_2068, w_073_2072, w_073_2074, w_073_2075, w_073_2076, w_073_2078, w_073_2080, w_073_2081, w_073_2083, w_073_2084, w_073_2085, w_073_2087, w_073_2088, w_073_2091, w_073_2094, w_073_2100, w_073_2101, w_073_2102, w_073_2103, w_073_2104, w_073_2105, w_073_2111, w_073_2115, w_073_2117, w_073_2118, w_073_2119, w_073_2120, w_073_2121, w_073_2122, w_073_2123, w_073_2125, w_073_2126, w_073_2131, w_073_2132, w_073_2135, w_073_2137, w_073_2144, w_073_2148, w_073_2150, w_073_2151, w_073_2155, w_073_2156, w_073_2159, w_073_2160, w_073_2163, w_073_2165, w_073_2167, w_073_2168, w_073_2169, w_073_2172, w_073_2173, w_073_2175, w_073_2178, w_073_2179, w_073_2180, w_073_2184, w_073_2185, w_073_2186, w_073_2187, w_073_2188, w_073_2190, w_073_2192, w_073_2193, w_073_2194, w_073_2195, w_073_2198, w_073_2199, w_073_2201, w_073_2202, w_073_2203, w_073_2204, w_073_2205, w_073_2206, w_073_2208, w_073_2211, w_073_2212, w_073_2214, w_073_2215, w_073_2218, w_073_2219, w_073_2223, w_073_2225, w_073_2226, w_073_2230, w_073_2233, w_073_2234, w_073_2236, w_073_2237, w_073_2238, w_073_2239, w_073_2240, w_073_2241, w_073_2242, w_073_2244, w_073_2246, w_073_2249, w_073_2250, w_073_2255, w_073_2263, w_073_2266, w_073_2267, w_073_2269, w_073_2270, w_073_2273, w_073_2275, w_073_2276, w_073_2277, w_073_2278, w_073_2279, w_073_2280, w_073_2282, w_073_2283, w_073_2284, w_073_2286, w_073_2287, w_073_2290, w_073_2291, w_073_2296, w_073_2299, w_073_2300, w_073_2301, w_073_2304, w_073_2305, w_073_2309, w_073_2310, w_073_2312, w_073_2315, w_073_2316, w_073_2317, w_073_2321, w_073_2326, w_073_2327, w_073_2328, w_073_2329, w_073_2331, w_073_2332, w_073_2335, w_073_2338, w_073_2339, w_073_2340, w_073_2341, w_073_2345, w_073_2346, w_073_2348, w_073_2350, w_073_2352, w_073_2355, w_073_2356, w_073_2357, w_073_2358, w_073_2359, w_073_2361, w_073_2362, w_073_2364, w_073_2367, w_073_2369, w_073_2370, w_073_2371, w_073_2373, w_073_2374, w_073_2376, w_073_2378, w_073_2381, w_073_2385, w_073_2386, w_073_2387, w_073_2388, w_073_2389, w_073_2390, w_073_2391, w_073_2393, w_073_2395, w_073_2397, w_073_2398, w_073_2399, w_073_2403, w_073_2404, w_073_2405, w_073_2406, w_073_2410, w_073_2414, w_073_2415, w_073_2420, w_073_2421, w_073_2422, w_073_2424, w_073_2427, w_073_2428, w_073_2430, w_073_2431, w_073_2433, w_073_2435, w_073_2436, w_073_2438, w_073_2440, w_073_2448, w_073_2451, w_073_2456, w_073_2459, w_073_2462, w_073_2464, w_073_2465, w_073_2469, w_073_2470, w_073_2471, w_073_2473, w_073_2474, w_073_2477, w_073_2480, w_073_2481, w_073_2486, w_073_2490, w_073_2491, w_073_2492, w_073_2493, w_073_2494, w_073_2495, w_073_2497, w_073_2498, w_073_2499, w_073_2500, w_073_2502, w_073_2503, w_073_2505, w_073_2506, w_073_2508, w_073_2509, w_073_2510, w_073_2511, w_073_2515, w_073_2517, w_073_2518, w_073_2522, w_073_2524, w_073_2526, w_073_2527, w_073_2529, w_073_2535, w_073_2539, w_073_2540, w_073_2542, w_073_2544, w_073_2545, w_073_2546, w_073_2547, w_073_2549, w_073_2550, w_073_2553, w_073_2556, w_073_2557, w_073_2559, w_073_2560, w_073_2563, w_073_2567, w_073_2568, w_073_2569, w_073_2572, w_073_2575, w_073_2576, w_073_2583, w_073_2584, w_073_2585, w_073_2586, w_073_2587, w_073_2589, w_073_2591, w_073_2593, w_073_2594, w_073_2596, w_073_2598, w_073_2599, w_073_2600, w_073_2602, w_073_2604, w_073_2608, w_073_2609, w_073_2610, w_073_2611, w_073_2612, w_073_2613, w_073_2614, w_073_2615, w_073_2617, w_073_2618, w_073_2621, w_073_2622, w_073_2627, w_073_2630, w_073_2632, w_073_2634, w_073_2637, w_073_2638, w_073_2640, w_073_2642, w_073_2643, w_073_2644, w_073_2645, w_073_2646, w_073_2651, w_073_2656, w_073_2658, w_073_2659, w_073_2664, w_073_2670, w_073_2671, w_073_2672, w_073_2674, w_073_2677, w_073_2679, w_073_2682, w_073_2684, w_073_2685, w_073_2686, w_073_2687, w_073_2690, w_073_2691, w_073_2695, w_073_2696, w_073_2697, w_073_2702, w_073_2703, w_073_2704, w_073_2709, w_073_2710, w_073_2712, w_073_2714, w_073_2715, w_073_2716, w_073_2717, w_073_2719, w_073_2720, w_073_2721, w_073_2725, w_073_2726, w_073_2727, w_073_2728, w_073_2731, w_073_2733, w_073_2734, w_073_2735, w_073_2736, w_073_2737, w_073_2739, w_073_2740, w_073_2743, w_073_2744, w_073_2745, w_073_2746, w_073_2747, w_073_2748, w_073_2749, w_073_2750, w_073_2751, w_073_2752, w_073_2753, w_073_2755, w_073_2756, w_073_2758, w_073_2759, w_073_2760, w_073_2763, w_073_2764, w_073_2766, w_073_2768, w_073_2770, w_073_2771, w_073_2772, w_073_2773, w_073_2774, w_073_2775, w_073_2776, w_073_2777, w_073_2779, w_073_2785, w_073_2786, w_073_2788, w_073_2793, w_073_2794, w_073_2795, w_073_2797, w_073_2798, w_073_2800, w_073_2801, w_073_2805, w_073_2807, w_073_2809, w_073_2812, w_073_2815, w_073_2816, w_073_2820, w_073_2821, w_073_2822, w_073_2824, w_073_2827, w_073_2829, w_073_2830, w_073_2831, w_073_2832, w_073_2835, w_073_2837, w_073_2838, w_073_2839, w_073_2842, w_073_2843, w_073_2844, w_073_2846, w_073_2852, w_073_2857, w_073_2861, w_073_2863, w_073_2869, w_073_2870, w_073_2871, w_073_2874, w_073_2876, w_073_2878, w_073_2879, w_073_2880, w_073_2881, w_073_2884, w_073_2885, w_073_2886, w_073_2887, w_073_2888, w_073_2889, w_073_2890, w_073_2891, w_073_2893, w_073_2897, w_073_2899, w_073_2900, w_073_2901, w_073_2902, w_073_2903, w_073_2904, w_073_2905, w_073_2906, w_073_2907, w_073_2912, w_073_2913, w_073_2914, w_073_2915, w_073_2917, w_073_2919, w_073_2920, w_073_2922, w_073_2923, w_073_2925, w_073_2929, w_073_2930, w_073_2934, w_073_2935, w_073_2936, w_073_2938, w_073_2939, w_073_2940, w_073_2941, w_073_2943, w_073_2945, w_073_2946, w_073_2947, w_073_2948, w_073_2949, w_073_2950, w_073_2951, w_073_2952, w_073_2953, w_073_2954, w_073_2955, w_073_2957, w_073_2958, w_073_2959, w_073_2963, w_073_2964, w_073_2965, w_073_2967, w_073_2969, w_073_2970, w_073_2972, w_073_2975, w_073_2976, w_073_2978, w_073_2981, w_073_2982, w_073_2983, w_073_2984, w_073_2985, w_073_2990, w_073_2991, w_073_2993, w_073_2995, w_073_2996, w_073_2998, w_073_3000, w_073_3001, w_073_3002, w_073_3003, w_073_3004, w_073_3006, w_073_3008, w_073_3009, w_073_3011, w_073_3013, w_073_3015, w_073_3017, w_073_3019, w_073_3021, w_073_3022, w_073_3024, w_073_3025, w_073_3026, w_073_3027, w_073_3033, w_073_3035, w_073_3036, w_073_3042, w_073_3043, w_073_3044, w_073_3050, w_073_3053, w_073_3054, w_073_3055, w_073_3058, w_073_3059, w_073_3061, w_073_3062, w_073_3067, w_073_3070, w_073_3071, w_073_3076, w_073_3077, w_073_3082, w_073_3083, w_073_3084, w_073_3086, w_073_3090, w_073_3091, w_073_3093, w_073_3094, w_073_3100, w_073_3102, w_073_3105, w_073_3106, w_073_3107, w_073_3108, w_073_3112, w_073_3113, w_073_3118, w_073_3122, w_073_3123, w_073_3124, w_073_3125, w_073_3126, w_073_3128, w_073_3131, w_073_3132, w_073_3134, w_073_3138, w_073_3141, w_073_3142, w_073_3144, w_073_3148, w_073_3149, w_073_3150, w_073_3151, w_073_3152, w_073_3153, w_073_3155, w_073_3156, w_073_3158, w_073_3161, w_073_3164, w_073_3165, w_073_3168, w_073_3169, w_073_3171, w_073_3174, w_073_3175, w_073_3181, w_073_3182, w_073_3184, w_073_3186, w_073_3189, w_073_3191, w_073_3193, w_073_3194, w_073_3195, w_073_3201, w_073_3204, w_073_3206, w_073_3207, w_073_3209, w_073_3212, w_073_3217, w_073_3218, w_073_3219, w_073_3221, w_073_3222, w_073_3227, w_073_3229, w_073_3230, w_073_3231, w_073_3234, w_073_3236, w_073_3238, w_073_3239, w_073_3240, w_073_3241, w_073_3242, w_073_3243, w_073_3244, w_073_3245, w_073_3248, w_073_3250, w_073_3251, w_073_3254, w_073_3255, w_073_3256, w_073_3258, w_073_3259, w_073_3260, w_073_3264, w_073_3265, w_073_3267, w_073_3268, w_073_3269, w_073_3274, w_073_3275, w_073_3276, w_073_3278, w_073_3279, w_073_3281, w_073_3282, w_073_3283, w_073_3284, w_073_3286, w_073_3288, w_073_3290, w_073_3291, w_073_3292, w_073_3293, w_073_3295, w_073_3297, w_073_3299, w_073_3300, w_073_3304, w_073_3306, w_073_3310, w_073_3311, w_073_3312, w_073_3313, w_073_3314, w_073_3316, w_073_3317, w_073_3320, w_073_3321, w_073_3326, w_073_3327, w_073_3328, w_073_3329, w_073_3330, w_073_3331, w_073_3333, w_073_3337, w_073_3338, w_073_3339, w_073_3340, w_073_3341, w_073_3342, w_073_3343, w_073_3348, w_073_3349, w_073_3351, w_073_3353, w_073_3354, w_073_3358, w_073_3360, w_073_3361, w_073_3362, w_073_3363, w_073_3364, w_073_3365, w_073_3367, w_073_3372, w_073_3377, w_073_3380, w_073_3383, w_073_3386, w_073_3387, w_073_3388, w_073_3389, w_073_3390, w_073_3391, w_073_3392, w_073_3393, w_073_3395, w_073_3397, w_073_3398, w_073_3399, w_073_3400, w_073_3401, w_073_3402, w_073_3403, w_073_3404, w_073_3406, w_073_3407, w_073_3408, w_073_3411, w_073_3413, w_073_3414, w_073_3415, w_073_3416, w_073_3419, w_073_3422, w_073_3423, w_073_3424, w_073_3425, w_073_3426, w_073_3427, w_073_3428, w_073_3430, w_073_3432, w_073_3434, w_073_3438, w_073_3439, w_073_3443, w_073_3445, w_073_3447, w_073_3448, w_073_3451, w_073_3456, w_073_3457, w_073_3458, w_073_3460, w_073_3461, w_073_3462, w_073_3466, w_073_3469, w_073_3470, w_073_3471, w_073_3474, w_073_3476, w_073_3477, w_073_3478, w_073_3481, w_073_3484, w_073_3486, w_073_3488, w_073_3489, w_073_3491, w_073_3492, w_073_3495, w_073_3496, w_073_3498, w_073_3502, w_073_3507, w_073_3508, w_073_3509, w_073_3510, w_073_3512, w_073_3513, w_073_3516, w_073_3517, w_073_3519, w_073_3525, w_073_3527, w_073_3528, w_073_3529, w_073_3530, w_073_3535, w_073_3537, w_073_3538, w_073_3539, w_073_3543, w_073_3544, w_073_3545, w_073_3546, w_073_3547, w_073_3548, w_073_3549, w_073_3552, w_073_3555, w_073_3558, w_073_3559, w_073_3562, w_073_3563, w_073_3564, w_073_3566, w_073_3567, w_073_3569, w_073_3570, w_073_3571, w_073_3575, w_073_3581, w_073_3584, w_073_3587, w_073_3592, w_073_3593, w_073_3594, w_073_3596, w_073_3597, w_073_3598, w_073_3600, w_073_3601, w_073_3602, w_073_3603, w_073_3606, w_073_3607, w_073_3609, w_073_3610, w_073_3611, w_073_3612, w_073_3615, w_073_3617, w_073_3621, w_073_3622, w_073_3627, w_073_3628, w_073_3629, w_073_3630, w_073_3631, w_073_3632, w_073_3634, w_073_3637, w_073_3638, w_073_3640, w_073_3642, w_073_3645, w_073_3646, w_073_3647, w_073_3648, w_073_3651, w_073_3652, w_073_3653, w_073_3654, w_073_3656, w_073_3657, w_073_3658, w_073_3661, w_073_3662, w_073_3664, w_073_3666, w_073_3667, w_073_3668, w_073_3669, w_073_3670, w_073_3672, w_073_3674, w_073_3675, w_073_3677, w_073_3679, w_073_3681, w_073_3682, w_073_3684, w_073_3686, w_073_3687, w_073_3688, w_073_3689, w_073_3691, w_073_3694, w_073_3695, w_073_3697, w_073_3700, w_073_3702, w_073_3703, w_073_3707, w_073_3708, w_073_3711, w_073_3716, w_073_3719, w_073_3721, w_073_3722, w_073_3723, w_073_3728, w_073_3730, w_073_3733, w_073_3736, w_073_3737, w_073_3738, w_073_3739, w_073_3740, w_073_3741, w_073_3743, w_073_3745, w_073_3746, w_073_3750, w_073_3754, w_073_3755, w_073_3756, w_073_3759, w_073_3760, w_073_3761, w_073_3762, w_073_3763, w_073_3765, w_073_3766, w_073_3767, w_073_3771, w_073_3772, w_073_3780, w_073_3782, w_073_3784, w_073_3788, w_073_3795, w_073_3796, w_073_3798, w_073_3799, w_073_3801, w_073_3802, w_073_3803, w_073_3804, w_073_3805, w_073_3806, w_073_3807, w_073_3808, w_073_3811, w_073_3813, w_073_3815, w_073_3816, w_073_3819, w_073_3820, w_073_3821, w_073_3822, w_073_3823, w_073_3825, w_073_3826, w_073_3827, w_073_3829, w_073_3832, w_073_3836, w_073_3838, w_073_3841, w_073_3843, w_073_3846, w_073_3848, w_073_3850, w_073_3851, w_073_3852, w_073_3855, w_073_3856, w_073_3857, w_073_3859, w_073_3860, w_073_3861, w_073_3862, w_073_3863, w_073_3865, w_073_3867, w_073_3871, w_073_3872, w_073_3874, w_073_3875, w_073_3876, w_073_3879, w_073_3880, w_073_3884, w_073_3885, w_073_3892, w_073_3893, w_073_3896, w_073_3898, w_073_3899, w_073_3900, w_073_3901, w_073_3903, w_073_3909, w_073_3911, w_073_3912, w_073_3914, w_073_3915, w_073_3920, w_073_3922, w_073_3927, w_073_3929, w_073_3933, w_073_3935, w_073_3936, w_073_3937, w_073_3938, w_073_3939, w_073_3941, w_073_3944, w_073_3946, w_073_3947, w_073_3950, w_073_3951, w_073_3952, w_073_3954, w_073_3956, w_073_3957, w_073_3959, w_073_3960, w_073_3962, w_073_3963, w_073_3964, w_073_3967, w_073_3969, w_073_3972, w_073_3974, w_073_3975, w_073_3976, w_073_3977, w_073_3981, w_073_3982, w_073_3983, w_073_3984, w_073_3986, w_073_3987, w_073_3988, w_073_3989, w_073_3990, w_073_3992, w_073_3993, w_073_3995, w_073_3996, w_073_3997, w_073_3998, w_073_3999, w_073_4008, w_073_4009, w_073_4013, w_073_4014, w_073_4024, w_073_4025, w_073_4029, w_073_4031, w_073_4032, w_073_4034, w_073_4037, w_073_4041, w_073_4050, w_073_4059, w_073_4077, w_073_4081, w_073_4087, w_073_4095, w_073_4099, w_073_4101, w_073_4104, w_073_4107, w_073_4108, w_073_4110, w_073_4113, w_073_4116, w_073_4117, w_073_4118, w_073_4119, w_073_4121, w_073_4125, w_073_4126, w_073_4135, w_073_4136, w_073_4144, w_073_4145, w_073_4148, w_073_4152, w_073_4154, w_073_4157, w_073_4159, w_073_4160, w_073_4162, w_073_4165, w_073_4170, w_073_4177, w_073_4180, w_073_4183, w_073_4184, w_073_4193, w_073_4200, w_073_4202, w_073_4204, w_073_4205, w_073_4210, w_073_4211, w_073_4213, w_073_4214, w_073_4219, w_073_4220, w_073_4221, w_073_4222, w_073_4223, w_073_4225, w_073_4231, w_073_4238, w_073_4242, w_073_4243, w_073_4244, w_073_4246, w_073_4247, w_073_4248, w_073_4255, w_073_4257, w_073_4259, w_073_4267, w_073_4273, w_073_4275, w_073_4280, w_073_4281, w_073_4286, w_073_4287, w_073_4289, w_073_4290, w_073_4292, w_073_4294, w_073_4296, w_073_4297, w_073_4300, w_073_4302, w_073_4305, w_073_4306, w_073_4308, w_073_4320, w_073_4323, w_073_4326, w_073_4327, w_073_4336, w_073_4340, w_073_4344, w_073_4348, w_073_4350, w_073_4351, w_073_4352, w_073_4365, w_073_4366, w_073_4368, w_073_4369, w_073_4370, w_073_4371, w_073_4373, w_073_4377, w_073_4381, w_073_4382, w_073_4388, w_073_4390, w_073_4392, w_073_4393, w_073_4399, w_073_4400, w_073_4402, w_073_4403, w_073_4405, w_073_4406, w_073_4407, w_073_4408, w_073_4409, w_073_4411, w_073_4412, w_073_4424, w_073_4425, w_073_4427, w_073_4430, w_073_4435, w_073_4439, w_073_4440, w_073_4441, w_073_4446, w_073_4448, w_073_4449, w_073_4457, w_073_4470, w_073_4471, w_073_4474, w_073_4479, w_073_4489, w_073_4491, w_073_4493, w_073_4496, w_073_4500, w_073_4501, w_073_4503, w_073_4508, w_073_4510, w_073_4517, w_073_4518, w_073_4519, w_073_4520, w_073_4521, w_073_4524, w_073_4525, w_073_4526, w_073_4529, w_073_4530, w_073_4531, w_073_4532, w_073_4536, w_073_4539, w_073_4543, w_073_4552, w_073_4553, w_073_4555, w_073_4559, w_073_4560, w_073_4561, w_073_4565, w_073_4578, w_073_4579, w_073_4583, w_073_4584, w_073_4590, w_073_4593, w_073_4596, w_073_4598, w_073_4599, w_073_4600, w_073_4603, w_073_4609, w_073_4613, w_073_4614, w_073_4620, w_073_4621, w_073_4622, w_073_4635, w_073_4636, w_073_4638, w_073_4646, w_073_4651, w_073_4653, w_073_4657, w_073_4662, w_073_4664, w_073_4665, w_073_4667, w_073_4668, w_073_4680, w_073_4682, w_073_4683, w_073_4685, w_073_4688, w_073_4690, w_073_4694, w_073_4701, w_073_4702, w_073_4710, w_073_4714, w_073_4715, w_073_4718, w_073_4720, w_073_4722, w_073_4727, w_073_4732, w_073_4733, w_073_4734, w_073_4738, w_073_4741, w_073_4742, w_073_4743, w_073_4744, w_073_4748, w_073_4749, w_073_4750, w_073_4752, w_073_4754, w_073_4758, w_073_4761, w_073_4765, w_073_4769, w_073_4770, w_073_4774, w_073_4775, w_073_4777, w_073_4782, w_073_4785, w_073_4786, w_073_4794, w_073_4798, w_073_4800, w_073_4802, w_073_4806, w_073_4812, w_073_4814, w_073_4815, w_073_4817, w_073_4818, w_073_4824, w_073_4826, w_073_4828, w_073_4830, w_073_4831, w_073_4833, w_073_4837, w_073_4838, w_073_4840, w_073_4844, w_073_4845, w_073_4847, w_073_4849, w_073_4852, w_073_4855, w_073_4856, w_073_4857, w_073_4859, w_073_4861, w_073_4865, w_073_4868, w_073_4869, w_073_4872, w_073_4875, w_073_4880, w_073_4889, w_073_4896, w_073_4899, w_073_4901, w_073_4903, w_073_4912, w_073_4915, w_073_4935, w_073_4936, w_073_4942, w_073_4946, w_073_4949, w_073_4951, w_073_4954, w_073_4955, w_073_4958, w_073_4959, w_073_4960, w_073_4967, w_073_4969, w_073_4970, w_073_4973, w_073_4975, w_073_4977, w_073_4979, w_073_4986, w_073_4988, w_073_4994, w_073_5002, w_073_5003, w_073_5007, w_073_5019, w_073_5020, w_073_5024, w_073_5026, w_073_5031, w_073_5041, w_073_5043, w_073_5044, w_073_5046, w_073_5051, w_073_5054, w_073_5060, w_073_5061, w_073_5076, w_073_5080, w_073_5083, w_073_5084, w_073_5085, w_073_5097, w_073_5098, w_073_5101, w_073_5102, w_073_5115, w_073_5119, w_073_5123, w_073_5124, w_073_5125, w_073_5130, w_073_5133, w_073_5142, w_073_5144, w_073_5148, w_073_5151, w_073_5153, w_073_5156, w_073_5157, w_073_5158, w_073_5159, w_073_5160, w_073_5162, w_073_5164, w_073_5167, w_073_5169, w_073_5170, w_073_5171, w_073_5173, w_073_5175, w_073_5177, w_073_5178, w_073_5179, w_073_5186, w_073_5188, w_073_5189, w_073_5194, w_073_5196, w_073_5198, w_073_5202, w_073_5207, w_073_5210, w_073_5213, w_073_5214, w_073_5217, w_073_5218, w_073_5222, w_073_5228, w_073_5229, w_073_5230, w_073_5233, w_073_5238, w_073_5240, w_073_5242, w_073_5246, w_073_5248, w_073_5250, w_073_5251, w_073_5255, w_073_5262, w_073_5267, w_073_5268, w_073_5269, w_073_5275, w_073_5276, w_073_5280, w_073_5289, w_073_5292, w_073_5293, w_073_5294, w_073_5299, w_073_5310, w_073_5311, w_073_5319, w_073_5328, w_073_5335, w_073_5336, w_073_5338, w_073_5339, w_073_5342, w_073_5349, w_073_5357, w_073_5359, w_073_5361, w_073_5364, w_073_5366, w_073_5367, w_073_5368, w_073_5369, w_073_5370, w_073_5372, w_073_5374, w_073_5376, w_073_5378, w_073_5380, w_073_5388, w_073_5391, w_073_5394, w_073_5396, w_073_5406, w_073_5413, w_073_5414, w_073_5416, w_073_5433, w_073_5437, w_073_5443, w_073_5444, w_073_5445, w_073_5447, w_073_5451, w_073_5453, w_073_5454, w_073_5463, w_073_5464, w_073_5465, w_073_5469, w_073_5470, w_073_5473, w_073_5479, w_073_5480, w_073_5482, w_073_5485, w_073_5488, w_073_5491, w_073_5495, w_073_5501, w_073_5503, w_073_5512, w_073_5516, w_073_5521, w_073_5525, w_073_5539, w_073_5542, w_073_5543, w_073_5544, w_073_5545, w_073_5546, w_073_5547, w_073_5553, w_073_5558, w_073_5559, w_073_5562, w_073_5563, w_073_5566, w_073_5567, w_073_5568, w_073_5569, w_073_5570, w_073_5574, w_073_5576, w_073_5577, w_073_5581, w_073_5583, w_073_5589, w_073_5591, w_073_5593, w_073_5594, w_073_5603, w_073_5608, w_073_5612, w_073_5613, w_073_5618, w_073_5619, w_073_5620, w_073_5621, w_073_5628, w_073_5635, w_073_5641, w_073_5643, w_073_5644, w_073_5651, w_073_5653, w_073_5656, w_073_5659, w_073_5665, w_073_5669, w_073_5671, w_073_5672, w_073_5673, w_073_5674, w_073_5675, w_073_5680, w_073_5686, w_073_5687, w_073_5691, w_073_5692, w_073_5697, w_073_5710, w_073_5711, w_073_5712, w_073_5713, w_073_5720, w_073_5721, w_073_5723, w_073_5725, w_073_5727, w_073_5729, w_073_5732, w_073_5733, w_073_5734, w_073_5739, w_073_5745, w_073_5752, w_073_5756, w_073_5757, w_073_5763, w_073_5768, w_073_5769, w_073_5772, w_073_5773, w_073_5774, w_073_5777, w_073_5786, w_073_5789, w_073_5791, w_073_5799, w_073_5803, w_073_5805, w_073_5806, w_073_5812, w_073_5814, w_073_5815, w_073_5816, w_073_5819, w_073_5832, w_073_5834, w_073_5835, w_073_5843, w_073_5851, w_073_5856, w_073_5857, w_073_5859, w_073_5863, w_073_5864, w_073_5865, w_073_5871, w_073_5872, w_073_5882, w_073_5884, w_073_5888, w_073_5895, w_073_5899, w_073_5906, w_073_5907, w_073_5908, w_073_5909, w_073_5912, w_073_5914, w_073_5915, w_073_5919, w_073_5921, w_073_5923, w_073_5924, w_073_5932, w_073_5933, w_073_5935, w_073_5936, w_073_5938, w_073_5944, w_073_5948, w_073_5949, w_073_5951, w_073_5954, w_073_5956, w_073_5957, w_073_5959, w_073_5962, w_073_5966, w_073_5969, w_073_5970, w_073_5973, w_073_5974, w_073_5975, w_073_5977;
  wire w_074_000, w_074_001, w_074_002, w_074_003, w_074_004, w_074_006, w_074_007, w_074_008, w_074_009, w_074_010, w_074_011, w_074_012, w_074_013, w_074_014, w_074_015, w_074_016, w_074_017, w_074_018, w_074_019, w_074_020, w_074_021, w_074_022, w_074_023, w_074_024, w_074_025, w_074_026, w_074_027, w_074_028, w_074_029, w_074_030, w_074_031, w_074_032, w_074_033, w_074_034, w_074_035, w_074_037, w_074_038, w_074_039, w_074_040, w_074_041, w_074_042, w_074_043, w_074_044, w_074_046, w_074_047, w_074_048, w_074_050, w_074_051, w_074_052, w_074_053, w_074_054, w_074_055, w_074_056, w_074_057, w_074_058, w_074_059, w_074_061, w_074_064, w_074_066, w_074_067, w_074_068, w_074_069, w_074_070, w_074_071, w_074_072, w_074_073, w_074_074, w_074_075, w_074_076, w_074_078, w_074_079, w_074_080, w_074_081, w_074_082, w_074_083, w_074_084, w_074_085, w_074_086, w_074_087, w_074_088, w_074_090, w_074_091, w_074_092, w_074_094, w_074_095, w_074_099, w_074_100, w_074_101, w_074_102, w_074_103, w_074_105, w_074_106, w_074_107, w_074_108, w_074_109, w_074_110, w_074_111, w_074_114, w_074_115, w_074_116, w_074_118, w_074_120, w_074_121, w_074_122, w_074_123, w_074_125, w_074_126, w_074_128, w_074_129, w_074_131, w_074_132, w_074_133, w_074_135, w_074_136, w_074_137, w_074_138, w_074_139, w_074_140, w_074_143, w_074_144, w_074_145, w_074_146, w_074_148, w_074_149, w_074_151, w_074_152, w_074_153, w_074_154, w_074_156, w_074_157, w_074_158, w_074_159, w_074_160, w_074_161, w_074_162, w_074_163, w_074_164, w_074_166, w_074_167, w_074_168, w_074_169, w_074_170, w_074_171, w_074_172, w_074_173, w_074_175, w_074_176, w_074_177, w_074_179, w_074_180, w_074_182, w_074_183, w_074_184, w_074_185, w_074_186, w_074_187, w_074_188, w_074_191, w_074_193, w_074_194, w_074_196, w_074_197, w_074_198, w_074_200, w_074_201, w_074_202, w_074_203, w_074_204, w_074_205, w_074_206, w_074_207, w_074_208, w_074_209, w_074_210, w_074_211, w_074_212, w_074_213, w_074_214, w_074_215, w_074_216, w_074_217, w_074_219, w_074_220, w_074_221, w_074_222, w_074_223, w_074_224, w_074_225, w_074_226, w_074_227, w_074_229, w_074_230, w_074_232, w_074_233, w_074_234, w_074_235, w_074_236, w_074_238, w_074_239, w_074_240, w_074_241, w_074_242, w_074_243, w_074_244, w_074_245, w_074_246, w_074_247, w_074_248, w_074_249, w_074_250, w_074_251, w_074_252, w_074_254, w_074_255, w_074_256, w_074_258, w_074_259, w_074_260, w_074_261, w_074_262, w_074_263, w_074_264, w_074_265, w_074_266, w_074_267, w_074_268, w_074_270, w_074_271, w_074_273, w_074_274, w_074_275, w_074_276, w_074_277, w_074_278, w_074_279, w_074_280, w_074_281, w_074_282, w_074_283, w_074_284, w_074_285, w_074_286, w_074_287, w_074_288, w_074_289, w_074_290, w_074_291, w_074_293, w_074_294, w_074_295, w_074_296, w_074_297, w_074_298, w_074_299, w_074_300, w_074_301, w_074_302, w_074_303, w_074_304, w_074_305, w_074_307, w_074_308, w_074_309, w_074_310, w_074_311, w_074_312, w_074_313, w_074_314, w_074_315, w_074_316, w_074_318, w_074_320, w_074_321, w_074_322, w_074_323, w_074_324, w_074_325, w_074_326, w_074_327, w_074_328, w_074_329, w_074_330, w_074_332, w_074_333, w_074_334, w_074_336, w_074_337, w_074_338, w_074_340, w_074_342, w_074_343, w_074_344, w_074_345, w_074_346, w_074_347, w_074_348, w_074_349, w_074_350, w_074_351, w_074_352, w_074_353, w_074_354, w_074_356, w_074_357, w_074_358, w_074_359, w_074_361, w_074_362, w_074_363, w_074_364, w_074_365, w_074_366, w_074_367, w_074_368, w_074_369, w_074_370, w_074_372, w_074_373, w_074_374, w_074_376, w_074_377, w_074_380, w_074_381, w_074_382, w_074_383, w_074_385, w_074_386, w_074_387, w_074_388, w_074_390, w_074_391, w_074_392, w_074_394, w_074_395, w_074_396, w_074_397, w_074_398, w_074_399, w_074_401, w_074_402, w_074_403, w_074_404, w_074_405, w_074_406, w_074_407, w_074_408, w_074_409, w_074_410, w_074_411, w_074_414, w_074_415, w_074_416, w_074_417, w_074_419, w_074_420, w_074_421, w_074_422, w_074_423, w_074_424, w_074_425, w_074_426, w_074_428, w_074_429, w_074_430, w_074_431, w_074_432, w_074_433, w_074_435, w_074_436, w_074_437, w_074_438, w_074_439, w_074_440, w_074_441, w_074_442, w_074_443, w_074_445, w_074_446, w_074_447, w_074_448, w_074_450, w_074_451, w_074_452, w_074_453, w_074_454, w_074_455, w_074_458, w_074_459, w_074_460, w_074_461, w_074_462, w_074_464, w_074_465, w_074_466, w_074_467, w_074_468, w_074_469, w_074_470, w_074_471, w_074_472, w_074_473, w_074_474, w_074_475, w_074_477, w_074_478, w_074_479, w_074_480, w_074_481, w_074_482, w_074_483, w_074_484, w_074_485, w_074_486, w_074_487, w_074_488, w_074_489, w_074_490, w_074_491, w_074_492, w_074_493, w_074_494, w_074_495, w_074_496, w_074_497, w_074_498, w_074_499, w_074_500, w_074_501, w_074_503, w_074_504, w_074_506, w_074_507, w_074_509, w_074_510, w_074_511, w_074_512, w_074_513, w_074_514, w_074_515, w_074_516, w_074_517, w_074_520, w_074_521, w_074_522, w_074_523, w_074_526, w_074_528, w_074_529, w_074_530, w_074_531, w_074_532, w_074_533, w_074_534, w_074_535, w_074_536, w_074_538, w_074_539, w_074_540, w_074_541, w_074_542, w_074_543, w_074_544, w_074_545, w_074_546, w_074_547, w_074_548, w_074_549, w_074_550, w_074_551, w_074_552, w_074_555, w_074_556, w_074_560, w_074_561, w_074_562, w_074_563, w_074_564, w_074_565, w_074_566, w_074_567, w_074_568, w_074_569, w_074_570, w_074_572, w_074_573, w_074_574, w_074_575, w_074_578, w_074_579, w_074_580, w_074_581, w_074_582, w_074_583, w_074_584, w_074_587, w_074_588, w_074_589, w_074_590, w_074_591, w_074_592, w_074_593, w_074_595, w_074_596, w_074_598, w_074_599, w_074_600, w_074_601, w_074_603, w_074_604, w_074_606, w_074_607, w_074_608, w_074_609, w_074_610, w_074_611, w_074_612, w_074_613, w_074_614, w_074_615, w_074_616, w_074_618, w_074_619, w_074_620, w_074_621, w_074_622, w_074_623, w_074_624, w_074_625, w_074_626, w_074_627, w_074_628, w_074_629, w_074_630, w_074_631, w_074_633, w_074_636, w_074_638, w_074_639, w_074_640, w_074_641, w_074_642, w_074_643, w_074_645, w_074_646, w_074_648, w_074_649, w_074_650, w_074_653, w_074_654, w_074_655, w_074_656, w_074_657, w_074_658, w_074_659, w_074_660, w_074_661, w_074_662, w_074_663, w_074_664, w_074_665, w_074_666, w_074_667, w_074_668, w_074_669, w_074_670, w_074_671, w_074_673, w_074_674, w_074_675, w_074_676, w_074_677, w_074_678, w_074_679, w_074_680, w_074_681, w_074_684, w_074_685, w_074_686, w_074_688, w_074_689, w_074_691, w_074_692, w_074_693, w_074_694, w_074_695, w_074_696, w_074_697, w_074_698, w_074_699, w_074_700, w_074_701, w_074_704, w_074_705, w_074_706, w_074_707, w_074_709, w_074_710, w_074_711, w_074_712, w_074_715, w_074_716, w_074_717, w_074_718, w_074_719, w_074_720, w_074_722, w_074_723, w_074_724, w_074_725, w_074_726, w_074_727, w_074_729, w_074_731, w_074_733, w_074_735, w_074_736, w_074_737, w_074_738, w_074_739, w_074_740, w_074_741, w_074_742, w_074_743, w_074_744, w_074_745, w_074_746, w_074_748, w_074_749, w_074_750, w_074_751, w_074_752, w_074_753, w_074_754, w_074_755, w_074_756, w_074_758, w_074_759, w_074_760, w_074_761, w_074_762, w_074_764, w_074_765, w_074_766, w_074_767, w_074_768, w_074_769, w_074_770, w_074_772, w_074_773, w_074_774, w_074_775, w_074_776, w_074_777, w_074_778, w_074_780, w_074_783, w_074_784, w_074_785, w_074_786, w_074_787, w_074_788, w_074_789, w_074_790, w_074_791, w_074_792, w_074_794, w_074_795, w_074_796, w_074_797, w_074_798, w_074_799, w_074_800, w_074_801, w_074_802, w_074_805, w_074_806, w_074_807, w_074_808, w_074_809, w_074_810, w_074_812, w_074_813, w_074_814, w_074_815, w_074_816, w_074_817, w_074_818, w_074_819, w_074_820, w_074_822, w_074_824, w_074_827, w_074_828, w_074_830, w_074_831, w_074_832, w_074_833, w_074_834, w_074_835, w_074_836, w_074_837, w_074_840, w_074_841, w_074_843, w_074_844, w_074_846, w_074_847, w_074_848, w_074_849, w_074_850, w_074_852, w_074_853, w_074_854, w_074_855, w_074_856, w_074_858, w_074_859, w_074_861, w_074_862, w_074_863, w_074_864, w_074_865, w_074_866, w_074_867, w_074_868, w_074_869, w_074_870, w_074_871, w_074_872, w_074_873, w_074_874, w_074_875, w_074_876, w_074_877, w_074_879, w_074_880, w_074_881, w_074_883, w_074_884, w_074_885, w_074_886, w_074_887, w_074_888, w_074_890, w_074_891, w_074_892, w_074_893, w_074_895, w_074_896, w_074_897, w_074_898, w_074_899, w_074_900, w_074_901, w_074_902, w_074_903, w_074_904, w_074_905, w_074_906, w_074_907, w_074_908, w_074_909, w_074_910, w_074_911, w_074_912, w_074_914, w_074_915, w_074_916, w_074_917, w_074_918, w_074_919, w_074_920, w_074_921, w_074_922, w_074_924, w_074_925, w_074_928, w_074_929, w_074_930, w_074_931, w_074_932, w_074_933, w_074_934, w_074_935, w_074_936, w_074_937, w_074_938, w_074_940, w_074_941, w_074_942, w_074_943, w_074_945, w_074_946, w_074_947, w_074_948, w_074_949, w_074_950, w_074_952, w_074_953, w_074_954, w_074_955, w_074_957, w_074_959, w_074_960, w_074_961, w_074_962, w_074_964, w_074_965, w_074_966, w_074_967, w_074_968, w_074_969, w_074_970, w_074_972, w_074_973, w_074_975, w_074_976, w_074_978, w_074_979, w_074_980, w_074_981, w_074_983, w_074_984, w_074_985, w_074_986, w_074_987, w_074_988, w_074_989, w_074_990, w_074_991, w_074_992, w_074_993, w_074_994, w_074_995, w_074_996, w_074_997, w_074_998, w_074_999, w_074_1000, w_074_1002, w_074_1003, w_074_1004, w_074_1005, w_074_1006, w_074_1007, w_074_1008, w_074_1010, w_074_1011, w_074_1012, w_074_1013, w_074_1014, w_074_1016, w_074_1017, w_074_1019, w_074_1020, w_074_1022, w_074_1023, w_074_1024, w_074_1025, w_074_1027, w_074_1028, w_074_1030, w_074_1031, w_074_1032, w_074_1033, w_074_1034, w_074_1035, w_074_1036, w_074_1037, w_074_1038, w_074_1039, w_074_1040, w_074_1041, w_074_1042, w_074_1043, w_074_1044, w_074_1045, w_074_1046, w_074_1047, w_074_1049, w_074_1050, w_074_1052, w_074_1053, w_074_1054, w_074_1055, w_074_1057, w_074_1058, w_074_1059, w_074_1060, w_074_1061, w_074_1062, w_074_1063, w_074_1064, w_074_1065, w_074_1066, w_074_1067, w_074_1068, w_074_1069, w_074_1070, w_074_1071, w_074_1072, w_074_1073, w_074_1076, w_074_1078, w_074_1080, w_074_1081, w_074_1082, w_074_1084, w_074_1087, w_074_1088, w_074_1089, w_074_1090, w_074_1092, w_074_1093, w_074_1094, w_074_1095, w_074_1096, w_074_1097, w_074_1098, w_074_1099, w_074_1101, w_074_1102, w_074_1103, w_074_1104, w_074_1105, w_074_1106, w_074_1107, w_074_1108, w_074_1109, w_074_1110, w_074_1111, w_074_1112, w_074_1114, w_074_1116, w_074_1117, w_074_1118, w_074_1119, w_074_1120, w_074_1121, w_074_1122, w_074_1123, w_074_1124, w_074_1126, w_074_1127, w_074_1128, w_074_1129, w_074_1130, w_074_1132, w_074_1133, w_074_1134, w_074_1135, w_074_1136, w_074_1137, w_074_1139, w_074_1140, w_074_1141, w_074_1142, w_074_1143, w_074_1144, w_074_1145, w_074_1147, w_074_1148, w_074_1150, w_074_1153, w_074_1154, w_074_1156, w_074_1157, w_074_1158, w_074_1159, w_074_1160, w_074_1163, w_074_1164, w_074_1165, w_074_1166, w_074_1167, w_074_1168, w_074_1169, w_074_1170, w_074_1171, w_074_1173, w_074_1174, w_074_1176, w_074_1177, w_074_1178, w_074_1179, w_074_1180, w_074_1181, w_074_1182, w_074_1183, w_074_1184, w_074_1185, w_074_1186, w_074_1187, w_074_1189, w_074_1190, w_074_1191, w_074_1193, w_074_1194, w_074_1196, w_074_1197, w_074_1199, w_074_1200, w_074_1201, w_074_1202, w_074_1203, w_074_1205, w_074_1206, w_074_1207, w_074_1209, w_074_1211, w_074_1212, w_074_1213, w_074_1214, w_074_1215, w_074_1217, w_074_1218, w_074_1219, w_074_1220, w_074_1222, w_074_1223, w_074_1224, w_074_1225, w_074_1226, w_074_1228, w_074_1230, w_074_1231, w_074_1232, w_074_1233, w_074_1234, w_074_1235, w_074_1236, w_074_1237, w_074_1238, w_074_1239, w_074_1240, w_074_1242, w_074_1243, w_074_1244, w_074_1245, w_074_1246, w_074_1247, w_074_1248, w_074_1249, w_074_1251, w_074_1253, w_074_1254, w_074_1255, w_074_1256, w_074_1258, w_074_1259, w_074_1260, w_074_1261, w_074_1262, w_074_1263, w_074_1264, w_074_1265, w_074_1267, w_074_1268, w_074_1269, w_074_1270, w_074_1271, w_074_1272, w_074_1273, w_074_1274, w_074_1275, w_074_1276, w_074_1277, w_074_1278, w_074_1279, w_074_1280, w_074_1281, w_074_1283, w_074_1284, w_074_1285, w_074_1287, w_074_1288, w_074_1290, w_074_1291, w_074_1292, w_074_1293, w_074_1294, w_074_1295, w_074_1296, w_074_1299, w_074_1300, w_074_1301, w_074_1303, w_074_1304, w_074_1305, w_074_1306, w_074_1307, w_074_1308, w_074_1309, w_074_1310, w_074_1313, w_074_1314, w_074_1315, w_074_1316, w_074_1318, w_074_1319, w_074_1320, w_074_1321, w_074_1322, w_074_1324, w_074_1325, w_074_1326, w_074_1327, w_074_1328, w_074_1329, w_074_1330, w_074_1332, w_074_1333, w_074_1334, w_074_1335, w_074_1336, w_074_1337, w_074_1339, w_074_1340, w_074_1341, w_074_1342, w_074_1343, w_074_1344, w_074_1345, w_074_1346, w_074_1347, w_074_1348, w_074_1349, w_074_1350, w_074_1351, w_074_1352, w_074_1353, w_074_1355, w_074_1356, w_074_1357, w_074_1358, w_074_1359, w_074_1360, w_074_1361, w_074_1362, w_074_1363, w_074_1364, w_074_1365, w_074_1366, w_074_1367, w_074_1368, w_074_1369, w_074_1370, w_074_1371, w_074_1373, w_074_1375, w_074_1376, w_074_1377, w_074_1379, w_074_1381, w_074_1382, w_074_1383, w_074_1384, w_074_1385, w_074_1386, w_074_1389, w_074_1390, w_074_1392, w_074_1393, w_074_1394, w_074_1395, w_074_1396, w_074_1397, w_074_1399, w_074_1400, w_074_1401, w_074_1402, w_074_1403, w_074_1404, w_074_1405, w_074_1408, w_074_1409, w_074_1410, w_074_1411, w_074_1412, w_074_1413, w_074_1414, w_074_1415, w_074_1416, w_074_1418, w_074_1419, w_074_1420, w_074_1422, w_074_1424, w_074_1425, w_074_1426, w_074_1428, w_074_1429, w_074_1431, w_074_1432, w_074_1433, w_074_1435, w_074_1436, w_074_1437, w_074_1438, w_074_1440, w_074_1441, w_074_1442, w_074_1443, w_074_1444, w_074_1446, w_074_1447, w_074_1448, w_074_1449, w_074_1450, w_074_1451, w_074_1452, w_074_1453, w_074_1455, w_074_1456, w_074_1457, w_074_1458, w_074_1459, w_074_1460, w_074_1461, w_074_1463, w_074_1464, w_074_1465, w_074_1466, w_074_1467, w_074_1469, w_074_1470, w_074_1471, w_074_1472, w_074_1473, w_074_1474, w_074_1476, w_074_1478, w_074_1479, w_074_1480, w_074_1481, w_074_1483, w_074_1484, w_074_1485, w_074_1486, w_074_1487, w_074_1488, w_074_1490, w_074_1491, w_074_1492, w_074_1493, w_074_1494, w_074_1495, w_074_1497, w_074_1498, w_074_1499, w_074_1500, w_074_1501, w_074_1503, w_074_1505, w_074_1507, w_074_1509, w_074_1510, w_074_1511, w_074_1512, w_074_1513, w_074_1515, w_074_1516, w_074_1517, w_074_1519, w_074_1520, w_074_1522, w_074_1523, w_074_1524, w_074_1525, w_074_1527, w_074_1530, w_074_1531, w_074_1533, w_074_1534, w_074_1535, w_074_1536, w_074_1537, w_074_1539, w_074_1541, w_074_1542, w_074_1543, w_074_1544, w_074_1545, w_074_1546, w_074_1548, w_074_1549, w_074_1550, w_074_1551, w_074_1552, w_074_1553, w_074_1554, w_074_1555, w_074_1556, w_074_1557, w_074_1559, w_074_1560, w_074_1561, w_074_1563, w_074_1564, w_074_1565, w_074_1566, w_074_1567, w_074_1568, w_074_1569, w_074_1570, w_074_1571, w_074_1572, w_074_1573, w_074_1574, w_074_1575, w_074_1576, w_074_1577, w_074_1578, w_074_1579, w_074_1580, w_074_1581, w_074_1582, w_074_1583, w_074_1584, w_074_1585, w_074_1586, w_074_1587, w_074_1588, w_074_1589, w_074_1591, w_074_1592, w_074_1593, w_074_1595, w_074_1597, w_074_1600, w_074_1601, w_074_1602, w_074_1603, w_074_1604, w_074_1605, w_074_1606, w_074_1607, w_074_1608, w_074_1609, w_074_1611, w_074_1612, w_074_1614, w_074_1615, w_074_1616, w_074_1617, w_074_1618, w_074_1619, w_074_1620, w_074_1621, w_074_1622, w_074_1624, w_074_1625, w_074_1626, w_074_1627, w_074_1628, w_074_1629, w_074_1630, w_074_1631, w_074_1632, w_074_1633, w_074_1634, w_074_1635, w_074_1636, w_074_1637, w_074_1638, w_074_1639, w_074_1640, w_074_1642, w_074_1643, w_074_1644, w_074_1645, w_074_1646, w_074_1647, w_074_1648, w_074_1649, w_074_1650, w_074_1651, w_074_1653, w_074_1654, w_074_1655, w_074_1656, w_074_1657, w_074_1658, w_074_1659, w_074_1661, w_074_1662, w_074_1663, w_074_1664, w_074_1665, w_074_1666, w_074_1667, w_074_1669, w_074_1670, w_074_1673, w_074_1674, w_074_1675, w_074_1676, w_074_1678, w_074_1679, w_074_1680, w_074_1681, w_074_1682, w_074_1683, w_074_1684, w_074_1685, w_074_1687, w_074_1688, w_074_1690, w_074_1691, w_074_1692, w_074_1693, w_074_1695, w_074_1696, w_074_1697, w_074_1699, w_074_1700, w_074_1701, w_074_1702, w_074_1703, w_074_1704, w_074_1707, w_074_1710, w_074_1711, w_074_1712, w_074_1713, w_074_1714, w_074_1716, w_074_1717, w_074_1718, w_074_1719, w_074_1720, w_074_1723, w_074_1724, w_074_1725, w_074_1726, w_074_1727, w_074_1728, w_074_1729, w_074_1730, w_074_1731, w_074_1733, w_074_1734, w_074_1735, w_074_1736, w_074_1737, w_074_1739, w_074_1740, w_074_1741, w_074_1742, w_074_1743, w_074_1744, w_074_1745, w_074_1749, w_074_1750, w_074_1751, w_074_1752, w_074_1753, w_074_1754, w_074_1755, w_074_1756, w_074_1757, w_074_1758, w_074_1759, w_074_1761, w_074_1762, w_074_1763, w_074_1764, w_074_1765, w_074_1766, w_074_1767, w_074_1769, w_074_1770, w_074_1772, w_074_1773, w_074_1774, w_074_1776, w_074_1777, w_074_1778, w_074_1779, w_074_1780, w_074_1781, w_074_1783, w_074_1784, w_074_1785, w_074_1786, w_074_1787, w_074_1788, w_074_1789, w_074_1790, w_074_1791, w_074_1792, w_074_1794, w_074_1795, w_074_1796, w_074_1797, w_074_1798, w_074_1799, w_074_1800, w_074_1802, w_074_1803, w_074_1804, w_074_1805, w_074_1806, w_074_1807, w_074_1809, w_074_1811, w_074_1812, w_074_1813, w_074_1814, w_074_1818, w_074_1819, w_074_1821, w_074_1822, w_074_1824, w_074_1825, w_074_1826, w_074_1828, w_074_1829, w_074_1830, w_074_1831, w_074_1832, w_074_1833, w_074_1834, w_074_1836, w_074_1838, w_074_1839, w_074_1840, w_074_1841, w_074_1842, w_074_1843, w_074_1844, w_074_1845, w_074_1846, w_074_1847, w_074_1848, w_074_1849, w_074_1850, w_074_1851, w_074_1852, w_074_1853, w_074_1854, w_074_1855, w_074_1856, w_074_1857, w_074_1858, w_074_1860, w_074_1861, w_074_1862, w_074_1863, w_074_1864, w_074_1865, w_074_1866, w_074_1867, w_074_1868, w_074_1869, w_074_1872, w_074_1874, w_074_1875, w_074_1876, w_074_1877, w_074_1878, w_074_1880, w_074_1881, w_074_1883, w_074_1885, w_074_1886, w_074_1887, w_074_1889, w_074_1891, w_074_1893, w_074_1894, w_074_1895, w_074_1896, w_074_1897, w_074_1898, w_074_1899, w_074_1900, w_074_1901, w_074_1902, w_074_1903, w_074_1904, w_074_1905, w_074_1906, w_074_1907, w_074_1909, w_074_1911, w_074_1912, w_074_1914, w_074_1915, w_074_1916, w_074_1917, w_074_1918, w_074_1919, w_074_1920, w_074_1921, w_074_1922, w_074_1923, w_074_1924, w_074_1925, w_074_1926, w_074_1927, w_074_1928, w_074_1929, w_074_1930, w_074_1931, w_074_1932, w_074_1933, w_074_1934, w_074_1935, w_074_1936, w_074_1937, w_074_1938, w_074_1939, w_074_1940, w_074_1942, w_074_1943, w_074_1944, w_074_1945, w_074_1946, w_074_1947, w_074_1948, w_074_1949, w_074_1950, w_074_1951, w_074_1953, w_074_1954, w_074_1955, w_074_1956, w_074_1957, w_074_1958, w_074_1959, w_074_1960, w_074_1961, w_074_1962, w_074_1964, w_074_1965, w_074_1966, w_074_1967, w_074_1970, w_074_1971, w_074_1972, w_074_1973, w_074_1974, w_074_1975, w_074_1976, w_074_1977, w_074_1978, w_074_1981, w_074_1983, w_074_1985, w_074_1986, w_074_1987, w_074_1988, w_074_1989, w_074_1990, w_074_1991, w_074_1993, w_074_1994, w_074_1996, w_074_1997, w_074_2000, w_074_2001;
  wire w_075_001, w_075_002, w_075_003, w_075_004, w_075_008, w_075_009, w_075_016, w_075_017, w_075_018, w_075_019, w_075_023, w_075_024, w_075_026, w_075_028, w_075_030, w_075_031, w_075_032, w_075_034, w_075_035, w_075_038, w_075_041, w_075_045, w_075_046, w_075_047, w_075_048, w_075_049, w_075_051, w_075_052, w_075_056, w_075_057, w_075_058, w_075_059, w_075_061, w_075_062, w_075_070, w_075_072, w_075_074, w_075_078, w_075_079, w_075_080, w_075_084, w_075_085, w_075_086, w_075_087, w_075_089, w_075_090, w_075_093, w_075_094, w_075_097, w_075_105, w_075_107, w_075_108, w_075_110, w_075_112, w_075_114, w_075_115, w_075_116, w_075_117, w_075_119, w_075_120, w_075_124, w_075_126, w_075_128, w_075_133, w_075_134, w_075_137, w_075_140, w_075_142, w_075_143, w_075_144, w_075_147, w_075_149, w_075_151, w_075_152, w_075_156, w_075_158, w_075_160, w_075_161, w_075_163, w_075_164, w_075_165, w_075_168, w_075_170, w_075_175, w_075_178, w_075_179, w_075_180, w_075_182, w_075_183, w_075_184, w_075_185, w_075_187, w_075_189, w_075_190, w_075_192, w_075_193, w_075_198, w_075_199, w_075_201, w_075_208, w_075_209, w_075_210, w_075_214, w_075_216, w_075_218, w_075_223, w_075_224, w_075_225, w_075_227, w_075_229, w_075_231, w_075_233, w_075_237, w_075_244, w_075_249, w_075_252, w_075_255, w_075_256, w_075_258, w_075_262, w_075_267, w_075_271, w_075_275, w_075_281, w_075_288, w_075_290, w_075_293, w_075_300, w_075_309, w_075_310, w_075_315, w_075_317, w_075_319, w_075_323, w_075_326, w_075_332, w_075_334, w_075_335, w_075_341, w_075_343, w_075_347, w_075_349, w_075_351, w_075_353, w_075_356, w_075_357, w_075_358, w_075_360, w_075_366, w_075_371, w_075_377, w_075_384, w_075_386, w_075_395, w_075_396, w_075_402, w_075_403, w_075_406, w_075_407, w_075_409, w_075_411, w_075_421, w_075_422, w_075_426, w_075_428, w_075_430, w_075_439, w_075_440, w_075_451, w_075_452, w_075_460, w_075_461, w_075_463, w_075_466, w_075_470, w_075_473, w_075_474, w_075_475, w_075_488, w_075_489, w_075_495, w_075_496, w_075_500, w_075_501, w_075_505, w_075_506, w_075_509, w_075_511, w_075_512, w_075_520, w_075_524, w_075_530, w_075_533, w_075_536, w_075_538, w_075_539, w_075_545, w_075_549, w_075_551, w_075_552, w_075_558, w_075_559, w_075_565, w_075_568, w_075_571, w_075_581, w_075_593, w_075_597, w_075_598, w_075_600, w_075_603, w_075_606, w_075_607, w_075_608, w_075_611, w_075_612, w_075_613, w_075_617, w_075_624, w_075_627, w_075_629, w_075_637, w_075_641, w_075_645, w_075_646, w_075_647, w_075_648, w_075_649, w_075_650, w_075_656, w_075_658, w_075_659, w_075_663, w_075_666, w_075_667, w_075_669, w_075_675, w_075_676, w_075_682, w_075_694, w_075_711, w_075_712, w_075_714, w_075_721, w_075_724, w_075_725, w_075_726, w_075_730, w_075_731, w_075_732, w_075_737, w_075_738, w_075_739, w_075_741, w_075_743, w_075_745, w_075_749, w_075_752, w_075_753, w_075_754, w_075_757, w_075_758, w_075_759, w_075_760, w_075_761, w_075_768, w_075_777, w_075_784, w_075_786, w_075_788, w_075_792, w_075_793, w_075_802, w_075_805, w_075_806, w_075_808, w_075_810, w_075_811, w_075_819, w_075_821, w_075_825, w_075_827, w_075_828, w_075_830, w_075_833, w_075_835, w_075_836, w_075_842, w_075_845, w_075_846, w_075_847, w_075_849, w_075_850, w_075_855, w_075_856, w_075_857, w_075_858, w_075_860, w_075_862, w_075_864, w_075_870, w_075_881, w_075_883, w_075_887, w_075_894, w_075_898, w_075_907, w_075_908, w_075_911, w_075_912, w_075_915, w_075_916, w_075_917, w_075_919, w_075_920, w_075_925, w_075_926, w_075_927, w_075_929, w_075_930, w_075_931, w_075_941, w_075_944, w_075_949, w_075_951, w_075_953, w_075_957, w_075_959, w_075_960, w_075_961, w_075_964, w_075_966, w_075_967, w_075_971, w_075_977, w_075_980, w_075_990, w_075_992, w_075_994, w_075_1002, w_075_1005, w_075_1006, w_075_1015, w_075_1018, w_075_1019, w_075_1030, w_075_1033, w_075_1036, w_075_1038, w_075_1039, w_075_1043, w_075_1044, w_075_1049, w_075_1051, w_075_1053, w_075_1057, w_075_1065, w_075_1066, w_075_1072, w_075_1074, w_075_1075, w_075_1077, w_075_1078, w_075_1079, w_075_1081, w_075_1085, w_075_1090, w_075_1092, w_075_1094, w_075_1101, w_075_1108, w_075_1109, w_075_1112, w_075_1113, w_075_1114, w_075_1118, w_075_1120, w_075_1121, w_075_1122, w_075_1125, w_075_1126, w_075_1132, w_075_1137, w_075_1139, w_075_1141, w_075_1143, w_075_1144, w_075_1146, w_075_1153, w_075_1154, w_075_1171, w_075_1178, w_075_1181, w_075_1183, w_075_1185, w_075_1187, w_075_1191, w_075_1192, w_075_1202, w_075_1209, w_075_1219, w_075_1225, w_075_1226, w_075_1228, w_075_1229, w_075_1231, w_075_1232, w_075_1236, w_075_1246, w_075_1250, w_075_1265, w_075_1266, w_075_1280, w_075_1281, w_075_1283, w_075_1286, w_075_1287, w_075_1288, w_075_1291, w_075_1294, w_075_1297, w_075_1298, w_075_1301, w_075_1302, w_075_1304, w_075_1305, w_075_1311, w_075_1314, w_075_1329, w_075_1339, w_075_1340, w_075_1344, w_075_1345, w_075_1351, w_075_1356, w_075_1357, w_075_1359, w_075_1360, w_075_1362, w_075_1363, w_075_1366, w_075_1367, w_075_1370, w_075_1372, w_075_1379, w_075_1381, w_075_1389, w_075_1391, w_075_1393, w_075_1395, w_075_1396, w_075_1400, w_075_1404, w_075_1411, w_075_1412, w_075_1415, w_075_1417, w_075_1418, w_075_1420, w_075_1422, w_075_1425, w_075_1426, w_075_1430, w_075_1434, w_075_1443, w_075_1447, w_075_1455, w_075_1460, w_075_1466, w_075_1467, w_075_1472, w_075_1474, w_075_1475, w_075_1481, w_075_1483, w_075_1489, w_075_1490, w_075_1495, w_075_1499, w_075_1501, w_075_1506, w_075_1509, w_075_1512, w_075_1518, w_075_1521, w_075_1525, w_075_1531, w_075_1532, w_075_1545, w_075_1546, w_075_1548, w_075_1560, w_075_1563, w_075_1572, w_075_1573, w_075_1578, w_075_1580, w_075_1583, w_075_1586, w_075_1592, w_075_1593, w_075_1594, w_075_1595, w_075_1596, w_075_1599, w_075_1600, w_075_1602, w_075_1610, w_075_1619, w_075_1624, w_075_1627, w_075_1632, w_075_1635, w_075_1643, w_075_1645, w_075_1648, w_075_1650, w_075_1655, w_075_1656, w_075_1658, w_075_1662, w_075_1668, w_075_1669, w_075_1674, w_075_1678, w_075_1679, w_075_1680, w_075_1681, w_075_1682, w_075_1683, w_075_1685, w_075_1687, w_075_1691, w_075_1694, w_075_1700, w_075_1701, w_075_1706, w_075_1707, w_075_1712, w_075_1714, w_075_1719, w_075_1721, w_075_1723, w_075_1724, w_075_1726, w_075_1733, w_075_1735, w_075_1744, w_075_1746, w_075_1749, w_075_1750, w_075_1753, w_075_1755, w_075_1756, w_075_1757, w_075_1762, w_075_1763, w_075_1768, w_075_1776, w_075_1784, w_075_1788, w_075_1793, w_075_1803, w_075_1809, w_075_1812, w_075_1816, w_075_1823, w_075_1826, w_075_1828, w_075_1830, w_075_1831, w_075_1834, w_075_1835, w_075_1836, w_075_1837, w_075_1841, w_075_1843, w_075_1847, w_075_1848, w_075_1850, w_075_1851, w_075_1859, w_075_1861, w_075_1862, w_075_1864, w_075_1871, w_075_1876, w_075_1877, w_075_1879, w_075_1883, w_075_1885, w_075_1888, w_075_1889, w_075_1896, w_075_1898, w_075_1899, w_075_1907, w_075_1912, w_075_1914, w_075_1916, w_075_1917, w_075_1924, w_075_1937, w_075_1940, w_075_1942, w_075_1944, w_075_1946, w_075_1949, w_075_1954, w_075_1958, w_075_1965, w_075_1968, w_075_1979, w_075_1980, w_075_1982, w_075_1984, w_075_1986, w_075_1988, w_075_1990, w_075_1994, w_075_1995, w_075_1996, w_075_2000, w_075_2003, w_075_2006, w_075_2009, w_075_2014, w_075_2019, w_075_2021, w_075_2025, w_075_2026, w_075_2029, w_075_2031, w_075_2033, w_075_2035, w_075_2041, w_075_2045, w_075_2046, w_075_2048, w_075_2051, w_075_2052, w_075_2056, w_075_2060, w_075_2065, w_075_2066, w_075_2071, w_075_2078, w_075_2083, w_075_2087, w_075_2088, w_075_2090, w_075_2096, w_075_2102, w_075_2111, w_075_2114, w_075_2118, w_075_2119, w_075_2123, w_075_2131, w_075_2134, w_075_2137, w_075_2141, w_075_2143, w_075_2146, w_075_2148, w_075_2149, w_075_2153, w_075_2158, w_075_2163, w_075_2166, w_075_2178, w_075_2183, w_075_2189, w_075_2193, w_075_2198, w_075_2199, w_075_2202, w_075_2214, w_075_2216, w_075_2217, w_075_2219, w_075_2226, w_075_2229, w_075_2230, w_075_2234, w_075_2237, w_075_2244, w_075_2251, w_075_2254, w_075_2255, w_075_2261, w_075_2269, w_075_2273, w_075_2282, w_075_2297, w_075_2303, w_075_2304, w_075_2305, w_075_2308, w_075_2309, w_075_2311, w_075_2312, w_075_2315, w_075_2316, w_075_2318, w_075_2319, w_075_2323, w_075_2325, w_075_2329, w_075_2330, w_075_2332, w_075_2337, w_075_2347, w_075_2361, w_075_2365, w_075_2367, w_075_2368, w_075_2373, w_075_2374, w_075_2376, w_075_2382, w_075_2384, w_075_2386, w_075_2389, w_075_2394, w_075_2395, w_075_2398, w_075_2407, w_075_2413, w_075_2415, w_075_2418, w_075_2419, w_075_2422, w_075_2424, w_075_2429, w_075_2430, w_075_2435, w_075_2439, w_075_2440, w_075_2441, w_075_2446, w_075_2448, w_075_2451, w_075_2454, w_075_2458, w_075_2459, w_075_2460, w_075_2471, w_075_2476, w_075_2481, w_075_2490, w_075_2492, w_075_2493, w_075_2495, w_075_2502, w_075_2503, w_075_2507, w_075_2508, w_075_2512, w_075_2515, w_075_2520, w_075_2521, w_075_2522, w_075_2529, w_075_2535, w_075_2538, w_075_2542, w_075_2543, w_075_2557, w_075_2559, w_075_2562, w_075_2564, w_075_2565, w_075_2569, w_075_2570, w_075_2575, w_075_2577, w_075_2581, w_075_2586, w_075_2587, w_075_2588, w_075_2592, w_075_2595, w_075_2598, w_075_2603, w_075_2605, w_075_2606, w_075_2608, w_075_2609, w_075_2613, w_075_2615, w_075_2619, w_075_2621, w_075_2627, w_075_2631, w_075_2632, w_075_2633, w_075_2636, w_075_2638, w_075_2639, w_075_2640, w_075_2644, w_075_2646, w_075_2647, w_075_2649, w_075_2651, w_075_2652, w_075_2653, w_075_2663, w_075_2664, w_075_2665, w_075_2668, w_075_2670, w_075_2681, w_075_2682, w_075_2684, w_075_2688, w_075_2691, w_075_2694, w_075_2697, w_075_2711, w_075_2712, w_075_2716, w_075_2720, w_075_2729, w_075_2730, w_075_2736, w_075_2741, w_075_2746, w_075_2749, w_075_2755, w_075_2761, w_075_2763, w_075_2764, w_075_2767, w_075_2776, w_075_2783, w_075_2785, w_075_2814, w_075_2815, w_075_2816, w_075_2817, w_075_2818, w_075_2819, w_075_2820, w_075_2821, w_075_2827, w_075_2828, w_075_2832, w_075_2834, w_075_2837, w_075_2838, w_075_2843, w_075_2848, w_075_2849, w_075_2857, w_075_2863, w_075_2870, w_075_2871, w_075_2875, w_075_2876, w_075_2881, w_075_2886, w_075_2890, w_075_2891, w_075_2894, w_075_2896, w_075_2903, w_075_2904, w_075_2912, w_075_2916, w_075_2919, w_075_2924, w_075_2926, w_075_2929, w_075_2931, w_075_2933, w_075_2939, w_075_2941, w_075_2944, w_075_2951, w_075_2955, w_075_2961, w_075_2964, w_075_2965, w_075_2966, w_075_2974, w_075_2975, w_075_2976, w_075_2978, w_075_2982, w_075_2985, w_075_2991, w_075_2992, w_075_2994, w_075_2997, w_075_3000, w_075_3001, w_075_3002, w_075_3010, w_075_3013, w_075_3015, w_075_3020, w_075_3025, w_075_3026, w_075_3038, w_075_3039, w_075_3041, w_075_3046, w_075_3048, w_075_3049, w_075_3050, w_075_3051, w_075_3057, w_075_3068, w_075_3071, w_075_3075, w_075_3076, w_075_3077, w_075_3082, w_075_3086, w_075_3090, w_075_3092, w_075_3097, w_075_3101, w_075_3105, w_075_3108, w_075_3112, w_075_3113, w_075_3115, w_075_3119, w_075_3126, w_075_3127, w_075_3132, w_075_3137, w_075_3139, w_075_3143, w_075_3146, w_075_3148, w_075_3153, w_075_3156, w_075_3163, w_075_3177, w_075_3183, w_075_3188, w_075_3190, w_075_3194, w_075_3197, w_075_3200, w_075_3201, w_075_3202, w_075_3205, w_075_3206, w_075_3207, w_075_3212, w_075_3214, w_075_3221, w_075_3222, w_075_3225, w_075_3236, w_075_3239, w_075_3240, w_075_3241, w_075_3242, w_075_3243, w_075_3245, w_075_3248, w_075_3253, w_075_3255, w_075_3258, w_075_3259, w_075_3260, w_075_3276, w_075_3279, w_075_3282, w_075_3283, w_075_3291, w_075_3292, w_075_3301, w_075_3305, w_075_3307, w_075_3310, w_075_3313, w_075_3314, w_075_3321, w_075_3322, w_075_3323, w_075_3328, w_075_3330, w_075_3348, w_075_3349, w_075_3350, w_075_3351, w_075_3355, w_075_3358, w_075_3361, w_075_3365, w_075_3372, w_075_3373, w_075_3376, w_075_3377, w_075_3380, w_075_3381, w_075_3382, w_075_3383, w_075_3385, w_075_3386, w_075_3391, w_075_3392, w_075_3393, w_075_3394, w_075_3395, w_075_3400, w_075_3406, w_075_3410, w_075_3414, w_075_3415, w_075_3420, w_075_3422, w_075_3431, w_075_3432, w_075_3433, w_075_3436, w_075_3438, w_075_3443, w_075_3448, w_075_3452, w_075_3453, w_075_3455, w_075_3460, w_075_3462, w_075_3465, w_075_3466, w_075_3467, w_075_3471, w_075_3472, w_075_3473, w_075_3474, w_075_3476, w_075_3483, w_075_3485, w_075_3488, w_075_3496, w_075_3501, w_075_3502, w_075_3505, w_075_3506, w_075_3507, w_075_3508, w_075_3510, w_075_3513, w_075_3515, w_075_3518, w_075_3521, w_075_3528, w_075_3530, w_075_3533, w_075_3536, w_075_3538, w_075_3556, w_075_3557, w_075_3561, w_075_3564, w_075_3565, w_075_3571, w_075_3574, w_075_3581, w_075_3589, w_075_3594, w_075_3595, w_075_3598, w_075_3600, w_075_3601, w_075_3606, w_075_3607, w_075_3608, w_075_3609, w_075_3614, w_075_3616, w_075_3624, w_075_3632, w_075_3633, w_075_3645, w_075_3646, w_075_3651, w_075_3652, w_075_3654, w_075_3657, w_075_3659, w_075_3660, w_075_3663, w_075_3665, w_075_3669, w_075_3670, w_075_3675, w_075_3676, w_075_3677, w_075_3680, w_075_3681, w_075_3683, w_075_3686, w_075_3688, w_075_3692, w_075_3694, w_075_3695, w_075_3698, w_075_3701, w_075_3703, w_075_3704, w_075_3705, w_075_3708, w_075_3713, w_075_3716, w_075_3717, w_075_3724, w_075_3728, w_075_3731, w_075_3738, w_075_3739, w_075_3741, w_075_3743, w_075_3748, w_075_3750, w_075_3761, w_075_3763, w_075_3764, w_075_3768, w_075_3769, w_075_3772, w_075_3777, w_075_3780, w_075_3781, w_075_3784, w_075_3795, w_075_3797, w_075_3799, w_075_3800, w_075_3803, w_075_3806, w_075_3809, w_075_3815, w_075_3820, w_075_3822, w_075_3823, w_075_3824, w_075_3829, w_075_3831, w_075_3832, w_075_3840, w_075_3845, w_075_3852, w_075_3858, w_075_3862, w_075_3864, w_075_3865, w_075_3870, w_075_3871, w_075_3875, w_075_3876, w_075_3884, w_075_3888, w_075_3889, w_075_3890, w_075_3894, w_075_3905, w_075_3907, w_075_3912, w_075_3917, w_075_3918, w_075_3919, w_075_3932, w_075_3933, w_075_3936, w_075_3937, w_075_3938, w_075_3950, w_075_3957, w_075_3958, w_075_3961, w_075_3964, w_075_3973, w_075_3974, w_075_3976, w_075_3978, w_075_3979, w_075_3980, w_075_3982, w_075_3988, w_075_3989, w_075_3990, w_075_3991, w_075_3995, w_075_4000, w_075_4010, w_075_4011, w_075_4015, w_075_4016, w_075_4017, w_075_4022, w_075_4030, w_075_4037, w_075_4046, w_075_4051, w_075_4052, w_075_4070, w_075_4077, w_075_4078, w_075_4083, w_075_4088, w_075_4091, w_075_4093, w_075_4096, w_075_4100, w_075_4101, w_075_4106, w_075_4115, w_075_4120, w_075_4121, w_075_4126, w_075_4128, w_075_4136, w_075_4137, w_075_4141, w_075_4142, w_075_4146, w_075_4149, w_075_4151, w_075_4157, w_075_4160, w_075_4161, w_075_4164, w_075_4166, w_075_4170, w_075_4174, w_075_4175, w_075_4180, w_075_4181, w_075_4188, w_075_4197, w_075_4198, w_075_4200, w_075_4201, w_075_4206, w_075_4213, w_075_4223, w_075_4236, w_075_4242, w_075_4247, w_075_4250, w_075_4255, w_075_4257, w_075_4261, w_075_4262, w_075_4263, w_075_4265, w_075_4278, w_075_4283, w_075_4288, w_075_4293, w_075_4294, w_075_4296, w_075_4297, w_075_4298, w_075_4300, w_075_4301, w_075_4303, w_075_4305, w_075_4309, w_075_4313, w_075_4317, w_075_4320, w_075_4322, w_075_4324, w_075_4326, w_075_4327, w_075_4329, w_075_4332, w_075_4336, w_075_4339, w_075_4341, w_075_4343, w_075_4345, w_075_4346, w_075_4348, w_075_4352, w_075_4355, w_075_4361, w_075_4364, w_075_4365, w_075_4367, w_075_4369, w_075_4385, w_075_4386, w_075_4391, w_075_4392, w_075_4395, w_075_4397, w_075_4401, w_075_4404, w_075_4408, w_075_4409, w_075_4410, w_075_4413, w_075_4415, w_075_4416, w_075_4418, w_075_4425, w_075_4430, w_075_4432, w_075_4435, w_075_4436, w_075_4437, w_075_4439, w_075_4443, w_075_4445, w_075_4447, w_075_4459, w_075_4461, w_075_4472, w_075_4473, w_075_4475, w_075_4477, w_075_4479, w_075_4483, w_075_4487, w_075_4488, w_075_4494, w_075_4499, w_075_4506, w_075_4512, w_075_4515, w_075_4516, w_075_4517, w_075_4518, w_075_4521, w_075_4523, w_075_4524, w_075_4529, w_075_4530, w_075_4534, w_075_4543, w_075_4546, w_075_4554, w_075_4557, w_075_4558, w_075_4566, w_075_4581, w_075_4583, w_075_4588, w_075_4589, w_075_4596, w_075_4600, w_075_4602, w_075_4603, w_075_4612, w_075_4614, w_075_4616, w_075_4620, w_075_4623, w_075_4630, w_075_4632, w_075_4635, w_075_4638, w_075_4643, w_075_4645, w_075_4654, w_075_4656, w_075_4666, w_075_4668, w_075_4670, w_075_4674, w_075_4682, w_075_4685, w_075_4689, w_075_4696, w_075_4699, w_075_4700, w_075_4709, w_075_4722, w_075_4735, w_075_4736, w_075_4737, w_075_4745, w_075_4746, w_075_4747, w_075_4750, w_075_4755, w_075_4756, w_075_4757, w_075_4759, w_075_4762, w_075_4765, w_075_4767, w_075_4773, w_075_4774, w_075_4775, w_075_4781, w_075_4783, w_075_4793, w_075_4795, w_075_4799, w_075_4801, w_075_4802, w_075_4807, w_075_4809, w_075_4813, w_075_4816, w_075_4826, w_075_4829, w_075_4830, w_075_4832, w_075_4839, w_075_4857, w_075_4878, w_075_4883, w_075_4889, w_075_4890, w_075_4892, w_075_4902, w_075_4903, w_075_4908, w_075_4915, w_075_4916, w_075_4923, w_075_4932, w_075_4933, w_075_4934, w_075_4938, w_075_4940, w_075_4943, w_075_4946, w_075_4948, w_075_4953, w_075_4956, w_075_4959, w_075_4961, w_075_4963, w_075_4967, w_075_4969, w_075_4970, w_075_4971, w_075_4973, w_075_4979, w_075_4980, w_075_4981, w_075_4989, w_075_4990, w_075_4992, w_075_4993, w_075_4997, w_075_5001, w_075_5003, w_075_5007, w_075_5009, w_075_5010, w_075_5014, w_075_5018, w_075_5020, w_075_5021, w_075_5026, w_075_5031, w_075_5032, w_075_5034, w_075_5041, w_075_5042, w_075_5053, w_075_5054, w_075_5058, w_075_5061, w_075_5064, w_075_5074, w_075_5078, w_075_5079, w_075_5087, w_075_5091, w_075_5094, w_075_5096, w_075_5103, w_075_5107, w_075_5109, w_075_5110, w_075_5116, w_075_5117, w_075_5119, w_075_5121, w_075_5129, w_075_5132, w_075_5133, w_075_5136, w_075_5138, w_075_5140, w_075_5142, w_075_5146, w_075_5147, w_075_5148, w_075_5149, w_075_5150, w_075_5151, w_075_5165, w_075_5168, w_075_5173, w_075_5178, w_075_5182, w_075_5183, w_075_5189, w_075_5190, w_075_5194, w_075_5195, w_075_5196, w_075_5209, w_075_5215, w_075_5216, w_075_5223, w_075_5226, w_075_5230, w_075_5232, w_075_5236, w_075_5246, w_075_5253, w_075_5256, w_075_5259, w_075_5262, w_075_5267, w_075_5280, w_075_5281, w_075_5284, w_075_5299, w_075_5305, w_075_5307, w_075_5309, w_075_5314, w_075_5316, w_075_5317, w_075_5318, w_075_5319, w_075_5324, w_075_5330, w_075_5332, w_075_5340, w_075_5344, w_075_5345, w_075_5346, w_075_5347, w_075_5349, w_075_5350, w_075_5352, w_075_5353, w_075_5355, w_075_5360, w_075_5361, w_075_5362, w_075_5366, w_075_5367, w_075_5368, w_075_5370, w_075_5377, w_075_5378, w_075_5379, w_075_5383, w_075_5387, w_075_5390, w_075_5397, w_075_5404, w_075_5407, w_075_5413, w_075_5416, w_075_5431, w_075_5432, w_075_5433, w_075_5434, w_075_5439, w_075_5444, w_075_5448, w_075_5449, w_075_5450, w_075_5460, w_075_5470, w_075_5487, w_075_5491, w_075_5492, w_075_5493, w_075_5494, w_075_5496, w_075_5497, w_075_5502, w_075_5504, w_075_5509, w_075_5516, w_075_5523, w_075_5527, w_075_5528, w_075_5531, w_075_5532, w_075_5543, w_075_5547, w_075_5552, w_075_5553, w_075_5554, w_075_5557, w_075_5562, w_075_5565, w_075_5570, w_075_5571, w_075_5573, w_075_5578, w_075_5581, w_075_5589, w_075_5593, w_075_5603, w_075_5604, w_075_5610, w_075_5617, w_075_5626, w_075_5628, w_075_5629, w_075_5633, w_075_5640, w_075_5644, w_075_5645, w_075_5647, w_075_5651, w_075_5654, w_075_5655, w_075_5657, w_075_5659, w_075_5660, w_075_5661, w_075_5663, w_075_5664, w_075_5667, w_075_5668, w_075_5671, w_075_5678, w_075_5679, w_075_5681, w_075_5683, w_075_5685, w_075_5687, w_075_5688, w_075_5689, w_075_5690, w_075_5696, w_075_5703, w_075_5704, w_075_5705, w_075_5706, w_075_5709, w_075_5711, w_075_5716, w_075_5717, w_075_5721, w_075_5723, w_075_5727, w_075_5733, w_075_5737, w_075_5738, w_075_5754, w_075_5756, w_075_5759, w_075_5761, w_075_5769, w_075_5770, w_075_5772, w_075_5773, w_075_5774, w_075_5776, w_075_5778, w_075_5780, w_075_5781, w_075_5784, w_075_5786, w_075_5788, w_075_5789, w_075_5797, w_075_5798, w_075_5803, w_075_5814, w_075_5819, w_075_5820, w_075_5821, w_075_5826, w_075_5831, w_075_5837, w_075_5838, w_075_5839, w_075_5840, w_075_5844, w_075_5850, w_075_5853, w_075_5855, w_075_5862, w_075_5863, w_075_5864, w_075_5866, w_075_5867, w_075_5869, w_075_5870, w_075_5875, w_075_5876, w_075_5877, w_075_5878, w_075_5881, w_075_5883, w_075_5886, w_075_5888, w_075_5889, w_075_5890, w_075_5894, w_075_5900, w_075_5901, w_075_5905, w_075_5907, w_075_5908, w_075_5909, w_075_5912, w_075_5913, w_075_5919, w_075_5921, w_075_5925, w_075_5927, w_075_5929, w_075_5931, w_075_5932, w_075_5933, w_075_5934, w_075_5940, w_075_5943, w_075_5947, w_075_5948, w_075_5956, w_075_5960, w_075_5961, w_075_5962, w_075_5965, w_075_5970, w_075_5972, w_075_5973, w_075_5975, w_075_5977, w_075_5979, w_075_5989, w_075_5990, w_075_5993, w_075_5994, w_075_5995, w_075_5996, w_075_6000, w_075_6002, w_075_6007, w_075_6009, w_075_6011, w_075_6012, w_075_6015, w_075_6016, w_075_6022, w_075_6029, w_075_6033, w_075_6037, w_075_6039, w_075_6042, w_075_6044, w_075_6049, w_075_6053, w_075_6054, w_075_6055, w_075_6056, w_075_6060, w_075_6064, w_075_6066, w_075_6069, w_075_6074, w_075_6079, w_075_6081, w_075_6084, w_075_6085, w_075_6090, w_075_6091, w_075_6105, w_075_6110, w_075_6117, w_075_6119, w_075_6120, w_075_6123, w_075_6131, w_075_6132, w_075_6136, w_075_6137, w_075_6139, w_075_6140, w_075_6143, w_075_6144, w_075_6146, w_075_6150, w_075_6152, w_075_6153, w_075_6159, w_075_6163, w_075_6168, w_075_6173, w_075_6174, w_075_6178, w_075_6180, w_075_6189, w_075_6210, w_075_6211, w_075_6215, w_075_6216, w_075_6218, w_075_6220, w_075_6222, w_075_6228, w_075_6231, w_075_6232, w_075_6234, w_075_6235, w_075_6236, w_075_6237, w_075_6242, w_075_6244, w_075_6245, w_075_6251, w_075_6257, w_075_6259, w_075_6262, w_075_6267, w_075_6269, w_075_6270, w_075_6273, w_075_6274, w_075_6277, w_075_6282, w_075_6284, w_075_6288, w_075_6300, w_075_6301, w_075_6303, w_075_6304, w_075_6305, w_075_6307, w_075_6309, w_075_6311, w_075_6324, w_075_6327, w_075_6336, w_075_6338, w_075_6340, w_075_6342, w_075_6346, w_075_6349, w_075_6357, w_075_6359, w_075_6371, w_075_6372, w_075_6376, w_075_6378, w_075_6381, w_075_6382, w_075_6388, w_075_6395, w_075_6400, w_075_6402, w_075_6403, w_075_6407, w_075_6413, w_075_6417, w_075_6423, w_075_6425, w_075_6432, w_075_6438, w_075_6440, w_075_6443, w_075_6449, w_075_6450, w_075_6452, w_075_6459, w_075_6460, w_075_6463, w_075_6468, w_075_6469, w_075_6471, w_075_6478, w_075_6484, w_075_6486, w_075_6489, w_075_6498, w_075_6503, w_075_6506, w_075_6509, w_075_6511, w_075_6515, w_075_6516, w_075_6519, w_075_6524, w_075_6533, w_075_6535, w_075_6536, w_075_6538, w_075_6539, w_075_6543, w_075_6546, w_075_6551, w_075_6552, w_075_6553, w_075_6554, w_075_6555, w_075_6556, w_075_6558, w_075_6572, w_075_6578, w_075_6580, w_075_6581, w_075_6582, w_075_6583, w_075_6586, w_075_6588, w_075_6589, w_075_6591, w_075_6593, w_075_6597, w_075_6601, w_075_6603, w_075_6607, w_075_6609, w_075_6610, w_075_6618, w_075_6620, w_075_6621, w_075_6623, w_075_6633, w_075_6644, w_075_6645, w_075_6649, w_075_6656, w_075_6658, w_075_6659, w_075_6660, w_075_6664, w_075_6666, w_075_6670, w_075_6671, w_075_6672, w_075_6673, w_075_6674, w_075_6678, w_075_6680, w_075_6683, w_075_6686, w_075_6692, w_075_6694, w_075_6697, w_075_6705, w_075_6707, w_075_6708, w_075_6714, w_075_6719, w_075_6721, w_075_6725, w_075_6728, w_075_6729, w_075_6732, w_075_6733, w_075_6734, w_075_6735, w_075_6737, w_075_6741, w_075_6742, w_075_6746, w_075_6753, w_075_6754, w_075_6763, w_075_6766, w_075_6769, w_075_6770, w_075_6771, w_075_6772, w_075_6773, w_075_6786, w_075_6802, w_075_6808, w_075_6809, w_075_6811, w_075_6813, w_075_6814, w_075_6817, w_075_6818, w_075_6819, w_075_6821, w_075_6822, w_075_6823, w_075_6825, w_075_6834, w_075_6836, w_075_6846, w_075_6850, w_075_6858, w_075_6861, w_075_6862, w_075_6863, w_075_6864, w_075_6869, w_075_6870, w_075_6872, w_075_6874, w_075_6875, w_075_6877, w_075_6879, w_075_6885, w_075_6886, w_075_6889, w_075_6892, w_075_6893, w_075_6894, w_075_6896, w_075_6897, w_075_6900, w_075_6901, w_075_6902, w_075_6906, w_075_6922, w_075_6923, w_075_6924, w_075_6937, w_075_6941, w_075_6944, w_075_6945, w_075_6946, w_075_6947, w_075_6949, w_075_6953, w_075_6954, w_075_6959, w_075_6963, w_075_6964, w_075_6965, w_075_6967, w_075_6970, w_075_6972, w_075_6975, w_075_6977, w_075_6984, w_075_6988, w_075_6994, w_075_6999, w_075_7002, w_075_7008, w_075_7010, w_075_7012, w_075_7013, w_075_7018, w_075_7022, w_075_7025, w_075_7030, w_075_7031, w_075_7032, w_075_7033, w_075_7040, w_075_7043, w_075_7048, w_075_7050, w_075_7057, w_075_7068, w_075_7077, w_075_7082, w_075_7083, w_075_7086, w_075_7087, w_075_7090, w_075_7091, w_075_7096, w_075_7097, w_075_7101, w_075_7102, w_075_7103, w_075_7104, w_075_7107, w_075_7110, w_075_7114, w_075_7115, w_075_7123, w_075_7134, w_075_7139, w_075_7141, w_075_7149, w_075_7154, w_075_7158, w_075_7159, w_075_7161, w_075_7163, w_075_7164, w_075_7173, w_075_7176, w_075_7178, w_075_7180, w_075_7183, w_075_7188, w_075_7190, w_075_7192, w_075_7193, w_075_7194, w_075_7196, w_075_7202, w_075_7204, w_075_7205, w_075_7207, w_075_7210, w_075_7211, w_075_7216, w_075_7217, w_075_7219, w_075_7223, w_075_7226, w_075_7229, w_075_7232, w_075_7233, w_075_7236, w_075_7237, w_075_7239, w_075_7242, w_075_7244, w_075_7246, w_075_7249, w_075_7251, w_075_7252, w_075_7256, w_075_7259, w_075_7265, w_075_7271, w_075_7272, w_075_7276, w_075_7279, w_075_7283, w_075_7284, w_075_7292, w_075_7295, w_075_7305, w_075_7306, w_075_7310, w_075_7314, w_075_7320, w_075_7323, w_075_7326, w_075_7331, w_075_7336, w_075_7340, w_075_7342, w_075_7346, w_075_7347, w_075_7348, w_075_7351, w_075_7353, w_075_7354, w_075_7355, w_075_7357, w_075_7361, w_075_7366, w_075_7367, w_075_7371, w_075_7375, w_075_7377, w_075_7381, w_075_7382, w_075_7383, w_075_7386, w_075_7398, w_075_7401, w_075_7412, w_075_7414, w_075_7415, w_075_7416, w_075_7419, w_075_7420, w_075_7422, w_075_7425, w_075_7429, w_075_7431, w_075_7434, w_075_7436, w_075_7438, w_075_7440, w_075_7443, w_075_7446, w_075_7452, w_075_7453, w_075_7454, w_075_7458, w_075_7469, w_075_7470, w_075_7472, w_075_7473, w_075_7476, w_075_7479, w_075_7480, w_075_7482, w_075_7486, w_075_7489, w_075_7498, w_075_7504, w_075_7505, w_075_7509, w_075_7513, w_075_7514, w_075_7518, w_075_7521, w_075_7528, w_075_7529, w_075_7530, w_075_7532, w_075_7533, w_075_7534, w_075_7535, w_075_7538, w_075_7542, w_075_7543, w_075_7544, w_075_7545, w_075_7550, w_075_7551, w_075_7552, w_075_7556, w_075_7569, w_075_7571, w_075_7585, w_075_7596, w_075_7597, w_075_7600, w_075_7602, w_075_7611, w_075_7615, w_075_7621, w_075_7640, w_075_7644, w_075_7646, w_075_7651, w_075_7653, w_075_7655, w_075_7660, w_075_7661, w_075_7664, w_075_7667, w_075_7671, w_075_7673, w_075_7674, w_075_7676, w_075_7684, w_075_7689, w_075_7691, w_075_7695, w_075_7699, w_075_7701, w_075_7706, w_075_7709, w_075_7713, w_075_7714, w_075_7717, w_075_7720, w_075_7725, w_075_7727, w_075_7732, w_075_7733, w_075_7737, w_075_7743, w_075_7745, w_075_7749, w_075_7750, w_075_7756, w_075_7758, w_075_7761, w_075_7766, w_075_7767, w_075_7775, w_075_7776, w_075_7777, w_075_7783, w_075_7786, w_075_7790, w_075_7794, w_075_7797, w_075_7802, w_075_7803, w_075_7805, w_075_7807, w_075_7812, w_075_7816, w_075_7818, w_075_7821, w_075_7827, w_075_7832, w_075_7839, w_075_7843, w_075_7845, w_075_7846, w_075_7849, w_075_7869, w_075_7882, w_075_7888, w_075_7890, w_075_7891, w_075_7901, w_075_7914, w_075_7919, w_075_7934, w_075_7937, w_075_7939, w_075_7941, w_075_7948, w_075_7954, w_075_7959, w_075_7961, w_075_7967, w_075_7971, w_075_7972, w_075_7978, w_075_7981, w_075_7985, w_075_7988, w_075_7989, w_075_7995, w_075_8004, w_075_8005, w_075_8006, w_075_8007, w_075_8008, w_075_8012, w_075_8014, w_075_8017, w_075_8021, w_075_8022, w_075_8024, w_075_8025, w_075_8026, w_075_8028, w_075_8029, w_075_8032, w_075_8039, w_075_8040, w_075_8044, w_075_8046, w_075_8047, w_075_8051, w_075_8052, w_075_8054, w_075_8065, w_075_8066, w_075_8070, w_075_8074, w_075_8075, w_075_8076, w_075_8078, w_075_8079, w_075_8090, w_075_8092, w_075_8095, w_075_8105, w_075_8108, w_075_8110, w_075_8112, w_075_8115, w_075_8120, w_075_8125, w_075_8133, w_075_8146, w_075_8152, w_075_8153, w_075_8154, w_075_8156, w_075_8157, w_075_8160, w_075_8165, w_075_8166, w_075_8167, w_075_8168, w_075_8174, w_075_8175, w_075_8179, w_075_8182, w_075_8184, w_075_8186, w_075_8187, w_075_8191, w_075_8200, w_075_8204, w_075_8208, w_075_8211, w_075_8213, w_075_8216, w_075_8225, w_075_8232, w_075_8233, w_075_8236, w_075_8238, w_075_8239, w_075_8241, w_075_8242, w_075_8250, w_075_8251, w_075_8252, w_075_8257, w_075_8260, w_075_8264, w_075_8267, w_075_8268, w_075_8280, w_075_8281, w_075_8286, w_075_8288, w_075_8294, w_075_8297, w_075_8298, w_075_8301, w_075_8308, w_075_8309, w_075_8311, w_075_8317, w_075_8319, w_075_8320, w_075_8325, w_075_8328, w_075_8334, w_075_8336, w_075_8338, w_075_8347, w_075_8348, w_075_8349, w_075_8352, w_075_8354, w_075_8357, w_075_8369, w_075_8372, w_075_8376, w_075_8381, w_075_8382, w_075_8383, w_075_8386, w_075_8391, w_075_8393, w_075_8398, w_075_8399, w_075_8400, w_075_8402, w_075_8411, w_075_8412, w_075_8415, w_075_8416, w_075_8425, w_075_8427, w_075_8433, w_075_8438, w_075_8440, w_075_8442, w_075_8444, w_075_8449, w_075_8451, w_075_8457, w_075_8458, w_075_8461, w_075_8467, w_075_8468, w_075_8469, w_075_8470, w_075_8472, w_075_8477, w_075_8480, w_075_8482, w_075_8484, w_075_8485, w_075_8488, w_075_8490, w_075_8491, w_075_8497, w_075_8502, w_075_8507, w_075_8508, w_075_8511, w_075_8514, w_075_8515, w_075_8516, w_075_8519, w_075_8521, w_075_8523, w_075_8526, w_075_8527, w_075_8529, w_075_8530, w_075_8531, w_075_8533, w_075_8536, w_075_8546, w_075_8549, w_075_8550, w_075_8553, w_075_8556, w_075_8558, w_075_8559, w_075_8563, w_075_8570, w_075_8572, w_075_8575, w_075_8576, w_075_8577, w_075_8580, w_075_8585, w_075_8586, w_075_8589, w_075_8591, w_075_8592, w_075_8593, w_075_8594, w_075_8596, w_075_8599, w_075_8601, w_075_8604, w_075_8605, w_075_8606, w_075_8609, w_075_8613, w_075_8614, w_075_8622, w_075_8625, w_075_8626, w_075_8628, w_075_8630, w_075_8631, w_075_8635, w_075_8641, w_075_8646, w_075_8651, w_075_8652, w_075_8653, w_075_8654, w_075_8658, w_075_8659, w_075_8662, w_075_8666, w_075_8668, w_075_8673, w_075_8676, w_075_8678, w_075_8680, w_075_8683, w_075_8687, w_075_8690, w_075_8691, w_075_8694, w_075_8698, w_075_8702, w_075_8706, w_075_8708, w_075_8715, w_075_8717, w_075_8719, w_075_8721, w_075_8722, w_075_8723, w_075_8727, w_075_8735, w_075_8740, w_075_8743, w_075_8744, w_075_8751, w_075_8754, w_075_8755, w_075_8756, w_075_8757, w_075_8758, w_075_8760, w_075_8761, w_075_8763, w_075_8767, w_075_8769, w_075_8770, w_075_8772, w_075_8774, w_075_8781, w_075_8785, w_075_8792, w_075_8793, w_075_8797, w_075_8798, w_075_8801, w_075_8803, w_075_8809, w_075_8810, w_075_8811, w_075_8819, w_075_8820, w_075_8821, w_075_8824, w_075_8826, w_075_8828, w_075_8829, w_075_8832, w_075_8833, w_075_8834, w_075_8837, w_075_8838, w_075_8839, w_075_8841, w_075_8842, w_075_8845, w_075_8847, w_075_8848, w_075_8850, w_075_8851, w_075_8852, w_075_8856, w_075_8858, w_075_8859, w_075_8864, w_075_8872, w_075_8874, w_075_8875, w_075_8877, w_075_8880, w_075_8892, w_075_8896, w_075_8898, w_075_8899, w_075_8900, w_075_8901, w_075_8906, w_075_8912, w_075_8914, w_075_8916, w_075_8917, w_075_8919, w_075_8925, w_075_8926, w_075_8927, w_075_8929, w_075_8930, w_075_8931, w_075_8937, w_075_8938, w_075_8939, w_075_8942, w_075_8950, w_075_8955, w_075_8959, w_075_8964, w_075_8966, w_075_8973, w_075_8975, w_075_8984, w_075_8985, w_075_8988, w_075_8990, w_075_8993, w_075_9007, w_075_9011, w_075_9021, w_075_9022, w_075_9023, w_075_9025, w_075_9026, w_075_9030, w_075_9033, w_075_9036, w_075_9037, w_075_9039, w_075_9040, w_075_9041, w_075_9048, w_075_9052, w_075_9057, w_075_9065, w_075_9071, w_075_9072, w_075_9073, w_075_9075, w_075_9076, w_075_9077, w_075_9079, w_075_9083, w_075_9084, w_075_9088, w_075_9089, w_075_9094, w_075_9097, w_075_9100, w_075_9104, w_075_9109, w_075_9110, w_075_9116, w_075_9118, w_075_9120, w_075_9125, w_075_9128, w_075_9131, w_075_9134, w_075_9135, w_075_9136, w_075_9140, w_075_9145, w_075_9154, w_075_9159, w_075_9168, w_075_9170, w_075_9171, w_075_9181, w_075_9184, w_075_9185, w_075_9189, w_075_9193, w_075_9196, w_075_9198, w_075_9199, w_075_9202, w_075_9205, w_075_9208, w_075_9209, w_075_9210, w_075_9211, w_075_9213, w_075_9214, w_075_9216, w_075_9217, w_075_9222, w_075_9223, w_075_9224, w_075_9225, w_075_9226, w_075_9227, w_075_9228, w_075_9232, w_075_9234, w_075_9237, w_075_9244, w_075_9245, w_075_9246, w_075_9247, w_075_9248, w_075_9252, w_075_9253, w_075_9257, w_075_9258, w_075_9262, w_075_9263, w_075_9265, w_075_9272, w_075_9274, w_075_9275, w_075_9291, w_075_9297, w_075_9300, w_075_9302, w_075_9303, w_075_9308, w_075_9309, w_075_9315, w_075_9319, w_075_9321, w_075_9322, w_075_9323, w_075_9326, w_075_9327, w_075_9328, w_075_9330, w_075_9332, w_075_9334, w_075_9338, w_075_9340, w_075_9342, w_075_9344, w_075_9346, w_075_9352, w_075_9353, w_075_9355, w_075_9357, w_075_9361, w_075_9364, w_075_9365, w_075_9367, w_075_9371, w_075_9374, w_075_9377, w_075_9379, w_075_9381, w_075_9389, w_075_9399, w_075_9405, w_075_9411, w_075_9414, w_075_9421, w_075_9428, w_075_9429, w_075_9433, w_075_9434, w_075_9436, w_075_9437, w_075_9438, w_075_9440, w_075_9441, w_075_9442, w_075_9443, w_075_9444, w_075_9445, w_075_9452, w_075_9456, w_075_9462, w_075_9469, w_075_9470, w_075_9471, w_075_9482, w_075_9486, w_075_9487, w_075_9489, w_075_9493, w_075_9496, w_075_9497, w_075_9498, w_075_9505, w_075_9506, w_075_9507, w_075_9517, w_075_9520, w_075_9522, w_075_9528, w_075_9530, w_075_9539, w_075_9543, w_075_9545, w_075_9552, w_075_9553, w_075_9554, w_075_9556, w_075_9564, w_075_9565, w_075_9567, w_075_9569, w_075_9571, w_075_9579, w_075_9582, w_075_9593, w_075_9595, w_075_9603, w_075_9604, w_075_9606, w_075_9609, w_075_9610, w_075_9611, w_075_9613, w_075_9619, w_075_9622, w_075_9623, w_075_9625, w_075_9631, w_075_9632, w_075_9638, w_075_9640, w_075_9644, w_075_9645, w_075_9646, w_075_9650, w_075_9654, w_075_9656, w_075_9670, w_075_9672, w_075_9678, w_075_9679, w_075_9680, w_075_9690, w_075_9694, w_075_9697, w_075_9699, w_075_9701, w_075_9703, w_075_9704, w_075_9705, w_075_9708, w_075_9709, w_075_9712, w_075_9715, w_075_9716, w_075_9723, w_075_9724, w_075_9725, w_075_9728, w_075_9729, w_075_9732, w_075_9733, w_075_9738, w_075_9744, w_075_9751, w_075_9756, w_075_9759, w_075_9760, w_075_9761, w_075_9762, w_075_9765, w_075_9768, w_075_9771, w_075_9773, w_075_9775, w_075_9776, w_075_9777, w_075_9780, w_075_9782, w_075_9783, w_075_9785, w_075_9788, w_075_9792, w_075_9797;
  wire w_076_000, w_076_001, w_076_004, w_076_005, w_076_006, w_076_008, w_076_009, w_076_010, w_076_011, w_076_012, w_076_013, w_076_014, w_076_016, w_076_017, w_076_018, w_076_022, w_076_023, w_076_024, w_076_025, w_076_026, w_076_027, w_076_030, w_076_033, w_076_035, w_076_036, w_076_038, w_076_041, w_076_043, w_076_044, w_076_045, w_076_046, w_076_047, w_076_049, w_076_050, w_076_052, w_076_056, w_076_060, w_076_061, w_076_067, w_076_070, w_076_071, w_076_073, w_076_074, w_076_076, w_076_077, w_076_083, w_076_084, w_076_086, w_076_088, w_076_089, w_076_092, w_076_093, w_076_094, w_076_095, w_076_097, w_076_098, w_076_101, w_076_102, w_076_104, w_076_105, w_076_106, w_076_107, w_076_108, w_076_111, w_076_112, w_076_113, w_076_114, w_076_115, w_076_116, w_076_118, w_076_119, w_076_120, w_076_123, w_076_124, w_076_125, w_076_126, w_076_137, w_076_138, w_076_143, w_076_144, w_076_146, w_076_147, w_076_149, w_076_150, w_076_154, w_076_156, w_076_157, w_076_160, w_076_162, w_076_163, w_076_166, w_076_167, w_076_177, w_076_178, w_076_180, w_076_181, w_076_184, w_076_186, w_076_188, w_076_189, w_076_192, w_076_194, w_076_195, w_076_198, w_076_201, w_076_205, w_076_210, w_076_212, w_076_216, w_076_218, w_076_220, w_076_228, w_076_231, w_076_236, w_076_243, w_076_245, w_076_246, w_076_247, w_076_250, w_076_255, w_076_256, w_076_258, w_076_262, w_076_265, w_076_267, w_076_268, w_076_270, w_076_273, w_076_276, w_076_277, w_076_278, w_076_279, w_076_283, w_076_287, w_076_289, w_076_295, w_076_297, w_076_298, w_076_300, w_076_301, w_076_302, w_076_303, w_076_304, w_076_306, w_076_309, w_076_311, w_076_312, w_076_317, w_076_323, w_076_324, w_076_327, w_076_328, w_076_330, w_076_331, w_076_332, w_076_333, w_076_335, w_076_336, w_076_341, w_076_343, w_076_344, w_076_348, w_076_349, w_076_352, w_076_353, w_076_354, w_076_357, w_076_358, w_076_360, w_076_362, w_076_363, w_076_366, w_076_370, w_076_371, w_076_372, w_076_376, w_076_377, w_076_382, w_076_383, w_076_384, w_076_386, w_076_388, w_076_390, w_076_401, w_076_403, w_076_404, w_076_406, w_076_408, w_076_409, w_076_410, w_076_411, w_076_413, w_076_414, w_076_417, w_076_418, w_076_419, w_076_420, w_076_423, w_076_429, w_076_430, w_076_433, w_076_434, w_076_436, w_076_437, w_076_439, w_076_442, w_076_445, w_076_448, w_076_452, w_076_453, w_076_455, w_076_456, w_076_462, w_076_463, w_076_466, w_076_470, w_076_472, w_076_474, w_076_476, w_076_481, w_076_483, w_076_484, w_076_485, w_076_486, w_076_488, w_076_489, w_076_490, w_076_494, w_076_495, w_076_497, w_076_499, w_076_500, w_076_501, w_076_502, w_076_503, w_076_506, w_076_508, w_076_512, w_076_513, w_076_514, w_076_516, w_076_517, w_076_524, w_076_529, w_076_530, w_076_531, w_076_532, w_076_533, w_076_534, w_076_538, w_076_539, w_076_540, w_076_543, w_076_544, w_076_548, w_076_550, w_076_553, w_076_555, w_076_557, w_076_563, w_076_564, w_076_565, w_076_566, w_076_567, w_076_568, w_076_570, w_076_571, w_076_572, w_076_573, w_076_576, w_076_583, w_076_586, w_076_587, w_076_588, w_076_590, w_076_593, w_076_594, w_076_597, w_076_598, w_076_603, w_076_605, w_076_608, w_076_609, w_076_615, w_076_617, w_076_619, w_076_622, w_076_623, w_076_625, w_076_626, w_076_628, w_076_629, w_076_631, w_076_634, w_076_636, w_076_637, w_076_638, w_076_639, w_076_642, w_076_643, w_076_644, w_076_645, w_076_646, w_076_653, w_076_655, w_076_656, w_076_657, w_076_658, w_076_659, w_076_662, w_076_664, w_076_665, w_076_667, w_076_668, w_076_670, w_076_671, w_076_673, w_076_674, w_076_675, w_076_684, w_076_685, w_076_688, w_076_689, w_076_690, w_076_691, w_076_692, w_076_694, w_076_695, w_076_697, w_076_699, w_076_702, w_076_705, w_076_706, w_076_707, w_076_708, w_076_709, w_076_710, w_076_713, w_076_714, w_076_715, w_076_719, w_076_720, w_076_725, w_076_727, w_076_729, w_076_730, w_076_731, w_076_732, w_076_735, w_076_736, w_076_737, w_076_739, w_076_741, w_076_749, w_076_751, w_076_754, w_076_755, w_076_756, w_076_758, w_076_759, w_076_763, w_076_764, w_076_766, w_076_767, w_076_768, w_076_769, w_076_771, w_076_772, w_076_775, w_076_777, w_076_778, w_076_782, w_076_783, w_076_784, w_076_787, w_076_788, w_076_790, w_076_791, w_076_792, w_076_793, w_076_794, w_076_795, w_076_796, w_076_798, w_076_799, w_076_800, w_076_802, w_076_804, w_076_805, w_076_813, w_076_815, w_076_817, w_076_819, w_076_820, w_076_821, w_076_823, w_076_825, w_076_826, w_076_827, w_076_828, w_076_829, w_076_834, w_076_835, w_076_840, w_076_847, w_076_848, w_076_849, w_076_850, w_076_853, w_076_855, w_076_856, w_076_858, w_076_861, w_076_862, w_076_869, w_076_872, w_076_873, w_076_874, w_076_876, w_076_878, w_076_881, w_076_883, w_076_885, w_076_887, w_076_891, w_076_892, w_076_894, w_076_895, w_076_896, w_076_897, w_076_900, w_076_904, w_076_906, w_076_907, w_076_911, w_076_912, w_076_913, w_076_914, w_076_917, w_076_918, w_076_919, w_076_920, w_076_921, w_076_924, w_076_925, w_076_926, w_076_933, w_076_934, w_076_937, w_076_938, w_076_939, w_076_940, w_076_942, w_076_943, w_076_945, w_076_952, w_076_953, w_076_954, w_076_956, w_076_959, w_076_961, w_076_962, w_076_963, w_076_966, w_076_970, w_076_972, w_076_973, w_076_975, w_076_977, w_076_979, w_076_980, w_076_982, w_076_983, w_076_984, w_076_989, w_076_990, w_076_992, w_076_995, w_076_996, w_076_998, w_076_1000, w_076_1001, w_076_1002, w_076_1004, w_076_1007, w_076_1008, w_076_1013, w_076_1019, w_076_1022, w_076_1023, w_076_1024, w_076_1025, w_076_1027, w_076_1032, w_076_1034, w_076_1036, w_076_1038, w_076_1039, w_076_1041, w_076_1042, w_076_1043, w_076_1047, w_076_1048, w_076_1051, w_076_1053, w_076_1054, w_076_1056, w_076_1057, w_076_1058, w_076_1060, w_076_1061, w_076_1063, w_076_1064, w_076_1067, w_076_1071, w_076_1072, w_076_1073, w_076_1074, w_076_1075, w_076_1077, w_076_1078, w_076_1079, w_076_1081, w_076_1083, w_076_1085, w_076_1086, w_076_1087, w_076_1094, w_076_1096, w_076_1098, w_076_1099, w_076_1101, w_076_1103, w_076_1104, w_076_1105, w_076_1106, w_076_1107, w_076_1108, w_076_1109, w_076_1116, w_076_1117, w_076_1118, w_076_1123, w_076_1124, w_076_1125, w_076_1127, w_076_1129, w_076_1132, w_076_1134, w_076_1135, w_076_1136, w_076_1141, w_076_1144, w_076_1145, w_076_1146, w_076_1147, w_076_1154, w_076_1155, w_076_1158, w_076_1161, w_076_1162, w_076_1163, w_076_1164, w_076_1165, w_076_1167, w_076_1168, w_076_1169, w_076_1177, w_076_1181, w_076_1184, w_076_1187, w_076_1189, w_076_1190, w_076_1192, w_076_1193, w_076_1194, w_076_1196, w_076_1197, w_076_1198, w_076_1199, w_076_1202, w_076_1204, w_076_1208, w_076_1209, w_076_1213, w_076_1214, w_076_1215, w_076_1216, w_076_1220, w_076_1221, w_076_1227, w_076_1228, w_076_1229, w_076_1230, w_076_1233, w_076_1234, w_076_1237, w_076_1240, w_076_1242, w_076_1244, w_076_1247, w_076_1250, w_076_1253, w_076_1255, w_076_1256, w_076_1257, w_076_1259, w_076_1260, w_076_1261, w_076_1263, w_076_1264, w_076_1268, w_076_1273, w_076_1275, w_076_1280, w_076_1281, w_076_1283, w_076_1286, w_076_1288, w_076_1290, w_076_1292, w_076_1293, w_076_1294, w_076_1295, w_076_1298, w_076_1299, w_076_1300, w_076_1301, w_076_1305, w_076_1306, w_076_1307, w_076_1308, w_076_1309, w_076_1310, w_076_1312, w_076_1313, w_076_1316, w_076_1317, w_076_1318, w_076_1320, w_076_1321, w_076_1322, w_076_1324, w_076_1325, w_076_1326, w_076_1327, w_076_1328, w_076_1335, w_076_1337, w_076_1338, w_076_1343, w_076_1345, w_076_1347, w_076_1349, w_076_1350, w_076_1354, w_076_1355, w_076_1358, w_076_1359, w_076_1360, w_076_1361, w_076_1362, w_076_1363, w_076_1366, w_076_1367, w_076_1370, w_076_1372, w_076_1373, w_076_1374, w_076_1376, w_076_1377, w_076_1379, w_076_1381, w_076_1382, w_076_1386, w_076_1388, w_076_1391, w_076_1393, w_076_1397, w_076_1398, w_076_1401, w_076_1405, w_076_1408, w_076_1409, w_076_1411, w_076_1413, w_076_1415, w_076_1416, w_076_1418, w_076_1423, w_076_1424, w_076_1425, w_076_1426, w_076_1427, w_076_1430, w_076_1433, w_076_1440, w_076_1443, w_076_1444, w_076_1446, w_076_1448, w_076_1449, w_076_1450, w_076_1455, w_076_1458, w_076_1459, w_076_1461, w_076_1462, w_076_1463, w_076_1465, w_076_1466, w_076_1468, w_076_1469, w_076_1470, w_076_1475, w_076_1479, w_076_1480, w_076_1481, w_076_1485, w_076_1488, w_076_1489, w_076_1491, w_076_1493, w_076_1494, w_076_1497, w_076_1499, w_076_1500, w_076_1502, w_076_1505, w_076_1506, w_076_1508, w_076_1509, w_076_1514, w_076_1515, w_076_1516, w_076_1517, w_076_1519, w_076_1525, w_076_1527, w_076_1528, w_076_1532, w_076_1534, w_076_1535, w_076_1537, w_076_1538, w_076_1540, w_076_1542, w_076_1543, w_076_1547, w_076_1549, w_076_1551, w_076_1554, w_076_1555, w_076_1556, w_076_1557, w_076_1560, w_076_1562, w_076_1563, w_076_1566, w_076_1569, w_076_1575, w_076_1577, w_076_1578, w_076_1581, w_076_1583, w_076_1585, w_076_1586, w_076_1587, w_076_1588, w_076_1589, w_076_1590, w_076_1592, w_076_1593, w_076_1595, w_076_1596, w_076_1598, w_076_1599, w_076_1600, w_076_1601, w_076_1605, w_076_1610, w_076_1612, w_076_1614, w_076_1615, w_076_1619, w_076_1621, w_076_1622, w_076_1623, w_076_1624, w_076_1625, w_076_1627, w_076_1632, w_076_1634, w_076_1639, w_076_1647, w_076_1648, w_076_1650, w_076_1651, w_076_1652, w_076_1654, w_076_1655, w_076_1657, w_076_1658, w_076_1661, w_076_1663, w_076_1664, w_076_1666, w_076_1667, w_076_1669, w_076_1672, w_076_1673, w_076_1675, w_076_1678, w_076_1686, w_076_1687, w_076_1688, w_076_1690, w_076_1693, w_076_1694, w_076_1697, w_076_1698, w_076_1699, w_076_1700, w_076_1701, w_076_1702, w_076_1705, w_076_1706, w_076_1710, w_076_1712, w_076_1713, w_076_1714, w_076_1718, w_076_1721, w_076_1725, w_076_1729, w_076_1736, w_076_1738, w_076_1739, w_076_1740, w_076_1748, w_076_1749, w_076_1752, w_076_1754, w_076_1756, w_076_1757, w_076_1760, w_076_1761, w_076_1762, w_076_1763, w_076_1764, w_076_1768, w_076_1769, w_076_1770, w_076_1773, w_076_1776, w_076_1778, w_076_1780, w_076_1781, w_076_1784, w_076_1786, w_076_1788, w_076_1789, w_076_1791, w_076_1794, w_076_1796, w_076_1798, w_076_1799, w_076_1800, w_076_1801, w_076_1804, w_076_1806, w_076_1808, w_076_1809, w_076_1811, w_076_1817, w_076_1818, w_076_1820, w_076_1821, w_076_1822, w_076_1824, w_076_1825, w_076_1827, w_076_1828, w_076_1833, w_076_1834, w_076_1835, w_076_1839, w_076_1840, w_076_1843, w_076_1846, w_076_1847, w_076_1856, w_076_1860, w_076_1862, w_076_1865, w_076_1874, w_076_1877, w_076_1880, w_076_1885, w_076_1886, w_076_1888, w_076_1889, w_076_1891, w_076_1892, w_076_1893, w_076_1894, w_076_1895, w_076_1898, w_076_1902, w_076_1903, w_076_1905, w_076_1906, w_076_1907, w_076_1908, w_076_1909, w_076_1912, w_076_1913, w_076_1914, w_076_1917, w_076_1918, w_076_1919, w_076_1920, w_076_1922, w_076_1925, w_076_1926, w_076_1927, w_076_1930, w_076_1931, w_076_1932, w_076_1933, w_076_1934, w_076_1935, w_076_1942, w_076_1943, w_076_1944, w_076_1946, w_076_1947, w_076_1952, w_076_1953, w_076_1954, w_076_1955, w_076_1958, w_076_1960, w_076_1963, w_076_1966, w_076_1973, w_076_1974, w_076_1975, w_076_1976, w_076_1977, w_076_1978, w_076_1979, w_076_1982, w_076_1983, w_076_1984, w_076_1987, w_076_1989, w_076_1996, w_076_1997, w_076_1999, w_076_2000, w_076_2002, w_076_2003, w_076_2004, w_076_2006, w_076_2007, w_076_2008, w_076_2009, w_076_2010, w_076_2011, w_076_2013, w_076_2014, w_076_2017, w_076_2021, w_076_2025, w_076_2026, w_076_2027, w_076_2028, w_076_2030, w_076_2032, w_076_2036, w_076_2040, w_076_2041, w_076_2046, w_076_2049, w_076_2052, w_076_2056, w_076_2057, w_076_2058, w_076_2060, w_076_2061, w_076_2062, w_076_2063, w_076_2064, w_076_2067, w_076_2072, w_076_2073, w_076_2076, w_076_2077, w_076_2078, w_076_2082, w_076_2086, w_076_2089, w_076_2090, w_076_2091, w_076_2092, w_076_2094, w_076_2095, w_076_2096, w_076_2097, w_076_2099, w_076_2100, w_076_2101, w_076_2102, w_076_2103, w_076_2109, w_076_2110, w_076_2114, w_076_2115, w_076_2116, w_076_2121, w_076_2124, w_076_2127, w_076_2131, w_076_2133, w_076_2134, w_076_2137, w_076_2138, w_076_2141, w_076_2142, w_076_2144, w_076_2145, w_076_2146, w_076_2149, w_076_2150, w_076_2151, w_076_2152, w_076_2153, w_076_2154, w_076_2157, w_076_2160, w_076_2162, w_076_2163, w_076_2164, w_076_2165, w_076_2166, w_076_2170, w_076_2172, w_076_2173, w_076_2174, w_076_2175, w_076_2176, w_076_2179, w_076_2181, w_076_2182, w_076_2183, w_076_2184, w_076_2185, w_076_2186, w_076_2187, w_076_2188, w_076_2189, w_076_2190, w_076_2191, w_076_2195, w_076_2196, w_076_2203, w_076_2204, w_076_2207, w_076_2208, w_076_2210, w_076_2211, w_076_2213, w_076_2214, w_076_2216, w_076_2219, w_076_2221, w_076_2228, w_076_2229, w_076_2231, w_076_2235, w_076_2238, w_076_2241, w_076_2242, w_076_2245, w_076_2246, w_076_2248, w_076_2250, w_076_2251, w_076_2252, w_076_2254, w_076_2255, w_076_2257, w_076_2258, w_076_2259, w_076_2263, w_076_2265, w_076_2266, w_076_2269, w_076_2273, w_076_2275, w_076_2278, w_076_2280, w_076_2281, w_076_2282, w_076_2285, w_076_2286, w_076_2287, w_076_2289, w_076_2293, w_076_2294, w_076_2298, w_076_2299, w_076_2300, w_076_2302, w_076_2304, w_076_2305, w_076_2307, w_076_2308, w_076_2310, w_076_2311, w_076_2315, w_076_2316, w_076_2317, w_076_2318, w_076_2320, w_076_2321, w_076_2323, w_076_2324, w_076_2325, w_076_2329, w_076_2330, w_076_2334, w_076_2339, w_076_2340, w_076_2341, w_076_2348, w_076_2349, w_076_2350, w_076_2351, w_076_2352, w_076_2353, w_076_2355, w_076_2356, w_076_2357, w_076_2359, w_076_2361, w_076_2362, w_076_2367, w_076_2368, w_076_2369, w_076_2372, w_076_2375, w_076_2376, w_076_2377, w_076_2382, w_076_2384, w_076_2385, w_076_2391, w_076_2392, w_076_2395, w_076_2396, w_076_2398, w_076_2405, w_076_2407, w_076_2408, w_076_2409, w_076_2410, w_076_2412, w_076_2413, w_076_2414, w_076_2415, w_076_2416, w_076_2417, w_076_2419, w_076_2420, w_076_2421, w_076_2422, w_076_2423, w_076_2425, w_076_2434, w_076_2435, w_076_2438, w_076_2440, w_076_2441, w_076_2443, w_076_2444, w_076_2446, w_076_2447, w_076_2448, w_076_2449, w_076_2450, w_076_2451, w_076_2453, w_076_2455, w_076_2456, w_076_2458, w_076_2460, w_076_2464, w_076_2465, w_076_2466, w_076_2467, w_076_2468, w_076_2469, w_076_2470, w_076_2474, w_076_2475, w_076_2476, w_076_2479, w_076_2483, w_076_2488, w_076_2489, w_076_2491, w_076_2495, w_076_2496, w_076_2497, w_076_2498, w_076_2499, w_076_2500, w_076_2501, w_076_2502, w_076_2503, w_076_2504, w_076_2505, w_076_2506, w_076_2507, w_076_2510, w_076_2511, w_076_2513, w_076_2514, w_076_2515, w_076_2520, w_076_2521, w_076_2523, w_076_2524, w_076_2525, w_076_2526, w_076_2528, w_076_2529, w_076_2530, w_076_2531, w_076_2534, w_076_2535, w_076_2537, w_076_2538, w_076_2543, w_076_2545, w_076_2546, w_076_2549, w_076_2550, w_076_2553, w_076_2555, w_076_2557, w_076_2558, w_076_2559, w_076_2560, w_076_2563, w_076_2564, w_076_2565, w_076_2568, w_076_2570, w_076_2571, w_076_2581, w_076_2582, w_076_2583, w_076_2587, w_076_2588, w_076_2589, w_076_2594, w_076_2595, w_076_2596, w_076_2598, w_076_2603, w_076_2604, w_076_2607, w_076_2608, w_076_2609, w_076_2610, w_076_2611, w_076_2614, w_076_2615, w_076_2618, w_076_2621, w_076_2624, w_076_2626, w_076_2627, w_076_2628, w_076_2631, w_076_2637, w_076_2642, w_076_2643, w_076_2646, w_076_2647, w_076_2660, w_076_2661, w_076_2662, w_076_2664, w_076_2666, w_076_2667, w_076_2668, w_076_2669, w_076_2670, w_076_2671, w_076_2672, w_076_2673, w_076_2674, w_076_2676, w_076_2677, w_076_2680, w_076_2683, w_076_2684, w_076_2686, w_076_2689, w_076_2691, w_076_2692, w_076_2693, w_076_2694, w_076_2695, w_076_2697, w_076_2698, w_076_2700, w_076_2703, w_076_2704, w_076_2706, w_076_2707, w_076_2710, w_076_2711, w_076_2716, w_076_2717, w_076_2719, w_076_2722, w_076_2725, w_076_2727, w_076_2728, w_076_2729, w_076_2731, w_076_2733, w_076_2734, w_076_2737, w_076_2740, w_076_2743, w_076_2747, w_076_2748, w_076_2749, w_076_2752, w_076_2753, w_076_2754, w_076_2762, w_076_2763, w_076_2765, w_076_2773, w_076_2779, w_076_2782, w_076_2783, w_076_2784, w_076_2786, w_076_2792, w_076_2795, w_076_2796, w_076_2799, w_076_2801, w_076_2806, w_076_2809, w_076_2811, w_076_2819, w_076_2824, w_076_2827, w_076_2830, w_076_2843, w_076_2844, w_076_2848, w_076_2850, w_076_2851, w_076_2852, w_076_2854, w_076_2859, w_076_2860, w_076_2863, w_076_2864, w_076_2869, w_076_2872, w_076_2874, w_076_2875, w_076_2877, w_076_2878, w_076_2879, w_076_2883, w_076_2889, w_076_2891, w_076_2895, w_076_2901, w_076_2906, w_076_2910, w_076_2912, w_076_2913, w_076_2915, w_076_2916, w_076_2918, w_076_2920, w_076_2921, w_076_2925, w_076_2931, w_076_2934, w_076_2937, w_076_2939, w_076_2940, w_076_2942, w_076_2944, w_076_2954, w_076_2955, w_076_2956, w_076_2958, w_076_2959, w_076_2962, w_076_2969, w_076_2971, w_076_2976, w_076_2978, w_076_2980, w_076_2986, w_076_2994, w_076_2998, w_076_3002, w_076_3004, w_076_3005, w_076_3008, w_076_3009, w_076_3010, w_076_3020, w_076_3021, w_076_3022, w_076_3027, w_076_3028, w_076_3032, w_076_3033, w_076_3034, w_076_3035, w_076_3041, w_076_3042, w_076_3044, w_076_3045, w_076_3050, w_076_3052, w_076_3062, w_076_3063, w_076_3065, w_076_3066, w_076_3070, w_076_3071, w_076_3081, w_076_3084, w_076_3087, w_076_3088, w_076_3089, w_076_3102, w_076_3109, w_076_3110, w_076_3111, w_076_3112, w_076_3116, w_076_3120, w_076_3121, w_076_3125, w_076_3133, w_076_3141, w_076_3142, w_076_3146, w_076_3147, w_076_3149, w_076_3150, w_076_3152, w_076_3154, w_076_3157, w_076_3161, w_076_3164, w_076_3180, w_076_3182, w_076_3184, w_076_3188, w_076_3192, w_076_3194, w_076_3195, w_076_3197, w_076_3200, w_076_3201, w_076_3203, w_076_3210, w_076_3211, w_076_3213, w_076_3218, w_076_3222, w_076_3225, w_076_3226, w_076_3227, w_076_3229, w_076_3230, w_076_3235, w_076_3240, w_076_3243, w_076_3244, w_076_3251, w_076_3253, w_076_3257, w_076_3259, w_076_3260, w_076_3263, w_076_3265, w_076_3267, w_076_3268, w_076_3279, w_076_3281, w_076_3288, w_076_3294, w_076_3299, w_076_3300, w_076_3310, w_076_3315, w_076_3324, w_076_3327, w_076_3329, w_076_3331, w_076_3333, w_076_3335, w_076_3336, w_076_3337, w_076_3338, w_076_3343, w_076_3346, w_076_3347, w_076_3349, w_076_3356, w_076_3361, w_076_3363, w_076_3366, w_076_3369, w_076_3384, w_076_3388, w_076_3391, w_076_3392, w_076_3393, w_076_3395, w_076_3398, w_076_3400, w_076_3401, w_076_3402, w_076_3409, w_076_3411, w_076_3416, w_076_3418, w_076_3420, w_076_3421, w_076_3423, w_076_3425, w_076_3428, w_076_3431, w_076_3434, w_076_3436, w_076_3439, w_076_3446, w_076_3455, w_076_3465, w_076_3468, w_076_3475, w_076_3477, w_076_3486, w_076_3487, w_076_3489, w_076_3496, w_076_3499, w_076_3503, w_076_3505, w_076_3510, w_076_3513, w_076_3514, w_076_3517, w_076_3523, w_076_3524, w_076_3527, w_076_3528, w_076_3530, w_076_3541, w_076_3543, w_076_3544, w_076_3547, w_076_3548, w_076_3550, w_076_3552, w_076_3556, w_076_3557, w_076_3558, w_076_3562, w_076_3565, w_076_3575, w_076_3577, w_076_3578, w_076_3580, w_076_3581, w_076_3582, w_076_3590, w_076_3592, w_076_3594, w_076_3597, w_076_3605, w_076_3607, w_076_3610, w_076_3614, w_076_3617, w_076_3620, w_076_3625, w_076_3629, w_076_3632, w_076_3636, w_076_3639, w_076_3640, w_076_3641, w_076_3644, w_076_3653, w_076_3655, w_076_3657, w_076_3658, w_076_3660, w_076_3664, w_076_3676, w_076_3681, w_076_3684, w_076_3685, w_076_3686, w_076_3688, w_076_3698, w_076_3700, w_076_3701, w_076_3702, w_076_3703, w_076_3705, w_076_3711, w_076_3720, w_076_3722, w_076_3727, w_076_3730, w_076_3735, w_076_3737, w_076_3740, w_076_3741, w_076_3742, w_076_3743, w_076_3745, w_076_3746, w_076_3747, w_076_3748, w_076_3751, w_076_3755, w_076_3763, w_076_3771, w_076_3774, w_076_3776, w_076_3782, w_076_3784, w_076_3786, w_076_3790, w_076_3791, w_076_3796, w_076_3799, w_076_3800, w_076_3801, w_076_3802, w_076_3804, w_076_3805, w_076_3806, w_076_3809, w_076_3818, w_076_3822, w_076_3826, w_076_3834, w_076_3836, w_076_3840, w_076_3841, w_076_3843, w_076_3844, w_076_3849, w_076_3850, w_076_3852, w_076_3862, w_076_3864, w_076_3865, w_076_3866, w_076_3875, w_076_3884, w_076_3886, w_076_3889, w_076_3890, w_076_3892, w_076_3895, w_076_3899, w_076_3900, w_076_3904, w_076_3912, w_076_3914, w_076_3918, w_076_3920, w_076_3921, w_076_3924, w_076_3925, w_076_3934, w_076_3936, w_076_3939, w_076_3941, w_076_3945, w_076_3948, w_076_3950, w_076_3951, w_076_3958, w_076_3959, w_076_3961, w_076_3964, w_076_3968, w_076_3971, w_076_3974, w_076_3975, w_076_3984, w_076_3985, w_076_3992, w_076_3995, w_076_3997, w_076_3998, w_076_4002, w_076_4004, w_076_4007, w_076_4010, w_076_4012, w_076_4032, w_076_4034, w_076_4035, w_076_4041, w_076_4044, w_076_4051, w_076_4063, w_076_4077, w_076_4079, w_076_4083, w_076_4086, w_076_4088, w_076_4089, w_076_4093, w_076_4095, w_076_4099, w_076_4104, w_076_4114, w_076_4118, w_076_4121, w_076_4122, w_076_4127, w_076_4128, w_076_4129, w_076_4130, w_076_4133, w_076_4134, w_076_4140, w_076_4141, w_076_4145, w_076_4151, w_076_4152, w_076_4154, w_076_4157, w_076_4159, w_076_4161, w_076_4164, w_076_4172, w_076_4173, w_076_4177, w_076_4180, w_076_4182, w_076_4190, w_076_4193, w_076_4196, w_076_4200, w_076_4209, w_076_4212, w_076_4213, w_076_4214, w_076_4216, w_076_4218, w_076_4221, w_076_4232, w_076_4234, w_076_4243, w_076_4247, w_076_4249, w_076_4251, w_076_4254, w_076_4262, w_076_4263, w_076_4264, w_076_4265, w_076_4268, w_076_4271, w_076_4275, w_076_4277, w_076_4282, w_076_4283, w_076_4285, w_076_4286, w_076_4287, w_076_4290, w_076_4292, w_076_4294, w_076_4298, w_076_4300, w_076_4301, w_076_4303, w_076_4304, w_076_4305, w_076_4310, w_076_4316, w_076_4322, w_076_4323, w_076_4325, w_076_4326, w_076_4327, w_076_4336, w_076_4337, w_076_4339, w_076_4342, w_076_4357, w_076_4362, w_076_4363, w_076_4367, w_076_4368, w_076_4369, w_076_4373, w_076_4377, w_076_4379, w_076_4380, w_076_4387, w_076_4389, w_076_4394, w_076_4400, w_076_4402, w_076_4407, w_076_4409, w_076_4412, w_076_4413, w_076_4416, w_076_4418, w_076_4421, w_076_4422, w_076_4425, w_076_4433, w_076_4434, w_076_4435, w_076_4446, w_076_4454, w_076_4461, w_076_4466, w_076_4469, w_076_4470, w_076_4471, w_076_4473, w_076_4475, w_076_4478, w_076_4484, w_076_4486, w_076_4488, w_076_4496, w_076_4500, w_076_4510, w_076_4514, w_076_4515, w_076_4518, w_076_4523, w_076_4524, w_076_4525, w_076_4530, w_076_4535, w_076_4539, w_076_4545, w_076_4546, w_076_4547, w_076_4549, w_076_4557, w_076_4559, w_076_4562, w_076_4563, w_076_4565, w_076_4575, w_076_4580, w_076_4585, w_076_4586, w_076_4590, w_076_4592, w_076_4600, w_076_4616, w_076_4618, w_076_4619, w_076_4623, w_076_4628, w_076_4633, w_076_4636, w_076_4639, w_076_4646, w_076_4651, w_076_4652, w_076_4653, w_076_4661, w_076_4664, w_076_4667, w_076_4668, w_076_4670, w_076_4673, w_076_4678, w_076_4685, w_076_4696, w_076_4701, w_076_4705, w_076_4709, w_076_4713, w_076_4715, w_076_4716, w_076_4720, w_076_4722, w_076_4726, w_076_4727, w_076_4731, w_076_4733, w_076_4734, w_076_4737, w_076_4749, w_076_4751, w_076_4752, w_076_4754, w_076_4755, w_076_4762, w_076_4769, w_076_4773, w_076_4774, w_076_4780, w_076_4791, w_076_4797, w_076_4799, w_076_4800, w_076_4805, w_076_4807, w_076_4811, w_076_4812, w_076_4813, w_076_4817, w_076_4819, w_076_4821, w_076_4822, w_076_4823, w_076_4827, w_076_4832, w_076_4835, w_076_4837, w_076_4838, w_076_4839, w_076_4842, w_076_4846, w_076_4851, w_076_4854, w_076_4855, w_076_4858, w_076_4860, w_076_4861, w_076_4862, w_076_4863, w_076_4864, w_076_4866, w_076_4867, w_076_4868, w_076_4870, w_076_4871, w_076_4873, w_076_4877, w_076_4879, w_076_4880, w_076_4892, w_076_4899, w_076_4902, w_076_4903, w_076_4912, w_076_4917, w_076_4921, w_076_4924, w_076_4927, w_076_4928, w_076_4931, w_076_4935, w_076_4936, w_076_4941, w_076_4945, w_076_4947, w_076_4949, w_076_4952, w_076_4953, w_076_4954, w_076_4959, w_076_4965, w_076_4966, w_076_4968, w_076_4970, w_076_4971, w_076_4975, w_076_4977, w_076_4979, w_076_4980, w_076_4985, w_076_4988, w_076_4989, w_076_4990, w_076_4992, w_076_5000, w_076_5005, w_076_5007, w_076_5009, w_076_5014, w_076_5015, w_076_5018, w_076_5025, w_076_5030, w_076_5036, w_076_5038, w_076_5047, w_076_5049, w_076_5055, w_076_5056, w_076_5061, w_076_5062, w_076_5063, w_076_5067, w_076_5068, w_076_5069, w_076_5071, w_076_5072, w_076_5077, w_076_5078, w_076_5082, w_076_5083, w_076_5086, w_076_5091, w_076_5092, w_076_5096, w_076_5097, w_076_5101, w_076_5105, w_076_5109, w_076_5111, w_076_5114, w_076_5115, w_076_5120, w_076_5123, w_076_5126, w_076_5128, w_076_5143, w_076_5147, w_076_5148, w_076_5150, w_076_5151, w_076_5162, w_076_5165, w_076_5169, w_076_5174, w_076_5176, w_076_5178, w_076_5181, w_076_5193, w_076_5194, w_076_5195, w_076_5201, w_076_5208, w_076_5211, w_076_5212, w_076_5219, w_076_5221, w_076_5228, w_076_5229, w_076_5239, w_076_5242, w_076_5244, w_076_5259, w_076_5275, w_076_5279, w_076_5281, w_076_5283, w_076_5289, w_076_5291, w_076_5293, w_076_5301, w_076_5303, w_076_5304, w_076_5305, w_076_5312, w_076_5314, w_076_5316, w_076_5320, w_076_5322, w_076_5328, w_076_5330, w_076_5335, w_076_5344, w_076_5356, w_076_5357, w_076_5361, w_076_5362, w_076_5365, w_076_5366, w_076_5369, w_076_5377, w_076_5378, w_076_5380, w_076_5384, w_076_5386, w_076_5389, w_076_5390, w_076_5392, w_076_5398, w_076_5401, w_076_5405, w_076_5406, w_076_5410, w_076_5413, w_076_5415, w_076_5419, w_076_5421, w_076_5426, w_076_5428, w_076_5433, w_076_5439, w_076_5442, w_076_5445, w_076_5447, w_076_5448, w_076_5450, w_076_5456, w_076_5460, w_076_5461, w_076_5467, w_076_5469, w_076_5470, w_076_5481, w_076_5482, w_076_5487, w_076_5489, w_076_5494, w_076_5502, w_076_5503, w_076_5508, w_076_5509, w_076_5511, w_076_5512, w_076_5516, w_076_5517, w_076_5520, w_076_5527, w_076_5532, w_076_5533, w_076_5535, w_076_5537, w_076_5541, w_076_5552, w_076_5556, w_076_5559, w_076_5561, w_076_5564, w_076_5566, w_076_5569, w_076_5576, w_076_5580, w_076_5590, w_076_5594, w_076_5595, w_076_5597, w_076_5601, w_076_5602, w_076_5604, w_076_5609, w_076_5611, w_076_5614, w_076_5623, w_076_5626, w_076_5627, w_076_5631, w_076_5633, w_076_5638, w_076_5639, w_076_5640, w_076_5641, w_076_5642, w_076_5643, w_076_5644, w_076_5647, w_076_5648, w_076_5650, w_076_5657, w_076_5659, w_076_5660, w_076_5669, w_076_5674, w_076_5675, w_076_5676, w_076_5677, w_076_5678, w_076_5680, w_076_5684, w_076_5688, w_076_5689, w_076_5692, w_076_5693, w_076_5694, w_076_5695, w_076_5697, w_076_5698, w_076_5701, w_076_5705, w_076_5712, w_076_5721, w_076_5723, w_076_5726, w_076_5729, w_076_5731, w_076_5735, w_076_5737, w_076_5738, w_076_5741, w_076_5748, w_076_5749, w_076_5760, w_076_5761, w_076_5762, w_076_5768, w_076_5784, w_076_5791, w_076_5792, w_076_5793, w_076_5796, w_076_5798, w_076_5802, w_076_5805, w_076_5806, w_076_5809, w_076_5811, w_076_5815, w_076_5819, w_076_5827, w_076_5832, w_076_5833, w_076_5837, w_076_5848, w_076_5853, w_076_5854, w_076_5856, w_076_5860, w_076_5862, w_076_5864, w_076_5873, w_076_5885, w_076_5886, w_076_5887, w_076_5891, w_076_5896, w_076_5897, w_076_5899, w_076_5905, w_076_5911, w_076_5916, w_076_5928, w_076_5930, w_076_5933, w_076_5934, w_076_5935, w_076_5941, w_076_5942, w_076_5959, w_076_5961, w_076_5964, w_076_5968, w_076_5970, w_076_5975, w_076_5982, w_076_5984, w_076_5985, w_076_5986, w_076_5987, w_076_5992, w_076_5993, w_076_5994, w_076_5997, w_076_5998, w_076_6006, w_076_6007, w_076_6008, w_076_6011, w_076_6014, w_076_6015, w_076_6023, w_076_6024, w_076_6032, w_076_6040, w_076_6041, w_076_6042, w_076_6044, w_076_6046, w_076_6048, w_076_6057, w_076_6059, w_076_6062, w_076_6064, w_076_6065, w_076_6068, w_076_6073, w_076_6075, w_076_6078, w_076_6079, w_076_6082, w_076_6083, w_076_6088, w_076_6090, w_076_6091, w_076_6092, w_076_6095, w_076_6097, w_076_6099, w_076_6103, w_076_6105, w_076_6108, w_076_6111, w_076_6115, w_076_6118, w_076_6122, w_076_6129, w_076_6138, w_076_6139, w_076_6142, w_076_6147, w_076_6149, w_076_6153, w_076_6158, w_076_6159, w_076_6162, w_076_6167, w_076_6168, w_076_6172, w_076_6173, w_076_6175, w_076_6177, w_076_6179, w_076_6183, w_076_6186, w_076_6187, w_076_6193, w_076_6200, w_076_6205, w_076_6221, w_076_6224, w_076_6233, w_076_6235, w_076_6236, w_076_6237, w_076_6240, w_076_6256, w_076_6261, w_076_6264, w_076_6270, w_076_6283, w_076_6284, w_076_6286, w_076_6290, w_076_6292, w_076_6297, w_076_6301, w_076_6305, w_076_6308, w_076_6309, w_076_6310, w_076_6329, w_076_6331, w_076_6340, w_076_6342, w_076_6343, w_076_6344, w_076_6345, w_076_6349, w_076_6350, w_076_6351, w_076_6352, w_076_6354, w_076_6358, w_076_6364, w_076_6367, w_076_6370, w_076_6372, w_076_6377, w_076_6380, w_076_6382, w_076_6386, w_076_6387, w_076_6388, w_076_6391, w_076_6393, w_076_6406, w_076_6408, w_076_6409, w_076_6410, w_076_6411, w_076_6412, w_076_6414, w_076_6421, w_076_6422, w_076_6423, w_076_6425, w_076_6426, w_076_6433, w_076_6439, w_076_6442, w_076_6443, w_076_6446, w_076_6447, w_076_6449, w_076_6450, w_076_6459, w_076_6460, w_076_6465, w_076_6466, w_076_6468, w_076_6469, w_076_6475, w_076_6477, w_076_6479, w_076_6484, w_076_6485, w_076_6490, w_076_6491, w_076_6493, w_076_6494, w_076_6496, w_076_6497, w_076_6503, w_076_6511, w_076_6512, w_076_6513, w_076_6517, w_076_6518, w_076_6519, w_076_6522, w_076_6532, w_076_6533, w_076_6540, w_076_6542, w_076_6544, w_076_6548, w_076_6552, w_076_6554, w_076_6556, w_076_6557, w_076_6562, w_076_6564, w_076_6576, w_076_6577, w_076_6588, w_076_6590, w_076_6600, w_076_6608, w_076_6610, w_076_6614, w_076_6618, w_076_6619, w_076_6620, w_076_6622, w_076_6624, w_076_6625, w_076_6628, w_076_6630, w_076_6634, w_076_6637, w_076_6640, w_076_6642, w_076_6646, w_076_6648, w_076_6655, w_076_6663, w_076_6666, w_076_6668, w_076_6670, w_076_6672, w_076_6673, w_076_6675, w_076_6676, w_076_6677, w_076_6678, w_076_6682, w_076_6684, w_076_6686, w_076_6690, w_076_6692, w_076_6693, w_076_6695, w_076_6698, w_076_6711, w_076_6713, w_076_6716, w_076_6719, w_076_6723, w_076_6726, w_076_6727, w_076_6728, w_076_6733, w_076_6745, w_076_6748, w_076_6749, w_076_6751, w_076_6758, w_076_6764, w_076_6765, w_076_6770, w_076_6772, w_076_6775, w_076_6785, w_076_6788, w_076_6789, w_076_6796, w_076_6798, w_076_6806, w_076_6808, w_076_6812, w_076_6813, w_076_6817, w_076_6819, w_076_6838, w_076_6840, w_076_6842, w_076_6845, w_076_6849, w_076_6850, w_076_6852, w_076_6855, w_076_6856, w_076_6857, w_076_6859, w_076_6864, w_076_6870, w_076_6876, w_076_6882, w_076_6883, w_076_6891, w_076_6892, w_076_6895, w_076_6896, w_076_6900, w_076_6901, w_076_6903, w_076_6908, w_076_6909, w_076_6911, w_076_6914, w_076_6916, w_076_6920, w_076_6923, w_076_6929, w_076_6931, w_076_6933, w_076_6939, w_076_6941, w_076_6942, w_076_6946, w_076_6948, w_076_6954, w_076_6956, w_076_6958, w_076_6959, w_076_6960, w_076_6963, w_076_6966, w_076_6970, w_076_6973, w_076_6974, w_076_6978, w_076_6983, w_076_6993, w_076_6994, w_076_6996, w_076_7005, w_076_7009, w_076_7013, w_076_7014, w_076_7026, w_076_7030, w_076_7032, w_076_7033, w_076_7034, w_076_7035, w_076_7036, w_076_7037, w_076_7041, w_076_7046, w_076_7051, w_076_7056, w_076_7057, w_076_7060, w_076_7061, w_076_7066, w_076_7073, w_076_7074, w_076_7075, w_076_7083, w_076_7093, w_076_7094, w_076_7095, w_076_7098, w_076_7099, w_076_7102, w_076_7109, w_076_7110, w_076_7116, w_076_7119, w_076_7131, w_076_7135, w_076_7136, w_076_7137, w_076_7138, w_076_7142, w_076_7144, w_076_7147, w_076_7149, w_076_7155, w_076_7157, w_076_7158, w_076_7165, w_076_7166, w_076_7171, w_076_7180, w_076_7183, w_076_7189, w_076_7190, w_076_7191, w_076_7193, w_076_7194, w_076_7195, w_076_7198, w_076_7203, w_076_7204, w_076_7212, w_076_7213, w_076_7214, w_076_7216, w_076_7217, w_076_7221, w_076_7224, w_076_7232, w_076_7235, w_076_7236, w_076_7239, w_076_7242;
  wire w_077_001, w_077_002, w_077_003, w_077_004, w_077_005, w_077_007, w_077_008, w_077_010, w_077_012, w_077_013, w_077_014, w_077_015, w_077_017, w_077_018, w_077_019, w_077_020, w_077_021, w_077_022, w_077_023, w_077_024, w_077_025, w_077_026, w_077_027, w_077_028, w_077_031, w_077_032, w_077_033, w_077_034, w_077_035, w_077_036, w_077_037, w_077_038, w_077_039, w_077_040, w_077_041, w_077_042, w_077_043, w_077_044, w_077_045, w_077_046, w_077_047, w_077_048, w_077_049, w_077_051, w_077_052, w_077_053, w_077_054, w_077_055, w_077_056, w_077_058, w_077_059, w_077_061, w_077_062, w_077_063, w_077_064, w_077_065, w_077_066, w_077_067, w_077_068, w_077_069, w_077_070, w_077_071, w_077_072, w_077_073, w_077_074, w_077_077, w_077_078, w_077_079, w_077_080, w_077_081, w_077_082, w_077_083, w_077_084, w_077_085, w_077_087, w_077_088, w_077_089, w_077_090, w_077_091, w_077_092, w_077_093, w_077_094, w_077_095, w_077_096, w_077_097, w_077_098, w_077_099, w_077_101, w_077_102, w_077_103, w_077_104, w_077_105, w_077_106, w_077_107, w_077_108, w_077_109, w_077_111, w_077_112, w_077_113, w_077_114, w_077_115, w_077_116, w_077_117, w_077_118, w_077_119, w_077_121, w_077_122, w_077_123, w_077_124, w_077_125, w_077_126, w_077_127, w_077_128, w_077_129, w_077_130, w_077_131, w_077_132, w_077_133, w_077_134, w_077_136, w_077_137, w_077_138, w_077_139, w_077_140, w_077_143, w_077_144, w_077_145, w_077_146, w_077_147, w_077_148, w_077_149, w_077_151, w_077_152, w_077_153, w_077_154, w_077_155, w_077_156, w_077_157, w_077_159, w_077_160, w_077_161, w_077_162, w_077_163, w_077_164, w_077_165, w_077_166, w_077_167, w_077_168, w_077_169, w_077_170, w_077_171, w_077_172, w_077_173, w_077_176, w_077_177, w_077_178, w_077_179, w_077_180, w_077_181, w_077_182, w_077_183, w_077_184, w_077_185, w_077_187, w_077_188, w_077_189, w_077_191, w_077_192, w_077_193, w_077_194, w_077_195, w_077_196, w_077_197, w_077_198, w_077_199, w_077_200, w_077_201, w_077_202, w_077_203, w_077_204, w_077_205, w_077_206, w_077_207, w_077_208, w_077_209, w_077_210, w_077_211, w_077_212, w_077_213, w_077_214, w_077_215, w_077_216, w_077_217, w_077_218, w_077_219, w_077_221, w_077_222, w_077_223, w_077_224, w_077_225, w_077_226, w_077_227, w_077_228, w_077_229, w_077_230, w_077_231, w_077_232, w_077_233, w_077_234, w_077_235, w_077_236, w_077_237, w_077_238, w_077_239, w_077_241, w_077_242, w_077_243, w_077_244, w_077_245, w_077_246, w_077_248, w_077_249, w_077_250, w_077_251, w_077_252, w_077_253, w_077_254, w_077_255, w_077_257, w_077_258, w_077_259, w_077_260, w_077_261, w_077_263, w_077_264, w_077_265, w_077_266, w_077_267, w_077_268, w_077_269, w_077_270, w_077_271, w_077_272, w_077_276, w_077_278, w_077_279, w_077_280, w_077_282, w_077_284, w_077_285, w_077_286, w_077_287, w_077_288, w_077_289, w_077_290, w_077_291, w_077_292, w_077_293, w_077_294, w_077_295, w_077_296, w_077_297, w_077_298, w_077_299, w_077_300, w_077_301, w_077_302, w_077_303, w_077_304, w_077_305, w_077_306, w_077_307, w_077_308, w_077_309, w_077_310, w_077_311, w_077_313, w_077_314, w_077_315, w_077_316, w_077_317, w_077_318, w_077_319, w_077_320, w_077_321, w_077_322, w_077_323, w_077_324, w_077_325, w_077_327, w_077_328, w_077_329, w_077_330, w_077_331, w_077_332, w_077_333, w_077_334, w_077_335, w_077_338, w_077_339, w_077_340, w_077_342, w_077_343, w_077_344, w_077_345, w_077_346, w_077_347, w_077_348, w_077_349, w_077_350, w_077_351, w_077_352, w_077_353, w_077_354, w_077_355, w_077_356, w_077_357, w_077_358, w_077_359, w_077_360, w_077_363, w_077_364, w_077_365, w_077_366, w_077_367, w_077_368, w_077_369, w_077_371, w_077_372, w_077_373, w_077_375, w_077_376, w_077_377, w_077_378, w_077_379, w_077_380, w_077_381, w_077_382, w_077_383, w_077_384, w_077_385, w_077_387, w_077_388, w_077_389, w_077_390, w_077_391, w_077_392, w_077_393, w_077_395, w_077_397, w_077_398, w_077_399, w_077_400, w_077_401, w_077_402, w_077_403, w_077_404, w_077_405, w_077_406, w_077_407, w_077_410, w_077_411, w_077_413, w_077_414, w_077_415, w_077_416, w_077_417, w_077_419, w_077_420, w_077_421, w_077_422, w_077_423, w_077_424, w_077_425, w_077_427, w_077_428, w_077_429, w_077_430, w_077_431, w_077_432, w_077_433, w_077_434, w_077_435, w_077_436, w_077_437, w_077_438, w_077_439, w_077_440, w_077_441, w_077_442, w_077_443, w_077_444, w_077_445, w_077_446, w_077_448, w_077_449, w_077_451, w_077_453, w_077_454, w_077_455, w_077_457, w_077_458, w_077_461, w_077_462, w_077_463, w_077_464, w_077_465, w_077_467, w_077_469, w_077_470, w_077_471, w_077_472, w_077_473, w_077_474, w_077_475, w_077_476, w_077_477, w_077_478, w_077_479, w_077_480, w_077_481, w_077_482, w_077_483, w_077_484, w_077_485, w_077_486, w_077_487, w_077_491, w_077_494, w_077_495, w_077_496, w_077_497, w_077_498, w_077_499, w_077_502, w_077_503, w_077_504, w_077_505, w_077_506, w_077_507, w_077_508, w_077_509, w_077_510, w_077_511, w_077_512, w_077_513, w_077_514, w_077_515, w_077_516, w_077_517, w_077_520, w_077_521, w_077_522, w_077_523, w_077_525, w_077_526, w_077_527, w_077_528, w_077_530, w_077_531, w_077_532, w_077_533, w_077_534, w_077_535, w_077_537, w_077_538, w_077_539, w_077_540, w_077_541, w_077_542, w_077_543, w_077_544, w_077_545, w_077_546, w_077_547, w_077_548, w_077_549, w_077_550, w_077_551, w_077_552, w_077_553, w_077_554, w_077_555, w_077_556, w_077_557, w_077_558, w_077_559, w_077_560, w_077_561, w_077_562, w_077_563, w_077_564, w_077_565, w_077_566, w_077_567, w_077_568, w_077_569, w_077_570, w_077_571, w_077_572, w_077_573, w_077_574, w_077_575, w_077_576, w_077_577, w_077_578, w_077_581, w_077_582, w_077_584, w_077_585, w_077_586, w_077_587, w_077_588, w_077_589, w_077_591, w_077_595, w_077_596, w_077_598, w_077_599, w_077_600, w_077_601, w_077_602, w_077_603, w_077_604, w_077_605, w_077_606, w_077_607, w_077_608, w_077_609, w_077_610, w_077_611, w_077_612, w_077_613, w_077_614, w_077_616, w_077_617, w_077_618, w_077_619, w_077_620, w_077_621, w_077_622, w_077_623, w_077_624, w_077_625, w_077_626, w_077_627, w_077_628, w_077_629, w_077_630, w_077_631, w_077_632, w_077_633, w_077_634, w_077_635, w_077_636, w_077_637, w_077_638, w_077_640, w_077_641, w_077_642, w_077_643, w_077_644, w_077_645, w_077_646, w_077_647, w_077_648, w_077_649, w_077_650, w_077_653, w_077_654, w_077_655, w_077_657, w_077_658, w_077_659, w_077_660, w_077_661, w_077_662, w_077_663, w_077_664, w_077_665, w_077_666, w_077_667, w_077_668, w_077_670, w_077_671, w_077_672, w_077_673, w_077_674, w_077_677, w_077_679, w_077_680, w_077_682, w_077_683, w_077_684, w_077_686, w_077_687, w_077_688, w_077_689, w_077_690, w_077_691, w_077_692, w_077_693, w_077_694, w_077_695, w_077_696, w_077_697, w_077_698, w_077_699, w_077_700, w_077_701, w_077_702, w_077_703, w_077_704, w_077_705, w_077_706, w_077_707, w_077_708, w_077_709, w_077_710, w_077_711, w_077_712, w_077_713, w_077_714, w_077_715, w_077_716, w_077_717, w_077_718, w_077_719, w_077_720, w_077_721, w_077_723, w_077_724, w_077_725, w_077_727, w_077_728, w_077_730, w_077_733, w_077_735, w_077_736, w_077_738, w_077_739, w_077_740, w_077_741, w_077_742, w_077_743, w_077_745, w_077_747, w_077_748, w_077_750, w_077_751, w_077_753, w_077_755, w_077_756, w_077_757, w_077_758, w_077_759, w_077_760, w_077_762, w_077_763, w_077_765, w_077_766, w_077_767, w_077_768, w_077_769, w_077_772, w_077_773, w_077_774, w_077_775, w_077_776, w_077_777, w_077_778, w_077_780, w_077_781, w_077_782, w_077_783, w_077_784, w_077_785, w_077_786, w_077_787, w_077_788, w_077_789, w_077_790, w_077_791, w_077_792, w_077_795, w_077_796, w_077_797, w_077_798, w_077_799, w_077_800, w_077_801, w_077_802, w_077_804, w_077_805, w_077_806, w_077_807, w_077_809, w_077_810, w_077_812, w_077_814, w_077_815, w_077_816, w_077_818, w_077_819, w_077_820, w_077_821, w_077_822, w_077_823, w_077_824, w_077_825, w_077_826, w_077_827, w_077_828, w_077_829, w_077_830, w_077_831, w_077_832, w_077_833, w_077_834, w_077_835, w_077_836, w_077_837, w_077_839, w_077_841, w_077_842, w_077_843, w_077_844, w_077_846, w_077_847, w_077_848, w_077_849, w_077_850, w_077_852, w_077_853, w_077_855, w_077_856, w_077_857, w_077_859, w_077_860, w_077_861, w_077_864, w_077_865, w_077_866, w_077_867, w_077_868, w_077_870, w_077_871, w_077_872, w_077_873, w_077_874, w_077_875, w_077_876, w_077_877, w_077_878, w_077_880, w_077_881, w_077_882, w_077_883, w_077_885, w_077_887, w_077_888, w_077_889, w_077_890, w_077_892, w_077_893, w_077_894, w_077_896, w_077_897, w_077_898, w_077_899, w_077_900, w_077_901, w_077_902, w_077_903, w_077_904, w_077_905, w_077_906, w_077_907, w_077_909, w_077_910, w_077_911, w_077_913, w_077_916, w_077_917, w_077_920, w_077_922, w_077_924, w_077_926, w_077_929, w_077_931, w_077_933, w_077_934, w_077_935, w_077_936, w_077_937, w_077_939, w_077_940, w_077_942, w_077_944, w_077_945, w_077_947, w_077_949, w_077_951, w_077_952, w_077_953, w_077_954, w_077_955, w_077_956, w_077_957, w_077_958, w_077_959, w_077_960, w_077_961, w_077_963, w_077_964, w_077_965, w_077_967, w_077_968, w_077_969, w_077_970, w_077_972, w_077_973, w_077_974, w_077_975, w_077_976, w_077_977, w_077_978, w_077_979, w_077_980, w_077_981, w_077_982, w_077_983, w_077_984, w_077_985, w_077_986, w_077_987, w_077_988, w_077_989, w_077_990, w_077_991, w_077_992, w_077_993, w_077_994, w_077_995, w_077_996, w_077_998, w_077_999, w_077_1000, w_077_1001, w_077_1002, w_077_1003, w_077_1004, w_077_1005, w_077_1006, w_077_1007, w_077_1008, w_077_1009, w_077_1010, w_077_1011, w_077_1012, w_077_1013, w_077_1014, w_077_1015, w_077_1016, w_077_1017, w_077_1019, w_077_1021, w_077_1023, w_077_1024, w_077_1025, w_077_1026, w_077_1027, w_077_1029, w_077_1030, w_077_1031, w_077_1032, w_077_1034, w_077_1035, w_077_1036, w_077_1037, w_077_1038, w_077_1040, w_077_1041, w_077_1043, w_077_1044, w_077_1045, w_077_1046, w_077_1047, w_077_1048, w_077_1049, w_077_1051, w_077_1053, w_077_1054, w_077_1055, w_077_1059, w_077_1060, w_077_1061, w_077_1062, w_077_1065, w_077_1066, w_077_1068, w_077_1069, w_077_1070, w_077_1071, w_077_1072, w_077_1073, w_077_1074, w_077_1075, w_077_1076, w_077_1077, w_077_1078, w_077_1079, w_077_1080, w_077_1081, w_077_1083, w_077_1084, w_077_1086, w_077_1087, w_077_1088, w_077_1091, w_077_1092, w_077_1093, w_077_1094, w_077_1096, w_077_1097, w_077_1098, w_077_1099, w_077_1100, w_077_1103, w_077_1104, w_077_1105, w_077_1106, w_077_1108, w_077_1109, w_077_1110, w_077_1112, w_077_1113, w_077_1116, w_077_1117, w_077_1118, w_077_1119, w_077_1120, w_077_1121, w_077_1122, w_077_1123, w_077_1124, w_077_1125, w_077_1127, w_077_1128, w_077_1129, w_077_1130, w_077_1132, w_077_1133, w_077_1134, w_077_1135, w_077_1136, w_077_1137, w_077_1138, w_077_1139, w_077_1140, w_077_1141, w_077_1143, w_077_1144, w_077_1145, w_077_1148, w_077_1151, w_077_1152, w_077_1154, w_077_1155, w_077_1159, w_077_1160, w_077_1162, w_077_1163, w_077_1164, w_077_1165, w_077_1166, w_077_1167, w_077_1168, w_077_1169, w_077_1170, w_077_1171, w_077_1173, w_077_1174, w_077_1175, w_077_1176, w_077_1177, w_077_1178, w_077_1179, w_077_1180, w_077_1181, w_077_1182, w_077_1183, w_077_1184, w_077_1185, w_077_1186, w_077_1187, w_077_1188, w_077_1189, w_077_1191, w_077_1192, w_077_1193, w_077_1194, w_077_1195, w_077_1196, w_077_1197, w_077_1198, w_077_1199, w_077_1200, w_077_1201, w_077_1202, w_077_1203, w_077_1204, w_077_1206, w_077_1208, w_077_1209, w_077_1210, w_077_1211, w_077_1212, w_077_1213, w_077_1214, w_077_1215, w_077_1216, w_077_1217, w_077_1218, w_077_1219, w_077_1220, w_077_1221, w_077_1222, w_077_1224, w_077_1225, w_077_1226, w_077_1227, w_077_1229, w_077_1231, w_077_1233, w_077_1234, w_077_1235, w_077_1237, w_077_1239, w_077_1240, w_077_1241, w_077_1242, w_077_1243, w_077_1244, w_077_1247, w_077_1248, w_077_1249, w_077_1250, w_077_1251, w_077_1253, w_077_1256, w_077_1257, w_077_1258, w_077_1259, w_077_1260, w_077_1262, w_077_1264, w_077_1266, w_077_1267, w_077_1269, w_077_1270, w_077_1271, w_077_1272, w_077_1273, w_077_1274, w_077_1277, w_077_1279, w_077_1280, w_077_1282, w_077_1283, w_077_1284, w_077_1285, w_077_1286, w_077_1287, w_077_1288, w_077_1289, w_077_1290, w_077_1291, w_077_1292, w_077_1293, w_077_1295, w_077_1296, w_077_1297, w_077_1299, w_077_1300, w_077_1301, w_077_1302, w_077_1303, w_077_1304, w_077_1305, w_077_1306, w_077_1307, w_077_1308, w_077_1309, w_077_1310, w_077_1311, w_077_1312, w_077_1314, w_077_1315, w_077_1317, w_077_1318, w_077_1319, w_077_1320, w_077_1321, w_077_1322, w_077_1323, w_077_1324, w_077_1325, w_077_1328, w_077_1329, w_077_1330, w_077_1331, w_077_1332, w_077_1333, w_077_1334, w_077_1336, w_077_1337, w_077_1338, w_077_1339, w_077_1340, w_077_1341, w_077_1342, w_077_1343, w_077_1344, w_077_1345, w_077_1346, w_077_1347, w_077_1348, w_077_1349, w_077_1350, w_077_1351, w_077_1352, w_077_1353, w_077_1354, w_077_1355, w_077_1356, w_077_1357, w_077_1358, w_077_1359, w_077_1360, w_077_1361, w_077_1362, w_077_1363, w_077_1364, w_077_1365, w_077_1366, w_077_1367, w_077_1368, w_077_1369, w_077_1370, w_077_1371, w_077_1372, w_077_1374, w_077_1375, w_077_1376, w_077_1377, w_077_1378, w_077_1379, w_077_1381, w_077_1382, w_077_1383, w_077_1385, w_077_1388, w_077_1389, w_077_1390, w_077_1391, w_077_1392, w_077_1393, w_077_1395, w_077_1396, w_077_1397, w_077_1398, w_077_1399, w_077_1400, w_077_1401, w_077_1402, w_077_1403, w_077_1404, w_077_1405, w_077_1406, w_077_1408, w_077_1409, w_077_1410, w_077_1411, w_077_1412, w_077_1414, w_077_1415, w_077_1416, w_077_1417, w_077_1418, w_077_1420, w_077_1421, w_077_1423, w_077_1425, w_077_1426, w_077_1428, w_077_1429, w_077_1430, w_077_1431, w_077_1432, w_077_1433, w_077_1434, w_077_1435, w_077_1436, w_077_1437, w_077_1438, w_077_1440, w_077_1441, w_077_1442, w_077_1444, w_077_1445, w_077_1446, w_077_1447, w_077_1448, w_077_1449, w_077_1450, w_077_1452, w_077_1453, w_077_1454, w_077_1455, w_077_1458, w_077_1459, w_077_1460, w_077_1461, w_077_1462, w_077_1463, w_077_1464, w_077_1465, w_077_1466, w_077_1467, w_077_1468, w_077_1469, w_077_1470, w_077_1471, w_077_1473, w_077_1474, w_077_1475, w_077_1476, w_077_1478, w_077_1479, w_077_1480, w_077_1481, w_077_1482, w_077_1483, w_077_1484, w_077_1485, w_077_1486, w_077_1488, w_077_1489, w_077_1490, w_077_1492, w_077_1496, w_077_1497, w_077_1498, w_077_1499, w_077_1501, w_077_1503, w_077_1505, w_077_1507, w_077_1508, w_077_1509, w_077_1510, w_077_1511, w_077_1512, w_077_1513, w_077_1514, w_077_1515, w_077_1516, w_077_1517, w_077_1518, w_077_1519, w_077_1520, w_077_1522, w_077_1523, w_077_1524, w_077_1525, w_077_1526, w_077_1527, w_077_1528, w_077_1529, w_077_1530, w_077_1531, w_077_1532, w_077_1534, w_077_1535, w_077_1536, w_077_1537, w_077_1539, w_077_1540, w_077_1541, w_077_1543, w_077_1545, w_077_1546, w_077_1547, w_077_1551, w_077_1552, w_077_1553, w_077_1555, w_077_1556, w_077_1557, w_077_1559, w_077_1561, w_077_1562, w_077_1563, w_077_1564, w_077_1565, w_077_1567, w_077_1568, w_077_1569, w_077_1570, w_077_1571, w_077_1572, w_077_1573, w_077_1574, w_077_1576, w_077_1577, w_077_1578, w_077_1579, w_077_1582, w_077_1583, w_077_1584, w_077_1585, w_077_1586, w_077_1587, w_077_1588, w_077_1590, w_077_1592, w_077_1593, w_077_1594, w_077_1595, w_077_1596, w_077_1597, w_077_1598, w_077_1599, w_077_1600, w_077_1601, w_077_1602, w_077_1603, w_077_1604, w_077_1605, w_077_1607, w_077_1608, w_077_1609, w_077_1610, w_077_1611, w_077_1612, w_077_1614, w_077_1615, w_077_1616, w_077_1617, w_077_1618, w_077_1619, w_077_1620, w_077_1621, w_077_1622, w_077_1623, w_077_1624, w_077_1625, w_077_1628, w_077_1629, w_077_1630, w_077_1631, w_077_1632, w_077_1633, w_077_1634, w_077_1635, w_077_1636, w_077_1637, w_077_1639, w_077_1640, w_077_1641, w_077_1642, w_077_1643, w_077_1644, w_077_1648, w_077_1649, w_077_1650, w_077_1651, w_077_1652, w_077_1654, w_077_1655, w_077_1657, w_077_1658, w_077_1659, w_077_1660, w_077_1661, w_077_1663, w_077_1664, w_077_1665, w_077_1666, w_077_1667, w_077_1668, w_077_1670, w_077_1671, w_077_1672, w_077_1673, w_077_1674, w_077_1675, w_077_1676, w_077_1677, w_077_1678, w_077_1680, w_077_1681, w_077_1684, w_077_1685, w_077_1686, w_077_1687, w_077_1688, w_077_1689, w_077_1690, w_077_1691, w_077_1692, w_077_1693, w_077_1694, w_077_1695, w_077_1696, w_077_1697, w_077_1698, w_077_1699, w_077_1700, w_077_1702, w_077_1703, w_077_1704, w_077_1706, w_077_1707, w_077_1708, w_077_1709, w_077_1711, w_077_1713, w_077_1714, w_077_1716, w_077_1718, w_077_1719, w_077_1720, w_077_1721, w_077_1722, w_077_1723, w_077_1724, w_077_1728, w_077_1729, w_077_1731, w_077_1732, w_077_1733, w_077_1734, w_077_1735, w_077_1736, w_077_1737, w_077_1738, w_077_1740, w_077_1741, w_077_1743, w_077_1744, w_077_1745, w_077_1746, w_077_1747, w_077_1748, w_077_1749, w_077_1750, w_077_1751, w_077_1752, w_077_1753, w_077_1754, w_077_1756, w_077_1757, w_077_1758, w_077_1759, w_077_1760, w_077_1761, w_077_1762, w_077_1763, w_077_1764, w_077_1765, w_077_1766, w_077_1768, w_077_1769, w_077_1771, w_077_1774, w_077_1776, w_077_1778, w_077_1780, w_077_1783, w_077_1784, w_077_1785, w_077_1786, w_077_1787, w_077_1788, w_077_1789, w_077_1790, w_077_1791, w_077_1793, w_077_1795, w_077_1796, w_077_1797, w_077_1798, w_077_1799, w_077_1800, w_077_1801, w_077_1802, w_077_1803, w_077_1804, w_077_1805, w_077_1806, w_077_1808, w_077_1812, w_077_1813, w_077_1814, w_077_1818, w_077_1819, w_077_1820, w_077_1823, w_077_1824, w_077_1826, w_077_1827, w_077_1828, w_077_1829, w_077_1830, w_077_1831, w_077_1833, w_077_1834, w_077_1835, w_077_1836, w_077_1837, w_077_1838, w_077_1839, w_077_1841, w_077_1842, w_077_1846, w_077_1847, w_077_1848, w_077_1849, w_077_1850, w_077_1851, w_077_1852, w_077_1853, w_077_1857, w_077_1858, w_077_1859, w_077_1860, w_077_1861, w_077_1863, w_077_1864, w_077_1865, w_077_1866, w_077_1867, w_077_1868, w_077_1869, w_077_1871, w_077_1872, w_077_1874, w_077_1875, w_077_1876, w_077_1878, w_077_1879, w_077_1880;
  wire w_078_000, w_078_001, w_078_002, w_078_003, w_078_004, w_078_005, w_078_006, w_078_007, w_078_008, w_078_009, w_078_010, w_078_011, w_078_012, w_078_013, w_078_014, w_078_015, w_078_016, w_078_018, w_078_019, w_078_021, w_078_022, w_078_024, w_078_025, w_078_026, w_078_027, w_078_028, w_078_029, w_078_030, w_078_031, w_078_033, w_078_034, w_078_035, w_078_036, w_078_037, w_078_038, w_078_039, w_078_040, w_078_041, w_078_042, w_078_043, w_078_044, w_078_045, w_078_046, w_078_047, w_078_048, w_078_049, w_078_050, w_078_051, w_078_052, w_078_053, w_078_054, w_078_055, w_078_056, w_078_057, w_078_058, w_078_059, w_078_060, w_078_061, w_078_062, w_078_063, w_078_064, w_078_065, w_078_066, w_078_067, w_078_068, w_078_069, w_078_070, w_078_071, w_078_072, w_078_073, w_078_074, w_078_075, w_078_076, w_078_077, w_078_078, w_078_079, w_078_080, w_078_081, w_078_082, w_078_083, w_078_084, w_078_085, w_078_086, w_078_087, w_078_088, w_078_089, w_078_090, w_078_091, w_078_092, w_078_093, w_078_094, w_078_095, w_078_096, w_078_097, w_078_098, w_078_099, w_078_100, w_078_101, w_078_102, w_078_103, w_078_104, w_078_105, w_078_106, w_078_107, w_078_108, w_078_109, w_078_110, w_078_111, w_078_113, w_078_114, w_078_115, w_078_116, w_078_117, w_078_118, w_078_119, w_078_120, w_078_121, w_078_122, w_078_123, w_078_124, w_078_125, w_078_126, w_078_127, w_078_128, w_078_129, w_078_130, w_078_131, w_078_132, w_078_133, w_078_134, w_078_135, w_078_136, w_078_137, w_078_138, w_078_140, w_078_141, w_078_142, w_078_143, w_078_144, w_078_145, w_078_146, w_078_147, w_078_148, w_078_149, w_078_150, w_078_151, w_078_152, w_078_153, w_078_154, w_078_155, w_078_156, w_078_157, w_078_158, w_078_159, w_078_160, w_078_161, w_078_162, w_078_163, w_078_164, w_078_165, w_078_166, w_078_167, w_078_168, w_078_169, w_078_170, w_078_171, w_078_172, w_078_173, w_078_174, w_078_175, w_078_176, w_078_177, w_078_178, w_078_179, w_078_180, w_078_181, w_078_182, w_078_183, w_078_184, w_078_185, w_078_186, w_078_187, w_078_188, w_078_189, w_078_190, w_078_191, w_078_192, w_078_193, w_078_194, w_078_195, w_078_196, w_078_197, w_078_198, w_078_200, w_078_201, w_078_202, w_078_203, w_078_204, w_078_205, w_078_206, w_078_207, w_078_208, w_078_209, w_078_210, w_078_211, w_078_212, w_078_213, w_078_214, w_078_215, w_078_216, w_078_217, w_078_218, w_078_219, w_078_220, w_078_221, w_078_222, w_078_223, w_078_224, w_078_225, w_078_226, w_078_227, w_078_228, w_078_229, w_078_230, w_078_231, w_078_232, w_078_233, w_078_234, w_078_235, w_078_236, w_078_237, w_078_238, w_078_239, w_078_240, w_078_241, w_078_242, w_078_243, w_078_244, w_078_245, w_078_246, w_078_247, w_078_248, w_078_249, w_078_250, w_078_251, w_078_252, w_078_253, w_078_254, w_078_255, w_078_256, w_078_257, w_078_258, w_078_259, w_078_260, w_078_261, w_078_262, w_078_263, w_078_264, w_078_265, w_078_266, w_078_267, w_078_268, w_078_269, w_078_270, w_078_271, w_078_272, w_078_273, w_078_274, w_078_275, w_078_276, w_078_277, w_078_278, w_078_279, w_078_280, w_078_281, w_078_282, w_078_284, w_078_285, w_078_286, w_078_287, w_078_288, w_078_289, w_078_290, w_078_291, w_078_292, w_078_293, w_078_294, w_078_295, w_078_296, w_078_297, w_078_298, w_078_299, w_078_300, w_078_301, w_078_302, w_078_303, w_078_304, w_078_305, w_078_308, w_078_309, w_078_310, w_078_311, w_078_312, w_078_313, w_078_314, w_078_315, w_078_316, w_078_317, w_078_318, w_078_319, w_078_320, w_078_321, w_078_323, w_078_324, w_078_325, w_078_326, w_078_327, w_078_328, w_078_329, w_078_330, w_078_331, w_078_332, w_078_333, w_078_334, w_078_335, w_078_336, w_078_337, w_078_338, w_078_339, w_078_340, w_078_341, w_078_342, w_078_343, w_078_344, w_078_345, w_078_346, w_078_347, w_078_348, w_078_349, w_078_350, w_078_351, w_078_353, w_078_354, w_078_355, w_078_356, w_078_357, w_078_358, w_078_359, w_078_360, w_078_361, w_078_362, w_078_363, w_078_364, w_078_365, w_078_366, w_078_367, w_078_369, w_078_370, w_078_371, w_078_372, w_078_373, w_078_374, w_078_375, w_078_376, w_078_377, w_078_378, w_078_379, w_078_380, w_078_381, w_078_382, w_078_383, w_078_384, w_078_385, w_078_386, w_078_387, w_078_388, w_078_390, w_078_391, w_078_392, w_078_393, w_078_394, w_078_395, w_078_396, w_078_397, w_078_398, w_078_399, w_078_400, w_078_401, w_078_402, w_078_403, w_078_404, w_078_405, w_078_406, w_078_407, w_078_408, w_078_409, w_078_410, w_078_411, w_078_412, w_078_413, w_078_414, w_078_415, w_078_416, w_078_417, w_078_418, w_078_419, w_078_420, w_078_421, w_078_422, w_078_423, w_078_424, w_078_426, w_078_427, w_078_429, w_078_430, w_078_431, w_078_432, w_078_433, w_078_434, w_078_435, w_078_436, w_078_437, w_078_438, w_078_440, w_078_442, w_078_443, w_078_444, w_078_445, w_078_446, w_078_447, w_078_448, w_078_449, w_078_450, w_078_451, w_078_452, w_078_453, w_078_454, w_078_455, w_078_456, w_078_457, w_078_458, w_078_459, w_078_460, w_078_461, w_078_462, w_078_464, w_078_465, w_078_466, w_078_467, w_078_468, w_078_469, w_078_470, w_078_471, w_078_472, w_078_473, w_078_474, w_078_475, w_078_476, w_078_478, w_078_479, w_078_481, w_078_482, w_078_483, w_078_484, w_078_485, w_078_486, w_078_487, w_078_488, w_078_489, w_078_490, w_078_492, w_078_493, w_078_494, w_078_495, w_078_496, w_078_497, w_078_498, w_078_499, w_078_500, w_078_501, w_078_502, w_078_503, w_078_504, w_078_505, w_078_506, w_078_507, w_078_508, w_078_509, w_078_510, w_078_511, w_078_512, w_078_513, w_078_514, w_078_515, w_078_516, w_078_518, w_078_519, w_078_520, w_078_521, w_078_522, w_078_523, w_078_524, w_078_525, w_078_526, w_078_527, w_078_528, w_078_529, w_078_530, w_078_531, w_078_532, w_078_533, w_078_534, w_078_535, w_078_536, w_078_537, w_078_538, w_078_539, w_078_540, w_078_541, w_078_542, w_078_543, w_078_544, w_078_545, w_078_546, w_078_548, w_078_549, w_078_550, w_078_551, w_078_552, w_078_553, w_078_554, w_078_555, w_078_556, w_078_557, w_078_558, w_078_559, w_078_560, w_078_561, w_078_562, w_078_563, w_078_564, w_078_565, w_078_566, w_078_567, w_078_568, w_078_569, w_078_570, w_078_571, w_078_572, w_078_573, w_078_574, w_078_575, w_078_576, w_078_577, w_078_578, w_078_579, w_078_580, w_078_581, w_078_582, w_078_583, w_078_584, w_078_585, w_078_586, w_078_587, w_078_588, w_078_589, w_078_590, w_078_591, w_078_592, w_078_593, w_078_594, w_078_595, w_078_596, w_078_597, w_078_598, w_078_599, w_078_600, w_078_601, w_078_602, w_078_603, w_078_604, w_078_605, w_078_606, w_078_607, w_078_608, w_078_609, w_078_610, w_078_611, w_078_612, w_078_613, w_078_614, w_078_615, w_078_616, w_078_617, w_078_618, w_078_619, w_078_620, w_078_621, w_078_622, w_078_623, w_078_624, w_078_625, w_078_626, w_078_627, w_078_628, w_078_629, w_078_630, w_078_631, w_078_632, w_078_633, w_078_634, w_078_635, w_078_636, w_078_637, w_078_638, w_078_640, w_078_641, w_078_642, w_078_643, w_078_644, w_078_645, w_078_646, w_078_647, w_078_648, w_078_649, w_078_650, w_078_651, w_078_652, w_078_653, w_078_654, w_078_655, w_078_656, w_078_657, w_078_658, w_078_659, w_078_660, w_078_661, w_078_662, w_078_663, w_078_665, w_078_666, w_078_667, w_078_668, w_078_669, w_078_670, w_078_672, w_078_673, w_078_674, w_078_675, w_078_676, w_078_677, w_078_678, w_078_679, w_078_680, w_078_682, w_078_683, w_078_684, w_078_685, w_078_686, w_078_687, w_078_688, w_078_689, w_078_690, w_078_691, w_078_692, w_078_693, w_078_694, w_078_695, w_078_696, w_078_697, w_078_698, w_078_699, w_078_700, w_078_701, w_078_702, w_078_703, w_078_704, w_078_705, w_078_706, w_078_708, w_078_709, w_078_710, w_078_711, w_078_712, w_078_713, w_078_714, w_078_716, w_078_717, w_078_718, w_078_719, w_078_720, w_078_721, w_078_722, w_078_724, w_078_725, w_078_726, w_078_727, w_078_728, w_078_729, w_078_732, w_078_733, w_078_734, w_078_736, w_078_737, w_078_738, w_078_739, w_078_740, w_078_741, w_078_742, w_078_743, w_078_744, w_078_745, w_078_746, w_078_747, w_078_748, w_078_749, w_078_750, w_078_751, w_078_752, w_078_753, w_078_754, w_078_755, w_078_756, w_078_757, w_078_758, w_078_759, w_078_760, w_078_761, w_078_762, w_078_763, w_078_764, w_078_765, w_078_766, w_078_767, w_078_768, w_078_769, w_078_770, w_078_771, w_078_772, w_078_773, w_078_774, w_078_775, w_078_776, w_078_777, w_078_778, w_078_779, w_078_780, w_078_781, w_078_782, w_078_784, w_078_785, w_078_786, w_078_787, w_078_788, w_078_789, w_078_790, w_078_791, w_078_792, w_078_793, w_078_794, w_078_795, w_078_796, w_078_798, w_078_799, w_078_800, w_078_801, w_078_802, w_078_804, w_078_805, w_078_806, w_078_807, w_078_808, w_078_809, w_078_810, w_078_811, w_078_812, w_078_813, w_078_814, w_078_815, w_078_816, w_078_817, w_078_818, w_078_819, w_078_821, w_078_822, w_078_823, w_078_825, w_078_826, w_078_827, w_078_828, w_078_829, w_078_830, w_078_831, w_078_832, w_078_833, w_078_834, w_078_836, w_078_837, w_078_838, w_078_839, w_078_840, w_078_841, w_078_842, w_078_843, w_078_844, w_078_845, w_078_846, w_078_847, w_078_848, w_078_849, w_078_850, w_078_852, w_078_853, w_078_854, w_078_856, w_078_857, w_078_858, w_078_859, w_078_860, w_078_861, w_078_862, w_078_863, w_078_864, w_078_865, w_078_866, w_078_867, w_078_868, w_078_869, w_078_871, w_078_872, w_078_873, w_078_874, w_078_875, w_078_876, w_078_877, w_078_878, w_078_879, w_078_880, w_078_881, w_078_882, w_078_883, w_078_884, w_078_885, w_078_886, w_078_887, w_078_889, w_078_890, w_078_891, w_078_892, w_078_893, w_078_894, w_078_895, w_078_896, w_078_897, w_078_898, w_078_899, w_078_900, w_078_901, w_078_902, w_078_903, w_078_904, w_078_905, w_078_906, w_078_907, w_078_908, w_078_909, w_078_910, w_078_911, w_078_912, w_078_913, w_078_914, w_078_915, w_078_916, w_078_917, w_078_918, w_078_919, w_078_920, w_078_921, w_078_922, w_078_923, w_078_924, w_078_925, w_078_927, w_078_928, w_078_929, w_078_932, w_078_933, w_078_934, w_078_935, w_078_937, w_078_939, w_078_940, w_078_941, w_078_942, w_078_943, w_078_944, w_078_945, w_078_946, w_078_947, w_078_948, w_078_949, w_078_950, w_078_951, w_078_952, w_078_953, w_078_954, w_078_955, w_078_956, w_078_957, w_078_958, w_078_959, w_078_960, w_078_961, w_078_962, w_078_963, w_078_964, w_078_965, w_078_966, w_078_967, w_078_968, w_078_969, w_078_970, w_078_971, w_078_972, w_078_973, w_078_974, w_078_975, w_078_976, w_078_978, w_078_979, w_078_980, w_078_981, w_078_982, w_078_983, w_078_984, w_078_985, w_078_986, w_078_988, w_078_989, w_078_990, w_078_991, w_078_992, w_078_993, w_078_994, w_078_995, w_078_996, w_078_997, w_078_998, w_078_999, w_078_1000, w_078_1001, w_078_1002, w_078_1003, w_078_1004, w_078_1005, w_078_1006, w_078_1008, w_078_1009, w_078_1010, w_078_1011, w_078_1012, w_078_1013, w_078_1015, w_078_1016, w_078_1017, w_078_1018, w_078_1019, w_078_1020, w_078_1021, w_078_1022, w_078_1023, w_078_1024, w_078_1025, w_078_1026, w_078_1027, w_078_1028, w_078_1029, w_078_1030, w_078_1031, w_078_1032, w_078_1033, w_078_1034, w_078_1035, w_078_1036, w_078_1037, w_078_1038, w_078_1039, w_078_1040, w_078_1041, w_078_1042, w_078_1044, w_078_1045, w_078_1047, w_078_1048, w_078_1049, w_078_1050, w_078_1051, w_078_1052, w_078_1053, w_078_1054, w_078_1055, w_078_1056, w_078_1057, w_078_1059, w_078_1060, w_078_1061, w_078_1062, w_078_1063, w_078_1064, w_078_1065, w_078_1066, w_078_1067, w_078_1068, w_078_1069, w_078_1070, w_078_1071, w_078_1072, w_078_1073, w_078_1074, w_078_1075, w_078_1076, w_078_1077, w_078_1078, w_078_1079, w_078_1080, w_078_1082, w_078_1083, w_078_1084, w_078_1085, w_078_1086, w_078_1087, w_078_1088, w_078_1089, w_078_1090, w_078_1091, w_078_1092, w_078_1093, w_078_1094, w_078_1095, w_078_1096, w_078_1097, w_078_1098, w_078_1099, w_078_1100, w_078_1101, w_078_1102, w_078_1103, w_078_1104, w_078_1105, w_078_1106, w_078_1107, w_078_1108, w_078_1109, w_078_1110, w_078_1111, w_078_1112, w_078_1113, w_078_1114, w_078_1115, w_078_1116, w_078_1117, w_078_1118, w_078_1119, w_078_1120, w_078_1121, w_078_1122, w_078_1123, w_078_1124, w_078_1126, w_078_1128, w_078_1129, w_078_1130, w_078_1131, w_078_1132, w_078_1133, w_078_1134, w_078_1135, w_078_1136, w_078_1137, w_078_1138, w_078_1139, w_078_1140, w_078_1141, w_078_1142, w_078_1143, w_078_1144, w_078_1145, w_078_1146, w_078_1147, w_078_1148;
  wire w_079_000, w_079_001, w_079_002, w_079_003, w_079_004, w_079_005, w_079_008, w_079_009, w_079_010, w_079_012, w_079_015, w_079_016, w_079_018, w_079_019, w_079_021, w_079_022, w_079_024, w_079_026, w_079_030, w_079_031, w_079_032, w_079_033, w_079_034, w_079_035, w_079_036, w_079_037, w_079_038, w_079_039, w_079_040, w_079_041, w_079_042, w_079_046, w_079_047, w_079_049, w_079_050, w_079_052, w_079_053, w_079_054, w_079_055, w_079_057, w_079_058, w_079_060, w_079_061, w_079_062, w_079_063, w_079_067, w_079_069, w_079_070, w_079_072, w_079_074, w_079_075, w_079_076, w_079_077, w_079_078, w_079_079, w_079_082, w_079_083, w_079_084, w_079_085, w_079_086, w_079_089, w_079_091, w_079_092, w_079_093, w_079_094, w_079_099, w_079_100, w_079_102, w_079_104, w_079_106, w_079_107, w_079_109, w_079_112, w_079_113, w_079_114, w_079_115, w_079_117, w_079_118, w_079_119, w_079_120, w_079_121, w_079_122, w_079_124, w_079_125, w_079_128, w_079_129, w_079_130, w_079_133, w_079_135, w_079_137, w_079_138, w_079_139, w_079_142, w_079_143, w_079_144, w_079_145, w_079_146, w_079_148, w_079_149, w_079_150, w_079_152, w_079_155, w_079_157, w_079_160, w_079_161, w_079_162, w_079_165, w_079_166, w_079_167, w_079_170, w_079_171, w_079_172, w_079_174, w_079_177, w_079_178, w_079_179, w_079_181, w_079_182, w_079_185, w_079_186, w_079_188, w_079_190, w_079_192, w_079_193, w_079_194, w_079_195, w_079_197, w_079_200, w_079_201, w_079_202, w_079_204, w_079_205, w_079_207, w_079_208, w_079_209, w_079_215, w_079_217, w_079_218, w_079_219, w_079_220, w_079_221, w_079_223, w_079_224, w_079_225, w_079_227, w_079_228, w_079_229, w_079_232, w_079_233, w_079_234, w_079_235, w_079_236, w_079_238, w_079_240, w_079_241, w_079_243, w_079_244, w_079_246, w_079_248, w_079_250, w_079_251, w_079_252, w_079_253, w_079_254, w_079_255, w_079_256, w_079_257, w_079_259, w_079_260, w_079_262, w_079_263, w_079_264, w_079_265, w_079_266, w_079_267, w_079_268, w_079_272, w_079_273, w_079_274, w_079_275, w_079_276, w_079_277, w_079_279, w_079_280, w_079_281, w_079_282, w_079_285, w_079_289, w_079_290, w_079_292, w_079_293, w_079_294, w_079_295, w_079_296, w_079_298, w_079_299, w_079_300, w_079_303, w_079_307, w_079_308, w_079_309, w_079_311, w_079_313, w_079_315, w_079_317, w_079_318, w_079_320, w_079_323, w_079_324, w_079_325, w_079_326, w_079_327, w_079_328, w_079_329, w_079_331, w_079_332, w_079_333, w_079_335, w_079_336, w_079_337, w_079_339, w_079_340, w_079_341, w_079_342, w_079_346, w_079_350, w_079_351, w_079_354, w_079_356, w_079_357, w_079_358, w_079_359, w_079_361, w_079_363, w_079_364, w_079_366, w_079_368, w_079_369, w_079_370, w_079_371, w_079_374, w_079_375, w_079_377, w_079_378, w_079_382, w_079_385, w_079_387, w_079_388, w_079_391, w_079_393, w_079_394, w_079_396, w_079_397, w_079_398, w_079_399, w_079_400, w_079_401, w_079_402, w_079_403, w_079_404, w_079_406, w_079_407, w_079_408, w_079_409, w_079_410, w_079_411, w_079_413, w_079_414, w_079_415, w_079_420, w_079_421, w_079_422, w_079_424, w_079_427, w_079_430, w_079_431, w_079_432, w_079_434, w_079_435, w_079_436, w_079_438, w_079_439, w_079_440, w_079_441, w_079_442, w_079_444, w_079_446, w_079_447, w_079_449, w_079_450, w_079_452, w_079_453, w_079_454, w_079_455, w_079_456, w_079_459, w_079_460, w_079_462, w_079_463, w_079_466, w_079_468, w_079_469, w_079_470, w_079_471, w_079_473, w_079_478, w_079_479, w_079_481, w_079_482, w_079_483, w_079_484, w_079_485, w_079_486, w_079_487, w_079_489, w_079_490, w_079_491, w_079_492, w_079_493, w_079_494, w_079_495, w_079_496, w_079_498, w_079_499, w_079_500, w_079_501, w_079_503, w_079_506, w_079_507, w_079_508, w_079_509, w_079_511, w_079_512, w_079_513, w_079_514, w_079_515, w_079_516, w_079_517, w_079_518, w_079_519, w_079_521, w_079_522, w_079_523, w_079_524, w_079_525, w_079_527, w_079_529, w_079_530, w_079_531, w_079_533, w_079_535, w_079_536, w_079_540, w_079_541, w_079_542, w_079_544, w_079_546, w_079_547, w_079_548, w_079_549, w_079_550, w_079_551, w_079_552, w_079_553, w_079_554, w_079_555, w_079_556, w_079_557, w_079_558, w_079_559, w_079_560, w_079_561, w_079_567, w_079_569, w_079_570, w_079_572, w_079_576, w_079_577, w_079_578, w_079_579, w_079_580, w_079_586, w_079_587, w_079_590, w_079_591, w_079_593, w_079_594, w_079_595, w_079_596, w_079_597, w_079_600, w_079_602, w_079_603, w_079_607, w_079_608, w_079_609, w_079_611, w_079_615, w_079_616, w_079_617, w_079_621, w_079_622, w_079_628, w_079_629, w_079_631, w_079_632, w_079_635, w_079_636, w_079_638, w_079_640, w_079_642, w_079_644, w_079_645, w_079_646, w_079_648, w_079_649, w_079_651, w_079_652, w_079_653, w_079_655, w_079_657, w_079_658, w_079_659, w_079_661, w_079_662, w_079_663, w_079_665, w_079_666, w_079_668, w_079_669, w_079_670, w_079_671, w_079_672, w_079_673, w_079_674, w_079_675, w_079_677, w_079_678, w_079_679, w_079_680, w_079_681, w_079_682, w_079_683, w_079_684, w_079_685, w_079_686, w_079_687, w_079_690, w_079_691, w_079_692, w_079_693, w_079_694, w_079_697, w_079_698, w_079_700, w_079_701, w_079_702, w_079_704, w_079_706, w_079_707, w_079_708, w_079_712, w_079_714, w_079_715, w_079_717, w_079_718, w_079_719, w_079_720, w_079_721, w_079_722, w_079_723, w_079_724, w_079_725, w_079_726, w_079_727, w_079_730, w_079_734, w_079_737, w_079_739, w_079_741, w_079_742, w_079_743, w_079_744, w_079_745, w_079_749, w_079_750, w_079_752, w_079_753, w_079_755, w_079_756, w_079_757, w_079_763, w_079_764, w_079_765, w_079_766, w_079_767, w_079_768, w_079_770, w_079_771, w_079_772, w_079_773, w_079_774, w_079_775, w_079_776, w_079_778, w_079_780, w_079_781, w_079_783, w_079_784, w_079_787, w_079_791, w_079_792, w_079_794, w_079_797, w_079_798, w_079_800, w_079_801, w_079_803, w_079_804, w_079_805, w_079_807, w_079_808, w_079_809, w_079_810, w_079_817, w_079_818, w_079_819, w_079_820, w_079_822, w_079_823, w_079_825, w_079_828, w_079_831, w_079_832, w_079_833, w_079_834, w_079_835, w_079_836, w_079_838, w_079_839, w_079_843, w_079_844, w_079_845, w_079_847, w_079_851, w_079_852, w_079_853, w_079_854, w_079_855, w_079_856, w_079_857, w_079_861, w_079_862, w_079_863, w_079_864, w_079_865, w_079_866, w_079_868, w_079_870, w_079_871, w_079_872, w_079_873, w_079_874, w_079_875, w_079_877, w_079_880, w_079_881, w_079_883, w_079_884, w_079_885, w_079_889, w_079_890, w_079_895, w_079_896, w_079_897, w_079_898, w_079_901, w_079_902, w_079_904, w_079_905, w_079_907, w_079_911, w_079_912, w_079_913, w_079_914, w_079_915, w_079_916, w_079_920, w_079_921, w_079_922, w_079_923, w_079_925, w_079_926, w_079_927, w_079_928, w_079_929, w_079_932, w_079_933, w_079_935, w_079_936, w_079_937, w_079_938, w_079_940, w_079_943, w_079_946, w_079_949, w_079_950, w_079_951, w_079_953, w_079_955, w_079_956, w_079_957, w_079_958, w_079_960, w_079_962, w_079_963, w_079_967, w_079_970, w_079_971, w_079_972, w_079_974, w_079_975, w_079_976, w_079_978, w_079_979, w_079_980, w_079_981, w_079_983, w_079_984, w_079_985, w_079_986, w_079_987, w_079_988, w_079_990, w_079_991, w_079_992, w_079_993, w_079_994, w_079_996, w_079_997, w_079_998, w_079_1000, w_079_1002, w_079_1003, w_079_1005, w_079_1006, w_079_1007, w_079_1009, w_079_1010, w_079_1011, w_079_1012, w_079_1015, w_079_1017, w_079_1024, w_079_1025, w_079_1026, w_079_1027, w_079_1028, w_079_1030, w_079_1034, w_079_1035, w_079_1039, w_079_1042, w_079_1043, w_079_1045, w_079_1050, w_079_1051, w_079_1055, w_079_1057, w_079_1059, w_079_1060, w_079_1064, w_079_1065, w_079_1066, w_079_1073, w_079_1077, w_079_1078, w_079_1081, w_079_1082, w_079_1083, w_079_1088, w_079_1089, w_079_1090, w_079_1091, w_079_1092, w_079_1094, w_079_1095, w_079_1100, w_079_1109, w_079_1111, w_079_1114, w_079_1116, w_079_1121, w_079_1123, w_079_1124, w_079_1127, w_079_1128, w_079_1129, w_079_1132, w_079_1133, w_079_1137, w_079_1139, w_079_1140, w_079_1142, w_079_1148, w_079_1149, w_079_1150, w_079_1155, w_079_1156, w_079_1161, w_079_1166, w_079_1168, w_079_1170, w_079_1171, w_079_1172, w_079_1173, w_079_1174, w_079_1176, w_079_1179, w_079_1180, w_079_1182, w_079_1184, w_079_1185, w_079_1187, w_079_1189, w_079_1191, w_079_1193, w_079_1195, w_079_1196, w_079_1197, w_079_1202, w_079_1203, w_079_1210, w_079_1212, w_079_1217, w_079_1219, w_079_1220, w_079_1221, w_079_1222, w_079_1225, w_079_1226, w_079_1229, w_079_1230, w_079_1231, w_079_1232, w_079_1233, w_079_1236, w_079_1237, w_079_1239, w_079_1240, w_079_1241, w_079_1243, w_079_1246, w_079_1247, w_079_1250, w_079_1251, w_079_1252, w_079_1254, w_079_1255, w_079_1257, w_079_1258, w_079_1259, w_079_1261, w_079_1268, w_079_1275, w_079_1277, w_079_1281, w_079_1283, w_079_1285, w_079_1286, w_079_1288, w_079_1289, w_079_1290, w_079_1291, w_079_1292, w_079_1293, w_079_1297, w_079_1298, w_079_1301, w_079_1303, w_079_1304, w_079_1306, w_079_1307, w_079_1308, w_079_1309, w_079_1311, w_079_1316, w_079_1318, w_079_1319, w_079_1321, w_079_1325, w_079_1326, w_079_1327, w_079_1331, w_079_1334, w_079_1338, w_079_1341, w_079_1343, w_079_1344, w_079_1345, w_079_1348, w_079_1349, w_079_1350, w_079_1354, w_079_1355, w_079_1357, w_079_1358, w_079_1364, w_079_1365, w_079_1368, w_079_1369, w_079_1371, w_079_1374, w_079_1377, w_079_1380, w_079_1381, w_079_1382, w_079_1385, w_079_1387, w_079_1388, w_079_1389, w_079_1391, w_079_1392, w_079_1393, w_079_1394, w_079_1395, w_079_1397, w_079_1399, w_079_1401, w_079_1403, w_079_1406, w_079_1407, w_079_1408, w_079_1409, w_079_1411, w_079_1413, w_079_1414, w_079_1419, w_079_1420, w_079_1422, w_079_1423, w_079_1424, w_079_1425, w_079_1426, w_079_1427, w_079_1429, w_079_1432, w_079_1433, w_079_1435, w_079_1436, w_079_1441, w_079_1443, w_079_1445, w_079_1447, w_079_1448, w_079_1450, w_079_1451, w_079_1454, w_079_1457, w_079_1458, w_079_1459, w_079_1460, w_079_1465, w_079_1466, w_079_1467, w_079_1468, w_079_1469, w_079_1471, w_079_1472, w_079_1474, w_079_1477, w_079_1480, w_079_1483, w_079_1484, w_079_1485, w_079_1487, w_079_1488, w_079_1492, w_079_1493, w_079_1494, w_079_1495, w_079_1496, w_079_1497, w_079_1498, w_079_1500, w_079_1505, w_079_1508, w_079_1509, w_079_1510, w_079_1511, w_079_1512, w_079_1513, w_079_1516, w_079_1517, w_079_1519, w_079_1520, w_079_1522, w_079_1524, w_079_1525, w_079_1526, w_079_1527, w_079_1528, w_079_1531, w_079_1533, w_079_1534, w_079_1540, w_079_1541, w_079_1543, w_079_1546, w_079_1547, w_079_1549, w_079_1552, w_079_1554, w_079_1555, w_079_1557, w_079_1559, w_079_1562, w_079_1564, w_079_1567, w_079_1568, w_079_1569, w_079_1570, w_079_1572, w_079_1573, w_079_1576, w_079_1578, w_079_1581, w_079_1583, w_079_1587, w_079_1589, w_079_1591, w_079_1597, w_079_1598, w_079_1602, w_079_1603, w_079_1605, w_079_1607, w_079_1608, w_079_1611, w_079_1612, w_079_1613, w_079_1616, w_079_1618, w_079_1623, w_079_1625, w_079_1626, w_079_1628, w_079_1631, w_079_1632, w_079_1633, w_079_1638, w_079_1640, w_079_1643, w_079_1646, w_079_1649, w_079_1651, w_079_1652, w_079_1655, w_079_1656, w_079_1657, w_079_1660, w_079_1663, w_079_1664, w_079_1665, w_079_1667, w_079_1668, w_079_1669, w_079_1670, w_079_1672, w_079_1675, w_079_1676, w_079_1677, w_079_1681, w_079_1684, w_079_1685, w_079_1686, w_079_1691, w_079_1692, w_079_1694, w_079_1696, w_079_1697, w_079_1698, w_079_1699, w_079_1701, w_079_1705, w_079_1706, w_079_1708, w_079_1710, w_079_1711, w_079_1714, w_079_1716, w_079_1717, w_079_1718, w_079_1720, w_079_1721, w_079_1722, w_079_1724, w_079_1725, w_079_1728, w_079_1730, w_079_1731, w_079_1732, w_079_1733, w_079_1734, w_079_1736, w_079_1739, w_079_1741, w_079_1743, w_079_1748, w_079_1751, w_079_1756, w_079_1757, w_079_1759, w_079_1760, w_079_1761, w_079_1763, w_079_1765, w_079_1766, w_079_1767, w_079_1768, w_079_1769, w_079_1772, w_079_1777, w_079_1779, w_079_1781, w_079_1783, w_079_1787, w_079_1789, w_079_1792, w_079_1794, w_079_1795, w_079_1796, w_079_1797, w_079_1800, w_079_1801, w_079_1802, w_079_1803, w_079_1805, w_079_1807, w_079_1808, w_079_1809, w_079_1810, w_079_1812, w_079_1816, w_079_1820, w_079_1821, w_079_1822, w_079_1824, w_079_1826, w_079_1827, w_079_1831, w_079_1833, w_079_1835, w_079_1837, w_079_1839, w_079_1841, w_079_1842, w_079_1843, w_079_1848, w_079_1850, w_079_1851, w_079_1854, w_079_1858, w_079_1860, w_079_1861, w_079_1863, w_079_1867, w_079_1868, w_079_1871, w_079_1873, w_079_1874, w_079_1875, w_079_1876, w_079_1878, w_079_1881, w_079_1883, w_079_1885, w_079_1886, w_079_1888, w_079_1891, w_079_1892, w_079_1893, w_079_1894, w_079_1898, w_079_1899, w_079_1900, w_079_1905, w_079_1906, w_079_1908, w_079_1910, w_079_1911, w_079_1914, w_079_1915, w_079_1916, w_079_1919, w_079_1921, w_079_1923, w_079_1927, w_079_1931, w_079_1934, w_079_1935, w_079_1938, w_079_1941, w_079_1946, w_079_1948, w_079_1950, w_079_1951, w_079_1954, w_079_1957, w_079_1958, w_079_1961, w_079_1962, w_079_1963, w_079_1966, w_079_1968, w_079_1969, w_079_1970, w_079_1971, w_079_1974, w_079_1975, w_079_1978, w_079_1990, w_079_1996, w_079_1997, w_079_1998, w_079_2000, w_079_2002, w_079_2003, w_079_2004, w_079_2007, w_079_2009, w_079_2013, w_079_2014, w_079_2015, w_079_2016, w_079_2021, w_079_2022, w_079_2023, w_079_2024, w_079_2025, w_079_2026, w_079_2027, w_079_2029, w_079_2033, w_079_2036, w_079_2038, w_079_2039, w_079_2040, w_079_2042, w_079_2043, w_079_2045, w_079_2046, w_079_2047, w_079_2052, w_079_2053, w_079_2054, w_079_2056, w_079_2061, w_079_2063, w_079_2065, w_079_2066, w_079_2069, w_079_2073, w_079_2074, w_079_2075, w_079_2076, w_079_2078, w_079_2081, w_079_2082, w_079_2083, w_079_2084, w_079_2087, w_079_2088, w_079_2089, w_079_2090, w_079_2091, w_079_2092, w_079_2093, w_079_2095, w_079_2099, w_079_2101, w_079_2103, w_079_2104, w_079_2106, w_079_2109, w_079_2111, w_079_2113, w_079_2115, w_079_2118, w_079_2120, w_079_2122, w_079_2123, w_079_2125, w_079_2126, w_079_2131, w_079_2133, w_079_2138, w_079_2139, w_079_2140, w_079_2141, w_079_2142, w_079_2145, w_079_2149, w_079_2150, w_079_2151, w_079_2152, w_079_2154, w_079_2155, w_079_2156, w_079_2158, w_079_2160, w_079_2161, w_079_2163, w_079_2165, w_079_2166, w_079_2167, w_079_2168, w_079_2169, w_079_2173, w_079_2174, w_079_2176, w_079_2177, w_079_2185, w_079_2188, w_079_2190, w_079_2192, w_079_2197, w_079_2198, w_079_2201, w_079_2202, w_079_2204, w_079_2206, w_079_2207, w_079_2210, w_079_2214, w_079_2215, w_079_2217, w_079_2218, w_079_2223, w_079_2225, w_079_2226, w_079_2229, w_079_2233, w_079_2234, w_079_2235, w_079_2238, w_079_2240, w_079_2241, w_079_2242, w_079_2244, w_079_2249, w_079_2252, w_079_2254, w_079_2256, w_079_2257, w_079_2259, w_079_2261, w_079_2264, w_079_2265, w_079_2266, w_079_2269, w_079_2272, w_079_2281, w_079_2282, w_079_2283, w_079_2286, w_079_2287, w_079_2290, w_079_2293, w_079_2294, w_079_2299, w_079_2301, w_079_2302, w_079_2303, w_079_2308, w_079_2309, w_079_2311, w_079_2313, w_079_2315, w_079_2316, w_079_2317, w_079_2320, w_079_2324, w_079_2325, w_079_2326, w_079_2328, w_079_2329, w_079_2331, w_079_2333, w_079_2336, w_079_2337, w_079_2338, w_079_2340, w_079_2343, w_079_2344, w_079_2345, w_079_2346, w_079_2347, w_079_2353, w_079_2354, w_079_2360, w_079_2362, w_079_2366, w_079_2367, w_079_2368, w_079_2371, w_079_2374, w_079_2382, w_079_2383, w_079_2386, w_079_2388, w_079_2390, w_079_2391, w_079_2392, w_079_2393, w_079_2394, w_079_2395, w_079_2399, w_079_2403, w_079_2404, w_079_2405, w_079_2406, w_079_2411, w_079_2412, w_079_2418, w_079_2419, w_079_2421, w_079_2422, w_079_2423, w_079_2424, w_079_2426, w_079_2430, w_079_2431, w_079_2434, w_079_2436, w_079_2439, w_079_2442, w_079_2445, w_079_2448, w_079_2449, w_079_2454, w_079_2459, w_079_2460, w_079_2461, w_079_2462, w_079_2469, w_079_2471, w_079_2472, w_079_2478, w_079_2482, w_079_2483, w_079_2484, w_079_2488, w_079_2489, w_079_2492, w_079_2494, w_079_2495, w_079_2496, w_079_2497, w_079_2499, w_079_2501, w_079_2503, w_079_2504, w_079_2505, w_079_2510, w_079_2512, w_079_2513, w_079_2514, w_079_2515, w_079_2517, w_079_2520, w_079_2521, w_079_2523, w_079_2524, w_079_2525, w_079_2527, w_079_2530, w_079_2531, w_079_2532, w_079_2534, w_079_2537, w_079_2542, w_079_2552, w_079_2555, w_079_2556, w_079_2557, w_079_2559, w_079_2560, w_079_2561, w_079_2562, w_079_2565, w_079_2566, w_079_2567, w_079_2571, w_079_2572, w_079_2574, w_079_2575, w_079_2580, w_079_2582, w_079_2586, w_079_2588, w_079_2589, w_079_2592, w_079_2595, w_079_2596, w_079_2597, w_079_2599, w_079_2601, w_079_2602, w_079_2604, w_079_2605, w_079_2607, w_079_2608, w_079_2609, w_079_2611, w_079_2612, w_079_2618, w_079_2622, w_079_2624, w_079_2627, w_079_2628, w_079_2631, w_079_2632, w_079_2633, w_079_2635, w_079_2636, w_079_2640, w_079_2641, w_079_2642, w_079_2643, w_079_2647, w_079_2648, w_079_2649, w_079_2651, w_079_2652, w_079_2654, w_079_2659, w_079_2662, w_079_2663, w_079_2664, w_079_2665, w_079_2666, w_079_2668, w_079_2670, w_079_2674, w_079_2679, w_079_2682, w_079_2683, w_079_2684, w_079_2685, w_079_2689, w_079_2690, w_079_2691, w_079_2692, w_079_2693, w_079_2697, w_079_2698, w_079_2699, w_079_2700, w_079_2708, w_079_2709, w_079_2710, w_079_2711, w_079_2712, w_079_2713, w_079_2714, w_079_2715, w_079_2720, w_079_2721, w_079_2725, w_079_2726, w_079_2727, w_079_2729, w_079_2730, w_079_2731, w_079_2733, w_079_2734, w_079_2735, w_079_2737, w_079_2738, w_079_2739, w_079_2740, w_079_2743, w_079_2746, w_079_2750, w_079_2752, w_079_2753, w_079_2755, w_079_2756, w_079_2757, w_079_2760, w_079_2761, w_079_2763, w_079_2764, w_079_2767, w_079_2769, w_079_2773, w_079_2775, w_079_2776, w_079_2777, w_079_2779, w_079_2781, w_079_2783, w_079_2789, w_079_2791, w_079_2792, w_079_2793, w_079_2795, w_079_2797, w_079_2800, w_079_2801, w_079_2802, w_079_2803, w_079_2804, w_079_2806, w_079_2809, w_079_2810, w_079_2813, w_079_2815, w_079_2816, w_079_2818, w_079_2824, w_079_2827, w_079_2832, w_079_2833, w_079_2834, w_079_2837, w_079_2838, w_079_2839, w_079_2840, w_079_2842, w_079_2848, w_079_2855, w_079_2856, w_079_2858, w_079_2862, w_079_2864, w_079_2866, w_079_2868, w_079_2870, w_079_2871, w_079_2872, w_079_2874, w_079_2879, w_079_2880, w_079_2882, w_079_2883, w_079_2884, w_079_2887, w_079_2888, w_079_2890, w_079_2891, w_079_2892, w_079_2893, w_079_2897, w_079_2899, w_079_2903, w_079_2904, w_079_2905, w_079_2906, w_079_2907, w_079_2910, w_079_2911, w_079_2913, w_079_2917, w_079_2919, w_079_2920, w_079_2926, w_079_2928, w_079_2932, w_079_2933, w_079_2936, w_079_2938, w_079_2939, w_079_2941, w_079_2946, w_079_2949, w_079_2950, w_079_2951, w_079_2956, w_079_2958, w_079_2961, w_079_2963, w_079_2966, w_079_2968, w_079_2970, w_079_2971, w_079_2972, w_079_2973, w_079_2975, w_079_2981, w_079_2983, w_079_2986, w_079_2988, w_079_2995, w_079_2998, w_079_2999, w_079_3005, w_079_3010, w_079_3011, w_079_3013, w_079_3015, w_079_3018, w_079_3019, w_079_3020, w_079_3021, w_079_3022, w_079_3023, w_079_3024, w_079_3026, w_079_3027, w_079_3028, w_079_3029, w_079_3031, w_079_3034, w_079_3035, w_079_3040, w_079_3042, w_079_3044, w_079_3045, w_079_3050, w_079_3052, w_079_3053, w_079_3054, w_079_3057, w_079_3061, w_079_3062, w_079_3065, w_079_3068, w_079_3076, w_079_3078, w_079_3079, w_079_3080, w_079_3083, w_079_3087, w_079_3091, w_079_3092, w_079_3093, w_079_3094, w_079_3095, w_079_3097, w_079_3102, w_079_3104, w_079_3106, w_079_3107, w_079_3110, w_079_3112, w_079_3114, w_079_3117, w_079_3118, w_079_3123, w_079_3124, w_079_3125, w_079_3129, w_079_3130, w_079_3133, w_079_3136, w_079_3138, w_079_3140, w_079_3141, w_079_3143, w_079_3144, w_079_3145, w_079_3146, w_079_3147, w_079_3148, w_079_3154, w_079_3156, w_079_3158, w_079_3159, w_079_3160, w_079_3162, w_079_3164, w_079_3166, w_079_3168, w_079_3173, w_079_3175, w_079_3177, w_079_3178, w_079_3179, w_079_3181, w_079_3182, w_079_3185, w_079_3189, w_079_3190, w_079_3192, w_079_3194, w_079_3196, w_079_3198, w_079_3199, w_079_3200, w_079_3202, w_079_3203, w_079_3207, w_079_3209, w_079_3210, w_079_3213, w_079_3214, w_079_3221, w_079_3224, w_079_3227, w_079_3228, w_079_3230, w_079_3231, w_079_3232, w_079_3233, w_079_3234, w_079_3236, w_079_3238, w_079_3239, w_079_3240, w_079_3244, w_079_3245, w_079_3248, w_079_3250, w_079_3252, w_079_3256, w_079_3257, w_079_3259, w_079_3260, w_079_3263, w_079_3268, w_079_3269, w_079_3270, w_079_3274, w_079_3279, w_079_3285, w_079_3288, w_079_3295, w_079_3299, w_079_3300, w_079_3303, w_079_3304, w_079_3307, w_079_3310, w_079_3312, w_079_3313, w_079_3314, w_079_3315, w_079_3316, w_079_3321, w_079_3325, w_079_3328, w_079_3333, w_079_3334, w_079_3335, w_079_3336, w_079_3337, w_079_3339, w_079_3341, w_079_3342, w_079_3344, w_079_3347, w_079_3348, w_079_3349, w_079_3355, w_079_3356, w_079_3359, w_079_3364, w_079_3366, w_079_3368, w_079_3370, w_079_3371, w_079_3372, w_079_3373, w_079_3374, w_079_3376, w_079_3377, w_079_3378, w_079_3386, w_079_3387, w_079_3388, w_079_3389, w_079_3390, w_079_3392, w_079_3395, w_079_3397, w_079_3398, w_079_3399, w_079_3405, w_079_3407, w_079_3408, w_079_3410, w_079_3411, w_079_3415, w_079_3416, w_079_3417, w_079_3420, w_079_3421, w_079_3422, w_079_3424, w_079_3425, w_079_3428, w_079_3429, w_079_3435, w_079_3440, w_079_3441, w_079_3442, w_079_3444, w_079_3445, w_079_3447, w_079_3449, w_079_3450, w_079_3451, w_079_3455, w_079_3457, w_079_3458, w_079_3459, w_079_3460, w_079_3461, w_079_3462, w_079_3465, w_079_3467, w_079_3469, w_079_3470, w_079_3471, w_079_3476, w_079_3479, w_079_3483, w_079_3484, w_079_3485, w_079_3486, w_079_3490, w_079_3492, w_079_3494, w_079_3495, w_079_3496, w_079_3498, w_079_3505, w_079_3506, w_079_3509, w_079_3510, w_079_3512, w_079_3514, w_079_3515, w_079_3517, w_079_3518, w_079_3519, w_079_3520, w_079_3521, w_079_3522, w_079_3523, w_079_3524, w_079_3527, w_079_3530, w_079_3531, w_079_3532, w_079_3533, w_079_3534, w_079_3539, w_079_3542, w_079_3544, w_079_3550, w_079_3553, w_079_3554, w_079_3557, w_079_3559, w_079_3561, w_079_3564, w_079_3566, w_079_3567, w_079_3570, w_079_3571, w_079_3574, w_079_3575, w_079_3577, w_079_3579, w_079_3581, w_079_3586, w_079_3589, w_079_3590, w_079_3592, w_079_3593, w_079_3594, w_079_3595, w_079_3599, w_079_3600, w_079_3602, w_079_3603, w_079_3605, w_079_3608, w_079_3610, w_079_3611, w_079_3612, w_079_3614, w_079_3616, w_079_3619, w_079_3620, w_079_3624, w_079_3626, w_079_3628, w_079_3629, w_079_3631, w_079_3632, w_079_3633, w_079_3634, w_079_3637, w_079_3639, w_079_3640, w_079_3645, w_079_3647, w_079_3648, w_079_3650, w_079_3652, w_079_3653, w_079_3656, w_079_3657, w_079_3658, w_079_3659, w_079_3664, w_079_3666, w_079_3668, w_079_3671, w_079_3674, w_079_3677, w_079_3679, w_079_3683, w_079_3684, w_079_3685, w_079_3686, w_079_3688, w_079_3690, w_079_3693, w_079_3695, w_079_3697, w_079_3698, w_079_3699, w_079_3700, w_079_3703, w_079_3704, w_079_3705, w_079_3706, w_079_3707, w_079_3711, w_079_3716, w_079_3720, w_079_3723, w_079_3725, w_079_3732, w_079_3736, w_079_3738, w_079_3740, w_079_3741, w_079_3746, w_079_3748, w_079_3750, w_079_3752, w_079_3758, w_079_3760, w_079_3763, w_079_3765, w_079_3766, w_079_3767, w_079_3768, w_079_3769, w_079_3771, w_079_3775, w_079_3776, w_079_3777, w_079_3779, w_079_3781, w_079_3784, w_079_3785, w_079_3790, w_079_3791, w_079_3792, w_079_3794, w_079_3797, w_079_3798, w_079_3799, w_079_3800, w_079_3801, w_079_3803, w_079_3804, w_079_3806, w_079_3808, w_079_3810, w_079_3811, w_079_3812, w_079_3813, w_079_3817, w_079_3819, w_079_3820, w_079_3822, w_079_3823, w_079_3824, w_079_3825, w_079_3826, w_079_3827, w_079_3829, w_079_3832, w_079_3834, w_079_3836, w_079_3839, w_079_3840, w_079_3841, w_079_3844, w_079_3845, w_079_3850, w_079_3851, w_079_3855, w_079_3856, w_079_3857, w_079_3859, w_079_3861, w_079_3863, w_079_3864, w_079_3870, w_079_3871, w_079_3872, w_079_3873, w_079_3874, w_079_3875, w_079_3876, w_079_3878, w_079_3880, w_079_3882, w_079_3884, w_079_3885, w_079_3886, w_079_3887, w_079_3888, w_079_3889, w_079_3894, w_079_3897, w_079_3901, w_079_3903, w_079_3905, w_079_3908, w_079_3915, w_079_3919, w_079_3922, w_079_3923, w_079_3924, w_079_3925, w_079_3928, w_079_3932, w_079_3933, w_079_3934, w_079_3935, w_079_3936, w_079_3938, w_079_3941, w_079_3943, w_079_3944, w_079_3947, w_079_3953, w_079_3954, w_079_3955, w_079_3957, w_079_3959, w_079_3961, w_079_3962, w_079_3966, w_079_3967, w_079_3968, w_079_3969, w_079_3972, w_079_3973, w_079_3974, w_079_3975, w_079_3976, w_079_3978, w_079_3983, w_079_3984, w_079_3986, w_079_3987, w_079_3989, w_079_3990, w_079_3992, w_079_3993, w_079_3994, w_079_3995, w_079_3997, w_079_3998, w_079_3999, w_079_4000, w_079_4001, w_079_4002, w_079_4003, w_079_4004, w_079_4006, w_079_4010, w_079_4011, w_079_4012, w_079_4013, w_079_4015, w_079_4018, w_079_4022, w_079_4025, w_079_4026, w_079_4030, w_079_4032, w_079_4034, w_079_4035, w_079_4036, w_079_4038, w_079_4039, w_079_4040, w_079_4042, w_079_4049, w_079_4052, w_079_4053, w_079_4058, w_079_4062, w_079_4064, w_079_4066, w_079_4068, w_079_4069, w_079_4070, w_079_4071, w_079_4072, w_079_4082, w_079_4083, w_079_4084, w_079_4085, w_079_4086, w_079_4087, w_079_4088, w_079_4089, w_079_4090, w_079_4091, w_079_4093, w_079_4097, w_079_4099, w_079_4102, w_079_4104, w_079_4107, w_079_4108, w_079_4112, w_079_4114, w_079_4115, w_079_4117, w_079_4118, w_079_4119, w_079_4122, w_079_4124, w_079_4126, w_079_4127, w_079_4128, w_079_4130, w_079_4134, w_079_4138, w_079_4139, w_079_4141, w_079_4143, w_079_4144, w_079_4147, w_079_4149, w_079_4151, w_079_4153, w_079_4156, w_079_4157, w_079_4160, w_079_4161, w_079_4162, w_079_4171, w_079_4172, w_079_4174, w_079_4175, w_079_4180, w_079_4181, w_079_4182, w_079_4183, w_079_4184, w_079_4191, w_079_4194, w_079_4197, w_079_4198, w_079_4199, w_079_4202, w_079_4208, w_079_4210, w_079_4214, w_079_4216, w_079_4218, w_079_4220, w_079_4222, w_079_4229, w_079_4233, w_079_4236, w_079_4237, w_079_4241, w_079_4243, w_079_4244, w_079_4245, w_079_4247, w_079_4248, w_079_4249, w_079_4251, w_079_4253, w_079_4254, w_079_4258, w_079_4262, w_079_4263, w_079_4265, w_079_4268, w_079_4269, w_079_4270, w_079_4271, w_079_4272, w_079_4273, w_079_4274, w_079_4279, w_079_4280, w_079_4282, w_079_4284, w_079_4285, w_079_4286, w_079_4287, w_079_4288, w_079_4290, w_079_4292, w_079_4294, w_079_4298, w_079_4299, w_079_4300, w_079_4302, w_079_4303, w_079_4304, w_079_4316, w_079_4318, w_079_4320, w_079_4322, w_079_4324, w_079_4328, w_079_4329, w_079_4333, w_079_4335, w_079_4336, w_079_4339, w_079_4341, w_079_4342, w_079_4346, w_079_4347, w_079_4350, w_079_4351, w_079_4355, w_079_4361, w_079_4363, w_079_4364, w_079_4366, w_079_4367, w_079_4368, w_079_4370, w_079_4372, w_079_4373, w_079_4374, w_079_4375, w_079_4376, w_079_4377, w_079_4381, w_079_4382, w_079_4383, w_079_4384, w_079_4385, w_079_4386, w_079_4387, w_079_4389, w_079_4391, w_079_4392, w_079_4396, w_079_4398, w_079_4400, w_079_4401, w_079_4404, w_079_4409, w_079_4413, w_079_4415, w_079_4417, w_079_4418, w_079_4424, w_079_4425, w_079_4426, w_079_4428, w_079_4429, w_079_4431, w_079_4432, w_079_4435, w_079_4437, w_079_4438, w_079_4440, w_079_4441, w_079_4443, w_079_4444, w_079_4445, w_079_4447, w_079_4450, w_079_4451, w_079_4452, w_079_4453, w_079_4454, w_079_4455, w_079_4456, w_079_4457, w_079_4459, w_079_4460, w_079_4464, w_079_4467, w_079_4470, w_079_4472, w_079_4474, w_079_4475, w_079_4477, w_079_4479, w_079_4483, w_079_4485, w_079_4486, w_079_4487;
  wire w_080_003, w_080_004, w_080_006, w_080_008, w_080_013, w_080_017, w_080_020, w_080_021, w_080_023, w_080_025, w_080_027, w_080_028, w_080_029, w_080_031, w_080_032, w_080_034, w_080_035, w_080_038, w_080_042, w_080_043, w_080_046, w_080_047, w_080_048, w_080_050, w_080_055, w_080_057, w_080_058, w_080_061, w_080_062, w_080_065, w_080_066, w_080_069, w_080_071, w_080_076, w_080_077, w_080_078, w_080_079, w_080_081, w_080_082, w_080_084, w_080_085, w_080_086, w_080_088, w_080_089, w_080_090, w_080_091, w_080_093, w_080_094, w_080_097, w_080_099, w_080_101, w_080_103, w_080_105, w_080_106, w_080_107, w_080_108, w_080_111, w_080_112, w_080_114, w_080_119, w_080_120, w_080_122, w_080_124, w_080_126, w_080_130, w_080_131, w_080_132, w_080_134, w_080_136, w_080_137, w_080_138, w_080_140, w_080_141, w_080_143, w_080_145, w_080_147, w_080_149, w_080_152, w_080_154, w_080_155, w_080_157, w_080_159, w_080_162, w_080_163, w_080_165, w_080_166, w_080_168, w_080_169, w_080_174, w_080_175, w_080_177, w_080_179, w_080_181, w_080_185, w_080_187, w_080_188, w_080_189, w_080_193, w_080_195, w_080_197, w_080_198, w_080_204, w_080_208, w_080_209, w_080_210, w_080_211, w_080_212, w_080_217, w_080_219, w_080_220, w_080_221, w_080_222, w_080_224, w_080_227, w_080_228, w_080_230, w_080_236, w_080_239, w_080_241, w_080_243, w_080_245, w_080_250, w_080_251, w_080_252, w_080_254, w_080_256, w_080_259, w_080_261, w_080_265, w_080_266, w_080_268, w_080_270, w_080_272, w_080_276, w_080_277, w_080_278, w_080_281, w_080_282, w_080_285, w_080_289, w_080_294, w_080_296, w_080_298, w_080_300, w_080_301, w_080_302, w_080_305, w_080_306, w_080_308, w_080_311, w_080_312, w_080_314, w_080_317, w_080_319, w_080_322, w_080_323, w_080_327, w_080_329, w_080_330, w_080_337, w_080_340, w_080_342, w_080_344, w_080_345, w_080_349, w_080_350, w_080_351, w_080_352, w_080_353, w_080_355, w_080_357, w_080_359, w_080_365, w_080_367, w_080_368, w_080_373, w_080_375, w_080_377, w_080_378, w_080_380, w_080_381, w_080_382, w_080_383, w_080_384, w_080_387, w_080_389, w_080_392, w_080_393, w_080_397, w_080_399, w_080_401, w_080_402, w_080_405, w_080_407, w_080_409, w_080_411, w_080_412, w_080_417, w_080_418, w_080_420, w_080_422, w_080_425, w_080_426, w_080_427, w_080_429, w_080_431, w_080_436, w_080_438, w_080_439, w_080_441, w_080_442, w_080_443, w_080_444, w_080_445, w_080_449, w_080_451, w_080_452, w_080_454, w_080_458, w_080_461, w_080_462, w_080_463, w_080_466, w_080_467, w_080_468, w_080_469, w_080_472, w_080_473, w_080_475, w_080_478, w_080_480, w_080_481, w_080_482, w_080_484, w_080_485, w_080_486, w_080_487, w_080_489, w_080_490, w_080_493, w_080_495, w_080_497, w_080_499, w_080_501, w_080_503, w_080_504, w_080_509, w_080_511, w_080_515, w_080_516, w_080_520, w_080_522, w_080_527, w_080_528, w_080_534, w_080_535, w_080_537, w_080_540, w_080_543, w_080_544, w_080_546, w_080_547, w_080_548, w_080_551, w_080_552, w_080_560, w_080_564, w_080_565, w_080_570, w_080_573, w_080_574, w_080_576, w_080_578, w_080_580, w_080_583, w_080_584, w_080_585, w_080_586, w_080_592, w_080_593, w_080_594, w_080_597, w_080_599, w_080_601, w_080_605, w_080_607, w_080_609, w_080_610, w_080_612, w_080_614, w_080_615, w_080_617, w_080_620, w_080_627, w_080_630, w_080_632, w_080_635, w_080_636, w_080_637, w_080_640, w_080_650, w_080_651, w_080_654, w_080_655, w_080_658, w_080_660, w_080_662, w_080_663, w_080_665, w_080_666, w_080_667, w_080_668, w_080_670, w_080_673, w_080_674, w_080_675, w_080_676, w_080_678, w_080_679, w_080_681, w_080_682, w_080_684, w_080_687, w_080_688, w_080_689, w_080_691, w_080_692, w_080_693, w_080_695, w_080_696, w_080_697, w_080_701, w_080_709, w_080_711, w_080_712, w_080_713, w_080_714, w_080_716, w_080_719, w_080_722, w_080_726, w_080_727, w_080_728, w_080_729, w_080_732, w_080_735, w_080_736, w_080_738, w_080_740, w_080_741, w_080_744, w_080_746, w_080_747, w_080_748, w_080_751, w_080_753, w_080_755, w_080_757, w_080_758, w_080_759, w_080_760, w_080_764, w_080_765, w_080_766, w_080_769, w_080_772, w_080_775, w_080_778, w_080_785, w_080_787, w_080_789, w_080_790, w_080_792, w_080_794, w_080_795, w_080_796, w_080_797, w_080_800, w_080_802, w_080_804, w_080_807, w_080_809, w_080_810, w_080_811, w_080_813, w_080_814, w_080_822, w_080_824, w_080_825, w_080_827, w_080_832, w_080_834, w_080_836, w_080_842, w_080_843, w_080_846, w_080_847, w_080_848, w_080_849, w_080_850, w_080_851, w_080_852, w_080_856, w_080_858, w_080_860, w_080_862, w_080_865, w_080_866, w_080_867, w_080_870, w_080_874, w_080_875, w_080_877, w_080_878, w_080_881, w_080_886, w_080_888, w_080_889, w_080_890, w_080_891, w_080_895, w_080_899, w_080_900, w_080_902, w_080_905, w_080_908, w_080_911, w_080_912, w_080_914, w_080_915, w_080_918, w_080_920, w_080_921, w_080_926, w_080_929, w_080_932, w_080_933, w_080_936, w_080_938, w_080_940, w_080_941, w_080_949, w_080_950, w_080_951, w_080_953, w_080_954, w_080_960, w_080_963, w_080_965, w_080_966, w_080_971, w_080_972, w_080_973, w_080_974, w_080_975, w_080_977, w_080_980, w_080_982, w_080_983, w_080_984, w_080_985, w_080_986, w_080_991, w_080_996, w_080_997, w_080_1000, w_080_1001, w_080_1003, w_080_1007, w_080_1008, w_080_1010, w_080_1012, w_080_1013, w_080_1015, w_080_1018, w_080_1019, w_080_1021, w_080_1023, w_080_1026, w_080_1028, w_080_1031, w_080_1033, w_080_1034, w_080_1039, w_080_1042, w_080_1043, w_080_1044, w_080_1045, w_080_1047, w_080_1048, w_080_1054, w_080_1055, w_080_1058, w_080_1061, w_080_1066, w_080_1067, w_080_1069, w_080_1071, w_080_1073, w_080_1074, w_080_1075, w_080_1076, w_080_1078, w_080_1079, w_080_1081, w_080_1082, w_080_1083, w_080_1084, w_080_1085, w_080_1086, w_080_1087, w_080_1088, w_080_1094, w_080_1095, w_080_1097, w_080_1098, w_080_1100, w_080_1101, w_080_1103, w_080_1104, w_080_1105, w_080_1107, w_080_1108, w_080_1109, w_080_1112, w_080_1118, w_080_1119, w_080_1127, w_080_1129, w_080_1131, w_080_1133, w_080_1134, w_080_1135, w_080_1139, w_080_1140, w_080_1141, w_080_1142, w_080_1144, w_080_1148, w_080_1149, w_080_1152, w_080_1153, w_080_1154, w_080_1155, w_080_1156, w_080_1158, w_080_1159, w_080_1160, w_080_1161, w_080_1166, w_080_1175, w_080_1179, w_080_1181, w_080_1187, w_080_1188, w_080_1189, w_080_1190, w_080_1192, w_080_1194, w_080_1197, w_080_1198, w_080_1202, w_080_1204, w_080_1205, w_080_1208, w_080_1210, w_080_1212, w_080_1215, w_080_1216, w_080_1217, w_080_1218, w_080_1220, w_080_1221, w_080_1222, w_080_1224, w_080_1225, w_080_1229, w_080_1231, w_080_1235, w_080_1236, w_080_1237, w_080_1238, w_080_1240, w_080_1241, w_080_1242, w_080_1243, w_080_1245, w_080_1246, w_080_1248, w_080_1249, w_080_1250, w_080_1252, w_080_1254, w_080_1258, w_080_1261, w_080_1263, w_080_1267, w_080_1268, w_080_1270, w_080_1271, w_080_1273, w_080_1275, w_080_1276, w_080_1277, w_080_1278, w_080_1279, w_080_1280, w_080_1283, w_080_1285, w_080_1286, w_080_1290, w_080_1292, w_080_1293, w_080_1294, w_080_1298, w_080_1301, w_080_1302, w_080_1303, w_080_1308, w_080_1310, w_080_1311, w_080_1312, w_080_1314, w_080_1315, w_080_1316, w_080_1319, w_080_1321, w_080_1323, w_080_1326, w_080_1327, w_080_1328, w_080_1330, w_080_1332, w_080_1333, w_080_1336, w_080_1337, w_080_1338, w_080_1339, w_080_1342, w_080_1343, w_080_1346, w_080_1347, w_080_1348, w_080_1349, w_080_1350, w_080_1353, w_080_1354, w_080_1356, w_080_1357, w_080_1360, w_080_1361, w_080_1365, w_080_1367, w_080_1368, w_080_1369, w_080_1370, w_080_1373, w_080_1375, w_080_1376, w_080_1378, w_080_1382, w_080_1384, w_080_1386, w_080_1394, w_080_1398, w_080_1399, w_080_1401, w_080_1402, w_080_1405, w_080_1406, w_080_1408, w_080_1409, w_080_1411, w_080_1413, w_080_1414, w_080_1415, w_080_1419, w_080_1420, w_080_1424, w_080_1429, w_080_1430, w_080_1431, w_080_1432, w_080_1434, w_080_1435, w_080_1437, w_080_1438, w_080_1439, w_080_1440, w_080_1442, w_080_1443, w_080_1446, w_080_1448, w_080_1449, w_080_1450, w_080_1453, w_080_1454, w_080_1456, w_080_1459, w_080_1461, w_080_1466, w_080_1467, w_080_1470, w_080_1476, w_080_1478, w_080_1480, w_080_1482, w_080_1483, w_080_1490, w_080_1492, w_080_1497, w_080_1498, w_080_1499, w_080_1500, w_080_1502, w_080_1503, w_080_1504, w_080_1508, w_080_1509, w_080_1514, w_080_1517, w_080_1518, w_080_1520, w_080_1522, w_080_1524, w_080_1525, w_080_1526, w_080_1528, w_080_1531, w_080_1533, w_080_1534, w_080_1535, w_080_1539, w_080_1541, w_080_1545, w_080_1548, w_080_1551, w_080_1552, w_080_1555, w_080_1556, w_080_1560, w_080_1563, w_080_1564, w_080_1566, w_080_1567, w_080_1568, w_080_1569, w_080_1570, w_080_1571, w_080_1576, w_080_1578, w_080_1580, w_080_1582, w_080_1583, w_080_1584, w_080_1585, w_080_1591, w_080_1595, w_080_1598, w_080_1599, w_080_1601, w_080_1602, w_080_1604, w_080_1605, w_080_1607, w_080_1611, w_080_1612, w_080_1614, w_080_1615, w_080_1617, w_080_1619, w_080_1620, w_080_1625, w_080_1626, w_080_1630, w_080_1632, w_080_1635, w_080_1643, w_080_1644, w_080_1645, w_080_1646, w_080_1648, w_080_1652, w_080_1657, w_080_1658, w_080_1663, w_080_1664, w_080_1667, w_080_1668, w_080_1669, w_080_1672, w_080_1675, w_080_1676, w_080_1677, w_080_1678, w_080_1681, w_080_1683, w_080_1684, w_080_1685, w_080_1686, w_080_1689, w_080_1690, w_080_1691, w_080_1692, w_080_1695, w_080_1698, w_080_1701, w_080_1702, w_080_1705, w_080_1707, w_080_1709, w_080_1711, w_080_1712, w_080_1713, w_080_1715, w_080_1720, w_080_1721, w_080_1727, w_080_1729, w_080_1730, w_080_1731, w_080_1733, w_080_1735, w_080_1738, w_080_1740, w_080_1743, w_080_1744, w_080_1745, w_080_1746, w_080_1749, w_080_1752, w_080_1754, w_080_1756, w_080_1757, w_080_1758, w_080_1765, w_080_1766, w_080_1767, w_080_1770, w_080_1771, w_080_1774, w_080_1775, w_080_1777, w_080_1778, w_080_1779, w_080_1780, w_080_1781, w_080_1782, w_080_1785, w_080_1786, w_080_1787, w_080_1790, w_080_1791, w_080_1792, w_080_1794, w_080_1796, w_080_1798, w_080_1799, w_080_1802, w_080_1806, w_080_1807, w_080_1810, w_080_1811, w_080_1815, w_080_1817, w_080_1818, w_080_1820, w_080_1821, w_080_1822, w_080_1823, w_080_1824, w_080_1825, w_080_1826, w_080_1828, w_080_1832, w_080_1833, w_080_1834, w_080_1836, w_080_1841, w_080_1842, w_080_1843, w_080_1844, w_080_1850, w_080_1852, w_080_1860, w_080_1861, w_080_1862, w_080_1863, w_080_1864, w_080_1865, w_080_1867, w_080_1868, w_080_1871, w_080_1873, w_080_1875, w_080_1877, w_080_1878, w_080_1881, w_080_1887, w_080_1888, w_080_1892, w_080_1897, w_080_1898, w_080_1899, w_080_1900, w_080_1903, w_080_1912, w_080_1914, w_080_1915, w_080_1918, w_080_1921, w_080_1922, w_080_1923, w_080_1924, w_080_1926, w_080_1929, w_080_1930, w_080_1932, w_080_1933, w_080_1935, w_080_1937, w_080_1938, w_080_1942, w_080_1943, w_080_1944, w_080_1949, w_080_1951, w_080_1953, w_080_1954, w_080_1958, w_080_1959, w_080_1960, w_080_1961, w_080_1962, w_080_1968, w_080_1969, w_080_1973, w_080_1975, w_080_1978, w_080_1980, w_080_1983, w_080_1984, w_080_1985, w_080_1989, w_080_1991, w_080_1992, w_080_1994, w_080_1999, w_080_2000, w_080_2002, w_080_2005, w_080_2007, w_080_2009, w_080_2011, w_080_2012, w_080_2014, w_080_2015, w_080_2017, w_080_2018, w_080_2019, w_080_2021, w_080_2022, w_080_2023, w_080_2025, w_080_2026, w_080_2029, w_080_2030, w_080_2034, w_080_2035, w_080_2037, w_080_2038, w_080_2039, w_080_2041, w_080_2042, w_080_2044, w_080_2045, w_080_2046, w_080_2047, w_080_2048, w_080_2050, w_080_2052, w_080_2054, w_080_2055, w_080_2058, w_080_2062, w_080_2064, w_080_2066, w_080_2067, w_080_2069, w_080_2070, w_080_2071, w_080_2072, w_080_2074, w_080_2077, w_080_2081, w_080_2082, w_080_2083, w_080_2085, w_080_2086, w_080_2088, w_080_2090, w_080_2092, w_080_2093, w_080_2094, w_080_2096, w_080_2098, w_080_2101, w_080_2104, w_080_2105, w_080_2107, w_080_2110, w_080_2112, w_080_2115, w_080_2116, w_080_2119, w_080_2120, w_080_2122, w_080_2126, w_080_2127, w_080_2130, w_080_2131, w_080_2134, w_080_2136, w_080_2137, w_080_2138, w_080_2139, w_080_2141, w_080_2142, w_080_2143, w_080_2145, w_080_2146, w_080_2147, w_080_2149, w_080_2151, w_080_2152, w_080_2153, w_080_2155, w_080_2159, w_080_2160, w_080_2162, w_080_2163, w_080_2167, w_080_2169, w_080_2173, w_080_2174, w_080_2175, w_080_2178, w_080_2179, w_080_2185, w_080_2186, w_080_2193, w_080_2194, w_080_2196, w_080_2197, w_080_2199, w_080_2200, w_080_2204, w_080_2205, w_080_2208, w_080_2210, w_080_2211, w_080_2214, w_080_2215, w_080_2220, w_080_2221, w_080_2225, w_080_2226, w_080_2227, w_080_2228, w_080_2229, w_080_2231, w_080_2234, w_080_2236, w_080_2239, w_080_2241, w_080_2242, w_080_2243, w_080_2244, w_080_2245, w_080_2246, w_080_2248, w_080_2249, w_080_2250, w_080_2253, w_080_2257, w_080_2258, w_080_2262, w_080_2263, w_080_2270, w_080_2273, w_080_2275, w_080_2277, w_080_2280, w_080_2283, w_080_2284, w_080_2285, w_080_2286, w_080_2293, w_080_2295, w_080_2300, w_080_2307, w_080_2309, w_080_2317, w_080_2319, w_080_2321, w_080_2329, w_080_2334, w_080_2336, w_080_2338, w_080_2339, w_080_2341, w_080_2343, w_080_2346, w_080_2353, w_080_2355, w_080_2358, w_080_2365, w_080_2370, w_080_2372, w_080_2374, w_080_2380, w_080_2383, w_080_2385, w_080_2386, w_080_2389, w_080_2390, w_080_2394, w_080_2395, w_080_2397, w_080_2402, w_080_2409, w_080_2410, w_080_2411, w_080_2412, w_080_2413, w_080_2415, w_080_2418, w_080_2420, w_080_2421, w_080_2425, w_080_2426, w_080_2442, w_080_2452, w_080_2454, w_080_2459, w_080_2461, w_080_2463, w_080_2465, w_080_2473, w_080_2475, w_080_2476, w_080_2481, w_080_2484, w_080_2485, w_080_2487, w_080_2489, w_080_2493, w_080_2500, w_080_2514, w_080_2517, w_080_2518, w_080_2521, w_080_2532, w_080_2533, w_080_2534, w_080_2537, w_080_2539, w_080_2547, w_080_2551, w_080_2552, w_080_2553, w_080_2560, w_080_2561, w_080_2562, w_080_2564, w_080_2572, w_080_2576, w_080_2579, w_080_2582, w_080_2584, w_080_2587, w_080_2589, w_080_2590, w_080_2592, w_080_2598, w_080_2600, w_080_2610, w_080_2611, w_080_2613, w_080_2615, w_080_2618, w_080_2626, w_080_2633, w_080_2642, w_080_2645, w_080_2648, w_080_2652, w_080_2654, w_080_2655, w_080_2660, w_080_2661, w_080_2662, w_080_2668, w_080_2676, w_080_2679, w_080_2680, w_080_2681, w_080_2684, w_080_2685, w_080_2690, w_080_2691, w_080_2700, w_080_2704, w_080_2709, w_080_2712, w_080_2724, w_080_2726, w_080_2731, w_080_2735, w_080_2738, w_080_2739, w_080_2740, w_080_2751, w_080_2752, w_080_2753, w_080_2759, w_080_2763, w_080_2764, w_080_2765, w_080_2770, w_080_2772, w_080_2773, w_080_2779, w_080_2780, w_080_2788, w_080_2791, w_080_2793, w_080_2797, w_080_2800, w_080_2801, w_080_2810, w_080_2813, w_080_2815, w_080_2818, w_080_2821, w_080_2825, w_080_2828, w_080_2833, w_080_2837, w_080_2838, w_080_2843, w_080_2845, w_080_2847, w_080_2848, w_080_2851, w_080_2852, w_080_2860, w_080_2862, w_080_2864, w_080_2866, w_080_2878, w_080_2883, w_080_2890, w_080_2900, w_080_2901, w_080_2905, w_080_2909, w_080_2911, w_080_2912, w_080_2921, w_080_2923, w_080_2927, w_080_2930, w_080_2934, w_080_2935, w_080_2938, w_080_2939, w_080_2940, w_080_2945, w_080_2947, w_080_2948, w_080_2949, w_080_2953, w_080_2954, w_080_2956, w_080_2959, w_080_2960, w_080_2962, w_080_2963, w_080_2964, w_080_2968, w_080_2974, w_080_2985, w_080_2986, w_080_2990, w_080_2991, w_080_2992, w_080_2995, w_080_2997, w_080_3010, w_080_3012, w_080_3016, w_080_3019, w_080_3023, w_080_3025, w_080_3027, w_080_3028, w_080_3032, w_080_3033, w_080_3039, w_080_3046, w_080_3050, w_080_3054, w_080_3056, w_080_3061, w_080_3066, w_080_3067, w_080_3069, w_080_3070, w_080_3072, w_080_3073, w_080_3076, w_080_3078, w_080_3081, w_080_3083, w_080_3084, w_080_3085, w_080_3090, w_080_3094, w_080_3095, w_080_3096, w_080_3103, w_080_3106, w_080_3110, w_080_3117, w_080_3120, w_080_3127, w_080_3131, w_080_3134, w_080_3138, w_080_3141, w_080_3143, w_080_3148, w_080_3150, w_080_3152, w_080_3154, w_080_3163, w_080_3165, w_080_3175, w_080_3176, w_080_3181, w_080_3187, w_080_3190, w_080_3191, w_080_3201, w_080_3202, w_080_3208, w_080_3219, w_080_3233, w_080_3237, w_080_3239, w_080_3247, w_080_3249, w_080_3250, w_080_3253, w_080_3254, w_080_3262, w_080_3264, w_080_3265, w_080_3271, w_080_3274, w_080_3276, w_080_3279, w_080_3280, w_080_3285, w_080_3286, w_080_3289, w_080_3292, w_080_3294, w_080_3295, w_080_3302, w_080_3303, w_080_3304, w_080_3306, w_080_3309, w_080_3312, w_080_3316, w_080_3317, w_080_3321, w_080_3324, w_080_3331, w_080_3335, w_080_3339, w_080_3342, w_080_3346, w_080_3347, w_080_3351, w_080_3360, w_080_3361, w_080_3363, w_080_3369, w_080_3375, w_080_3376, w_080_3383, w_080_3384, w_080_3389, w_080_3390, w_080_3391, w_080_3392, w_080_3393, w_080_3396, w_080_3398, w_080_3405, w_080_3407, w_080_3409, w_080_3412, w_080_3415, w_080_3418, w_080_3424, w_080_3425, w_080_3428, w_080_3430, w_080_3437, w_080_3444, w_080_3445, w_080_3446, w_080_3447, w_080_3451, w_080_3456, w_080_3459, w_080_3461, w_080_3474, w_080_3475, w_080_3476, w_080_3480, w_080_3481, w_080_3482, w_080_3484, w_080_3485, w_080_3486, w_080_3495, w_080_3499, w_080_3508, w_080_3509, w_080_3510, w_080_3512, w_080_3523, w_080_3529, w_080_3530, w_080_3531, w_080_3532, w_080_3534, w_080_3535, w_080_3541, w_080_3542, w_080_3549, w_080_3550, w_080_3555, w_080_3561, w_080_3562, w_080_3563, w_080_3568, w_080_3569, w_080_3570, w_080_3581, w_080_3582, w_080_3589, w_080_3590, w_080_3598, w_080_3601, w_080_3602, w_080_3606, w_080_3608, w_080_3616, w_080_3617, w_080_3622, w_080_3626, w_080_3627, w_080_3630, w_080_3631, w_080_3637, w_080_3638, w_080_3639, w_080_3640, w_080_3647, w_080_3650, w_080_3651, w_080_3652, w_080_3654, w_080_3662, w_080_3666, w_080_3667, w_080_3672, w_080_3676, w_080_3677, w_080_3682, w_080_3684, w_080_3685, w_080_3686, w_080_3691, w_080_3711, w_080_3712, w_080_3721, w_080_3725, w_080_3731, w_080_3740, w_080_3743, w_080_3746, w_080_3749, w_080_3754, w_080_3765, w_080_3770, w_080_3772, w_080_3773, w_080_3774, w_080_3775, w_080_3778, w_080_3786, w_080_3789, w_080_3790, w_080_3807, w_080_3812, w_080_3813, w_080_3819, w_080_3820, w_080_3822, w_080_3833, w_080_3834, w_080_3835, w_080_3836, w_080_3839, w_080_3840, w_080_3842, w_080_3847, w_080_3849, w_080_3851, w_080_3856, w_080_3858, w_080_3861, w_080_3870, w_080_3873, w_080_3877, w_080_3883, w_080_3884, w_080_3886, w_080_3891, w_080_3895, w_080_3897, w_080_3902, w_080_3905, w_080_3907, w_080_3909, w_080_3910, w_080_3911, w_080_3912, w_080_3918, w_080_3919, w_080_3920, w_080_3922, w_080_3926, w_080_3931, w_080_3933, w_080_3934, w_080_3935, w_080_3937, w_080_3941, w_080_3942, w_080_3943, w_080_3944, w_080_3945, w_080_3950, w_080_3954, w_080_3957, w_080_3959, w_080_3962, w_080_3965, w_080_3966, w_080_3970, w_080_3977, w_080_3982, w_080_3988, w_080_3994, w_080_3997, w_080_3999, w_080_4000, w_080_4001, w_080_4002, w_080_4007, w_080_4013, w_080_4016, w_080_4019, w_080_4023, w_080_4024, w_080_4028, w_080_4036, w_080_4040, w_080_4043, w_080_4044, w_080_4050, w_080_4057, w_080_4058, w_080_4059, w_080_4060, w_080_4061, w_080_4063, w_080_4064, w_080_4065, w_080_4069, w_080_4073, w_080_4077, w_080_4078, w_080_4080, w_080_4087, w_080_4092, w_080_4093, w_080_4095, w_080_4097, w_080_4099, w_080_4106, w_080_4107, w_080_4112, w_080_4120, w_080_4121, w_080_4126, w_080_4135, w_080_4136, w_080_4137, w_080_4138, w_080_4141, w_080_4145, w_080_4154, w_080_4156, w_080_4161, w_080_4165, w_080_4167, w_080_4169, w_080_4176, w_080_4177, w_080_4179, w_080_4190, w_080_4196, w_080_4201, w_080_4202, w_080_4206, w_080_4211, w_080_4216, w_080_4220, w_080_4223, w_080_4225, w_080_4226, w_080_4230, w_080_4233, w_080_4235, w_080_4236, w_080_4242, w_080_4243, w_080_4245, w_080_4249, w_080_4251, w_080_4256, w_080_4260, w_080_4261, w_080_4267, w_080_4272, w_080_4273, w_080_4274, w_080_4294, w_080_4299, w_080_4301, w_080_4302, w_080_4305, w_080_4308, w_080_4314, w_080_4315, w_080_4317, w_080_4320, w_080_4324, w_080_4325, w_080_4333, w_080_4334, w_080_4338, w_080_4348, w_080_4355, w_080_4363, w_080_4364, w_080_4368, w_080_4370, w_080_4390, w_080_4391, w_080_4392, w_080_4393, w_080_4394, w_080_4395, w_080_4401, w_080_4403, w_080_4404, w_080_4405, w_080_4409, w_080_4411, w_080_4412, w_080_4421, w_080_4423, w_080_4429, w_080_4430, w_080_4432, w_080_4436, w_080_4437, w_080_4440, w_080_4443, w_080_4444, w_080_4450, w_080_4451, w_080_4455, w_080_4458, w_080_4463, w_080_4464, w_080_4468, w_080_4472, w_080_4474, w_080_4476, w_080_4480, w_080_4484, w_080_4485, w_080_4490, w_080_4491, w_080_4497, w_080_4506, w_080_4509, w_080_4518, w_080_4520, w_080_4524, w_080_4527, w_080_4540, w_080_4544, w_080_4548, w_080_4549, w_080_4552, w_080_4554, w_080_4556, w_080_4559, w_080_4560, w_080_4563, w_080_4567, w_080_4570, w_080_4571, w_080_4574, w_080_4577, w_080_4581, w_080_4583, w_080_4584, w_080_4590, w_080_4593, w_080_4599, w_080_4600, w_080_4607, w_080_4611, w_080_4615, w_080_4619, w_080_4620, w_080_4621, w_080_4627, w_080_4635, w_080_4644, w_080_4646, w_080_4647, w_080_4648, w_080_4651, w_080_4652, w_080_4656, w_080_4663, w_080_4665, w_080_4667, w_080_4671, w_080_4678, w_080_4679, w_080_4685, w_080_4686, w_080_4687, w_080_4688, w_080_4694, w_080_4695, w_080_4696, w_080_4698, w_080_4702, w_080_4704, w_080_4706, w_080_4707, w_080_4708, w_080_4712, w_080_4723, w_080_4726, w_080_4743, w_080_4744, w_080_4745, w_080_4752, w_080_4756, w_080_4760, w_080_4765, w_080_4767, w_080_4771, w_080_4776, w_080_4779, w_080_4784, w_080_4793, w_080_4795, w_080_4799, w_080_4804, w_080_4805, w_080_4806, w_080_4808, w_080_4811, w_080_4816, w_080_4820, w_080_4821, w_080_4823, w_080_4826, w_080_4829, w_080_4830, w_080_4831, w_080_4832, w_080_4837, w_080_4840, w_080_4842, w_080_4844, w_080_4848, w_080_4849, w_080_4863, w_080_4866, w_080_4867, w_080_4868, w_080_4870, w_080_4874, w_080_4875, w_080_4876, w_080_4877, w_080_4880, w_080_4883, w_080_4886, w_080_4889, w_080_4890, w_080_4896, w_080_4899, w_080_4900, w_080_4901, w_080_4902, w_080_4906, w_080_4907, w_080_4908, w_080_4914, w_080_4915, w_080_4916, w_080_4917, w_080_4929, w_080_4932, w_080_4933, w_080_4937, w_080_4938, w_080_4946, w_080_4954, w_080_4960, w_080_4962, w_080_4963, w_080_4967, w_080_4971, w_080_4975, w_080_4976, w_080_4988, w_080_4990, w_080_4991, w_080_4994, w_080_4998, w_080_5004, w_080_5010, w_080_5014, w_080_5017, w_080_5018, w_080_5025, w_080_5028, w_080_5037, w_080_5049, w_080_5051, w_080_5054, w_080_5058, w_080_5060, w_080_5064, w_080_5066, w_080_5070, w_080_5072, w_080_5073, w_080_5074, w_080_5076, w_080_5079, w_080_5083, w_080_5084, w_080_5086, w_080_5087, w_080_5089, w_080_5093, w_080_5094, w_080_5099, w_080_5107, w_080_5108, w_080_5112, w_080_5114, w_080_5115, w_080_5118, w_080_5121, w_080_5122, w_080_5125, w_080_5126, w_080_5133, w_080_5137, w_080_5138, w_080_5150, w_080_5159, w_080_5165, w_080_5171, w_080_5174, w_080_5176, w_080_5177, w_080_5178, w_080_5179, w_080_5180, w_080_5186, w_080_5188, w_080_5189, w_080_5191, w_080_5196, w_080_5198, w_080_5202, w_080_5208, w_080_5214, w_080_5217, w_080_5219, w_080_5224, w_080_5228, w_080_5230, w_080_5237, w_080_5242, w_080_5245, w_080_5249, w_080_5256, w_080_5264, w_080_5268, w_080_5269, w_080_5280, w_080_5285, w_080_5286, w_080_5290, w_080_5309, w_080_5313, w_080_5315, w_080_5317, w_080_5319, w_080_5323, w_080_5325, w_080_5327, w_080_5329, w_080_5331, w_080_5335, w_080_5337, w_080_5343, w_080_5344, w_080_5350, w_080_5356, w_080_5365, w_080_5366, w_080_5371, w_080_5376, w_080_5379, w_080_5385, w_080_5393, w_080_5394, w_080_5395, w_080_5397, w_080_5398, w_080_5399, w_080_5402, w_080_5404, w_080_5405, w_080_5406, w_080_5407, w_080_5412, w_080_5413, w_080_5419, w_080_5421, w_080_5428, w_080_5429, w_080_5430, w_080_5432, w_080_5434, w_080_5447, w_080_5448, w_080_5451, w_080_5452, w_080_5455, w_080_5457, w_080_5459, w_080_5460, w_080_5466, w_080_5468, w_080_5473, w_080_5474, w_080_5476, w_080_5481, w_080_5486, w_080_5491, w_080_5498, w_080_5503, w_080_5506, w_080_5509, w_080_5516, w_080_5521, w_080_5535, w_080_5538, w_080_5539, w_080_5555, w_080_5558, w_080_5560, w_080_5561, w_080_5568, w_080_5571, w_080_5574, w_080_5580, w_080_5581, w_080_5587, w_080_5588, w_080_5589, w_080_5592, w_080_5597, w_080_5602, w_080_5603, w_080_5606, w_080_5610, w_080_5613, w_080_5616, w_080_5618, w_080_5619, w_080_5627, w_080_5628, w_080_5630, w_080_5632, w_080_5635, w_080_5638, w_080_5643, w_080_5646, w_080_5647, w_080_5650, w_080_5653, w_080_5654, w_080_5663, w_080_5664, w_080_5665, w_080_5670, w_080_5673, w_080_5676, w_080_5679, w_080_5681, w_080_5686, w_080_5690, w_080_5692, w_080_5693, w_080_5695, w_080_5697, w_080_5703, w_080_5704, w_080_5708, w_080_5709, w_080_5714, w_080_5716, w_080_5717, w_080_5720, w_080_5721, w_080_5725, w_080_5727, w_080_5730, w_080_5733, w_080_5742, w_080_5744, w_080_5748, w_080_5750, w_080_5752, w_080_5753, w_080_5758, w_080_5763, w_080_5764, w_080_5773, w_080_5787, w_080_5789, w_080_5792, w_080_5794, w_080_5796, w_080_5797, w_080_5799, w_080_5800, w_080_5801, w_080_5805, w_080_5807, w_080_5810, w_080_5818, w_080_5820, w_080_5824, w_080_5825, w_080_5826, w_080_5836, w_080_5838, w_080_5839, w_080_5840, w_080_5843, w_080_5850, w_080_5853, w_080_5855, w_080_5856, w_080_5861, w_080_5870, w_080_5871, w_080_5872, w_080_5873, w_080_5874, w_080_5875, w_080_5877, w_080_5884, w_080_5889, w_080_5890, w_080_5898, w_080_5904, w_080_5910, w_080_5913, w_080_5914, w_080_5915, w_080_5917, w_080_5920, w_080_5930, w_080_5932, w_080_5933, w_080_5934, w_080_5936, w_080_5937, w_080_5939, w_080_5941, w_080_5942, w_080_5944, w_080_5958, w_080_5969, w_080_5972, w_080_5973, w_080_5974, w_080_5980, w_080_5981, w_080_5990, w_080_5991, w_080_6002, w_080_6004, w_080_6005, w_080_6006, w_080_6009, w_080_6016, w_080_6027, w_080_6031, w_080_6033, w_080_6038, w_080_6039, w_080_6041, w_080_6045, w_080_6048, w_080_6052, w_080_6057, w_080_6058, w_080_6063, w_080_6064, w_080_6065, w_080_6073, w_080_6075, w_080_6076, w_080_6084, w_080_6087, w_080_6088, w_080_6090, w_080_6094, w_080_6098, w_080_6103, w_080_6106, w_080_6107, w_080_6108, w_080_6112, w_080_6120, w_080_6125, w_080_6128, w_080_6131, w_080_6136, w_080_6159, w_080_6161, w_080_6165, w_080_6169, w_080_6172, w_080_6174, w_080_6183, w_080_6184, w_080_6186, w_080_6193, w_080_6197, w_080_6200, w_080_6203, w_080_6204, w_080_6205, w_080_6213, w_080_6216, w_080_6219, w_080_6220, w_080_6222, w_080_6229, w_080_6235, w_080_6243, w_080_6245, w_080_6250, w_080_6254, w_080_6255, w_080_6257, w_080_6262, w_080_6263, w_080_6264, w_080_6268, w_080_6271, w_080_6275, w_080_6278, w_080_6281, w_080_6283, w_080_6286, w_080_6288, w_080_6290, w_080_6291, w_080_6292, w_080_6293, w_080_6294, w_080_6295, w_080_6302, w_080_6310, w_080_6312, w_080_6314, w_080_6316, w_080_6320, w_080_6325, w_080_6327, w_080_6330, w_080_6345, w_080_6349, w_080_6352, w_080_6356, w_080_6359, w_080_6360, w_080_6361, w_080_6365, w_080_6372, w_080_6381, w_080_6386, w_080_6387, w_080_6389, w_080_6391, w_080_6393, w_080_6397, w_080_6399, w_080_6404, w_080_6405, w_080_6407, w_080_6414, w_080_6417, w_080_6419, w_080_6420, w_080_6421, w_080_6425, w_080_6429, w_080_6434, w_080_6436, w_080_6445, w_080_6448, w_080_6450, w_080_6456, w_080_6457, w_080_6463, w_080_6465, w_080_6468, w_080_6472, w_080_6481, w_080_6482, w_080_6483, w_080_6485, w_080_6486, w_080_6490, w_080_6491, w_080_6492, w_080_6493, w_080_6496, w_080_6504, w_080_6510, w_080_6515, w_080_6519, w_080_6521, w_080_6531, w_080_6532, w_080_6535, w_080_6536, w_080_6538, w_080_6541, w_080_6548, w_080_6549, w_080_6552, w_080_6554, w_080_6561, w_080_6562, w_080_6563, w_080_6566, w_080_6568, w_080_6570, w_080_6578, w_080_6581, w_080_6583, w_080_6585, w_080_6588, w_080_6590, w_080_6591, w_080_6593, w_080_6601, w_080_6603, w_080_6604, w_080_6612, w_080_6613, w_080_6614, w_080_6617, w_080_6618, w_080_6620, w_080_6621, w_080_6624, w_080_6628, w_080_6629, w_080_6633, w_080_6635, w_080_6641, w_080_6644, w_080_6645, w_080_6648, w_080_6649, w_080_6655, w_080_6656, w_080_6657, w_080_6660, w_080_6662, w_080_6681, w_080_6688, w_080_6701, w_080_6709, w_080_6713, w_080_6716, w_080_6719, w_080_6721, w_080_6724, w_080_6725, w_080_6726, w_080_6731, w_080_6732, w_080_6735, w_080_6737, w_080_6743, w_080_6749, w_080_6754, w_080_6760, w_080_6763, w_080_6772, w_080_6774, w_080_6781, w_080_6782, w_080_6787, w_080_6788, w_080_6791, w_080_6796, w_080_6797, w_080_6801, w_080_6803, w_080_6811, w_080_6812, w_080_6815, w_080_6817, w_080_6826, w_080_6834, w_080_6838, w_080_6839, w_080_6841, w_080_6842, w_080_6848, w_080_6851, w_080_6853, w_080_6854, w_080_6855, w_080_6856, w_080_6858, w_080_6862, w_080_6863, w_080_6866, w_080_6868, w_080_6869, w_080_6870, w_080_6871, w_080_6872, w_080_6874, w_080_6876, w_080_6882, w_080_6886, w_080_6898, w_080_6900, w_080_6901, w_080_6907, w_080_6912, w_080_6914, w_080_6919, w_080_6923, w_080_6926, w_080_6927, w_080_6933, w_080_6935, w_080_6943, w_080_6944, w_080_6953, w_080_6955, w_080_6958, w_080_6962, w_080_6963, w_080_6966, w_080_6967, w_080_6968, w_080_6971, w_080_6975, w_080_6981, w_080_6985, w_080_6988, w_080_6991, w_080_6992, w_080_6994, w_080_6996, w_080_6998, w_080_7000, w_080_7003, w_080_7016, w_080_7017, w_080_7021, w_080_7022, w_080_7023, w_080_7026, w_080_7031, w_080_7045, w_080_7048, w_080_7049, w_080_7050, w_080_7053, w_080_7058, w_080_7059, w_080_7064, w_080_7068, w_080_7070, w_080_7071, w_080_7073, w_080_7075, w_080_7079, w_080_7083, w_080_7088, w_080_7091, w_080_7096, w_080_7098, w_080_7105, w_080_7108, w_080_7109, w_080_7115, w_080_7117, w_080_7121, w_080_7124, w_080_7127, w_080_7132, w_080_7135, w_080_7138, w_080_7142, w_080_7143, w_080_7147, w_080_7150, w_080_7151, w_080_7154, w_080_7160, w_080_7164, w_080_7166, w_080_7171, w_080_7172, w_080_7175, w_080_7185, w_080_7195, w_080_7196, w_080_7202, w_080_7204, w_080_7206, w_080_7213, w_080_7221, w_080_7224, w_080_7232, w_080_7240, w_080_7243, w_080_7246, w_080_7248, w_080_7254, w_080_7257, w_080_7258, w_080_7262, w_080_7263, w_080_7270, w_080_7271, w_080_7273, w_080_7275, w_080_7279, w_080_7284, w_080_7288, w_080_7290, w_080_7291, w_080_7296, w_080_7302, w_080_7308, w_080_7310, w_080_7312, w_080_7314, w_080_7316, w_080_7318, w_080_7323, w_080_7326, w_080_7330, w_080_7334, w_080_7339, w_080_7340, w_080_7343, w_080_7345, w_080_7356, w_080_7361, w_080_7367, w_080_7368, w_080_7371, w_080_7374, w_080_7381, w_080_7385, w_080_7387, w_080_7388, w_080_7389, w_080_7390, w_080_7391, w_080_7392, w_080_7396, w_080_7398, w_080_7399, w_080_7402, w_080_7403, w_080_7405, w_080_7409, w_080_7414, w_080_7419, w_080_7420, w_080_7424, w_080_7431, w_080_7433, w_080_7434, w_080_7435, w_080_7436, w_080_7438, w_080_7440, w_080_7441, w_080_7442, w_080_7444, w_080_7445, w_080_7458, w_080_7460, w_080_7479, w_080_7481, w_080_7483, w_080_7487, w_080_7488, w_080_7490, w_080_7493, w_080_7496, w_080_7497, w_080_7501, w_080_7503, w_080_7505, w_080_7506, w_080_7508, w_080_7525, w_080_7531, w_080_7536, w_080_7539, w_080_7543, w_080_7546, w_080_7550, w_080_7551, w_080_7552, w_080_7555, w_080_7560, w_080_7571, w_080_7574, w_080_7575, w_080_7581, w_080_7582, w_080_7587, w_080_7588, w_080_7592, w_080_7599, w_080_7600, w_080_7602, w_080_7603, w_080_7607, w_080_7613, w_080_7615, w_080_7624, w_080_7628, w_080_7631, w_080_7634, w_080_7636, w_080_7640, w_080_7641, w_080_7646, w_080_7649, w_080_7650, w_080_7651, w_080_7652, w_080_7654, w_080_7655, w_080_7656, w_080_7657, w_080_7660, w_080_7663, w_080_7667, w_080_7675, w_080_7678, w_080_7680, w_080_7684, w_080_7691, w_080_7693, w_080_7694, w_080_7695, w_080_7696, w_080_7700, w_080_7703, w_080_7705, w_080_7712;
  wire w_081_001, w_081_002, w_081_003, w_081_004, w_081_006, w_081_008, w_081_011, w_081_012, w_081_015, w_081_016, w_081_018, w_081_022, w_081_023, w_081_024, w_081_026, w_081_027, w_081_028, w_081_029, w_081_034, w_081_035, w_081_037, w_081_039, w_081_040, w_081_041, w_081_042, w_081_043, w_081_050, w_081_054, w_081_061, w_081_062, w_081_065, w_081_066, w_081_067, w_081_071, w_081_072, w_081_075, w_081_076, w_081_077, w_081_078, w_081_080, w_081_087, w_081_088, w_081_089, w_081_091, w_081_093, w_081_094, w_081_095, w_081_096, w_081_097, w_081_100, w_081_102, w_081_104, w_081_106, w_081_107, w_081_111, w_081_112, w_081_114, w_081_115, w_081_118, w_081_120, w_081_121, w_081_122, w_081_123, w_081_124, w_081_125, w_081_127, w_081_137, w_081_142, w_081_143, w_081_146, w_081_147, w_081_148, w_081_152, w_081_153, w_081_155, w_081_156, w_081_159, w_081_160, w_081_161, w_081_162, w_081_163, w_081_165, w_081_167, w_081_169, w_081_171, w_081_172, w_081_175, w_081_181, w_081_182, w_081_184, w_081_186, w_081_187, w_081_189, w_081_192, w_081_197, w_081_200, w_081_201, w_081_204, w_081_205, w_081_206, w_081_208, w_081_210, w_081_212, w_081_213, w_081_214, w_081_217, w_081_221, w_081_225, w_081_232, w_081_235, w_081_237, w_081_238, w_081_239, w_081_242, w_081_244, w_081_245, w_081_247, w_081_249, w_081_250, w_081_251, w_081_252, w_081_253, w_081_255, w_081_256, w_081_259, w_081_261, w_081_263, w_081_264, w_081_265, w_081_266, w_081_270, w_081_272, w_081_275, w_081_277, w_081_278, w_081_279, w_081_280, w_081_282, w_081_283, w_081_285, w_081_287, w_081_293, w_081_295, w_081_296, w_081_297, w_081_298, w_081_299, w_081_303, w_081_305, w_081_308, w_081_310, w_081_312, w_081_314, w_081_316, w_081_318, w_081_319, w_081_321, w_081_322, w_081_324, w_081_332, w_081_334, w_081_335, w_081_336, w_081_337, w_081_338, w_081_345, w_081_348, w_081_351, w_081_352, w_081_353, w_081_356, w_081_357, w_081_358, w_081_360, w_081_362, w_081_363, w_081_365, w_081_368, w_081_374, w_081_376, w_081_377, w_081_379, w_081_382, w_081_383, w_081_384, w_081_387, w_081_388, w_081_392, w_081_397, w_081_400, w_081_402, w_081_404, w_081_405, w_081_410, w_081_411, w_081_413, w_081_418, w_081_422, w_081_424, w_081_425, w_081_427, w_081_428, w_081_429, w_081_430, w_081_431, w_081_434, w_081_436, w_081_437, w_081_438, w_081_440, w_081_441, w_081_443, w_081_444, w_081_445, w_081_446, w_081_447, w_081_449, w_081_450, w_081_452, w_081_454, w_081_455, w_081_456, w_081_464, w_081_467, w_081_468, w_081_475, w_081_477, w_081_480, w_081_481, w_081_483, w_081_484, w_081_486, w_081_490, w_081_491, w_081_492, w_081_493, w_081_495, w_081_497, w_081_498, w_081_500, w_081_501, w_081_502, w_081_503, w_081_505, w_081_506, w_081_507, w_081_509, w_081_513, w_081_514, w_081_515, w_081_522, w_081_524, w_081_526, w_081_527, w_081_528, w_081_534, w_081_537, w_081_538, w_081_543, w_081_549, w_081_550, w_081_552, w_081_554, w_081_556, w_081_559, w_081_561, w_081_563, w_081_566, w_081_567, w_081_568, w_081_569, w_081_570, w_081_574, w_081_577, w_081_579, w_081_581, w_081_583, w_081_586, w_081_587, w_081_590, w_081_591, w_081_592, w_081_597, w_081_599, w_081_602, w_081_604, w_081_605, w_081_606, w_081_610, w_081_611, w_081_612, w_081_613, w_081_614, w_081_615, w_081_617, w_081_619, w_081_621, w_081_623, w_081_624, w_081_626, w_081_629, w_081_630, w_081_633, w_081_634, w_081_636, w_081_643, w_081_644, w_081_645, w_081_647, w_081_649, w_081_650, w_081_655, w_081_657, w_081_660, w_081_661, w_081_663, w_081_664, w_081_667, w_081_670, w_081_672, w_081_677, w_081_678, w_081_679, w_081_680, w_081_681, w_081_683, w_081_685, w_081_687, w_081_688, w_081_689, w_081_690, w_081_692, w_081_693, w_081_699, w_081_702, w_081_704, w_081_705, w_081_707, w_081_708, w_081_709, w_081_710, w_081_712, w_081_713, w_081_714, w_081_717, w_081_720, w_081_722, w_081_723, w_081_725, w_081_727, w_081_732, w_081_734, w_081_735, w_081_742, w_081_745, w_081_746, w_081_747, w_081_749, w_081_751, w_081_754, w_081_755, w_081_756, w_081_758, w_081_759, w_081_760, w_081_762, w_081_763, w_081_767, w_081_768, w_081_769, w_081_772, w_081_773, w_081_775, w_081_776, w_081_783, w_081_790, w_081_791, w_081_792, w_081_793, w_081_796, w_081_799, w_081_803, w_081_804, w_081_808, w_081_809, w_081_810, w_081_815, w_081_818, w_081_821, w_081_827, w_081_828, w_081_831, w_081_832, w_081_833, w_081_834, w_081_836, w_081_837, w_081_839, w_081_842, w_081_844, w_081_848, w_081_852, w_081_856, w_081_857, w_081_858, w_081_859, w_081_862, w_081_863, w_081_864, w_081_867, w_081_872, w_081_873, w_081_875, w_081_876, w_081_884, w_081_886, w_081_888, w_081_892, w_081_893, w_081_896, w_081_898, w_081_901, w_081_902, w_081_903, w_081_905, w_081_906, w_081_909, w_081_910, w_081_911, w_081_912, w_081_914, w_081_915, w_081_916, w_081_918, w_081_919, w_081_922, w_081_923, w_081_927, w_081_928, w_081_933, w_081_934, w_081_937, w_081_939, w_081_942, w_081_945, w_081_947, w_081_948, w_081_949, w_081_950, w_081_955, w_081_956, w_081_957, w_081_960, w_081_961, w_081_964, w_081_965, w_081_966, w_081_969, w_081_970, w_081_971, w_081_972, w_081_973, w_081_974, w_081_978, w_081_980, w_081_986, w_081_988, w_081_989, w_081_990, w_081_991, w_081_992, w_081_994, w_081_996, w_081_997, w_081_998, w_081_999, w_081_1000, w_081_1002, w_081_1006, w_081_1007, w_081_1008, w_081_1010, w_081_1011, w_081_1012, w_081_1014, w_081_1015, w_081_1017, w_081_1019, w_081_1020, w_081_1023, w_081_1025, w_081_1026, w_081_1027, w_081_1030, w_081_1034, w_081_1039, w_081_1042, w_081_1043, w_081_1045, w_081_1046, w_081_1047, w_081_1049, w_081_1055, w_081_1058, w_081_1060, w_081_1066, w_081_1069, w_081_1073, w_081_1075, w_081_1078, w_081_1080, w_081_1081, w_081_1084, w_081_1088, w_081_1089, w_081_1093, w_081_1096, w_081_1097, w_081_1098, w_081_1099, w_081_1100, w_081_1107, w_081_1108, w_081_1109, w_081_1113, w_081_1114, w_081_1118, w_081_1119, w_081_1120, w_081_1121, w_081_1122, w_081_1123, w_081_1124, w_081_1127, w_081_1132, w_081_1135, w_081_1136, w_081_1137, w_081_1139, w_081_1141, w_081_1142, w_081_1143, w_081_1145, w_081_1146, w_081_1150, w_081_1151, w_081_1152, w_081_1153, w_081_1154, w_081_1156, w_081_1159, w_081_1160, w_081_1161, w_081_1164, w_081_1165, w_081_1167, w_081_1169, w_081_1170, w_081_1173, w_081_1174, w_081_1175, w_081_1176, w_081_1178, w_081_1179, w_081_1181, w_081_1183, w_081_1185, w_081_1189, w_081_1190, w_081_1194, w_081_1195, w_081_1196, w_081_1197, w_081_1199, w_081_1200, w_081_1202, w_081_1203, w_081_1206, w_081_1208, w_081_1211, w_081_1213, w_081_1214, w_081_1215, w_081_1216, w_081_1218, w_081_1220, w_081_1221, w_081_1222, w_081_1223, w_081_1225, w_081_1226, w_081_1229, w_081_1231, w_081_1234, w_081_1235, w_081_1237, w_081_1238, w_081_1239, w_081_1241, w_081_1242, w_081_1243, w_081_1244, w_081_1246, w_081_1247, w_081_1249, w_081_1251, w_081_1254, w_081_1255, w_081_1256, w_081_1259, w_081_1260, w_081_1261, w_081_1263, w_081_1266, w_081_1269, w_081_1271, w_081_1273, w_081_1276, w_081_1277, w_081_1282, w_081_1283, w_081_1286, w_081_1287, w_081_1288, w_081_1289, w_081_1290, w_081_1291, w_081_1292, w_081_1293, w_081_1296, w_081_1299, w_081_1300, w_081_1302, w_081_1304, w_081_1305, w_081_1306, w_081_1307, w_081_1312, w_081_1313, w_081_1315, w_081_1316, w_081_1317, w_081_1319, w_081_1323, w_081_1325, w_081_1327, w_081_1328, w_081_1330, w_081_1333, w_081_1338, w_081_1340, w_081_1343, w_081_1344, w_081_1345, w_081_1346, w_081_1347, w_081_1350, w_081_1352, w_081_1355, w_081_1356, w_081_1357, w_081_1360, w_081_1362, w_081_1364, w_081_1365, w_081_1369, w_081_1370, w_081_1372, w_081_1378, w_081_1379, w_081_1380, w_081_1381, w_081_1383, w_081_1386, w_081_1387, w_081_1389, w_081_1390, w_081_1395, w_081_1396, w_081_1398, w_081_1400, w_081_1402, w_081_1403, w_081_1404, w_081_1406, w_081_1410, w_081_1412, w_081_1413, w_081_1415, w_081_1416, w_081_1417, w_081_1423, w_081_1432, w_081_1435, w_081_1437, w_081_1442, w_081_1443, w_081_1447, w_081_1450, w_081_1452, w_081_1455, w_081_1456, w_081_1459, w_081_1463, w_081_1466, w_081_1467, w_081_1468, w_081_1469, w_081_1471, w_081_1473, w_081_1474, w_081_1476, w_081_1477, w_081_1479, w_081_1482, w_081_1483, w_081_1484, w_081_1486, w_081_1490, w_081_1491, w_081_1492, w_081_1495, w_081_1498, w_081_1499, w_081_1501, w_081_1504, w_081_1506, w_081_1507, w_081_1509, w_081_1511, w_081_1513, w_081_1514, w_081_1516, w_081_1517, w_081_1521, w_081_1523, w_081_1525, w_081_1526, w_081_1529, w_081_1530, w_081_1533, w_081_1535, w_081_1538, w_081_1540, w_081_1541, w_081_1544, w_081_1547, w_081_1549, w_081_1552, w_081_1555, w_081_1557, w_081_1561, w_081_1562, w_081_1563, w_081_1564, w_081_1565, w_081_1567, w_081_1571, w_081_1572, w_081_1574, w_081_1576, w_081_1579, w_081_1580, w_081_1581, w_081_1582, w_081_1589, w_081_1591, w_081_1592, w_081_1593, w_081_1594, w_081_1598, w_081_1599, w_081_1601, w_081_1604, w_081_1605, w_081_1607, w_081_1610, w_081_1612, w_081_1613, w_081_1614, w_081_1616, w_081_1619, w_081_1622, w_081_1625, w_081_1626, w_081_1627, w_081_1630, w_081_1633, w_081_1637, w_081_1638, w_081_1640, w_081_1642, w_081_1643, w_081_1645, w_081_1647, w_081_1648, w_081_1649, w_081_1653, w_081_1656, w_081_1658, w_081_1659, w_081_1660, w_081_1661, w_081_1664, w_081_1670, w_081_1673, w_081_1674, w_081_1677, w_081_1680, w_081_1681, w_081_1684, w_081_1685, w_081_1689, w_081_1692, w_081_1696, w_081_1697, w_081_1700, w_081_1701, w_081_1705, w_081_1707, w_081_1708, w_081_1709, w_081_1713, w_081_1715, w_081_1716, w_081_1717, w_081_1719, w_081_1723, w_081_1727, w_081_1729, w_081_1732, w_081_1738, w_081_1739, w_081_1742, w_081_1743, w_081_1744, w_081_1745, w_081_1746, w_081_1747, w_081_1749, w_081_1751, w_081_1753, w_081_1755, w_081_1760, w_081_1761, w_081_1762, w_081_1764, w_081_1766, w_081_1767, w_081_1768, w_081_1769, w_081_1771, w_081_1772, w_081_1773, w_081_1774, w_081_1778, w_081_1780, w_081_1781, w_081_1782, w_081_1783, w_081_1784, w_081_1786, w_081_1787, w_081_1795, w_081_1796, w_081_1797, w_081_1798, w_081_1804, w_081_1806, w_081_1807, w_081_1808, w_081_1810, w_081_1812, w_081_1816, w_081_1819, w_081_1821, w_081_1827, w_081_1828, w_081_1829, w_081_1831, w_081_1833, w_081_1834, w_081_1835, w_081_1840, w_081_1841, w_081_1844, w_081_1847, w_081_1852, w_081_1853, w_081_1854, w_081_1856, w_081_1858, w_081_1863, w_081_1865, w_081_1866, w_081_1869, w_081_1870, w_081_1872, w_081_1873, w_081_1874, w_081_1876, w_081_1878, w_081_1879, w_081_1880, w_081_1882, w_081_1883, w_081_1884, w_081_1888, w_081_1891, w_081_1892, w_081_1893, w_081_1894, w_081_1896, w_081_1899, w_081_1900, w_081_1901, w_081_1902, w_081_1903, w_081_1905, w_081_1906, w_081_1910, w_081_1912, w_081_1916, w_081_1917, w_081_1919, w_081_1920, w_081_1925, w_081_1926, w_081_1927, w_081_1930, w_081_1931, w_081_1932, w_081_1939, w_081_1941, w_081_1942, w_081_1944, w_081_1945, w_081_1947, w_081_1950, w_081_1955, w_081_1957, w_081_1958, w_081_1959, w_081_1960, w_081_1961, w_081_1962, w_081_1963, w_081_1966, w_081_1969, w_081_1970, w_081_1973, w_081_1976, w_081_1979, w_081_1981, w_081_1982, w_081_1984, w_081_1988, w_081_1990, w_081_1991, w_081_1994, w_081_1995, w_081_1999, w_081_2000, w_081_2001, w_081_2004, w_081_2006, w_081_2008, w_081_2009, w_081_2010, w_081_2012, w_081_2013, w_081_2015, w_081_2017, w_081_2018, w_081_2019, w_081_2020, w_081_2023, w_081_2027, w_081_2033, w_081_2034, w_081_2036, w_081_2037, w_081_2038, w_081_2040, w_081_2042, w_081_2043, w_081_2048, w_081_2049, w_081_2051, w_081_2053, w_081_2054, w_081_2056, w_081_2058, w_081_2059, w_081_2062, w_081_2064, w_081_2065, w_081_2066, w_081_2068, w_081_2070, w_081_2071, w_081_2073, w_081_2074, w_081_2075, w_081_2076, w_081_2077, w_081_2078, w_081_2081, w_081_2083, w_081_2084, w_081_2087, w_081_2088, w_081_2092, w_081_2096, w_081_2097, w_081_2098, w_081_2100, w_081_2102, w_081_2106, w_081_2107, w_081_2110, w_081_2112, w_081_2114, w_081_2115, w_081_2116, w_081_2117, w_081_2119, w_081_2122, w_081_2124, w_081_2125, w_081_2128, w_081_2129, w_081_2130, w_081_2131, w_081_2132, w_081_2134, w_081_2137, w_081_2140, w_081_2141, w_081_2142, w_081_2143, w_081_2148, w_081_2151, w_081_2153, w_081_2155, w_081_2157, w_081_2159, w_081_2161, w_081_2162, w_081_2163, w_081_2167, w_081_2169, w_081_2170, w_081_2173, w_081_2175, w_081_2176, w_081_2186, w_081_2188, w_081_2190, w_081_2192, w_081_2193, w_081_2199, w_081_2200, w_081_2202, w_081_2205, w_081_2206, w_081_2208, w_081_2213, w_081_2217, w_081_2218, w_081_2219, w_081_2221, w_081_2224, w_081_2226, w_081_2227, w_081_2228, w_081_2229, w_081_2235, w_081_2238, w_081_2242, w_081_2246, w_081_2250, w_081_2251, w_081_2252, w_081_2253, w_081_2254, w_081_2255, w_081_2260, w_081_2263, w_081_2264, w_081_2267, w_081_2271, w_081_2272, w_081_2273, w_081_2274, w_081_2275, w_081_2276, w_081_2277, w_081_2279, w_081_2283, w_081_2285, w_081_2286, w_081_2288, w_081_2293, w_081_2294, w_081_2297, w_081_2300, w_081_2302, w_081_2303, w_081_2304, w_081_2305, w_081_2307, w_081_2308, w_081_2309, w_081_2311, w_081_2313, w_081_2316, w_081_2320, w_081_2321, w_081_2323, w_081_2324, w_081_2325, w_081_2327, w_081_2331, w_081_2334, w_081_2337, w_081_2338, w_081_2339, w_081_2340, w_081_2341, w_081_2343, w_081_2349, w_081_2352, w_081_2356, w_081_2362, w_081_2364, w_081_2365, w_081_2366, w_081_2367, w_081_2372, w_081_2374, w_081_2375, w_081_2377, w_081_2379, w_081_2380, w_081_2381, w_081_2387, w_081_2390, w_081_2391, w_081_2392, w_081_2393, w_081_2395, w_081_2396, w_081_2397, w_081_2401, w_081_2403, w_081_2404, w_081_2406, w_081_2409, w_081_2410, w_081_2413, w_081_2414, w_081_2415, w_081_2416, w_081_2418, w_081_2419, w_081_2420, w_081_2421, w_081_2424, w_081_2428, w_081_2432, w_081_2433, w_081_2434, w_081_2436, w_081_2437, w_081_2438, w_081_2440, w_081_2441, w_081_2442, w_081_2443, w_081_2446, w_081_2447, w_081_2450, w_081_2452, w_081_2454, w_081_2455, w_081_2457, w_081_2462, w_081_2463, w_081_2467, w_081_2468, w_081_2469, w_081_2473, w_081_2476, w_081_2477, w_081_2480, w_081_2485, w_081_2487, w_081_2488, w_081_2490, w_081_2492, w_081_2494, w_081_2496, w_081_2497, w_081_2498, w_081_2499, w_081_2501, w_081_2505, w_081_2508, w_081_2509, w_081_2510, w_081_2512, w_081_2513, w_081_2516, w_081_2517, w_081_2518, w_081_2519, w_081_2520, w_081_2524, w_081_2525, w_081_2528, w_081_2529, w_081_2531, w_081_2534, w_081_2535, w_081_2537, w_081_2538, w_081_2542, w_081_2545, w_081_2548, w_081_2551, w_081_2552, w_081_2554, w_081_2557, w_081_2560, w_081_2563, w_081_2568, w_081_2569, w_081_2571, w_081_2572, w_081_2573, w_081_2574, w_081_2575, w_081_2584, w_081_2586, w_081_2587, w_081_2588, w_081_2589, w_081_2590, w_081_2591, w_081_2592, w_081_2594, w_081_2598, w_081_2599, w_081_2601, w_081_2603, w_081_2606, w_081_2609, w_081_2612, w_081_2614, w_081_2617, w_081_2623, w_081_2627, w_081_2632, w_081_2635, w_081_2636, w_081_2637, w_081_2641, w_081_2642, w_081_2643, w_081_2645, w_081_2646, w_081_2650, w_081_2653, w_081_2654, w_081_2655, w_081_2658, w_081_2660, w_081_2663, w_081_2666, w_081_2667, w_081_2668, w_081_2670, w_081_2671, w_081_2673, w_081_2674, w_081_2676, w_081_2677, w_081_2682, w_081_2684, w_081_2686, w_081_2689, w_081_2690, w_081_2691, w_081_2692, w_081_2694, w_081_2697, w_081_2698, w_081_2699, w_081_2700, w_081_2701, w_081_2702, w_081_2703, w_081_2707, w_081_2711, w_081_2713, w_081_2714, w_081_2717, w_081_2719, w_081_2720, w_081_2722, w_081_2723, w_081_2729, w_081_2730, w_081_2731, w_081_2732, w_081_2734, w_081_2736, w_081_2737, w_081_2742, w_081_2743, w_081_2748, w_081_2749, w_081_2750, w_081_2753, w_081_2755, w_081_2757, w_081_2763, w_081_2766, w_081_2768, w_081_2770, w_081_2772, w_081_2775, w_081_2776, w_081_2777, w_081_2779, w_081_2781, w_081_2782, w_081_2785, w_081_2786, w_081_2787, w_081_2788, w_081_2791, w_081_2793, w_081_2794, w_081_2795, w_081_2798, w_081_2799, w_081_2800, w_081_2801, w_081_2802, w_081_2806, w_081_2808, w_081_2809, w_081_2810, w_081_2811, w_081_2813, w_081_2815, w_081_2817, w_081_2818, w_081_2819, w_081_2820, w_081_2821, w_081_2829, w_081_2831, w_081_2833, w_081_2834, w_081_2835, w_081_2836, w_081_2837, w_081_2838, w_081_2839, w_081_2844, w_081_2845, w_081_2848, w_081_2852, w_081_2853, w_081_2854, w_081_2855, w_081_2856, w_081_2857, w_081_2859, w_081_2862, w_081_2865, w_081_2867, w_081_2868, w_081_2869, w_081_2870, w_081_2872, w_081_2873, w_081_2876, w_081_2878, w_081_2882, w_081_2884, w_081_2888, w_081_2892, w_081_2894, w_081_2895, w_081_2899, w_081_2901, w_081_2905, w_081_2908, w_081_2912, w_081_2913, w_081_2914, w_081_2920, w_081_2924, w_081_2926, w_081_2927, w_081_2928, w_081_2929, w_081_2931, w_081_2934, w_081_2935, w_081_2936, w_081_2937, w_081_2938, w_081_2939, w_081_2942, w_081_2943, w_081_2944, w_081_2945, w_081_2948, w_081_2949, w_081_2950, w_081_2951, w_081_2953, w_081_2954, w_081_2957, w_081_2959, w_081_2960, w_081_2961, w_081_2963, w_081_2964, w_081_2965, w_081_2970, w_081_2971, w_081_2972, w_081_2983, w_081_2993, w_081_2995, w_081_2999, w_081_3002, w_081_3004, w_081_3007, w_081_3011, w_081_3014, w_081_3016, w_081_3017, w_081_3018, w_081_3019, w_081_3021, w_081_3022, w_081_3023, w_081_3029, w_081_3030, w_081_3032, w_081_3037, w_081_3038, w_081_3039, w_081_3044, w_081_3047, w_081_3048, w_081_3049, w_081_3051, w_081_3053, w_081_3054, w_081_3056, w_081_3057, w_081_3058, w_081_3059, w_081_3061, w_081_3062, w_081_3064, w_081_3066, w_081_3067, w_081_3068, w_081_3069, w_081_3073, w_081_3074, w_081_3077, w_081_3078, w_081_3082, w_081_3083, w_081_3084, w_081_3085, w_081_3088, w_081_3090, w_081_3091, w_081_3096, w_081_3098, w_081_3099, w_081_3106, w_081_3108, w_081_3109, w_081_3110, w_081_3112, w_081_3113, w_081_3117, w_081_3118, w_081_3120, w_081_3122, w_081_3124, w_081_3125, w_081_3127, w_081_3130, w_081_3134, w_081_3135, w_081_3140, w_081_3141, w_081_3143, w_081_3145, w_081_3146, w_081_3148, w_081_3151, w_081_3152, w_081_3162, w_081_3163, w_081_3164, w_081_3166, w_081_3171, w_081_3172, w_081_3176, w_081_3178, w_081_3179, w_081_3180, w_081_3186, w_081_3187, w_081_3191, w_081_3192, w_081_3193, w_081_3194, w_081_3201, w_081_3204, w_081_3205, w_081_3207, w_081_3209, w_081_3212, w_081_3214, w_081_3215, w_081_3216, w_081_3217, w_081_3218, w_081_3219, w_081_3222, w_081_3223, w_081_3225, w_081_3226, w_081_3230, w_081_3233, w_081_3234, w_081_3235, w_081_3236, w_081_3237, w_081_3239, w_081_3240, w_081_3242, w_081_3248, w_081_3250, w_081_3254, w_081_3255, w_081_3256, w_081_3257, w_081_3259, w_081_3260, w_081_3261, w_081_3265, w_081_3266, w_081_3268, w_081_3273, w_081_3277, w_081_3278, w_081_3279, w_081_3284, w_081_3285, w_081_3286, w_081_3288, w_081_3295, w_081_3298, w_081_3300, w_081_3301, w_081_3304, w_081_3307, w_081_3308, w_081_3309, w_081_3313, w_081_3314, w_081_3315, w_081_3317, w_081_3318, w_081_3320, w_081_3324, w_081_3327, w_081_3330, w_081_3331, w_081_3332, w_081_3336, w_081_3338, w_081_3339, w_081_3340, w_081_3341, w_081_3342, w_081_3343, w_081_3345, w_081_3347, w_081_3348, w_081_3349, w_081_3350, w_081_3353, w_081_3354, w_081_3356, w_081_3360, w_081_3361, w_081_3364, w_081_3368, w_081_3372, w_081_3374, w_081_3375, w_081_3376, w_081_3378, w_081_3379, w_081_3381, w_081_3382, w_081_3383, w_081_3385, w_081_3386, w_081_3387, w_081_3388, w_081_3389, w_081_3390, w_081_3391, w_081_3392, w_081_3394, w_081_3395, w_081_3396, w_081_3400, w_081_3402, w_081_3406, w_081_3410, w_081_3414, w_081_3415, w_081_3418, w_081_3419, w_081_3422, w_081_3423, w_081_3425, w_081_3427, w_081_3428, w_081_3431, w_081_3433, w_081_3434, w_081_3435, w_081_3437, w_081_3439, w_081_3442, w_081_3448, w_081_3450, w_081_3451, w_081_3454, w_081_3460, w_081_3462, w_081_3465, w_081_3466, w_081_3468, w_081_3469, w_081_3470, w_081_3474, w_081_3477, w_081_3479, w_081_3480, w_081_3482, w_081_3483, w_081_3490, w_081_3492, w_081_3494, w_081_3495, w_081_3499, w_081_3500, w_081_3501, w_081_3502, w_081_3504, w_081_3505, w_081_3506, w_081_3509, w_081_3510, w_081_3512, w_081_3513, w_081_3516, w_081_3518, w_081_3522, w_081_3525, w_081_3532, w_081_3533, w_081_3536, w_081_3539, w_081_3540, w_081_3541, w_081_3542, w_081_3543, w_081_3544, w_081_3546, w_081_3548, w_081_3549, w_081_3551, w_081_3552, w_081_3553, w_081_3554, w_081_3555, w_081_3560, w_081_3562, w_081_3567, w_081_3568, w_081_3569, w_081_3570, w_081_3571, w_081_3572, w_081_3575, w_081_3577, w_081_3580, w_081_3582, w_081_3584, w_081_3585, w_081_3586, w_081_3587, w_081_3588, w_081_3593, w_081_3596, w_081_3597, w_081_3598, w_081_3599, w_081_3601, w_081_3602, w_081_3603, w_081_3605, w_081_3606, w_081_3607, w_081_3610, w_081_3611, w_081_3612, w_081_3613, w_081_3617, w_081_3618, w_081_3620, w_081_3621, w_081_3623, w_081_3626, w_081_3632, w_081_3637, w_081_3638, w_081_3639, w_081_3640, w_081_3650, w_081_3654, w_081_3655, w_081_3656, w_081_3660, w_081_3662, w_081_3665, w_081_3668, w_081_3670, w_081_3673, w_081_3679, w_081_3680, w_081_3682, w_081_3683, w_081_3686, w_081_3688, w_081_3689, w_081_3690, w_081_3691, w_081_3692, w_081_3693, w_081_3698, w_081_3701, w_081_3704, w_081_3705, w_081_3708, w_081_3709, w_081_3710, w_081_3714, w_081_3715, w_081_3716, w_081_3718, w_081_3719, w_081_3720, w_081_3724, w_081_3725, w_081_3726, w_081_3728, w_081_3733, w_081_3734, w_081_3735, w_081_3736, w_081_3737, w_081_3738, w_081_3739, w_081_3740, w_081_3741, w_081_3746, w_081_3748, w_081_3751, w_081_3756, w_081_3757, w_081_3759, w_081_3762, w_081_3764, w_081_3766, w_081_3767, w_081_3769, w_081_3771, w_081_3778, w_081_3779, w_081_3782, w_081_3784, w_081_3787, w_081_3788, w_081_3790, w_081_3791, w_081_3794, w_081_3796, w_081_3798, w_081_3801, w_081_3804, w_081_3805, w_081_3806, w_081_3807, w_081_3814, w_081_3816, w_081_3817, w_081_3819, w_081_3820, w_081_3821, w_081_3822, w_081_3823, w_081_3824, w_081_3825, w_081_3826, w_081_3831, w_081_3832, w_081_3833, w_081_3835, w_081_3836, w_081_3837, w_081_3843, w_081_3844, w_081_3845, w_081_3848, w_081_3849, w_081_3855, w_081_3857, w_081_3864, w_081_3865, w_081_3867, w_081_3869, w_081_3872, w_081_3873, w_081_3875, w_081_3878, w_081_3879, w_081_3880, w_081_3881, w_081_3883, w_081_3884, w_081_3887, w_081_3888, w_081_3894, w_081_3895, w_081_3898, w_081_3899, w_081_3900, w_081_3901, w_081_3902, w_081_3905, w_081_3907, w_081_3908, w_081_3912, w_081_3914, w_081_3915, w_081_3916, w_081_3918, w_081_3919, w_081_3927, w_081_3934, w_081_3936, w_081_3938, w_081_3940, w_081_3944, w_081_3945, w_081_3946, w_081_3947, w_081_3948, w_081_3949, w_081_3952, w_081_3955, w_081_3957, w_081_3958, w_081_3959, w_081_3961, w_081_3962, w_081_3963, w_081_3967, w_081_3968, w_081_3969, w_081_3970, w_081_3971, w_081_3972, w_081_3976, w_081_3977, w_081_3980, w_081_3983, w_081_3987, w_081_3989, w_081_3990, w_081_3991, w_081_3992, w_081_3993, w_081_3994, w_081_3995, w_081_3997, w_081_4005, w_081_4008, w_081_4013, w_081_4015, w_081_4016, w_081_4022, w_081_4023, w_081_4025, w_081_4026, w_081_4028, w_081_4031, w_081_4033, w_081_4038, w_081_4040, w_081_4042, w_081_4045, w_081_4048, w_081_4050, w_081_4052, w_081_4056, w_081_4057, w_081_4059, w_081_4060, w_081_4061, w_081_4062, w_081_4063, w_081_4065, w_081_4066, w_081_4067, w_081_4070, w_081_4072, w_081_4073, w_081_4075, w_081_4076, w_081_4077, w_081_4078, w_081_4082, w_081_4083, w_081_4084, w_081_4087, w_081_4088, w_081_4091, w_081_4093, w_081_4095, w_081_4097, w_081_4106, w_081_4107, w_081_4108, w_081_4112, w_081_4116, w_081_4119, w_081_4120, w_081_4121, w_081_4123, w_081_4125, w_081_4127, w_081_4129, w_081_4132, w_081_4134, w_081_4135, w_081_4137, w_081_4140, w_081_4141, w_081_4145, w_081_4147, w_081_4149, w_081_4150, w_081_4151, w_081_4152, w_081_4154, w_081_4158, w_081_4161, w_081_4163, w_081_4164, w_081_4168, w_081_4171, w_081_4172, w_081_4173, w_081_4175, w_081_4176, w_081_4179, w_081_4180, w_081_4181, w_081_4185, w_081_4186, w_081_4187, w_081_4190, w_081_4194, w_081_4195, w_081_4197, w_081_4198, w_081_4199, w_081_4200, w_081_4203, w_081_4205, w_081_4207, w_081_4208, w_081_4211, w_081_4213, w_081_4215, w_081_4216, w_081_4220, w_081_4221, w_081_4223, w_081_4224, w_081_4226, w_081_4227, w_081_4229, w_081_4230, w_081_4232, w_081_4236, w_081_4237, w_081_4239, w_081_4247, w_081_4248, w_081_4253, w_081_4254, w_081_4255, w_081_4258, w_081_4260, w_081_4261, w_081_4263, w_081_4264, w_081_4266, w_081_4267, w_081_4268, w_081_4270, w_081_4271, w_081_4273, w_081_4275, w_081_4276, w_081_4279, w_081_4280, w_081_4281, w_081_4282, w_081_4283, w_081_4284, w_081_4285, w_081_4287, w_081_4288, w_081_4289, w_081_4294, w_081_4295, w_081_4296, w_081_4299, w_081_4300, w_081_4301, w_081_4302, w_081_4305, w_081_4307, w_081_4310, w_081_4315, w_081_4321, w_081_4324, w_081_4326, w_081_4329, w_081_4330, w_081_4335, w_081_4336, w_081_4340, w_081_4341, w_081_4342, w_081_4348, w_081_4350, w_081_4353, w_081_4355, w_081_4357, w_081_4358, w_081_4361, w_081_4362, w_081_4363, w_081_4367, w_081_4369, w_081_4371, w_081_4373, w_081_4377, w_081_4379, w_081_4382, w_081_4386, w_081_4390, w_081_4391, w_081_4394, w_081_4396, w_081_4399, w_081_4404, w_081_4406, w_081_4407, w_081_4412, w_081_4414, w_081_4415, w_081_4417, w_081_4418, w_081_4424, w_081_4426, w_081_4428, w_081_4429, w_081_4430, w_081_4431, w_081_4432, w_081_4434, w_081_4437, w_081_4438, w_081_4442, w_081_4443, w_081_4444, w_081_4446, w_081_4447, w_081_4450, w_081_4452, w_081_4456, w_081_4457, w_081_4460, w_081_4461, w_081_4468, w_081_4472, w_081_4475, w_081_4476, w_081_4477, w_081_4478, w_081_4482, w_081_4486, w_081_4489, w_081_4490, w_081_4491, w_081_4493, w_081_4495, w_081_4496, w_081_4497, w_081_4498, w_081_4499, w_081_4500, w_081_4502, w_081_4503, w_081_4504, w_081_4505, w_081_4506, w_081_4507, w_081_4509, w_081_4512, w_081_4513, w_081_4518, w_081_4519, w_081_4520, w_081_4521, w_081_4522, w_081_4523, w_081_4524, w_081_4533, w_081_4534, w_081_4535, w_081_4537, w_081_4538, w_081_4539, w_081_4540, w_081_4541, w_081_4546, w_081_4547, w_081_4553, w_081_4554, w_081_4556, w_081_4557, w_081_4559, w_081_4562, w_081_4563, w_081_4565, w_081_4568, w_081_4573, w_081_4574, w_081_4575, w_081_4579, w_081_4580, w_081_4582, w_081_4588, w_081_4591, w_081_4592, w_081_4595, w_081_4597, w_081_4601, w_081_4603, w_081_4605, w_081_4606, w_081_4607, w_081_4608, w_081_4611, w_081_4612, w_081_4613, w_081_4615, w_081_4620, w_081_4621, w_081_4626, w_081_4627, w_081_4628, w_081_4629, w_081_4634, w_081_4638, w_081_4651, w_081_4654, w_081_4656, w_081_4657, w_081_4658, w_081_4659, w_081_4664, w_081_4668, w_081_4674, w_081_4675, w_081_4678, w_081_4679, w_081_4680, w_081_4687, w_081_4690, w_081_4691, w_081_4693, w_081_4695, w_081_4699, w_081_4700, w_081_4712, w_081_4714, w_081_4720, w_081_4722, w_081_4724, w_081_4726, w_081_4728, w_081_4732, w_081_4733, w_081_4744, w_081_4749, w_081_4751, w_081_4755, w_081_4762, w_081_4770, w_081_4772, w_081_4774, w_081_4775, w_081_4780, w_081_4788, w_081_4793, w_081_4796, w_081_4806, w_081_4812, w_081_4822, w_081_4827, w_081_4828, w_081_4830, w_081_4833, w_081_4834, w_081_4835, w_081_4838, w_081_4839, w_081_4840, w_081_4843, w_081_4851, w_081_4853, w_081_4854, w_081_4856, w_081_4857, w_081_4862, w_081_4865, w_081_4866, w_081_4870, w_081_4879, w_081_4882, w_081_4888, w_081_4896, w_081_4899, w_081_4904, w_081_4905, w_081_4906, w_081_4907, w_081_4910, w_081_4913, w_081_4914, w_081_4916, w_081_4917, w_081_4921, w_081_4922, w_081_4926, w_081_4927, w_081_4945, w_081_4949, w_081_4952, w_081_4959, w_081_4963, w_081_4968, w_081_4977, w_081_4978, w_081_4979, w_081_4980, w_081_4986, w_081_4987, w_081_4989, w_081_4994, w_081_4997, w_081_5000, w_081_5001, w_081_5004, w_081_5005, w_081_5008, w_081_5012, w_081_5014, w_081_5019, w_081_5020, w_081_5025, w_081_5027, w_081_5029, w_081_5031, w_081_5035, w_081_5036, w_081_5037, w_081_5039, w_081_5040, w_081_5041, w_081_5043, w_081_5045, w_081_5052, w_081_5053, w_081_5056, w_081_5058, w_081_5059, w_081_5063, w_081_5067, w_081_5078, w_081_5083, w_081_5095, w_081_5096, w_081_5103, w_081_5106, w_081_5112, w_081_5115, w_081_5118, w_081_5119, w_081_5120, w_081_5128, w_081_5129, w_081_5130, w_081_5132, w_081_5134, w_081_5136, w_081_5147, w_081_5148, w_081_5149, w_081_5154, w_081_5157, w_081_5158, w_081_5164, w_081_5169, w_081_5175, w_081_5181, w_081_5182, w_081_5183, w_081_5186, w_081_5193, w_081_5195, w_081_5207, w_081_5213, w_081_5220, w_081_5221, w_081_5230, w_081_5232, w_081_5240, w_081_5241, w_081_5243, w_081_5256, w_081_5257, w_081_5260, w_081_5261, w_081_5266, w_081_5271, w_081_5273, w_081_5285, w_081_5288, w_081_5291, w_081_5292, w_081_5294, w_081_5299, w_081_5301, w_081_5308, w_081_5310, w_081_5312, w_081_5315, w_081_5327, w_081_5333, w_081_5336, w_081_5337, w_081_5340, w_081_5341, w_081_5344, w_081_5351, w_081_5352, w_081_5353, w_081_5356, w_081_5361, w_081_5362, w_081_5365, w_081_5369, w_081_5373, w_081_5377, w_081_5381, w_081_5383;
  wire w_082_000, w_082_001, w_082_002, w_082_003, w_082_005, w_082_010, w_082_011, w_082_013, w_082_014, w_082_016, w_082_017, w_082_020, w_082_023, w_082_025, w_082_026, w_082_028, w_082_029, w_082_032, w_082_036, w_082_038, w_082_044, w_082_045, w_082_048, w_082_049, w_082_050, w_082_053, w_082_054, w_082_061, w_082_062, w_082_071, w_082_074, w_082_075, w_082_077, w_082_078, w_082_079, w_082_080, w_082_081, w_082_082, w_082_083, w_082_084, w_082_087, w_082_088, w_082_091, w_082_094, w_082_095, w_082_096, w_082_098, w_082_099, w_082_102, w_082_105, w_082_107, w_082_108, w_082_110, w_082_111, w_082_112, w_082_114, w_082_115, w_082_117, w_082_118, w_082_119, w_082_121, w_082_122, w_082_123, w_082_124, w_082_127, w_082_132, w_082_133, w_082_134, w_082_135, w_082_137, w_082_138, w_082_140, w_082_141, w_082_144, w_082_145, w_082_146, w_082_147, w_082_149, w_082_153, w_082_156, w_082_157, w_082_158, w_082_160, w_082_161, w_082_163, w_082_164, w_082_165, w_082_166, w_082_167, w_082_168, w_082_170, w_082_172, w_082_174, w_082_180, w_082_181, w_082_182, w_082_183, w_082_185, w_082_186, w_082_187, w_082_190, w_082_191, w_082_192, w_082_194, w_082_196, w_082_199, w_082_200, w_082_201, w_082_204, w_082_205, w_082_206, w_082_208, w_082_210, w_082_211, w_082_212, w_082_214, w_082_215, w_082_216, w_082_217, w_082_220, w_082_224, w_082_225, w_082_226, w_082_227, w_082_229, w_082_231, w_082_233, w_082_235, w_082_237, w_082_239, w_082_240, w_082_243, w_082_245, w_082_246, w_082_247, w_082_248, w_082_249, w_082_250, w_082_252, w_082_253, w_082_255, w_082_256, w_082_257, w_082_258, w_082_261, w_082_262, w_082_263, w_082_264, w_082_266, w_082_267, w_082_268, w_082_269, w_082_272, w_082_273, w_082_274, w_082_276, w_082_278, w_082_279, w_082_283, w_082_284, w_082_285, w_082_286, w_082_287, w_082_289, w_082_290, w_082_293, w_082_295, w_082_296, w_082_297, w_082_298, w_082_299, w_082_300, w_082_301, w_082_302, w_082_305, w_082_307, w_082_308, w_082_310, w_082_311, w_082_313, w_082_316, w_082_317, w_082_319, w_082_322, w_082_323, w_082_324, w_082_325, w_082_327, w_082_330, w_082_332, w_082_333, w_082_340, w_082_341, w_082_342, w_082_344, w_082_347, w_082_348, w_082_349, w_082_350, w_082_354, w_082_355, w_082_357, w_082_358, w_082_359, w_082_360, w_082_361, w_082_362, w_082_365, w_082_367, w_082_368, w_082_369, w_082_370, w_082_371, w_082_375, w_082_376, w_082_378, w_082_379, w_082_380, w_082_381, w_082_382, w_082_386, w_082_387, w_082_388, w_082_391, w_082_392, w_082_393, w_082_394, w_082_395, w_082_397, w_082_399, w_082_400, w_082_401, w_082_402, w_082_408, w_082_409, w_082_410, w_082_414, w_082_416, w_082_417, w_082_418, w_082_421, w_082_422, w_082_424, w_082_426, w_082_428, w_082_429, w_082_430, w_082_432, w_082_434, w_082_435, w_082_437, w_082_439, w_082_440, w_082_442, w_082_443, w_082_445, w_082_447, w_082_449, w_082_450, w_082_452, w_082_454, w_082_455, w_082_456, w_082_460, w_082_462, w_082_464, w_082_465, w_082_468, w_082_471, w_082_472, w_082_473, w_082_475, w_082_477, w_082_479, w_082_482, w_082_484, w_082_486, w_082_487, w_082_488, w_082_489, w_082_492, w_082_494, w_082_496, w_082_497, w_082_498, w_082_501, w_082_502, w_082_503, w_082_504, w_082_505, w_082_507, w_082_509, w_082_510, w_082_512, w_082_513, w_082_514, w_082_515, w_082_516, w_082_519, w_082_521, w_082_523, w_082_524, w_082_525, w_082_526, w_082_528, w_082_529, w_082_530, w_082_531, w_082_533, w_082_535, w_082_536, w_082_538, w_082_539, w_082_540, w_082_541, w_082_544, w_082_545, w_082_547, w_082_550, w_082_552, w_082_553, w_082_554, w_082_555, w_082_556, w_082_560, w_082_562, w_082_563, w_082_565, w_082_566, w_082_567, w_082_568, w_082_569, w_082_570, w_082_571, w_082_572, w_082_573, w_082_574, w_082_575, w_082_579, w_082_584, w_082_585, w_082_586, w_082_587, w_082_588, w_082_590, w_082_591, w_082_592, w_082_595, w_082_599, w_082_600, w_082_602, w_082_605, w_082_607, w_082_609, w_082_613, w_082_615, w_082_616, w_082_617, w_082_619, w_082_620, w_082_623, w_082_624, w_082_625, w_082_626, w_082_630, w_082_631, w_082_633, w_082_635, w_082_636, w_082_637, w_082_638, w_082_641, w_082_642, w_082_643, w_082_644, w_082_645, w_082_647, w_082_649, w_082_650, w_082_651, w_082_653, w_082_654, w_082_655, w_082_656, w_082_658, w_082_662, w_082_664, w_082_666, w_082_667, w_082_668, w_082_670, w_082_672, w_082_673, w_082_674, w_082_675, w_082_676, w_082_677, w_082_678, w_082_680, w_082_682, w_082_683, w_082_684, w_082_685, w_082_686, w_082_687, w_082_688, w_082_689, w_082_692, w_082_693, w_082_696, w_082_697, w_082_698, w_082_700, w_082_701, w_082_704, w_082_706, w_082_707, w_082_712, w_082_715, w_082_716, w_082_717, w_082_720, w_082_722, w_082_723, w_082_724, w_082_726, w_082_730, w_082_733, w_082_736, w_082_738, w_082_739, w_082_740, w_082_742, w_082_743, w_082_744, w_082_746, w_082_747, w_082_749, w_082_752, w_082_753, w_082_754, w_082_756, w_082_757, w_082_759, w_082_760, w_082_764, w_082_765, w_082_766, w_082_767, w_082_769, w_082_771, w_082_773, w_082_774, w_082_775, w_082_777, w_082_779, w_082_783, w_082_784, w_082_785, w_082_788, w_082_789, w_082_790, w_082_792, w_082_793, w_082_796, w_082_798, w_082_799, w_082_800, w_082_802, w_082_804, w_082_806, w_082_807, w_082_808, w_082_809, w_082_812, w_082_813, w_082_814, w_082_818, w_082_819, w_082_821, w_082_823, w_082_824, w_082_825, w_082_827, w_082_828, w_082_830, w_082_832, w_082_833, w_082_834, w_082_838, w_082_839, w_082_840, w_082_842, w_082_844, w_082_845, w_082_846, w_082_847, w_082_853, w_082_855, w_082_856, w_082_858, w_082_860, w_082_861, w_082_866, w_082_867, w_082_868, w_082_870, w_082_873, w_082_874, w_082_875, w_082_879, w_082_881, w_082_883, w_082_884, w_082_885, w_082_886, w_082_890, w_082_891, w_082_892, w_082_894, w_082_898, w_082_900, w_082_905, w_082_907, w_082_909, w_082_912, w_082_915, w_082_916, w_082_917, w_082_919, w_082_921, w_082_922, w_082_924, w_082_926, w_082_927, w_082_930, w_082_931, w_082_932, w_082_934, w_082_935, w_082_939, w_082_940, w_082_942, w_082_946, w_082_947, w_082_948, w_082_949, w_082_950, w_082_954, w_082_955, w_082_958, w_082_959, w_082_960, w_082_961, w_082_964, w_082_966, w_082_967, w_082_968, w_082_971, w_082_973, w_082_975, w_082_976, w_082_977, w_082_978, w_082_981, w_082_983, w_082_984, w_082_985, w_082_986, w_082_987, w_082_988, w_082_990, w_082_991, w_082_994, w_082_995, w_082_996, w_082_997, w_082_998, w_082_999, w_082_1001, w_082_1002, w_082_1003, w_082_1004, w_082_1010, w_082_1014, w_082_1016, w_082_1018, w_082_1019, w_082_1020, w_082_1021, w_082_1022, w_082_1023, w_082_1024, w_082_1026, w_082_1028, w_082_1029, w_082_1030, w_082_1031, w_082_1032, w_082_1033, w_082_1034, w_082_1035, w_082_1037, w_082_1038, w_082_1042, w_082_1043, w_082_1044, w_082_1045, w_082_1046, w_082_1047, w_082_1048, w_082_1050, w_082_1051, w_082_1052, w_082_1056, w_082_1057, w_082_1059, w_082_1064, w_082_1065, w_082_1066, w_082_1067, w_082_1068, w_082_1069, w_082_1070, w_082_1073, w_082_1076, w_082_1078, w_082_1079, w_082_1080, w_082_1081, w_082_1084, w_082_1088, w_082_1092, w_082_1093, w_082_1095, w_082_1098, w_082_1100, w_082_1101, w_082_1103, w_082_1104, w_082_1105, w_082_1106, w_082_1107, w_082_1110, w_082_1112, w_082_1113, w_082_1114, w_082_1116, w_082_1117, w_082_1118, w_082_1121, w_082_1126, w_082_1130, w_082_1132, w_082_1133, w_082_1134, w_082_1135, w_082_1139, w_082_1141, w_082_1142, w_082_1145, w_082_1150, w_082_1152, w_082_1157, w_082_1159, w_082_1164, w_082_1165, w_082_1167, w_082_1168, w_082_1170, w_082_1173, w_082_1183, w_082_1185, w_082_1186, w_082_1190, w_082_1192, w_082_1195, w_082_1196, w_082_1197, w_082_1200, w_082_1202, w_082_1204, w_082_1206, w_082_1207, w_082_1209, w_082_1210, w_082_1211, w_082_1212, w_082_1216, w_082_1218, w_082_1221, w_082_1222, w_082_1224, w_082_1229, w_082_1230, w_082_1232, w_082_1233, w_082_1235, w_082_1236, w_082_1237, w_082_1242, w_082_1243, w_082_1245, w_082_1249, w_082_1252, w_082_1253, w_082_1254, w_082_1257, w_082_1258, w_082_1259, w_082_1260, w_082_1263, w_082_1267, w_082_1269, w_082_1271, w_082_1274, w_082_1275, w_082_1276, w_082_1279, w_082_1280, w_082_1283, w_082_1285, w_082_1286, w_082_1290, w_082_1291, w_082_1294, w_082_1295, w_082_1296, w_082_1298, w_082_1299, w_082_1300, w_082_1302, w_082_1307, w_082_1311, w_082_1313, w_082_1314, w_082_1316, w_082_1318, w_082_1320, w_082_1322, w_082_1323, w_082_1327, w_082_1329, w_082_1332, w_082_1333, w_082_1334, w_082_1335, w_082_1336, w_082_1338, w_082_1342, w_082_1343, w_082_1344, w_082_1346, w_082_1347, w_082_1348, w_082_1349, w_082_1350, w_082_1351, w_082_1352, w_082_1355, w_082_1359, w_082_1360, w_082_1362, w_082_1363, w_082_1364, w_082_1367, w_082_1368, w_082_1375, w_082_1379, w_082_1381, w_082_1382, w_082_1383, w_082_1384, w_082_1386, w_082_1389, w_082_1392, w_082_1394, w_082_1398, w_082_1399, w_082_1400, w_082_1401, w_082_1404, w_082_1405, w_082_1409, w_082_1412, w_082_1414, w_082_1417, w_082_1418, w_082_1423, w_082_1424, w_082_1425, w_082_1429, w_082_1431, w_082_1432, w_082_1433, w_082_1436, w_082_1437, w_082_1438, w_082_1448, w_082_1449, w_082_1451, w_082_1452, w_082_1456, w_082_1457, w_082_1461, w_082_1464, w_082_1470, w_082_1475, w_082_1478, w_082_1480, w_082_1481, w_082_1490, w_082_1491, w_082_1492, w_082_1493, w_082_1494, w_082_1495, w_082_1497, w_082_1498, w_082_1500, w_082_1502, w_082_1503, w_082_1505, w_082_1510, w_082_1511, w_082_1512, w_082_1513, w_082_1515, w_082_1516, w_082_1517, w_082_1518, w_082_1519, w_082_1520, w_082_1522, w_082_1525, w_082_1528, w_082_1530, w_082_1531, w_082_1532, w_082_1533, w_082_1538, w_082_1540, w_082_1541, w_082_1542, w_082_1545, w_082_1546, w_082_1547, w_082_1548, w_082_1549, w_082_1550, w_082_1551, w_082_1553, w_082_1557, w_082_1559, w_082_1560, w_082_1561, w_082_1565, w_082_1566, w_082_1569, w_082_1570, w_082_1573, w_082_1575, w_082_1577, w_082_1578, w_082_1582, w_082_1583, w_082_1587, w_082_1589, w_082_1591, w_082_1593, w_082_1594, w_082_1595, w_082_1596, w_082_1597, w_082_1598, w_082_1600, w_082_1603, w_082_1604, w_082_1606, w_082_1607, w_082_1608, w_082_1613, w_082_1614, w_082_1618, w_082_1619, w_082_1622, w_082_1626, w_082_1630, w_082_1631, w_082_1632, w_082_1633, w_082_1635, w_082_1638, w_082_1643, w_082_1647, w_082_1648, w_082_1651, w_082_1652, w_082_1656, w_082_1657, w_082_1659, w_082_1660, w_082_1661, w_082_1662, w_082_1666, w_082_1667, w_082_1668, w_082_1669, w_082_1670, w_082_1671, w_082_1672, w_082_1674, w_082_1676, w_082_1678, w_082_1679, w_082_1680, w_082_1681, w_082_1685, w_082_1687, w_082_1688, w_082_1689, w_082_1691, w_082_1692, w_082_1696, w_082_1697, w_082_1700, w_082_1701, w_082_1702, w_082_1709, w_082_1714, w_082_1716, w_082_1719, w_082_1724, w_082_1725, w_082_1728, w_082_1730, w_082_1731, w_082_1732, w_082_1733, w_082_1735, w_082_1736, w_082_1740, w_082_1744, w_082_1745, w_082_1746, w_082_1747, w_082_1748, w_082_1749, w_082_1750, w_082_1752, w_082_1753, w_082_1756, w_082_1758, w_082_1761, w_082_1762, w_082_1763, w_082_1764, w_082_1765, w_082_1766, w_082_1767, w_082_1771, w_082_1774, w_082_1777, w_082_1779, w_082_1783, w_082_1784, w_082_1788, w_082_1789, w_082_1791, w_082_1792, w_082_1794, w_082_1795, w_082_1796, w_082_1799, w_082_1800, w_082_1803, w_082_1804, w_082_1807, w_082_1811, w_082_1815, w_082_1817, w_082_1818, w_082_1821, w_082_1822, w_082_1825, w_082_1834, w_082_1835, w_082_1836, w_082_1841, w_082_1843, w_082_1844, w_082_1846, w_082_1848, w_082_1849, w_082_1852, w_082_1854, w_082_1855, w_082_1857, w_082_1858, w_082_1862, w_082_1864, w_082_1865, w_082_1866, w_082_1868, w_082_1870, w_082_1871, w_082_1872, w_082_1875, w_082_1880, w_082_1881, w_082_1882, w_082_1883, w_082_1884, w_082_1885, w_082_1887, w_082_1888, w_082_1890, w_082_1891, w_082_1893, w_082_1896, w_082_1898, w_082_1902, w_082_1903, w_082_1907, w_082_1908, w_082_1911, w_082_1912, w_082_1914, w_082_1916, w_082_1921, w_082_1922, w_082_1923, w_082_1927, w_082_1932, w_082_1937, w_082_1939, w_082_1940, w_082_1942, w_082_1946, w_082_1951, w_082_1952, w_082_1953, w_082_1954, w_082_1955, w_082_1959, w_082_1961, w_082_1962, w_082_1963, w_082_1970, w_082_1973, w_082_1974, w_082_1979, w_082_1980, w_082_1982, w_082_1983, w_082_1987, w_082_1988, w_082_1990, w_082_1992, w_082_1993, w_082_1994, w_082_1996, w_082_1998, w_082_1999, w_082_2001, w_082_2003, w_082_2006, w_082_2007, w_082_2011, w_082_2012, w_082_2017, w_082_2019, w_082_2020, w_082_2021, w_082_2022, w_082_2024, w_082_2028, w_082_2030, w_082_2031, w_082_2035, w_082_2037, w_082_2038, w_082_2040, w_082_2041, w_082_2043, w_082_2044, w_082_2047, w_082_2049, w_082_2050, w_082_2051, w_082_2054, w_082_2057, w_082_2058, w_082_2059, w_082_2060, w_082_2061, w_082_2065, w_082_2068, w_082_2071, w_082_2072, w_082_2076, w_082_2079, w_082_2084, w_082_2085, w_082_2088, w_082_2090, w_082_2091, w_082_2092, w_082_2095, w_082_2096, w_082_2099, w_082_2107, w_082_2108, w_082_2110, w_082_2114, w_082_2117, w_082_2119, w_082_2120, w_082_2121, w_082_2122, w_082_2123, w_082_2126, w_082_2132, w_082_2136, w_082_2137, w_082_2138, w_082_2139, w_082_2140, w_082_2141, w_082_2142, w_082_2143, w_082_2145, w_082_2149, w_082_2150, w_082_2152, w_082_2154, w_082_2155, w_082_2156, w_082_2158, w_082_2160, w_082_2165, w_082_2167, w_082_2168, w_082_2171, w_082_2172, w_082_2173, w_082_2175, w_082_2179, w_082_2185, w_082_2187, w_082_2191, w_082_2193, w_082_2197, w_082_2198, w_082_2201, w_082_2206, w_082_2209, w_082_2211, w_082_2214, w_082_2216, w_082_2220, w_082_2225, w_082_2226, w_082_2227, w_082_2228, w_082_2230, w_082_2231, w_082_2234, w_082_2235, w_082_2236, w_082_2238, w_082_2239, w_082_2241, w_082_2244, w_082_2245, w_082_2247, w_082_2250, w_082_2251, w_082_2252, w_082_2253, w_082_2256, w_082_2258, w_082_2260, w_082_2263, w_082_2264, w_082_2273, w_082_2274, w_082_2275, w_082_2277, w_082_2278, w_082_2279, w_082_2283, w_082_2284, w_082_2286, w_082_2287, w_082_2291, w_082_2294, w_082_2295, w_082_2296, w_082_2301, w_082_2303, w_082_2305, w_082_2306, w_082_2307, w_082_2308, w_082_2312, w_082_2315, w_082_2316, w_082_2317, w_082_2324, w_082_2327, w_082_2329, w_082_2330, w_082_2332, w_082_2334, w_082_2335, w_082_2336, w_082_2340, w_082_2342, w_082_2343, w_082_2351, w_082_2353, w_082_2354, w_082_2357, w_082_2358, w_082_2359, w_082_2360, w_082_2361, w_082_2362, w_082_2367, w_082_2368, w_082_2370, w_082_2371, w_082_2373, w_082_2376, w_082_2379, w_082_2383, w_082_2384, w_082_2386, w_082_2388, w_082_2389, w_082_2390, w_082_2393, w_082_2396, w_082_2400, w_082_2401, w_082_2402, w_082_2403, w_082_2405, w_082_2406, w_082_2408, w_082_2409, w_082_2410, w_082_2412, w_082_2416, w_082_2418, w_082_2419, w_082_2420, w_082_2421, w_082_2422, w_082_2427, w_082_2432, w_082_2433, w_082_2437, w_082_2438, w_082_2440, w_082_2442, w_082_2443, w_082_2444, w_082_2447, w_082_2449, w_082_2454, w_082_2455, w_082_2456, w_082_2458, w_082_2459, w_082_2460, w_082_2462, w_082_2463, w_082_2466, w_082_2467, w_082_2472, w_082_2473, w_082_2474, w_082_2482, w_082_2483, w_082_2484, w_082_2486, w_082_2489, w_082_2493, w_082_2494, w_082_2498, w_082_2500, w_082_2501, w_082_2509, w_082_2511, w_082_2512, w_082_2513, w_082_2514, w_082_2515, w_082_2518, w_082_2519, w_082_2521, w_082_2523, w_082_2525, w_082_2529, w_082_2531, w_082_2537, w_082_2539, w_082_2540, w_082_2542, w_082_2543, w_082_2546, w_082_2547, w_082_2549, w_082_2550, w_082_2551, w_082_2552, w_082_2555, w_082_2561, w_082_2563, w_082_2565, w_082_2566, w_082_2567, w_082_2569, w_082_2572, w_082_2574, w_082_2576, w_082_2580, w_082_2584, w_082_2587, w_082_2588, w_082_2590, w_082_2592, w_082_2594, w_082_2596, w_082_2597, w_082_2598, w_082_2602, w_082_2607, w_082_2608, w_082_2609, w_082_2612, w_082_2616, w_082_2617, w_082_2619, w_082_2621, w_082_2622, w_082_2623, w_082_2624, w_082_2625, w_082_2626, w_082_2628, w_082_2630, w_082_2631, w_082_2632, w_082_2636, w_082_2638, w_082_2640, w_082_2646, w_082_2648, w_082_2650, w_082_2651, w_082_2655, w_082_2657, w_082_2659, w_082_2660, w_082_2661, w_082_2662, w_082_2664, w_082_2666, w_082_2667, w_082_2676, w_082_2678, w_082_2679, w_082_2681, w_082_2682, w_082_2683, w_082_2685, w_082_2688, w_082_2691, w_082_2692, w_082_2693, w_082_2694, w_082_2695, w_082_2698, w_082_2699, w_082_2700, w_082_2703, w_082_2704, w_082_2713, w_082_2718, w_082_2719, w_082_2720, w_082_2722, w_082_2723, w_082_2726, w_082_2728, w_082_2729, w_082_2731, w_082_2733, w_082_2734, w_082_2737, w_082_2741, w_082_2742, w_082_2743, w_082_2747, w_082_2748, w_082_2750, w_082_2753, w_082_2754, w_082_2755, w_082_2757, w_082_2760, w_082_2763, w_082_2765, w_082_2766, w_082_2767, w_082_2768, w_082_2774, w_082_2776, w_082_2779, w_082_2780, w_082_2782, w_082_2785, w_082_2790, w_082_2793, w_082_2794, w_082_2795, w_082_2803, w_082_2804, w_082_2806, w_082_2807, w_082_2809, w_082_2810, w_082_2811, w_082_2813, w_082_2815, w_082_2816, w_082_2818, w_082_2820, w_082_2821, w_082_2822, w_082_2823, w_082_2828, w_082_2829, w_082_2832, w_082_2835, w_082_2838, w_082_2840, w_082_2842, w_082_2844, w_082_2846, w_082_2851, w_082_2859, w_082_2860, w_082_2864, w_082_2868, w_082_2871, w_082_2874, w_082_2876, w_082_2878, w_082_2879, w_082_2886, w_082_2887, w_082_2890, w_082_2891, w_082_2892, w_082_2894, w_082_2895, w_082_2896, w_082_2898, w_082_2899, w_082_2900, w_082_2903, w_082_2904, w_082_2905, w_082_2909, w_082_2911, w_082_2912, w_082_2915, w_082_2916, w_082_2919, w_082_2921, w_082_2922, w_082_2923, w_082_2926, w_082_2927, w_082_2928, w_082_2929, w_082_2930, w_082_2931, w_082_2932, w_082_2938, w_082_2939, w_082_2942, w_082_2944, w_082_2947, w_082_2949, w_082_2951, w_082_2952, w_082_2955, w_082_2956, w_082_2957, w_082_2958, w_082_2960, w_082_2961, w_082_2962, w_082_2964, w_082_2966, w_082_2967, w_082_2968, w_082_2970, w_082_2974, w_082_2979, w_082_2980, w_082_2981, w_082_2984, w_082_2990, w_082_2991, w_082_2994, w_082_2997, w_082_3001, w_082_3002, w_082_3003, w_082_3004, w_082_3011, w_082_3014, w_082_3015, w_082_3016, w_082_3020, w_082_3026, w_082_3027, w_082_3029, w_082_3030, w_082_3032, w_082_3035, w_082_3036, w_082_3039, w_082_3042, w_082_3043, w_082_3044, w_082_3045, w_082_3046, w_082_3054, w_082_3055, w_082_3056, w_082_3058, w_082_3061, w_082_3064, w_082_3066, w_082_3068, w_082_3069, w_082_3071, w_082_3074, w_082_3075, w_082_3076, w_082_3082, w_082_3084, w_082_3085, w_082_3092, w_082_3093, w_082_3095, w_082_3096, w_082_3098, w_082_3100, w_082_3101, w_082_3102, w_082_3103, w_082_3105, w_082_3107, w_082_3109, w_082_3111, w_082_3112, w_082_3115, w_082_3116, w_082_3119, w_082_3120, w_082_3124, w_082_3126, w_082_3132, w_082_3134, w_082_3137, w_082_3139, w_082_3140, w_082_3141, w_082_3144, w_082_3146, w_082_3147, w_082_3149, w_082_3153, w_082_3155, w_082_3158, w_082_3162, w_082_3163, w_082_3165, w_082_3167, w_082_3171, w_082_3173, w_082_3176, w_082_3177, w_082_3178, w_082_3180, w_082_3185, w_082_3186, w_082_3191, w_082_3193, w_082_3195, w_082_3196, w_082_3197, w_082_3198, w_082_3200, w_082_3201, w_082_3205, w_082_3207, w_082_3208, w_082_3209, w_082_3211, w_082_3214, w_082_3218, w_082_3219, w_082_3220, w_082_3221, w_082_3225, w_082_3226, w_082_3231, w_082_3232, w_082_3233, w_082_3234, w_082_3235, w_082_3242, w_082_3244, w_082_3245, w_082_3246, w_082_3247, w_082_3252, w_082_3253, w_082_3256, w_082_3258, w_082_3260, w_082_3261, w_082_3262, w_082_3264, w_082_3267, w_082_3272, w_082_3276, w_082_3277, w_082_3280, w_082_3281, w_082_3282, w_082_3283, w_082_3289, w_082_3290, w_082_3294, w_082_3295, w_082_3297, w_082_3298, w_082_3301, w_082_3302, w_082_3303, w_082_3305, w_082_3306, w_082_3307, w_082_3311, w_082_3314, w_082_3315, w_082_3316, w_082_3318, w_082_3319, w_082_3320, w_082_3321, w_082_3323, w_082_3324, w_082_3325, w_082_3326, w_082_3331, w_082_3332, w_082_3333, w_082_3336, w_082_3337, w_082_3340, w_082_3342, w_082_3346, w_082_3352, w_082_3354, w_082_3359, w_082_3361, w_082_3363, w_082_3366, w_082_3367, w_082_3372, w_082_3374, w_082_3378, w_082_3379, w_082_3380, w_082_3383, w_082_3386, w_082_3387, w_082_3394, w_082_3395, w_082_3396, w_082_3398, w_082_3400, w_082_3405, w_082_3406, w_082_3407, w_082_3409, w_082_3410, w_082_3411, w_082_3416, w_082_3418, w_082_3421, w_082_3423, w_082_3424, w_082_3425, w_082_3428, w_082_3430, w_082_3431, w_082_3432, w_082_3435, w_082_3436, w_082_3439, w_082_3440, w_082_3443, w_082_3444, w_082_3451, w_082_3452, w_082_3455, w_082_3457, w_082_3459, w_082_3460, w_082_3462, w_082_3464, w_082_3466, w_082_3467, w_082_3469, w_082_3470, w_082_3471, w_082_3475, w_082_3476, w_082_3477, w_082_3479, w_082_3481, w_082_3482, w_082_3483, w_082_3491, w_082_3492, w_082_3494, w_082_3498, w_082_3499, w_082_3501, w_082_3503, w_082_3506, w_082_3516, w_082_3519, w_082_3523, w_082_3524, w_082_3531, w_082_3535, w_082_3537, w_082_3540, w_082_3541, w_082_3542, w_082_3545, w_082_3546, w_082_3548, w_082_3549, w_082_3550, w_082_3553, w_082_3554, w_082_3558, w_082_3561, w_082_3564, w_082_3566, w_082_3568, w_082_3569, w_082_3570, w_082_3571, w_082_3572, w_082_3573, w_082_3578, w_082_3580, w_082_3584, w_082_3585, w_082_3586, w_082_3587, w_082_3589, w_082_3590, w_082_3591, w_082_3594, w_082_3596, w_082_3597, w_082_3598, w_082_3599, w_082_3600, w_082_3602, w_082_3606, w_082_3607, w_082_3610, w_082_3612, w_082_3613, w_082_3614, w_082_3615, w_082_3625, w_082_3626, w_082_3628, w_082_3629, w_082_3631, w_082_3633, w_082_3634, w_082_3638, w_082_3640, w_082_3641, w_082_3642, w_082_3643, w_082_3647, w_082_3654, w_082_3656, w_082_3658, w_082_3659, w_082_3662, w_082_3663, w_082_3666, w_082_3669, w_082_3672, w_082_3673, w_082_3679, w_082_3680, w_082_3682, w_082_3688, w_082_3690, w_082_3691, w_082_3694, w_082_3696, w_082_3702, w_082_3708, w_082_3714, w_082_3716, w_082_3717, w_082_3721, w_082_3722, w_082_3723, w_082_3725, w_082_3726, w_082_3727, w_082_3729, w_082_3730, w_082_3731, w_082_3732, w_082_3734, w_082_3736, w_082_3739, w_082_3743, w_082_3746, w_082_3747, w_082_3748, w_082_3749, w_082_3754, w_082_3756, w_082_3758, w_082_3759, w_082_3760, w_082_3762, w_082_3763, w_082_3769, w_082_3771, w_082_3772, w_082_3773, w_082_3774, w_082_3776, w_082_3780, w_082_3786, w_082_3787, w_082_3788, w_082_3789, w_082_3791, w_082_3794, w_082_3798, w_082_3799, w_082_3800, w_082_3801, w_082_3805, w_082_3807, w_082_3810, w_082_3811, w_082_3814, w_082_3815, w_082_3819, w_082_3820, w_082_3821, w_082_3824, w_082_3825, w_082_3826, w_082_3827, w_082_3829, w_082_3830, w_082_3832, w_082_3833, w_082_3834, w_082_3839, w_082_3844, w_082_3845, w_082_3848, w_082_3852, w_082_3854, w_082_3856, w_082_3857, w_082_3858, w_082_3860, w_082_3861, w_082_3863, w_082_3864, w_082_3869, w_082_3871, w_082_3872, w_082_3873, w_082_3874, w_082_3877, w_082_3884, w_082_3887, w_082_3888, w_082_3895, w_082_3898, w_082_3907, w_082_3908, w_082_3909, w_082_3910, w_082_3911, w_082_3915, w_082_3917, w_082_3920, w_082_3922, w_082_3924, w_082_3925, w_082_3928, w_082_3929, w_082_3930, w_082_3932, w_082_3939, w_082_3940, w_082_3942, w_082_3945, w_082_3946, w_082_3948, w_082_3952, w_082_3953, w_082_3956, w_082_3960, w_082_3961, w_082_3968, w_082_3972, w_082_3976, w_082_3977, w_082_3979, w_082_3981, w_082_3984, w_082_3987, w_082_3993, w_082_3997, w_082_3999, w_082_4000, w_082_4001, w_082_4002, w_082_4007, w_082_4008, w_082_4010, w_082_4011, w_082_4013, w_082_4014, w_082_4015, w_082_4017, w_082_4020, w_082_4022, w_082_4027, w_082_4029, w_082_4030, w_082_4031, w_082_4032, w_082_4035, w_082_4036, w_082_4037, w_082_4038, w_082_4040, w_082_4041, w_082_4043, w_082_4047, w_082_4049, w_082_4050, w_082_4054, w_082_4057, w_082_4058, w_082_4059, w_082_4060, w_082_4064, w_082_4065, w_082_4066, w_082_4071, w_082_4073, w_082_4077, w_082_4081, w_082_4084, w_082_4085, w_082_4086, w_082_4087, w_082_4092, w_082_4093, w_082_4096, w_082_4098, w_082_4099, w_082_4102, w_082_4104, w_082_4105, w_082_4109, w_082_4110, w_082_4116, w_082_4118, w_082_4119, w_082_4121, w_082_4126, w_082_4127, w_082_4128, w_082_4130, w_082_4132, w_082_4134, w_082_4135, w_082_4139, w_082_4143, w_082_4144, w_082_4146, w_082_4147, w_082_4152, w_082_4153, w_082_4163, w_082_4165, w_082_4171, w_082_4172, w_082_4176, w_082_4177, w_082_4183, w_082_4184, w_082_4185, w_082_4186, w_082_4188, w_082_4189, w_082_4190, w_082_4192, w_082_4193, w_082_4195, w_082_4197, w_082_4198, w_082_4199, w_082_4201, w_082_4202, w_082_4205, w_082_4207, w_082_4208, w_082_4211, w_082_4215, w_082_4216, w_082_4218, w_082_4220, w_082_4221, w_082_4222, w_082_4223, w_082_4224, w_082_4226, w_082_4228, w_082_4232, w_082_4234, w_082_4239, w_082_4241, w_082_4242, w_082_4243, w_082_4248, w_082_4250, w_082_4254, w_082_4256, w_082_4257, w_082_4259, w_082_4260, w_082_4264, w_082_4265, w_082_4266, w_082_4268, w_082_4269, w_082_4270, w_082_4271, w_082_4272, w_082_4273, w_082_4274, w_082_4277, w_082_4278, w_082_4279, w_082_4282, w_082_4285, w_082_4287, w_082_4288, w_082_4289, w_082_4291, w_082_4292, w_082_4293, w_082_4295, w_082_4296, w_082_4298, w_082_4299, w_082_4300, w_082_4303, w_082_4304, w_082_4309, w_082_4310, w_082_4313, w_082_4314, w_082_4315, w_082_4316, w_082_4319, w_082_4321, w_082_4322, w_082_4324, w_082_4327, w_082_4329, w_082_4332, w_082_4340, w_082_4341, w_082_4342, w_082_4344, w_082_4346, w_082_4348, w_082_4349, w_082_4350, w_082_4351, w_082_4353, w_082_4354, w_082_4355, w_082_4357, w_082_4360, w_082_4362, w_082_4363, w_082_4366, w_082_4370, w_082_4372, w_082_4373, w_082_4376, w_082_4378, w_082_4380, w_082_4381, w_082_4382, w_082_4384, w_082_4390, w_082_4391, w_082_4393, w_082_4394, w_082_4396, w_082_4399, w_082_4400, w_082_4401, w_082_4402, w_082_4403, w_082_4405, w_082_4407, w_082_4414, w_082_4416, w_082_4419, w_082_4421, w_082_4422, w_082_4423, w_082_4424, w_082_4427, w_082_4430, w_082_4431, w_082_4435, w_082_4438;
  wire w_083_002, w_083_003, w_083_004, w_083_005, w_083_007, w_083_009, w_083_011, w_083_016, w_083_017, w_083_021, w_083_022, w_083_023, w_083_025, w_083_026, w_083_028, w_083_029, w_083_030, w_083_031, w_083_033, w_083_037, w_083_046, w_083_048, w_083_051, w_083_054, w_083_057, w_083_058, w_083_067, w_083_068, w_083_070, w_083_071, w_083_074, w_083_077, w_083_078, w_083_079, w_083_081, w_083_083, w_083_086, w_083_089, w_083_090, w_083_091, w_083_092, w_083_093, w_083_094, w_083_095, w_083_097, w_083_100, w_083_101, w_083_102, w_083_106, w_083_107, w_083_109, w_083_111, w_083_113, w_083_115, w_083_126, w_083_129, w_083_132, w_083_135, w_083_137, w_083_139, w_083_140, w_083_142, w_083_143, w_083_144, w_083_146, w_083_150, w_083_153, w_083_156, w_083_157, w_083_159, w_083_160, w_083_163, w_083_165, w_083_166, w_083_169, w_083_171, w_083_172, w_083_173, w_083_174, w_083_177, w_083_178, w_083_182, w_083_183, w_083_185, w_083_186, w_083_189, w_083_190, w_083_191, w_083_192, w_083_196, w_083_197, w_083_200, w_083_203, w_083_204, w_083_205, w_083_206, w_083_207, w_083_209, w_083_210, w_083_211, w_083_214, w_083_216, w_083_218, w_083_221, w_083_222, w_083_226, w_083_228, w_083_230, w_083_235, w_083_241, w_083_243, w_083_245, w_083_247, w_083_249, w_083_250, w_083_256, w_083_263, w_083_265, w_083_266, w_083_268, w_083_270, w_083_271, w_083_273, w_083_274, w_083_278, w_083_280, w_083_281, w_083_282, w_083_285, w_083_286, w_083_287, w_083_289, w_083_290, w_083_291, w_083_294, w_083_296, w_083_299, w_083_300, w_083_301, w_083_302, w_083_304, w_083_307, w_083_308, w_083_315, w_083_317, w_083_320, w_083_321, w_083_326, w_083_327, w_083_328, w_083_329, w_083_334, w_083_335, w_083_337, w_083_340, w_083_341, w_083_343, w_083_344, w_083_347, w_083_348, w_083_350, w_083_355, w_083_359, w_083_361, w_083_362, w_083_364, w_083_366, w_083_367, w_083_368, w_083_369, w_083_373, w_083_376, w_083_378, w_083_379, w_083_381, w_083_382, w_083_383, w_083_384, w_083_387, w_083_392, w_083_400, w_083_402, w_083_403, w_083_404, w_083_405, w_083_407, w_083_408, w_083_409, w_083_410, w_083_411, w_083_412, w_083_415, w_083_417, w_083_418, w_083_419, w_083_420, w_083_423, w_083_424, w_083_429, w_083_431, w_083_434, w_083_435, w_083_437, w_083_439, w_083_440, w_083_443, w_083_444, w_083_446, w_083_447, w_083_449, w_083_450, w_083_451, w_083_453, w_083_455, w_083_456, w_083_457, w_083_459, w_083_460, w_083_463, w_083_464, w_083_465, w_083_469, w_083_470, w_083_471, w_083_472, w_083_478, w_083_482, w_083_484, w_083_486, w_083_488, w_083_489, w_083_492, w_083_493, w_083_494, w_083_495, w_083_500, w_083_503, w_083_505, w_083_506, w_083_509, w_083_511, w_083_514, w_083_515, w_083_518, w_083_519, w_083_520, w_083_521, w_083_522, w_083_523, w_083_525, w_083_527, w_083_528, w_083_529, w_083_531, w_083_534, w_083_535, w_083_537, w_083_538, w_083_542, w_083_543, w_083_544, w_083_546, w_083_549, w_083_557, w_083_558, w_083_560, w_083_561, w_083_562, w_083_565, w_083_573, w_083_575, w_083_576, w_083_579, w_083_581, w_083_583, w_083_584, w_083_585, w_083_587, w_083_590, w_083_591, w_083_593, w_083_598, w_083_599, w_083_601, w_083_602, w_083_610, w_083_619, w_083_621, w_083_622, w_083_625, w_083_626, w_083_628, w_083_630, w_083_633, w_083_636, w_083_639, w_083_642, w_083_643, w_083_645, w_083_646, w_083_652, w_083_655, w_083_658, w_083_659, w_083_664, w_083_666, w_083_670, w_083_673, w_083_676, w_083_677, w_083_679, w_083_680, w_083_681, w_083_683, w_083_684, w_083_685, w_083_687, w_083_691, w_083_692, w_083_693, w_083_694, w_083_696, w_083_697, w_083_701, w_083_702, w_083_703, w_083_705, w_083_706, w_083_708, w_083_710, w_083_714, w_083_718, w_083_722, w_083_724, w_083_726, w_083_727, w_083_731, w_083_732, w_083_733, w_083_735, w_083_736, w_083_737, w_083_738, w_083_739, w_083_740, w_083_742, w_083_743, w_083_749, w_083_750, w_083_751, w_083_752, w_083_753, w_083_754, w_083_755, w_083_759, w_083_760, w_083_763, w_083_766, w_083_770, w_083_771, w_083_772, w_083_774, w_083_775, w_083_782, w_083_783, w_083_787, w_083_788, w_083_790, w_083_792, w_083_795, w_083_796, w_083_798, w_083_801, w_083_804, w_083_805, w_083_806, w_083_807, w_083_808, w_083_809, w_083_810, w_083_816, w_083_817, w_083_820, w_083_821, w_083_822, w_083_823, w_083_824, w_083_825, w_083_828, w_083_835, w_083_838, w_083_839, w_083_840, w_083_841, w_083_847, w_083_848, w_083_849, w_083_850, w_083_851, w_083_852, w_083_853, w_083_854, w_083_858, w_083_860, w_083_864, w_083_865, w_083_867, w_083_868, w_083_869, w_083_870, w_083_875, w_083_876, w_083_877, w_083_879, w_083_885, w_083_886, w_083_887, w_083_888, w_083_889, w_083_890, w_083_891, w_083_892, w_083_893, w_083_895, w_083_896, w_083_898, w_083_901, w_083_909, w_083_910, w_083_912, w_083_913, w_083_915, w_083_916, w_083_917, w_083_918, w_083_922, w_083_923, w_083_924, w_083_925, w_083_927, w_083_928, w_083_930, w_083_933, w_083_934, w_083_936, w_083_937, w_083_938, w_083_942, w_083_943, w_083_947, w_083_949, w_083_951, w_083_952, w_083_955, w_083_958, w_083_960, w_083_961, w_083_962, w_083_966, w_083_967, w_083_969, w_083_971, w_083_973, w_083_974, w_083_976, w_083_977, w_083_980, w_083_981, w_083_982, w_083_987, w_083_988, w_083_989, w_083_990, w_083_995, w_083_997, w_083_998, w_083_999, w_083_1000, w_083_1004, w_083_1007, w_083_1008, w_083_1013, w_083_1014, w_083_1015, w_083_1018, w_083_1020, w_083_1021, w_083_1025, w_083_1026, w_083_1029, w_083_1030, w_083_1031, w_083_1032, w_083_1033, w_083_1036, w_083_1038, w_083_1041, w_083_1044, w_083_1045, w_083_1047, w_083_1049, w_083_1051, w_083_1053, w_083_1054, w_083_1056, w_083_1058, w_083_1061, w_083_1063, w_083_1064, w_083_1065, w_083_1066, w_083_1067, w_083_1068, w_083_1071, w_083_1074, w_083_1076, w_083_1077, w_083_1080, w_083_1081, w_083_1083, w_083_1084, w_083_1085, w_083_1087, w_083_1088, w_083_1090, w_083_1091, w_083_1092, w_083_1095, w_083_1096, w_083_1100, w_083_1101, w_083_1102, w_083_1108, w_083_1110, w_083_1113, w_083_1117, w_083_1118, w_083_1119, w_083_1120, w_083_1122, w_083_1123, w_083_1127, w_083_1128, w_083_1129, w_083_1133, w_083_1137, w_083_1141, w_083_1148, w_083_1153, w_083_1156, w_083_1158, w_083_1162, w_083_1163, w_083_1164, w_083_1165, w_083_1166, w_083_1167, w_083_1170, w_083_1171, w_083_1175, w_083_1178, w_083_1181, w_083_1184, w_083_1185, w_083_1190, w_083_1191, w_083_1192, w_083_1193, w_083_1195, w_083_1196, w_083_1198, w_083_1199, w_083_1200, w_083_1203, w_083_1205, w_083_1206, w_083_1207, w_083_1211, w_083_1212, w_083_1216, w_083_1219, w_083_1220, w_083_1224, w_083_1226, w_083_1228, w_083_1233, w_083_1235, w_083_1237, w_083_1238, w_083_1239, w_083_1240, w_083_1241, w_083_1243, w_083_1244, w_083_1246, w_083_1247, w_083_1249, w_083_1251, w_083_1252, w_083_1261, w_083_1262, w_083_1265, w_083_1268, w_083_1271, w_083_1272, w_083_1276, w_083_1278, w_083_1283, w_083_1284, w_083_1288, w_083_1289, w_083_1291, w_083_1293, w_083_1295, w_083_1297, w_083_1301, w_083_1302, w_083_1305, w_083_1307, w_083_1309, w_083_1310, w_083_1311, w_083_1312, w_083_1314, w_083_1316, w_083_1318, w_083_1321, w_083_1323, w_083_1328, w_083_1329, w_083_1331, w_083_1332, w_083_1333, w_083_1335, w_083_1336, w_083_1337, w_083_1338, w_083_1339, w_083_1350, w_083_1351, w_083_1352, w_083_1353, w_083_1357, w_083_1358, w_083_1361, w_083_1363, w_083_1376, w_083_1379, w_083_1381, w_083_1384, w_083_1387, w_083_1388, w_083_1390, w_083_1393, w_083_1394, w_083_1396, w_083_1399, w_083_1400, w_083_1402, w_083_1403, w_083_1406, w_083_1408, w_083_1414, w_083_1417, w_083_1419, w_083_1421, w_083_1423, w_083_1425, w_083_1427, w_083_1431, w_083_1433, w_083_1434, w_083_1435, w_083_1436, w_083_1438, w_083_1448, w_083_1450, w_083_1454, w_083_1455, w_083_1457, w_083_1462, w_083_1465, w_083_1466, w_083_1469, w_083_1471, w_083_1472, w_083_1473, w_083_1483, w_083_1485, w_083_1493, w_083_1496, w_083_1498, w_083_1499, w_083_1500, w_083_1501, w_083_1502, w_083_1504, w_083_1505, w_083_1507, w_083_1510, w_083_1516, w_083_1517, w_083_1519, w_083_1522, w_083_1527, w_083_1529, w_083_1530, w_083_1531, w_083_1535, w_083_1538, w_083_1541, w_083_1548, w_083_1549, w_083_1550, w_083_1551, w_083_1554, w_083_1558, w_083_1559, w_083_1562, w_083_1569, w_083_1572, w_083_1573, w_083_1578, w_083_1581, w_083_1582, w_083_1584, w_083_1585, w_083_1586, w_083_1588, w_083_1591, w_083_1594, w_083_1596, w_083_1599, w_083_1600, w_083_1604, w_083_1605, w_083_1606, w_083_1607, w_083_1609, w_083_1611, w_083_1615, w_083_1618, w_083_1623, w_083_1625, w_083_1626, w_083_1627, w_083_1628, w_083_1629, w_083_1633, w_083_1638, w_083_1639, w_083_1641, w_083_1642, w_083_1643, w_083_1644, w_083_1646, w_083_1647, w_083_1649, w_083_1653, w_083_1655, w_083_1659, w_083_1660, w_083_1661, w_083_1665, w_083_1666, w_083_1667, w_083_1668, w_083_1669, w_083_1670, w_083_1675, w_083_1677, w_083_1678, w_083_1684, w_083_1686, w_083_1687, w_083_1688, w_083_1689, w_083_1694, w_083_1696, w_083_1700, w_083_1701, w_083_1705, w_083_1707, w_083_1708, w_083_1710, w_083_1711, w_083_1712, w_083_1717, w_083_1721, w_083_1724, w_083_1725, w_083_1726, w_083_1730, w_083_1731, w_083_1732, w_083_1735, w_083_1738, w_083_1740, w_083_1741, w_083_1742, w_083_1743, w_083_1744, w_083_1747, w_083_1749, w_083_1751, w_083_1753, w_083_1757, w_083_1758, w_083_1759, w_083_1762, w_083_1764, w_083_1766, w_083_1768, w_083_1769, w_083_1771, w_083_1772, w_083_1774, w_083_1776, w_083_1777, w_083_1779, w_083_1781, w_083_1782, w_083_1783, w_083_1784, w_083_1786, w_083_1787, w_083_1789, w_083_1792, w_083_1796, w_083_1798, w_083_1801, w_083_1804, w_083_1805, w_083_1806, w_083_1807, w_083_1808, w_083_1811, w_083_1812, w_083_1813, w_083_1814, w_083_1815, w_083_1816, w_083_1821, w_083_1823, w_083_1825, w_083_1827, w_083_1828, w_083_1830, w_083_1832, w_083_1833, w_083_1835, w_083_1836, w_083_1839, w_083_1841, w_083_1842, w_083_1843, w_083_1844, w_083_1850, w_083_1851, w_083_1854, w_083_1856, w_083_1858, w_083_1861, w_083_1862, w_083_1863, w_083_1865, w_083_1868, w_083_1869, w_083_1871, w_083_1872, w_083_1873, w_083_1881, w_083_1882, w_083_1886, w_083_1888, w_083_1893, w_083_1894, w_083_1895, w_083_1896, w_083_1897, w_083_1898, w_083_1900, w_083_1901, w_083_1905, w_083_1906, w_083_1908, w_083_1911, w_083_1913, w_083_1919, w_083_1921, w_083_1924, w_083_1925, w_083_1926, w_083_1929, w_083_1930, w_083_1934, w_083_1937, w_083_1939, w_083_1941, w_083_1942, w_083_1944, w_083_1945, w_083_1946, w_083_1950, w_083_1951, w_083_1957, w_083_1960, w_083_1963, w_083_1964, w_083_1965, w_083_1966, w_083_1968, w_083_1970, w_083_1972, w_083_1973, w_083_1974, w_083_1977, w_083_1978, w_083_1979, w_083_1980, w_083_1981, w_083_1985, w_083_1987, w_083_1991, w_083_1992, w_083_1994, w_083_1995, w_083_1997, w_083_1999, w_083_2000, w_083_2005, w_083_2006, w_083_2011, w_083_2014, w_083_2018, w_083_2020, w_083_2021, w_083_2024, w_083_2029, w_083_2031, w_083_2032, w_083_2033, w_083_2034, w_083_2036, w_083_2037, w_083_2038, w_083_2040, w_083_2041, w_083_2044, w_083_2045, w_083_2046, w_083_2049, w_083_2052, w_083_2055, w_083_2058, w_083_2060, w_083_2061, w_083_2062, w_083_2064, w_083_2067, w_083_2068, w_083_2069, w_083_2070, w_083_2072, w_083_2074, w_083_2077, w_083_2080, w_083_2083, w_083_2087, w_083_2088, w_083_2090, w_083_2091, w_083_2096, w_083_2098, w_083_2101, w_083_2102, w_083_2105, w_083_2112, w_083_2114, w_083_2115, w_083_2116, w_083_2118, w_083_2121, w_083_2123, w_083_2125, w_083_2126, w_083_2128, w_083_2133, w_083_2135, w_083_2137, w_083_2138, w_083_2141, w_083_2142, w_083_2146, w_083_2147, w_083_2148, w_083_2149, w_083_2151, w_083_2153, w_083_2154, w_083_2157, w_083_2158, w_083_2161, w_083_2162, w_083_2164, w_083_2167, w_083_2169, w_083_2170, w_083_2172, w_083_2174, w_083_2177, w_083_2179, w_083_2181, w_083_2182, w_083_2183, w_083_2187, w_083_2189, w_083_2190, w_083_2191, w_083_2192, w_083_2195, w_083_2196, w_083_2201, w_083_2205, w_083_2206, w_083_2208, w_083_2209, w_083_2211, w_083_2212, w_083_2213, w_083_2214, w_083_2220, w_083_2222, w_083_2226, w_083_2227, w_083_2228, w_083_2236, w_083_2239, w_083_2242, w_083_2243, w_083_2251, w_083_2253, w_083_2258, w_083_2259, w_083_2260, w_083_2261, w_083_2262, w_083_2266, w_083_2268, w_083_2271, w_083_2274, w_083_2277, w_083_2278, w_083_2282, w_083_2284, w_083_2285, w_083_2287, w_083_2288, w_083_2291, w_083_2295, w_083_2297, w_083_2298, w_083_2299, w_083_2302, w_083_2303, w_083_2308, w_083_2311, w_083_2312, w_083_2315, w_083_2316, w_083_2318, w_083_2321, w_083_2322, w_083_2324, w_083_2327, w_083_2328, w_083_2332, w_083_2334, w_083_2339, w_083_2341, w_083_2345, w_083_2346, w_083_2347, w_083_2349, w_083_2350, w_083_2351, w_083_2354, w_083_2355, w_083_2358, w_083_2360, w_083_2363, w_083_2365, w_083_2374, w_083_2375, w_083_2376, w_083_2382, w_083_2389, w_083_2390, w_083_2395, w_083_2398, w_083_2407, w_083_2408, w_083_2415, w_083_2422, w_083_2424, w_083_2428, w_083_2429, w_083_2433, w_083_2434, w_083_2435, w_083_2438, w_083_2441, w_083_2449, w_083_2450, w_083_2452, w_083_2458, w_083_2459, w_083_2460, w_083_2464, w_083_2467, w_083_2471, w_083_2472, w_083_2477, w_083_2489, w_083_2491, w_083_2492, w_083_2504, w_083_2507, w_083_2524, w_083_2529, w_083_2532, w_083_2535, w_083_2538, w_083_2548, w_083_2563, w_083_2567, w_083_2568, w_083_2571, w_083_2580, w_083_2583, w_083_2591, w_083_2592, w_083_2596, w_083_2597, w_083_2600, w_083_2609, w_083_2611, w_083_2620, w_083_2622, w_083_2626, w_083_2627, w_083_2629, w_083_2630, w_083_2634, w_083_2636, w_083_2641, w_083_2644, w_083_2645, w_083_2650, w_083_2652, w_083_2653, w_083_2654, w_083_2655, w_083_2656, w_083_2663, w_083_2664, w_083_2684, w_083_2685, w_083_2687, w_083_2690, w_083_2691, w_083_2692, w_083_2693, w_083_2705, w_083_2710, w_083_2711, w_083_2713, w_083_2714, w_083_2723, w_083_2730, w_083_2737, w_083_2740, w_083_2745, w_083_2750, w_083_2752, w_083_2753, w_083_2756, w_083_2763, w_083_2776, w_083_2780, w_083_2781, w_083_2783, w_083_2784, w_083_2785, w_083_2788, w_083_2791, w_083_2796, w_083_2797, w_083_2798, w_083_2799, w_083_2801, w_083_2803, w_083_2807, w_083_2823, w_083_2829, w_083_2830, w_083_2838, w_083_2840, w_083_2843, w_083_2844, w_083_2847, w_083_2859, w_083_2860, w_083_2864, w_083_2867, w_083_2869, w_083_2880, w_083_2881, w_083_2882, w_083_2885, w_083_2889, w_083_2901, w_083_2904, w_083_2905, w_083_2906, w_083_2909, w_083_2912, w_083_2913, w_083_2915, w_083_2916, w_083_2921, w_083_2927, w_083_2929, w_083_2937, w_083_2943, w_083_2944, w_083_2946, w_083_2948, w_083_2950, w_083_2953, w_083_2958, w_083_2964, w_083_2967, w_083_2972, w_083_2978, w_083_2979, w_083_2985, w_083_2988, w_083_2996, w_083_3001, w_083_3004, w_083_3005, w_083_3007, w_083_3010, w_083_3014, w_083_3024, w_083_3027, w_083_3034, w_083_3038, w_083_3041, w_083_3042, w_083_3043, w_083_3051, w_083_3054, w_083_3057, w_083_3061, w_083_3068, w_083_3071, w_083_3072, w_083_3074, w_083_3079, w_083_3080, w_083_3081, w_083_3089, w_083_3091, w_083_3096, w_083_3103, w_083_3105, w_083_3115, w_083_3117, w_083_3120, w_083_3122, w_083_3123, w_083_3129, w_083_3131, w_083_3136, w_083_3143, w_083_3147, w_083_3148, w_083_3149, w_083_3156, w_083_3160, w_083_3162, w_083_3174, w_083_3176, w_083_3177, w_083_3182, w_083_3197, w_083_3203, w_083_3204, w_083_3215, w_083_3222, w_083_3225, w_083_3231, w_083_3241, w_083_3243, w_083_3244, w_083_3248, w_083_3252, w_083_3260, w_083_3262, w_083_3266, w_083_3272, w_083_3275, w_083_3278, w_083_3279, w_083_3280, w_083_3281, w_083_3284, w_083_3288, w_083_3299, w_083_3301, w_083_3303, w_083_3307, w_083_3310, w_083_3311, w_083_3312, w_083_3319, w_083_3321, w_083_3329, w_083_3341, w_083_3355, w_083_3358, w_083_3365, w_083_3374, w_083_3376, w_083_3380, w_083_3381, w_083_3382, w_083_3386, w_083_3388, w_083_3397, w_083_3398, w_083_3405, w_083_3411, w_083_3419, w_083_3425, w_083_3426, w_083_3429, w_083_3433, w_083_3441, w_083_3448, w_083_3453, w_083_3455, w_083_3456, w_083_3461, w_083_3462, w_083_3474, w_083_3485, w_083_3490, w_083_3491, w_083_3506, w_083_3510, w_083_3515, w_083_3517, w_083_3519, w_083_3522, w_083_3524, w_083_3526, w_083_3531, w_083_3540, w_083_3543, w_083_3545, w_083_3552, w_083_3553, w_083_3555, w_083_3563, w_083_3565, w_083_3568, w_083_3569, w_083_3572, w_083_3573, w_083_3574, w_083_3576, w_083_3583, w_083_3584, w_083_3586, w_083_3589, w_083_3599, w_083_3603, w_083_3607, w_083_3609, w_083_3611, w_083_3612, w_083_3614, w_083_3621, w_083_3625, w_083_3633, w_083_3635, w_083_3639, w_083_3641, w_083_3644, w_083_3648, w_083_3649, w_083_3655, w_083_3656, w_083_3657, w_083_3662, w_083_3671, w_083_3679, w_083_3680, w_083_3681, w_083_3683, w_083_3684, w_083_3689, w_083_3693, w_083_3700, w_083_3702, w_083_3704, w_083_3705, w_083_3707, w_083_3709, w_083_3711, w_083_3712, w_083_3716, w_083_3720, w_083_3727, w_083_3730, w_083_3733, w_083_3743, w_083_3745, w_083_3746, w_083_3753, w_083_3755, w_083_3758, w_083_3760, w_083_3764, w_083_3765, w_083_3775, w_083_3776, w_083_3787, w_083_3791, w_083_3794, w_083_3798, w_083_3803, w_083_3806, w_083_3807, w_083_3809, w_083_3810, w_083_3817, w_083_3822, w_083_3830, w_083_3831, w_083_3833, w_083_3839, w_083_3841, w_083_3847, w_083_3853, w_083_3854, w_083_3859, w_083_3865, w_083_3868, w_083_3870, w_083_3877, w_083_3882, w_083_3889, w_083_3894, w_083_3895, w_083_3902, w_083_3904, w_083_3912, w_083_3914, w_083_3915, w_083_3918, w_083_3919, w_083_3920, w_083_3922, w_083_3930, w_083_3933, w_083_3936, w_083_3944, w_083_3949, w_083_3956, w_083_3963, w_083_3964, w_083_3966, w_083_3968, w_083_3972, w_083_3978, w_083_3984, w_083_3986, w_083_3987, w_083_3990, w_083_3992, w_083_3995, w_083_3997, w_083_4000, w_083_4002, w_083_4006, w_083_4015, w_083_4018, w_083_4022, w_083_4024, w_083_4029, w_083_4031, w_083_4032, w_083_4036, w_083_4039, w_083_4045, w_083_4047, w_083_4048, w_083_4050, w_083_4054, w_083_4056, w_083_4067, w_083_4072, w_083_4073, w_083_4078, w_083_4080, w_083_4082, w_083_4087, w_083_4092, w_083_4099, w_083_4103, w_083_4112, w_083_4115, w_083_4119, w_083_4132, w_083_4134, w_083_4135, w_083_4137, w_083_4139, w_083_4145, w_083_4154, w_083_4157, w_083_4158, w_083_4159, w_083_4171, w_083_4174, w_083_4179, w_083_4182, w_083_4187, w_083_4188, w_083_4189, w_083_4197, w_083_4201, w_083_4211, w_083_4216, w_083_4217, w_083_4222, w_083_4223, w_083_4224, w_083_4228, w_083_4229, w_083_4234, w_083_4241, w_083_4245, w_083_4247, w_083_4252, w_083_4255, w_083_4279, w_083_4282, w_083_4284, w_083_4286, w_083_4287, w_083_4288, w_083_4295, w_083_4296, w_083_4297, w_083_4302, w_083_4306, w_083_4307, w_083_4308, w_083_4309, w_083_4311, w_083_4318, w_083_4319, w_083_4321, w_083_4325, w_083_4328, w_083_4331, w_083_4337, w_083_4340, w_083_4343, w_083_4355, w_083_4362, w_083_4366, w_083_4368, w_083_4374, w_083_4376, w_083_4378, w_083_4381, w_083_4392, w_083_4395, w_083_4409, w_083_4414, w_083_4415, w_083_4419, w_083_4420, w_083_4431, w_083_4432, w_083_4439, w_083_4443, w_083_4447, w_083_4449, w_083_4457, w_083_4458, w_083_4460, w_083_4464, w_083_4465, w_083_4466, w_083_4468, w_083_4472, w_083_4475, w_083_4482, w_083_4484, w_083_4485, w_083_4494, w_083_4496, w_083_4497, w_083_4500, w_083_4501, w_083_4504, w_083_4505, w_083_4506, w_083_4507, w_083_4511, w_083_4516, w_083_4524, w_083_4528, w_083_4533, w_083_4536, w_083_4539, w_083_4542, w_083_4546, w_083_4551, w_083_4554, w_083_4555, w_083_4556, w_083_4563, w_083_4567, w_083_4569, w_083_4570, w_083_4575, w_083_4577, w_083_4581, w_083_4584, w_083_4586, w_083_4587, w_083_4591, w_083_4592, w_083_4597, w_083_4601, w_083_4602, w_083_4603, w_083_4609, w_083_4611, w_083_4613, w_083_4616, w_083_4617, w_083_4619, w_083_4624, w_083_4626, w_083_4629, w_083_4630, w_083_4631, w_083_4633, w_083_4637, w_083_4639, w_083_4640, w_083_4645, w_083_4646, w_083_4648, w_083_4657, w_083_4658, w_083_4662, w_083_4663, w_083_4667, w_083_4674, w_083_4682, w_083_4694, w_083_4700, w_083_4702, w_083_4707, w_083_4708, w_083_4716, w_083_4718, w_083_4720, w_083_4721, w_083_4729, w_083_4731, w_083_4734, w_083_4738, w_083_4739, w_083_4741, w_083_4744, w_083_4746, w_083_4762, w_083_4763, w_083_4765, w_083_4766, w_083_4768, w_083_4770, w_083_4773, w_083_4774, w_083_4775, w_083_4781, w_083_4786, w_083_4793, w_083_4798, w_083_4806, w_083_4810, w_083_4811, w_083_4813, w_083_4819, w_083_4822, w_083_4824, w_083_4831, w_083_4833, w_083_4836, w_083_4838, w_083_4839, w_083_4847, w_083_4848, w_083_4853, w_083_4858, w_083_4863, w_083_4865, w_083_4868, w_083_4870, w_083_4873, w_083_4883, w_083_4884, w_083_4887, w_083_4889, w_083_4890, w_083_4898, w_083_4900, w_083_4904, w_083_4908, w_083_4909, w_083_4916, w_083_4922, w_083_4928, w_083_4935, w_083_4937, w_083_4938, w_083_4941, w_083_4942, w_083_4953, w_083_4955, w_083_4961, w_083_4962, w_083_4965, w_083_4969, w_083_4972, w_083_4979, w_083_4981, w_083_4985, w_083_4989, w_083_4991, w_083_5003, w_083_5008, w_083_5025, w_083_5028, w_083_5032, w_083_5036, w_083_5038, w_083_5045, w_083_5067, w_083_5068, w_083_5072, w_083_5083, w_083_5085, w_083_5088, w_083_5093, w_083_5098, w_083_5099, w_083_5102, w_083_5104, w_083_5106, w_083_5114, w_083_5121, w_083_5130, w_083_5132, w_083_5136, w_083_5142, w_083_5144, w_083_5145, w_083_5147, w_083_5156, w_083_5157, w_083_5165, w_083_5166, w_083_5167, w_083_5170, w_083_5171, w_083_5175, w_083_5177, w_083_5178, w_083_5181, w_083_5182, w_083_5183, w_083_5190, w_083_5193, w_083_5194, w_083_5198, w_083_5200, w_083_5206, w_083_5209, w_083_5211, w_083_5212, w_083_5213, w_083_5217, w_083_5219, w_083_5220, w_083_5222, w_083_5226, w_083_5229, w_083_5233, w_083_5234, w_083_5236, w_083_5241, w_083_5246, w_083_5254, w_083_5255, w_083_5261, w_083_5264, w_083_5270, w_083_5271, w_083_5272, w_083_5278, w_083_5290, w_083_5298, w_083_5302, w_083_5308, w_083_5317, w_083_5321, w_083_5322, w_083_5324, w_083_5326, w_083_5335, w_083_5336, w_083_5339, w_083_5340, w_083_5342, w_083_5345, w_083_5346, w_083_5348, w_083_5351, w_083_5353, w_083_5355, w_083_5356, w_083_5358, w_083_5363, w_083_5366, w_083_5380, w_083_5384, w_083_5392, w_083_5394, w_083_5395, w_083_5397, w_083_5404, w_083_5408, w_083_5409, w_083_5410, w_083_5412, w_083_5413, w_083_5416, w_083_5417, w_083_5418, w_083_5424, w_083_5428, w_083_5431, w_083_5433, w_083_5436, w_083_5442, w_083_5443, w_083_5448, w_083_5452, w_083_5454, w_083_5456, w_083_5457, w_083_5459, w_083_5467, w_083_5469, w_083_5470, w_083_5474, w_083_5480, w_083_5483, w_083_5496, w_083_5501, w_083_5503, w_083_5504, w_083_5512, w_083_5514, w_083_5519, w_083_5521, w_083_5524, w_083_5532, w_083_5536, w_083_5539, w_083_5546, w_083_5547, w_083_5552, w_083_5555, w_083_5559, w_083_5560, w_083_5563, w_083_5572, w_083_5574, w_083_5578, w_083_5590, w_083_5593, w_083_5594, w_083_5596, w_083_5607, w_083_5610, w_083_5611, w_083_5616, w_083_5618, w_083_5620, w_083_5626, w_083_5628, w_083_5647, w_083_5651, w_083_5654, w_083_5656, w_083_5659, w_083_5662, w_083_5664, w_083_5665, w_083_5666, w_083_5667, w_083_5670, w_083_5672, w_083_5677, w_083_5679, w_083_5690, w_083_5693, w_083_5694, w_083_5695, w_083_5702, w_083_5706, w_083_5708, w_083_5710, w_083_5712, w_083_5713, w_083_5717, w_083_5719, w_083_5720, w_083_5722, w_083_5737, w_083_5743, w_083_5745, w_083_5753, w_083_5757, w_083_5758, w_083_5762, w_083_5769, w_083_5772, w_083_5774, w_083_5777, w_083_5778, w_083_5779, w_083_5784, w_083_5795, w_083_5798, w_083_5801, w_083_5804, w_083_5808, w_083_5809, w_083_5816, w_083_5817, w_083_5820, w_083_5826, w_083_5834, w_083_5835, w_083_5843, w_083_5844, w_083_5848, w_083_5850, w_083_5865, w_083_5869, w_083_5873, w_083_5879, w_083_5883, w_083_5886, w_083_5888, w_083_5890, w_083_5891, w_083_5895, w_083_5897, w_083_5901, w_083_5903, w_083_5906, w_083_5908, w_083_5909, w_083_5910, w_083_5913, w_083_5917, w_083_5921, w_083_5923, w_083_5924, w_083_5926, w_083_5930, w_083_5931, w_083_5934, w_083_5940, w_083_5945, w_083_5946, w_083_5950, w_083_5961, w_083_5962, w_083_5963, w_083_5966, w_083_5979, w_083_5986, w_083_5996, w_083_6001, w_083_6002, w_083_6006, w_083_6007, w_083_6009, w_083_6010, w_083_6016, w_083_6018, w_083_6020, w_083_6022, w_083_6023, w_083_6032, w_083_6037, w_083_6044, w_083_6051, w_083_6054, w_083_6056, w_083_6057, w_083_6058, w_083_6062, w_083_6065, w_083_6067, w_083_6069, w_083_6070, w_083_6074, w_083_6075, w_083_6083, w_083_6087, w_083_6100, w_083_6101, w_083_6103, w_083_6123, w_083_6127, w_083_6129, w_083_6133, w_083_6137, w_083_6144, w_083_6145, w_083_6147, w_083_6150, w_083_6153, w_083_6154, w_083_6155, w_083_6159, w_083_6162, w_083_6164, w_083_6167, w_083_6172, w_083_6173, w_083_6177, w_083_6178, w_083_6183, w_083_6185, w_083_6197, w_083_6215, w_083_6216, w_083_6223, w_083_6224, w_083_6227, w_083_6230, w_083_6231, w_083_6238, w_083_6243, w_083_6244, w_083_6249, w_083_6250, w_083_6251, w_083_6258, w_083_6263, w_083_6265, w_083_6271, w_083_6272, w_083_6273, w_083_6277, w_083_6278, w_083_6279, w_083_6285, w_083_6287, w_083_6288, w_083_6291, w_083_6296, w_083_6302, w_083_6303, w_083_6304, w_083_6305, w_083_6309, w_083_6311, w_083_6312, w_083_6314, w_083_6316, w_083_6317, w_083_6318, w_083_6319, w_083_6320, w_083_6328, w_083_6329, w_083_6332, w_083_6337, w_083_6339, w_083_6343, w_083_6354, w_083_6356, w_083_6357, w_083_6358, w_083_6360, w_083_6361, w_083_6362, w_083_6366, w_083_6368, w_083_6374, w_083_6380, w_083_6390, w_083_6392, w_083_6396, w_083_6399, w_083_6403, w_083_6404, w_083_6405, w_083_6407, w_083_6409, w_083_6411, w_083_6413, w_083_6420, w_083_6422, w_083_6425, w_083_6427, w_083_6430, w_083_6432, w_083_6435, w_083_6441, w_083_6446, w_083_6451, w_083_6455, w_083_6456, w_083_6457, w_083_6460, w_083_6464, w_083_6466, w_083_6469, w_083_6476, w_083_6481, w_083_6483, w_083_6486, w_083_6490, w_083_6493, w_083_6500, w_083_6505, w_083_6510, w_083_6519, w_083_6520, w_083_6526, w_083_6530, w_083_6532, w_083_6534, w_083_6540, w_083_6544, w_083_6549, w_083_6553, w_083_6555, w_083_6558, w_083_6560, w_083_6561, w_083_6565, w_083_6569, w_083_6571, w_083_6575, w_083_6577, w_083_6582, w_083_6586, w_083_6591, w_083_6593, w_083_6598, w_083_6599, w_083_6611, w_083_6616, w_083_6628, w_083_6630, w_083_6634, w_083_6646, w_083_6650, w_083_6655, w_083_6656, w_083_6657, w_083_6658, w_083_6662, w_083_6665, w_083_6669, w_083_6674, w_083_6675, w_083_6678, w_083_6683, w_083_6690, w_083_6695, w_083_6701, w_083_6702, w_083_6704, w_083_6709, w_083_6711, w_083_6713, w_083_6715, w_083_6716, w_083_6717, w_083_6718, w_083_6720, w_083_6725, w_083_6727, w_083_6731, w_083_6732, w_083_6736, w_083_6744, w_083_6745, w_083_6750, w_083_6755, w_083_6756, w_083_6759, w_083_6764, w_083_6771, w_083_6772, w_083_6775, w_083_6777, w_083_6778, w_083_6783, w_083_6787, w_083_6796, w_083_6797, w_083_6800, w_083_6801, w_083_6803, w_083_6812, w_083_6816, w_083_6817, w_083_6818, w_083_6819, w_083_6820, w_083_6834, w_083_6836, w_083_6839, w_083_6842, w_083_6848, w_083_6852, w_083_6860, w_083_6863, w_083_6865, w_083_6866, w_083_6867, w_083_6868, w_083_6875, w_083_6876, w_083_6880, w_083_6884, w_083_6885, w_083_6889, w_083_6891, w_083_6892, w_083_6895, w_083_6897, w_083_6902, w_083_6903, w_083_6911, w_083_6917, w_083_6921, w_083_6922, w_083_6923, w_083_6924, w_083_6927, w_083_6928, w_083_6936, w_083_6937, w_083_6942, w_083_6947, w_083_6948, w_083_6950, w_083_6951, w_083_6952, w_083_6953, w_083_6955, w_083_6959, w_083_6972, w_083_6974, w_083_6983, w_083_6984, w_083_6986, w_083_6990, w_083_6992, w_083_6995, w_083_6996, w_083_6997, w_083_7006, w_083_7007, w_083_7009, w_083_7010, w_083_7012, w_083_7015, w_083_7016, w_083_7025, w_083_7028, w_083_7029, w_083_7031, w_083_7032, w_083_7035, w_083_7038, w_083_7040, w_083_7043, w_083_7045, w_083_7050, w_083_7052, w_083_7053, w_083_7056, w_083_7059, w_083_7061, w_083_7064, w_083_7065, w_083_7068, w_083_7073, w_083_7082, w_083_7083, w_083_7084, w_083_7100, w_083_7101, w_083_7102, w_083_7104, w_083_7106, w_083_7111, w_083_7112, w_083_7115, w_083_7117, w_083_7120, w_083_7123, w_083_7137, w_083_7142, w_083_7152, w_083_7160, w_083_7162, w_083_7169, w_083_7172, w_083_7176, w_083_7177, w_083_7181, w_083_7184, w_083_7192, w_083_7197, w_083_7198, w_083_7209, w_083_7210, w_083_7212, w_083_7215, w_083_7216, w_083_7219, w_083_7222, w_083_7226, w_083_7228, w_083_7229, w_083_7231, w_083_7237, w_083_7244, w_083_7249, w_083_7251, w_083_7255, w_083_7264, w_083_7266, w_083_7270, w_083_7272, w_083_7274, w_083_7276, w_083_7283, w_083_7286, w_083_7290, w_083_7291, w_083_7293, w_083_7297, w_083_7298, w_083_7301, w_083_7302, w_083_7304, w_083_7306, w_083_7307, w_083_7310, w_083_7311, w_083_7316, w_083_7319, w_083_7323, w_083_7324, w_083_7325, w_083_7328, w_083_7335, w_083_7345, w_083_7346, w_083_7349, w_083_7350, w_083_7354, w_083_7355, w_083_7356, w_083_7357, w_083_7359, w_083_7361, w_083_7363, w_083_7367, w_083_7370, w_083_7372, w_083_7374, w_083_7378, w_083_7382, w_083_7383, w_083_7390, w_083_7392, w_083_7393, w_083_7397, w_083_7407, w_083_7421, w_083_7425, w_083_7428, w_083_7438, w_083_7440, w_083_7441, w_083_7446, w_083_7449, w_083_7450, w_083_7462, w_083_7465, w_083_7469, w_083_7471, w_083_7478, w_083_7479, w_083_7488, w_083_7489, w_083_7495, w_083_7501, w_083_7502, w_083_7508, w_083_7516, w_083_7519, w_083_7520, w_083_7525, w_083_7526, w_083_7527, w_083_7530, w_083_7531, w_083_7534, w_083_7537, w_083_7540, w_083_7549, w_083_7550, w_083_7555, w_083_7557, w_083_7559, w_083_7561, w_083_7568, w_083_7569, w_083_7571, w_083_7572, w_083_7577, w_083_7578, w_083_7588, w_083_7589, w_083_7590, w_083_7593, w_083_7595, w_083_7596, w_083_7599, w_083_7600, w_083_7603, w_083_7604, w_083_7608, w_083_7610, w_083_7613, w_083_7623, w_083_7629, w_083_7631, w_083_7632, w_083_7639, w_083_7644;
  wire w_084_000, w_084_001, w_084_003, w_084_004, w_084_006, w_084_007, w_084_008, w_084_010, w_084_011, w_084_014, w_084_015, w_084_016, w_084_017, w_084_020, w_084_021, w_084_022, w_084_023, w_084_025, w_084_026, w_084_027, w_084_028, w_084_029, w_084_030, w_084_032, w_084_034, w_084_035, w_084_036, w_084_037, w_084_038, w_084_039, w_084_042, w_084_043, w_084_044, w_084_045, w_084_046, w_084_047, w_084_048, w_084_049, w_084_050, w_084_051, w_084_052, w_084_053, w_084_054, w_084_055, w_084_056, w_084_057, w_084_058, w_084_059, w_084_060, w_084_061, w_084_062, w_084_063, w_084_064, w_084_065, w_084_066, w_084_068, w_084_069, w_084_070, w_084_073, w_084_074, w_084_075, w_084_077, w_084_078, w_084_079, w_084_081, w_084_082, w_084_085, w_084_086, w_084_087, w_084_088, w_084_089, w_084_090, w_084_091, w_084_093, w_084_095, w_084_096, w_084_097, w_084_098, w_084_100, w_084_101, w_084_102, w_084_103, w_084_104, w_084_105, w_084_106, w_084_107, w_084_108, w_084_109, w_084_110, w_084_111, w_084_112, w_084_113, w_084_114, w_084_115, w_084_116, w_084_117, w_084_118, w_084_119, w_084_120, w_084_122, w_084_123, w_084_124, w_084_125, w_084_126, w_084_127, w_084_128, w_084_129, w_084_130, w_084_131, w_084_132, w_084_133, w_084_134, w_084_136, w_084_137, w_084_138, w_084_140, w_084_141, w_084_142, w_084_143, w_084_145, w_084_146, w_084_147, w_084_148, w_084_150, w_084_151, w_084_152, w_084_153, w_084_154, w_084_155, w_084_156, w_084_157, w_084_158, w_084_159, w_084_161, w_084_162, w_084_163, w_084_164, w_084_165, w_084_167, w_084_168, w_084_169, w_084_170, w_084_172, w_084_173, w_084_174, w_084_175, w_084_177, w_084_178, w_084_179, w_084_182, w_084_183, w_084_184, w_084_185, w_084_186, w_084_187, w_084_188, w_084_190, w_084_191, w_084_193, w_084_194, w_084_195, w_084_196, w_084_198, w_084_199, w_084_200, w_084_202, w_084_203, w_084_204, w_084_205, w_084_206, w_084_207, w_084_208, w_084_210, w_084_211, w_084_212, w_084_213, w_084_214, w_084_215, w_084_216, w_084_218, w_084_219, w_084_220, w_084_221, w_084_222, w_084_223, w_084_224, w_084_227, w_084_228, w_084_229, w_084_230, w_084_231, w_084_232, w_084_233, w_084_234, w_084_235, w_084_236, w_084_237, w_084_239, w_084_240, w_084_241, w_084_242, w_084_243, w_084_244, w_084_245, w_084_246, w_084_247, w_084_248, w_084_249, w_084_250, w_084_251, w_084_252, w_084_253, w_084_254, w_084_256, w_084_258, w_084_259, w_084_260, w_084_261, w_084_262, w_084_263, w_084_264, w_084_265, w_084_266, w_084_267, w_084_268, w_084_269, w_084_270, w_084_271, w_084_272, w_084_274, w_084_275, w_084_276, w_084_277, w_084_279, w_084_281, w_084_282, w_084_284, w_084_285, w_084_287, w_084_289, w_084_290, w_084_291, w_084_293, w_084_294, w_084_295, w_084_296, w_084_298, w_084_299, w_084_300, w_084_301, w_084_302, w_084_303, w_084_304, w_084_305, w_084_306, w_084_307, w_084_308, w_084_309, w_084_310, w_084_311, w_084_312, w_084_313, w_084_314, w_084_316, w_084_317, w_084_318, w_084_319, w_084_320, w_084_321, w_084_322, w_084_323, w_084_326, w_084_327, w_084_328, w_084_329, w_084_330, w_084_331, w_084_332, w_084_333, w_084_334, w_084_335, w_084_336, w_084_338, w_084_339, w_084_340, w_084_341, w_084_342, w_084_343, w_084_344, w_084_345, w_084_346, w_084_347, w_084_348, w_084_349, w_084_350, w_084_351, w_084_352, w_084_354, w_084_355, w_084_356, w_084_357, w_084_358, w_084_359, w_084_360, w_084_361, w_084_362, w_084_363, w_084_364, w_084_365, w_084_366, w_084_367, w_084_371, w_084_372, w_084_373, w_084_375, w_084_376, w_084_378, w_084_379, w_084_380, w_084_381, w_084_382, w_084_383, w_084_385, w_084_386, w_084_387, w_084_388, w_084_389, w_084_390, w_084_391, w_084_392, w_084_393, w_084_394, w_084_395, w_084_396, w_084_397, w_084_398, w_084_399, w_084_400, w_084_401, w_084_402, w_084_403, w_084_404, w_084_405, w_084_406, w_084_407, w_084_408, w_084_409, w_084_410, w_084_412, w_084_413, w_084_414, w_084_415, w_084_416, w_084_417, w_084_418, w_084_419, w_084_420, w_084_421, w_084_422, w_084_423, w_084_424, w_084_425, w_084_426, w_084_427, w_084_430, w_084_431, w_084_432, w_084_433, w_084_435, w_084_436, w_084_437, w_084_438, w_084_439, w_084_441, w_084_442, w_084_443, w_084_445, w_084_446, w_084_447, w_084_448, w_084_449, w_084_450, w_084_451, w_084_452, w_084_453, w_084_454, w_084_455, w_084_456, w_084_457, w_084_459, w_084_460, w_084_461, w_084_463, w_084_464, w_084_465, w_084_466, w_084_468, w_084_469, w_084_470, w_084_472, w_084_473, w_084_476, w_084_477, w_084_478, w_084_479, w_084_480, w_084_481, w_084_483, w_084_484, w_084_485, w_084_486, w_084_488, w_084_489, w_084_490, w_084_491, w_084_492, w_084_493, w_084_494, w_084_495, w_084_496, w_084_497, w_084_498, w_084_499, w_084_500, w_084_501, w_084_502, w_084_503, w_084_505, w_084_508, w_084_509, w_084_510, w_084_511, w_084_512, w_084_513, w_084_515, w_084_516, w_084_517, w_084_519, w_084_520, w_084_521, w_084_522, w_084_523, w_084_524, w_084_525, w_084_526, w_084_528, w_084_529, w_084_531, w_084_532, w_084_533, w_084_534, w_084_535, w_084_536, w_084_539, w_084_540, w_084_541, w_084_542, w_084_543, w_084_544, w_084_545, w_084_546, w_084_547, w_084_548, w_084_549, w_084_550, w_084_551, w_084_552, w_084_553, w_084_554, w_084_555, w_084_556, w_084_557, w_084_558, w_084_560, w_084_561, w_084_562, w_084_563, w_084_564, w_084_565, w_084_566, w_084_568, w_084_569, w_084_570, w_084_571, w_084_572, w_084_573, w_084_575, w_084_576, w_084_577, w_084_578, w_084_580, w_084_581, w_084_583, w_084_584, w_084_585, w_084_587, w_084_588, w_084_589, w_084_590, w_084_591, w_084_592, w_084_593, w_084_594, w_084_595, w_084_596, w_084_598, w_084_599, w_084_600, w_084_601, w_084_602, w_084_603, w_084_604, w_084_605, w_084_606, w_084_608, w_084_609, w_084_610, w_084_611, w_084_612, w_084_613, w_084_614, w_084_615, w_084_616, w_084_617, w_084_618, w_084_620, w_084_621, w_084_622, w_084_623, w_084_624, w_084_625, w_084_626, w_084_628, w_084_629, w_084_630, w_084_631, w_084_632, w_084_634, w_084_635, w_084_636, w_084_637, w_084_638, w_084_640, w_084_641, w_084_642, w_084_643, w_084_644, w_084_645, w_084_646, w_084_647, w_084_649, w_084_650, w_084_651, w_084_652, w_084_653, w_084_654, w_084_655, w_084_656, w_084_657, w_084_659, w_084_660, w_084_661, w_084_663, w_084_664, w_084_665, w_084_666, w_084_667, w_084_669, w_084_670, w_084_671, w_084_672, w_084_673, w_084_674, w_084_675, w_084_676, w_084_677, w_084_679, w_084_680, w_084_681, w_084_682, w_084_683, w_084_684, w_084_685, w_084_686, w_084_687, w_084_688, w_084_689, w_084_690, w_084_691, w_084_692, w_084_693, w_084_694, w_084_696, w_084_697, w_084_699, w_084_700, w_084_701, w_084_702, w_084_703, w_084_704, w_084_706, w_084_707, w_084_708, w_084_709, w_084_710, w_084_711, w_084_712, w_084_713, w_084_715, w_084_716, w_084_717, w_084_718, w_084_720, w_084_721, w_084_722, w_084_723, w_084_724, w_084_725, w_084_726, w_084_729, w_084_731, w_084_733, w_084_734, w_084_735, w_084_736, w_084_737, w_084_738, w_084_739, w_084_740, w_084_742, w_084_743, w_084_745, w_084_746, w_084_747, w_084_748, w_084_749, w_084_750, w_084_751, w_084_753, w_084_754, w_084_755, w_084_756, w_084_758, w_084_759, w_084_760, w_084_761, w_084_762, w_084_763, w_084_764, w_084_766, w_084_768, w_084_769, w_084_770, w_084_771, w_084_772, w_084_773, w_084_774, w_084_775, w_084_776, w_084_777, w_084_778, w_084_781, w_084_782, w_084_784, w_084_785, w_084_786, w_084_787, w_084_788, w_084_789, w_084_790, w_084_792, w_084_793, w_084_794, w_084_795, w_084_796, w_084_797, w_084_798, w_084_799, w_084_800, w_084_801, w_084_802, w_084_803, w_084_804, w_084_805, w_084_806, w_084_807, w_084_808, w_084_809, w_084_810, w_084_811, w_084_812, w_084_813, w_084_814, w_084_815, w_084_816, w_084_817, w_084_818, w_084_819, w_084_820, w_084_821, w_084_822, w_084_824, w_084_825, w_084_826, w_084_827, w_084_828, w_084_829, w_084_830, w_084_831, w_084_832, w_084_833, w_084_834, w_084_835, w_084_836, w_084_837, w_084_838, w_084_839, w_084_840, w_084_841, w_084_842, w_084_843, w_084_844, w_084_845, w_084_846, w_084_847, w_084_848, w_084_849, w_084_850, w_084_851, w_084_852, w_084_853, w_084_854, w_084_856, w_084_857, w_084_858, w_084_859, w_084_861, w_084_862, w_084_864, w_084_865, w_084_867, w_084_868, w_084_869, w_084_870, w_084_871, w_084_872, w_084_873, w_084_874, w_084_875, w_084_876, w_084_877, w_084_879, w_084_882, w_084_883, w_084_884, w_084_885, w_084_886, w_084_887, w_084_888, w_084_889, w_084_890, w_084_891, w_084_892, w_084_893, w_084_894, w_084_895, w_084_896, w_084_897, w_084_900, w_084_901, w_084_902, w_084_903, w_084_904, w_084_905, w_084_906, w_084_907, w_084_909, w_084_911, w_084_912, w_084_913, w_084_915, w_084_916, w_084_917, w_084_918, w_084_919, w_084_921, w_084_922, w_084_923, w_084_925, w_084_926, w_084_927, w_084_928, w_084_929, w_084_931, w_084_933, w_084_934, w_084_935, w_084_936, w_084_937, w_084_938, w_084_940, w_084_941, w_084_942, w_084_943, w_084_944, w_084_945, w_084_946, w_084_947, w_084_948, w_084_949, w_084_950, w_084_951, w_084_952, w_084_953, w_084_955, w_084_956, w_084_957, w_084_958, w_084_959, w_084_960, w_084_961, w_084_962, w_084_963, w_084_964, w_084_965, w_084_966, w_084_967, w_084_968, w_084_969, w_084_970, w_084_971, w_084_972, w_084_974, w_084_975, w_084_976, w_084_977, w_084_978, w_084_979, w_084_981, w_084_982, w_084_983, w_084_984, w_084_985, w_084_986, w_084_987, w_084_988, w_084_989, w_084_990, w_084_992, w_084_993, w_084_994, w_084_995, w_084_996, w_084_997, w_084_998, w_084_999, w_084_1000, w_084_1002, w_084_1003, w_084_1004, w_084_1005, w_084_1006, w_084_1007, w_084_1008, w_084_1009, w_084_1010, w_084_1012, w_084_1014, w_084_1015, w_084_1016, w_084_1017, w_084_1018, w_084_1019, w_084_1020, w_084_1022, w_084_1023, w_084_1025, w_084_1027, w_084_1028, w_084_1029, w_084_1030, w_084_1031, w_084_1032, w_084_1033, w_084_1034, w_084_1035, w_084_1036, w_084_1037, w_084_1038, w_084_1040, w_084_1041, w_084_1043, w_084_1044, w_084_1045, w_084_1046, w_084_1047, w_084_1048, w_084_1049, w_084_1050, w_084_1051, w_084_1053, w_084_1054, w_084_1055, w_084_1056, w_084_1057, w_084_1058, w_084_1059, w_084_1060, w_084_1063, w_084_1064, w_084_1065, w_084_1067, w_084_1068, w_084_1069, w_084_1070, w_084_1071, w_084_1075, w_084_1077, w_084_1078, w_084_1079, w_084_1080, w_084_1081, w_084_1082, w_084_1083, w_084_1084, w_084_1085, w_084_1086, w_084_1087, w_084_1088, w_084_1089, w_084_1090, w_084_1091, w_084_1093, w_084_1094, w_084_1095, w_084_1096, w_084_1097, w_084_1098, w_084_1099, w_084_1100, w_084_1101, w_084_1102, w_084_1103, w_084_1104, w_084_1105, w_084_1106, w_084_1107, w_084_1108, w_084_1109, w_084_1110, w_084_1112, w_084_1114, w_084_1116, w_084_1117, w_084_1118, w_084_1119, w_084_1120, w_084_1122, w_084_1123, w_084_1124, w_084_1125, w_084_1126, w_084_1127, w_084_1128, w_084_1129, w_084_1130, w_084_1132, w_084_1133, w_084_1134, w_084_1136, w_084_1137, w_084_1138, w_084_1139, w_084_1140, w_084_1141, w_084_1143, w_084_1144, w_084_1145, w_084_1146, w_084_1147, w_084_1148, w_084_1149, w_084_1152, w_084_1153, w_084_1154, w_084_1155, w_084_1156, w_084_1157, w_084_1158, w_084_1159, w_084_1160, w_084_1161, w_084_1163, w_084_1166, w_084_1167, w_084_1168, w_084_1172, w_084_1173, w_084_1174, w_084_1175, w_084_1176, w_084_1178, w_084_1180, w_084_1182, w_084_1184, w_084_1185, w_084_1186, w_084_1187, w_084_1188, w_084_1189, w_084_1190, w_084_1191, w_084_1192, w_084_1195, w_084_1196, w_084_1197, w_084_1199, w_084_1203, w_084_1206, w_084_1207, w_084_1208, w_084_1209, w_084_1210, w_084_1211, w_084_1212, w_084_1213, w_084_1214, w_084_1215, w_084_1216, w_084_1217, w_084_1218, w_084_1220, w_084_1221, w_084_1222, w_084_1223, w_084_1224, w_084_1225, w_084_1226, w_084_1227, w_084_1228, w_084_1229, w_084_1230, w_084_1231, w_084_1232, w_084_1234, w_084_1235, w_084_1236, w_084_1237, w_084_1238, w_084_1239, w_084_1240, w_084_1241, w_084_1242, w_084_1243, w_084_1244, w_084_1246, w_084_1247, w_084_1248, w_084_1249, w_084_1251, w_084_1252, w_084_1254, w_084_1256, w_084_1257, w_084_1259, w_084_1260, w_084_1261, w_084_1262, w_084_1263, w_084_1264, w_084_1265, w_084_1268, w_084_1270, w_084_1271, w_084_1272, w_084_1274, w_084_1276, w_084_1277, w_084_1278, w_084_1279, w_084_1280, w_084_1282, w_084_1283, w_084_1284, w_084_1285, w_084_1287, w_084_1289, w_084_1290, w_084_1291, w_084_1294, w_084_1295, w_084_1296, w_084_1297, w_084_1300, w_084_1302, w_084_1303, w_084_1304, w_084_1305, w_084_1306, w_084_1307, w_084_1309, w_084_1310, w_084_1311, w_084_1312, w_084_1313, w_084_1315, w_084_1316, w_084_1317, w_084_1318, w_084_1319, w_084_1320, w_084_1321, w_084_1322, w_084_1323, w_084_1324, w_084_1325, w_084_1326, w_084_1327, w_084_1328, w_084_1329, w_084_1332, w_084_1333, w_084_1335, w_084_1336, w_084_1338, w_084_1340, w_084_1341, w_084_1342, w_084_1343, w_084_1345, w_084_1346, w_084_1347, w_084_1348, w_084_1350, w_084_1351, w_084_1353, w_084_1354, w_084_1356, w_084_1357, w_084_1358, w_084_1360, w_084_1361, w_084_1362, w_084_1364, w_084_1366, w_084_1367, w_084_1368, w_084_1369, w_084_1370, w_084_1371, w_084_1373, w_084_1375, w_084_1376, w_084_1377, w_084_1378, w_084_1379, w_084_1380, w_084_1381, w_084_1383, w_084_1384, w_084_1385, w_084_1386, w_084_1387, w_084_1388, w_084_1389, w_084_1390, w_084_1392, w_084_1393, w_084_1394, w_084_1395, w_084_1397, w_084_1398, w_084_1400, w_084_1401, w_084_1402, w_084_1403, w_084_1404, w_084_1405, w_084_1407, w_084_1408, w_084_1409, w_084_1410, w_084_1411, w_084_1412, w_084_1413, w_084_1414, w_084_1415, w_084_1416, w_084_1417, w_084_1418, w_084_1420, w_084_1421, w_084_1422, w_084_1423, w_084_1425, w_084_1426, w_084_1427, w_084_1428, w_084_1429, w_084_1430, w_084_1432, w_084_1433, w_084_1434, w_084_1436, w_084_1437, w_084_1438, w_084_1440, w_084_1441, w_084_1442, w_084_1443, w_084_1444, w_084_1445, w_084_1447, w_084_1448, w_084_1449, w_084_1450, w_084_1452, w_084_1453, w_084_1454, w_084_1455, w_084_1456, w_084_1457, w_084_1458, w_084_1461, w_084_1462, w_084_1465, w_084_1467, w_084_1469, w_084_1470, w_084_1471, w_084_1472, w_084_1473, w_084_1474, w_084_1475, w_084_1476, w_084_1477, w_084_1479, w_084_1480, w_084_1481, w_084_1482, w_084_1483, w_084_1484, w_084_1485, w_084_1486, w_084_1489, w_084_1490, w_084_1493, w_084_1494, w_084_1497, w_084_1498, w_084_1499, w_084_1500, w_084_1501, w_084_1502, w_084_1503, w_084_1505, w_084_1506, w_084_1507, w_084_1508, w_084_1510, w_084_1511, w_084_1512, w_084_1514, w_084_1515, w_084_1516, w_084_1517, w_084_1519, w_084_1520, w_084_1521, w_084_1522, w_084_1523, w_084_1525, w_084_1526, w_084_1527, w_084_1529, w_084_1531, w_084_1532, w_084_1534, w_084_1536, w_084_1537, w_084_1538, w_084_1539, w_084_1540, w_084_1541, w_084_1542, w_084_1544, w_084_1545, w_084_1549, w_084_1551, w_084_1552, w_084_1553, w_084_1554, w_084_1555, w_084_1558, w_084_1559, w_084_1561, w_084_1562, w_084_1563, w_084_1564, w_084_1565, w_084_1567, w_084_1568, w_084_1569, w_084_1570, w_084_1571, w_084_1572, w_084_1573, w_084_1574, w_084_1575, w_084_1576, w_084_1577, w_084_1578, w_084_1579, w_084_1580, w_084_1581, w_084_1582, w_084_1583, w_084_1584, w_084_1585, w_084_1588, w_084_1589, w_084_1590, w_084_1591, w_084_1592, w_084_1593, w_084_1594, w_084_1595, w_084_1596, w_084_1597, w_084_1598, w_084_1599, w_084_1600, w_084_1602, w_084_1603, w_084_1604, w_084_1608, w_084_1609, w_084_1611, w_084_1612, w_084_1614, w_084_1615, w_084_1616, w_084_1617, w_084_1618, w_084_1619, w_084_1622, w_084_1623, w_084_1624, w_084_1627, w_084_1629, w_084_1630, w_084_1631, w_084_1632, w_084_1633, w_084_1634, w_084_1635, w_084_1636, w_084_1637, w_084_1638, w_084_1639, w_084_1641, w_084_1642, w_084_1643, w_084_1644, w_084_1645, w_084_1646, w_084_1647, w_084_1649, w_084_1650, w_084_1651, w_084_1652, w_084_1653, w_084_1654, w_084_1655, w_084_1656, w_084_1657, w_084_1660, w_084_1661, w_084_1662, w_084_1665, w_084_1667, w_084_1668, w_084_1669, w_084_1670, w_084_1671, w_084_1672, w_084_1673, w_084_1674, w_084_1675, w_084_1676, w_084_1677, w_084_1678, w_084_1679, w_084_1680, w_084_1681, w_084_1682, w_084_1683, w_084_1684, w_084_1685, w_084_1686, w_084_1688, w_084_1690, w_084_1691, w_084_1692, w_084_1693, w_084_1694, w_084_1696, w_084_1699, w_084_1700, w_084_1703, w_084_1704, w_084_1705, w_084_1706, w_084_1707, w_084_1709, w_084_1710, w_084_1711, w_084_1712, w_084_1713, w_084_1714, w_084_1715, w_084_1716, w_084_1717, w_084_1718, w_084_1719, w_084_1721, w_084_1723, w_084_1724, w_084_1725, w_084_1726, w_084_1727, w_084_1728, w_084_1729, w_084_1730, w_084_1731, w_084_1734, w_084_1735, w_084_1737, w_084_1738, w_084_1739, w_084_1740, w_084_1743, w_084_1744, w_084_1745, w_084_1747, w_084_1748, w_084_1749, w_084_1750, w_084_1751, w_084_1753, w_084_1755, w_084_1757, w_084_1758, w_084_1759, w_084_1761;
  wire w_085_001, w_085_003, w_085_004, w_085_007, w_085_010, w_085_012, w_085_013, w_085_016, w_085_017, w_085_018, w_085_019, w_085_023, w_085_025, w_085_028, w_085_029, w_085_030, w_085_031, w_085_032, w_085_033, w_085_035, w_085_036, w_085_037, w_085_038, w_085_040, w_085_041, w_085_045, w_085_048, w_085_049, w_085_050, w_085_051, w_085_052, w_085_053, w_085_055, w_085_056, w_085_057, w_085_059, w_085_061, w_085_063, w_085_064, w_085_065, w_085_067, w_085_068, w_085_073, w_085_074, w_085_083, w_085_088, w_085_089, w_085_100, w_085_103, w_085_108, w_085_110, w_085_112, w_085_113, w_085_116, w_085_117, w_085_119, w_085_120, w_085_123, w_085_129, w_085_130, w_085_137, w_085_139, w_085_141, w_085_142, w_085_143, w_085_144, w_085_145, w_085_150, w_085_151, w_085_154, w_085_158, w_085_165, w_085_166, w_085_167, w_085_169, w_085_171, w_085_172, w_085_173, w_085_174, w_085_176, w_085_178, w_085_180, w_085_182, w_085_185, w_085_190, w_085_191, w_085_192, w_085_194, w_085_195, w_085_197, w_085_198, w_085_203, w_085_204, w_085_205, w_085_208, w_085_211, w_085_213, w_085_214, w_085_218, w_085_219, w_085_222, w_085_223, w_085_226, w_085_227, w_085_228, w_085_229, w_085_233, w_085_234, w_085_235, w_085_236, w_085_239, w_085_240, w_085_244, w_085_250, w_085_255, w_085_256, w_085_257, w_085_258, w_085_261, w_085_262, w_085_265, w_085_266, w_085_267, w_085_269, w_085_271, w_085_272, w_085_276, w_085_277, w_085_279, w_085_285, w_085_287, w_085_288, w_085_291, w_085_292, w_085_294, w_085_296, w_085_299, w_085_300, w_085_301, w_085_303, w_085_306, w_085_307, w_085_318, w_085_320, w_085_321, w_085_326, w_085_328, w_085_329, w_085_331, w_085_339, w_085_344, w_085_345, w_085_346, w_085_347, w_085_348, w_085_349, w_085_350, w_085_351, w_085_354, w_085_356, w_085_357, w_085_358, w_085_362, w_085_363, w_085_367, w_085_369, w_085_371, w_085_375, w_085_376, w_085_378, w_085_379, w_085_380, w_085_384, w_085_388, w_085_396, w_085_400, w_085_401, w_085_404, w_085_406, w_085_409, w_085_410, w_085_412, w_085_414, w_085_415, w_085_416, w_085_417, w_085_418, w_085_420, w_085_425, w_085_426, w_085_428, w_085_430, w_085_433, w_085_436, w_085_444, w_085_446, w_085_448, w_085_450, w_085_451, w_085_452, w_085_453, w_085_457, w_085_459, w_085_461, w_085_462, w_085_466, w_085_469, w_085_472, w_085_477, w_085_480, w_085_481, w_085_482, w_085_483, w_085_489, w_085_490, w_085_491, w_085_494, w_085_495, w_085_497, w_085_498, w_085_499, w_085_501, w_085_505, w_085_506, w_085_507, w_085_511, w_085_512, w_085_513, w_085_514, w_085_515, w_085_516, w_085_517, w_085_518, w_085_522, w_085_524, w_085_525, w_085_526, w_085_527, w_085_531, w_085_533, w_085_534, w_085_543, w_085_546, w_085_547, w_085_551, w_085_552, w_085_556, w_085_559, w_085_560, w_085_561, w_085_566, w_085_567, w_085_568, w_085_571, w_085_576, w_085_577, w_085_578, w_085_580, w_085_581, w_085_583, w_085_587, w_085_592, w_085_594, w_085_595, w_085_596, w_085_598, w_085_599, w_085_602, w_085_603, w_085_605, w_085_609, w_085_611, w_085_614, w_085_615, w_085_618, w_085_620, w_085_623, w_085_624, w_085_628, w_085_630, w_085_632, w_085_633, w_085_634, w_085_635, w_085_639, w_085_642, w_085_646, w_085_648, w_085_652, w_085_653, w_085_657, w_085_660, w_085_662, w_085_664, w_085_666, w_085_667, w_085_669, w_085_670, w_085_671, w_085_673, w_085_674, w_085_676, w_085_677, w_085_678, w_085_679, w_085_683, w_085_685, w_085_686, w_085_687, w_085_690, w_085_691, w_085_692, w_085_694, w_085_695, w_085_696, w_085_698, w_085_702, w_085_706, w_085_707, w_085_711, w_085_712, w_085_715, w_085_716, w_085_718, w_085_724, w_085_725, w_085_727, w_085_728, w_085_729, w_085_732, w_085_734, w_085_735, w_085_738, w_085_739, w_085_740, w_085_741, w_085_744, w_085_745, w_085_747, w_085_750, w_085_753, w_085_754, w_085_757, w_085_759, w_085_760, w_085_764, w_085_765, w_085_767, w_085_770, w_085_775, w_085_776, w_085_779, w_085_781, w_085_782, w_085_783, w_085_784, w_085_786, w_085_787, w_085_789, w_085_790, w_085_794, w_085_795, w_085_798, w_085_800, w_085_803, w_085_806, w_085_807, w_085_810, w_085_812, w_085_817, w_085_818, w_085_821, w_085_822, w_085_823, w_085_825, w_085_828, w_085_835, w_085_837, w_085_838, w_085_840, w_085_841, w_085_845, w_085_850, w_085_851, w_085_856, w_085_858, w_085_860, w_085_862, w_085_866, w_085_867, w_085_871, w_085_873, w_085_878, w_085_880, w_085_881, w_085_884, w_085_888, w_085_890, w_085_892, w_085_893, w_085_895, w_085_896, w_085_905, w_085_908, w_085_911, w_085_915, w_085_917, w_085_920, w_085_921, w_085_922, w_085_923, w_085_925, w_085_929, w_085_930, w_085_932, w_085_934, w_085_936, w_085_937, w_085_940, w_085_941, w_085_944, w_085_947, w_085_948, w_085_949, w_085_950, w_085_951, w_085_952, w_085_953, w_085_955, w_085_957, w_085_960, w_085_964, w_085_966, w_085_968, w_085_969, w_085_971, w_085_974, w_085_977, w_085_978, w_085_979, w_085_983, w_085_988, w_085_989, w_085_990, w_085_992, w_085_993, w_085_997, w_085_999, w_085_1000, w_085_1001, w_085_1003, w_085_1005, w_085_1006, w_085_1009, w_085_1010, w_085_1011, w_085_1012, w_085_1015, w_085_1017, w_085_1018, w_085_1024, w_085_1025, w_085_1026, w_085_1028, w_085_1029, w_085_1032, w_085_1033, w_085_1034, w_085_1039, w_085_1040, w_085_1041, w_085_1042, w_085_1043, w_085_1045, w_085_1046, w_085_1047, w_085_1050, w_085_1051, w_085_1052, w_085_1054, w_085_1057, w_085_1058, w_085_1059, w_085_1064, w_085_1065, w_085_1066, w_085_1067, w_085_1073, w_085_1076, w_085_1077, w_085_1079, w_085_1081, w_085_1087, w_085_1092, w_085_1093, w_085_1094, w_085_1098, w_085_1099, w_085_1104, w_085_1106, w_085_1108, w_085_1109, w_085_1110, w_085_1111, w_085_1116, w_085_1120, w_085_1121, w_085_1122, w_085_1124, w_085_1127, w_085_1129, w_085_1135, w_085_1142, w_085_1143, w_085_1145, w_085_1147, w_085_1148, w_085_1149, w_085_1150, w_085_1152, w_085_1154, w_085_1155, w_085_1158, w_085_1159, w_085_1161, w_085_1163, w_085_1166, w_085_1167, w_085_1169, w_085_1171, w_085_1173, w_085_1175, w_085_1178, w_085_1179, w_085_1181, w_085_1182, w_085_1185, w_085_1186, w_085_1187, w_085_1192, w_085_1196, w_085_1198, w_085_1201, w_085_1204, w_085_1209, w_085_1211, w_085_1213, w_085_1215, w_085_1217, w_085_1218, w_085_1219, w_085_1220, w_085_1222, w_085_1223, w_085_1225, w_085_1227, w_085_1232, w_085_1233, w_085_1236, w_085_1237, w_085_1241, w_085_1243, w_085_1245, w_085_1246, w_085_1247, w_085_1251, w_085_1255, w_085_1256, w_085_1257, w_085_1258, w_085_1260, w_085_1263, w_085_1264, w_085_1265, w_085_1267, w_085_1270, w_085_1272, w_085_1276, w_085_1279, w_085_1284, w_085_1287, w_085_1290, w_085_1293, w_085_1297, w_085_1300, w_085_1302, w_085_1308, w_085_1311, w_085_1314, w_085_1316, w_085_1319, w_085_1321, w_085_1323, w_085_1325, w_085_1326, w_085_1327, w_085_1329, w_085_1332, w_085_1333, w_085_1334, w_085_1335, w_085_1338, w_085_1339, w_085_1340, w_085_1341, w_085_1342, w_085_1343, w_085_1346, w_085_1347, w_085_1348, w_085_1350, w_085_1353, w_085_1354, w_085_1356, w_085_1357, w_085_1361, w_085_1362, w_085_1364, w_085_1365, w_085_1369, w_085_1372, w_085_1379, w_085_1380, w_085_1381, w_085_1382, w_085_1383, w_085_1385, w_085_1386, w_085_1389, w_085_1392, w_085_1393, w_085_1394, w_085_1396, w_085_1397, w_085_1398, w_085_1403, w_085_1407, w_085_1410, w_085_1415, w_085_1420, w_085_1423, w_085_1424, w_085_1425, w_085_1427, w_085_1431, w_085_1436, w_085_1438, w_085_1441, w_085_1445, w_085_1446, w_085_1448, w_085_1449, w_085_1450, w_085_1452, w_085_1453, w_085_1454, w_085_1456, w_085_1459, w_085_1460, w_085_1464, w_085_1465, w_085_1466, w_085_1467, w_085_1469, w_085_1470, w_085_1471, w_085_1472, w_085_1482, w_085_1484, w_085_1486, w_085_1487, w_085_1489, w_085_1491, w_085_1493, w_085_1494, w_085_1496, w_085_1497, w_085_1498, w_085_1503, w_085_1505, w_085_1507, w_085_1511, w_085_1512, w_085_1514, w_085_1517, w_085_1528, w_085_1530, w_085_1533, w_085_1535, w_085_1538, w_085_1539, w_085_1543, w_085_1545, w_085_1549, w_085_1550, w_085_1551, w_085_1553, w_085_1557, w_085_1558, w_085_1560, w_085_1561, w_085_1564, w_085_1565, w_085_1566, w_085_1567, w_085_1569, w_085_1570, w_085_1571, w_085_1573, w_085_1574, w_085_1575, w_085_1582, w_085_1583, w_085_1584, w_085_1587, w_085_1590, w_085_1594, w_085_1598, w_085_1601, w_085_1604, w_085_1609, w_085_1610, w_085_1613, w_085_1617, w_085_1621, w_085_1622, w_085_1624, w_085_1625, w_085_1627, w_085_1629, w_085_1633, w_085_1636, w_085_1638, w_085_1639, w_085_1643, w_085_1644, w_085_1647, w_085_1652, w_085_1653, w_085_1654, w_085_1655, w_085_1659, w_085_1660, w_085_1661, w_085_1663, w_085_1665, w_085_1668, w_085_1671, w_085_1673, w_085_1676, w_085_1681, w_085_1682, w_085_1685, w_085_1687, w_085_1689, w_085_1692, w_085_1693, w_085_1698, w_085_1699, w_085_1703, w_085_1707, w_085_1710, w_085_1712, w_085_1713, w_085_1717, w_085_1718, w_085_1720, w_085_1721, w_085_1722, w_085_1723, w_085_1724, w_085_1725, w_085_1727, w_085_1728, w_085_1730, w_085_1731, w_085_1732, w_085_1733, w_085_1734, w_085_1735, w_085_1736, w_085_1737, w_085_1738, w_085_1741, w_085_1743, w_085_1746, w_085_1751, w_085_1755, w_085_1756, w_085_1757, w_085_1758, w_085_1760, w_085_1761, w_085_1763, w_085_1764, w_085_1765, w_085_1766, w_085_1767, w_085_1769, w_085_1770, w_085_1772, w_085_1773, w_085_1775, w_085_1777, w_085_1780, w_085_1781, w_085_1786, w_085_1788, w_085_1789, w_085_1790, w_085_1791, w_085_1792, w_085_1793, w_085_1798, w_085_1799, w_085_1800, w_085_1801, w_085_1808, w_085_1809, w_085_1810, w_085_1812, w_085_1813, w_085_1816, w_085_1817, w_085_1819, w_085_1824, w_085_1827, w_085_1828, w_085_1830, w_085_1831, w_085_1832, w_085_1833, w_085_1834, w_085_1836, w_085_1837, w_085_1840, w_085_1842, w_085_1843, w_085_1844, w_085_1845, w_085_1847, w_085_1849, w_085_1856, w_085_1858, w_085_1860, w_085_1861, w_085_1862, w_085_1863, w_085_1868, w_085_1869, w_085_1870, w_085_1871, w_085_1873, w_085_1876, w_085_1882, w_085_1883, w_085_1886, w_085_1887, w_085_1889, w_085_1890, w_085_1893, w_085_1896, w_085_1897, w_085_1898, w_085_1899, w_085_1901, w_085_1904, w_085_1907, w_085_1908, w_085_1909, w_085_1911, w_085_1914, w_085_1915, w_085_1917, w_085_1918, w_085_1919, w_085_1922, w_085_1924, w_085_1926, w_085_1931, w_085_1933, w_085_1937, w_085_1943, w_085_1947, w_085_1949, w_085_1951, w_085_1955, w_085_1956, w_085_1960, w_085_1963, w_085_1967, w_085_1968, w_085_1970, w_085_1973, w_085_1974, w_085_1977, w_085_1983, w_085_1987, w_085_1988, w_085_1989, w_085_1992, w_085_1993, w_085_1994, w_085_1995, w_085_1996, w_085_1997, w_085_1999, w_085_2001, w_085_2004, w_085_2005, w_085_2013, w_085_2014, w_085_2017, w_085_2018, w_085_2019, w_085_2026, w_085_2031, w_085_2032, w_085_2033, w_085_2034, w_085_2036, w_085_2038, w_085_2041, w_085_2043, w_085_2044, w_085_2045, w_085_2046, w_085_2047, w_085_2049, w_085_2051, w_085_2052, w_085_2054, w_085_2058, w_085_2059, w_085_2062, w_085_2065, w_085_2066, w_085_2068, w_085_2069, w_085_2075, w_085_2077, w_085_2079, w_085_2086, w_085_2088, w_085_2089, w_085_2090, w_085_2092, w_085_2096, w_085_2098, w_085_2099, w_085_2100, w_085_2104, w_085_2105, w_085_2106, w_085_2110, w_085_2111, w_085_2112, w_085_2119, w_085_2121, w_085_2122, w_085_2123, w_085_2125, w_085_2126, w_085_2131, w_085_2133, w_085_2134, w_085_2135, w_085_2136, w_085_2137, w_085_2143, w_085_2146, w_085_2150, w_085_2152, w_085_2153, w_085_2155, w_085_2156, w_085_2158, w_085_2162, w_085_2163, w_085_2166, w_085_2168, w_085_2170, w_085_2172, w_085_2173, w_085_2175, w_085_2176, w_085_2177, w_085_2178, w_085_2179, w_085_2180, w_085_2183, w_085_2185, w_085_2187, w_085_2188, w_085_2189, w_085_2190, w_085_2191, w_085_2194, w_085_2200, w_085_2201, w_085_2202, w_085_2204, w_085_2206, w_085_2209, w_085_2210, w_085_2213, w_085_2214, w_085_2215, w_085_2218, w_085_2220, w_085_2223, w_085_2226, w_085_2227, w_085_2228, w_085_2229, w_085_2235, w_085_2236, w_085_2239, w_085_2242, w_085_2246, w_085_2250, w_085_2251, w_085_2252, w_085_2253, w_085_2254, w_085_2255, w_085_2257, w_085_2259, w_085_2260, w_085_2262, w_085_2265, w_085_2266, w_085_2267, w_085_2268, w_085_2269, w_085_2271, w_085_2273, w_085_2274, w_085_2275, w_085_2280, w_085_2282, w_085_2284, w_085_2285, w_085_2286, w_085_2288, w_085_2289, w_085_2290, w_085_2291, w_085_2293, w_085_2295, w_085_2297, w_085_2298, w_085_2305, w_085_2306, w_085_2307, w_085_2309, w_085_2316, w_085_2321, w_085_2322, w_085_2324, w_085_2326, w_085_2328, w_085_2329, w_085_2332, w_085_2335, w_085_2338, w_085_2341, w_085_2343, w_085_2345, w_085_2347, w_085_2348, w_085_2349, w_085_2350, w_085_2351, w_085_2352, w_085_2355, w_085_2356, w_085_2360, w_085_2361, w_085_2364, w_085_2365, w_085_2366, w_085_2367, w_085_2374, w_085_2375, w_085_2377, w_085_2379, w_085_2380, w_085_2381, w_085_2383, w_085_2385, w_085_2388, w_085_2389, w_085_2390, w_085_2391, w_085_2393, w_085_2397, w_085_2398, w_085_2401, w_085_2403, w_085_2405, w_085_2407, w_085_2411, w_085_2412, w_085_2413, w_085_2415, w_085_2416, w_085_2418, w_085_2419, w_085_2420, w_085_2421, w_085_2423, w_085_2424, w_085_2435, w_085_2439, w_085_2441, w_085_2444, w_085_2445, w_085_2446, w_085_2447, w_085_2449, w_085_2450, w_085_2451, w_085_2454, w_085_2455, w_085_2457, w_085_2460, w_085_2461, w_085_2463, w_085_2464, w_085_2465, w_085_2466, w_085_2470, w_085_2471, w_085_2472, w_085_2473, w_085_2475, w_085_2476, w_085_2479, w_085_2485, w_085_2487, w_085_2490, w_085_2492, w_085_2493, w_085_2496, w_085_2499, w_085_2500, w_085_2501, w_085_2503, w_085_2504, w_085_2509, w_085_2510, w_085_2512, w_085_2513, w_085_2518, w_085_2520, w_085_2521, w_085_2522, w_085_2523, w_085_2533, w_085_2534, w_085_2535, w_085_2537, w_085_2538, w_085_2542, w_085_2543, w_085_2546, w_085_2548, w_085_2553, w_085_2554, w_085_2555, w_085_2556, w_085_2557, w_085_2558, w_085_2561, w_085_2563, w_085_2564, w_085_2567, w_085_2568, w_085_2570, w_085_2571, w_085_2573, w_085_2580, w_085_2583, w_085_2585, w_085_2590, w_085_2592, w_085_2594, w_085_2595, w_085_2597, w_085_2598, w_085_2599, w_085_2604, w_085_2605, w_085_2608, w_085_2612, w_085_2613, w_085_2614, w_085_2615, w_085_2619, w_085_2620, w_085_2621, w_085_2622, w_085_2625, w_085_2627, w_085_2631, w_085_2637, w_085_2638, w_085_2641, w_085_2644, w_085_2648, w_085_2649, w_085_2652, w_085_2654, w_085_2659, w_085_2660, w_085_2662, w_085_2666, w_085_2668, w_085_2670, w_085_2671, w_085_2672, w_085_2674, w_085_2676, w_085_2680, w_085_2681, w_085_2684, w_085_2686, w_085_2690, w_085_2691, w_085_2692, w_085_2693, w_085_2695, w_085_2698, w_085_2700, w_085_2702, w_085_2708, w_085_2709, w_085_2711, w_085_2714, w_085_2716, w_085_2717, w_085_2719, w_085_2721, w_085_2724, w_085_2728, w_085_2729, w_085_2731, w_085_2734, w_085_2736, w_085_2738, w_085_2739, w_085_2740, w_085_2742, w_085_2743, w_085_2745, w_085_2746, w_085_2747, w_085_2750, w_085_2753, w_085_2756, w_085_2759, w_085_2760, w_085_2761, w_085_2768, w_085_2772, w_085_2776, w_085_2778, w_085_2779, w_085_2783, w_085_2788, w_085_2789, w_085_2790, w_085_2794, w_085_2795, w_085_2796, w_085_2797, w_085_2799, w_085_2800, w_085_2801, w_085_2803, w_085_2805, w_085_2806, w_085_2809, w_085_2810, w_085_2814, w_085_2816, w_085_2821, w_085_2828, w_085_2833, w_085_2834, w_085_2835, w_085_2836, w_085_2837, w_085_2841, w_085_2848, w_085_2849, w_085_2850, w_085_2851, w_085_2852, w_085_2854, w_085_2855, w_085_2857, w_085_2859, w_085_2860, w_085_2862, w_085_2863, w_085_2864, w_085_2866, w_085_2869, w_085_2871, w_085_2876, w_085_2880, w_085_2883, w_085_2884, w_085_2885, w_085_2886, w_085_2890, w_085_2896, w_085_2898, w_085_2899, w_085_2901, w_085_2903, w_085_2909, w_085_2910, w_085_2911, w_085_2915, w_085_2916, w_085_2917, w_085_2919, w_085_2920, w_085_2921, w_085_2922, w_085_2923, w_085_2924, w_085_2926, w_085_2927, w_085_2931, w_085_2934, w_085_2935, w_085_2939, w_085_2942, w_085_2945, w_085_2948, w_085_2949, w_085_2952, w_085_2953, w_085_2954, w_085_2955, w_085_2957, w_085_2959, w_085_2961, w_085_2962, w_085_2963, w_085_2964, w_085_2967, w_085_2969, w_085_2973, w_085_2974, w_085_2975, w_085_2976, w_085_2977, w_085_2978, w_085_2979, w_085_2984, w_085_2986, w_085_2988, w_085_2989, w_085_2991, w_085_2993, w_085_2994, w_085_2996, w_085_3001, w_085_3004, w_085_3005, w_085_3008, w_085_3009, w_085_3014, w_085_3018, w_085_3023, w_085_3026, w_085_3029, w_085_3030, w_085_3031, w_085_3033, w_085_3034, w_085_3037, w_085_3045, w_085_3046, w_085_3047, w_085_3049, w_085_3050, w_085_3051, w_085_3052, w_085_3062, w_085_3064, w_085_3065, w_085_3069, w_085_3074, w_085_3075, w_085_3079, w_085_3082, w_085_3085, w_085_3086, w_085_3088, w_085_3090, w_085_3092, w_085_3093, w_085_3096, w_085_3097, w_085_3099, w_085_3101, w_085_3102, w_085_3106, w_085_3108, w_085_3111, w_085_3112, w_085_3113, w_085_3115, w_085_3117, w_085_3118, w_085_3120, w_085_3123, w_085_3124, w_085_3126, w_085_3127, w_085_3129, w_085_3133, w_085_3140, w_085_3143, w_085_3146, w_085_3147, w_085_3150, w_085_3151, w_085_3153, w_085_3154, w_085_3157, w_085_3158, w_085_3164, w_085_3168, w_085_3169, w_085_3178, w_085_3180, w_085_3183, w_085_3184, w_085_3186, w_085_3187, w_085_3189, w_085_3190, w_085_3192, w_085_3193, w_085_3196, w_085_3200, w_085_3201, w_085_3203, w_085_3212, w_085_3213, w_085_3214, w_085_3217, w_085_3220, w_085_3221, w_085_3222, w_085_3225, w_085_3226, w_085_3230, w_085_3232, w_085_3237, w_085_3240, w_085_3242, w_085_3243, w_085_3245, w_085_3246, w_085_3247, w_085_3249, w_085_3253, w_085_3255, w_085_3256, w_085_3258, w_085_3260, w_085_3261, w_085_3263, w_085_3264, w_085_3265, w_085_3269, w_085_3271, w_085_3273, w_085_3275, w_085_3279, w_085_3282, w_085_3283, w_085_3284, w_085_3288, w_085_3291, w_085_3295, w_085_3297, w_085_3300, w_085_3302, w_085_3303, w_085_3304, w_085_3305, w_085_3307, w_085_3311, w_085_3313, w_085_3318, w_085_3321, w_085_3323, w_085_3325, w_085_3327, w_085_3328, w_085_3329, w_085_3335, w_085_3336, w_085_3343, w_085_3344, w_085_3346, w_085_3347, w_085_3348, w_085_3349, w_085_3350, w_085_3354, w_085_3355, w_085_3359, w_085_3362, w_085_3363, w_085_3366, w_085_3367, w_085_3368, w_085_3369, w_085_3373, w_085_3374, w_085_3378, w_085_3380, w_085_3383, w_085_3384, w_085_3389, w_085_3393, w_085_3395, w_085_3400, w_085_3402, w_085_3403, w_085_3404, w_085_3405, w_085_3408, w_085_3409, w_085_3411, w_085_3412, w_085_3416, w_085_3418, w_085_3419, w_085_3420, w_085_3424, w_085_3425, w_085_3426, w_085_3427, w_085_3429, w_085_3430, w_085_3432, w_085_3433, w_085_3435, w_085_3439, w_085_3441, w_085_3442, w_085_3446, w_085_3447, w_085_3451, w_085_3453, w_085_3456, w_085_3457, w_085_3458, w_085_3459, w_085_3461, w_085_3462, w_085_3463, w_085_3465, w_085_3466, w_085_3472, w_085_3473, w_085_3474, w_085_3477, w_085_3483, w_085_3485, w_085_3487, w_085_3491, w_085_3494, w_085_3495, w_085_3497, w_085_3499, w_085_3500, w_085_3504, w_085_3505, w_085_3508, w_085_3510, w_085_3511, w_085_3512, w_085_3515, w_085_3517, w_085_3520, w_085_3522, w_085_3524, w_085_3526, w_085_3527, w_085_3531, w_085_3532, w_085_3535, w_085_3539, w_085_3544, w_085_3545, w_085_3546, w_085_3548, w_085_3549, w_085_3550, w_085_3551, w_085_3553, w_085_3556, w_085_3562, w_085_3564, w_085_3566, w_085_3567, w_085_3568, w_085_3576, w_085_3578, w_085_3582, w_085_3585, w_085_3588, w_085_3592, w_085_3593, w_085_3594, w_085_3595, w_085_3597, w_085_3598, w_085_3599, w_085_3600, w_085_3603, w_085_3604, w_085_3606, w_085_3607, w_085_3608, w_085_3611, w_085_3613, w_085_3614, w_085_3615, w_085_3616, w_085_3617, w_085_3618, w_085_3619, w_085_3623, w_085_3627, w_085_3628, w_085_3629, w_085_3630, w_085_3631, w_085_3632, w_085_3633, w_085_3634, w_085_3635, w_085_3636, w_085_3637, w_085_3645, w_085_3647, w_085_3650, w_085_3651, w_085_3655, w_085_3657, w_085_3658, w_085_3659, w_085_3661, w_085_3662, w_085_3664, w_085_3666, w_085_3667, w_085_3669, w_085_3672, w_085_3675, w_085_3683, w_085_3686, w_085_3690, w_085_3692, w_085_3693, w_085_3694, w_085_3701, w_085_3703, w_085_3706, w_085_3709, w_085_3710, w_085_3711, w_085_3714, w_085_3716, w_085_3718, w_085_3719, w_085_3720, w_085_3721, w_085_3724, w_085_3726, w_085_3729, w_085_3733, w_085_3739, w_085_3742, w_085_3745, w_085_3746, w_085_3747, w_085_3748, w_085_3749, w_085_3752, w_085_3756, w_085_3758, w_085_3760, w_085_3762, w_085_3763, w_085_3765, w_085_3766, w_085_3767, w_085_3768, w_085_3771, w_085_3774, w_085_3775, w_085_3778, w_085_3779, w_085_3781, w_085_3782, w_085_3783, w_085_3786, w_085_3789, w_085_3791, w_085_3792, w_085_3794, w_085_3796, w_085_3799, w_085_3801, w_085_3804, w_085_3807, w_085_3809, w_085_3810, w_085_3812, w_085_3815, w_085_3821, w_085_3827, w_085_3828, w_085_3829, w_085_3830, w_085_3835, w_085_3836, w_085_3839, w_085_3840, w_085_3841, w_085_3846, w_085_3847, w_085_3849, w_085_3850, w_085_3852, w_085_3853, w_085_3855, w_085_3856, w_085_3858, w_085_3859, w_085_3861, w_085_3864, w_085_3865, w_085_3866, w_085_3868, w_085_3869, w_085_3870, w_085_3872, w_085_3874, w_085_3876, w_085_3881, w_085_3883, w_085_3884, w_085_3885, w_085_3888, w_085_3889, w_085_3894, w_085_3895, w_085_3899, w_085_3900, w_085_3901, w_085_3902, w_085_3905, w_085_3906, w_085_3907, w_085_3909, w_085_3911, w_085_3913, w_085_3916, w_085_3918, w_085_3922, w_085_3924, w_085_3925, w_085_3929, w_085_3933, w_085_3939, w_085_3943, w_085_3944, w_085_3945, w_085_3947, w_085_3948, w_085_3949, w_085_3951, w_085_3952, w_085_3962, w_085_3965, w_085_3968, w_085_3972, w_085_3973, w_085_3978, w_085_3979, w_085_3980, w_085_3981, w_085_3983, w_085_3986, w_085_3991, w_085_3994, w_085_3995, w_085_3996, w_085_3997, w_085_3998, w_085_3999, w_085_4000, w_085_4001, w_085_4005, w_085_4008, w_085_4010, w_085_4011, w_085_4012, w_085_4013, w_085_4018, w_085_4019, w_085_4023, w_085_4029, w_085_4030, w_085_4031, w_085_4032, w_085_4035, w_085_4038, w_085_4039, w_085_4040, w_085_4043, w_085_4046, w_085_4048, w_085_4049, w_085_4050, w_085_4053, w_085_4054, w_085_4058, w_085_4059, w_085_4061, w_085_4062, w_085_4067, w_085_4068, w_085_4069, w_085_4071, w_085_4072, w_085_4074, w_085_4075, w_085_4079, w_085_4080, w_085_4081, w_085_4084, w_085_4087, w_085_4088, w_085_4089, w_085_4092, w_085_4093, w_085_4094, w_085_4095, w_085_4097, w_085_4098, w_085_4099, w_085_4101, w_085_4102, w_085_4105, w_085_4107, w_085_4110, w_085_4111, w_085_4114, w_085_4119, w_085_4120, w_085_4122, w_085_4124, w_085_4127, w_085_4128, w_085_4129, w_085_4130, w_085_4134, w_085_4138, w_085_4145, w_085_4146, w_085_4150, w_085_4152, w_085_4153, w_085_4154, w_085_4156, w_085_4162, w_085_4163, w_085_4164, w_085_4165, w_085_4167, w_085_4168, w_085_4170, w_085_4173, w_085_4174, w_085_4175, w_085_4177, w_085_4178, w_085_4180, w_085_4183, w_085_4185, w_085_4186, w_085_4189, w_085_4190, w_085_4191, w_085_4194, w_085_4195, w_085_4196, w_085_4202, w_085_4204, w_085_4205, w_085_4210, w_085_4211, w_085_4214, w_085_4215, w_085_4217, w_085_4219, w_085_4222, w_085_4223, w_085_4224, w_085_4225, w_085_4227, w_085_4228, w_085_4231, w_085_4232, w_085_4233, w_085_4234, w_085_4235, w_085_4236, w_085_4237, w_085_4242, w_085_4246, w_085_4250, w_085_4252, w_085_4256, w_085_4257, w_085_4258, w_085_4260, w_085_4263, w_085_4264, w_085_4266, w_085_4267, w_085_4268, w_085_4271, w_085_4273, w_085_4275, w_085_4276, w_085_4277, w_085_4278, w_085_4279, w_085_4281, w_085_4282, w_085_4286, w_085_4289, w_085_4290, w_085_4291, w_085_4292, w_085_4293, w_085_4294, w_085_4296, w_085_4299, w_085_4300, w_085_4303, w_085_4306, w_085_4307, w_085_4310, w_085_4314, w_085_4316, w_085_4317, w_085_4321, w_085_4328, w_085_4331, w_085_4334, w_085_4335, w_085_4337, w_085_4338, w_085_4342, w_085_4343, w_085_4344, w_085_4347, w_085_4350, w_085_4358, w_085_4359, w_085_4362, w_085_4364, w_085_4366, w_085_4371, w_085_4375, w_085_4376, w_085_4378, w_085_4379, w_085_4380, w_085_4381, w_085_4385, w_085_4389, w_085_4391, w_085_4393, w_085_4395, w_085_4398, w_085_4400, w_085_4402, w_085_4403, w_085_4404, w_085_4406, w_085_4408, w_085_4409, w_085_4410, w_085_4413, w_085_4414, w_085_4417, w_085_4426, w_085_4428, w_085_4429, w_085_4431, w_085_4432, w_085_4434, w_085_4436, w_085_4442, w_085_4445, w_085_4446, w_085_4447, w_085_4448, w_085_4449, w_085_4450, w_085_4452, w_085_4455, w_085_4456, w_085_4463, w_085_4464, w_085_4467, w_085_4468, w_085_4469, w_085_4470, w_085_4471, w_085_4476, w_085_4478, w_085_4479, w_085_4480, w_085_4481, w_085_4482, w_085_4483, w_085_4484, w_085_4487, w_085_4490, w_085_4491, w_085_4493, w_085_4495, w_085_4498, w_085_4500, w_085_4502, w_085_4503, w_085_4504, w_085_4506, w_085_4512, w_085_4513, w_085_4516, w_085_4521, w_085_4522, w_085_4523, w_085_4530, w_085_4531, w_085_4532, w_085_4538, w_085_4540, w_085_4543, w_085_4545, w_085_4546, w_085_4547, w_085_4549, w_085_4552, w_085_4553, w_085_4554, w_085_4556, w_085_4559, w_085_4560, w_085_4562, w_085_4564, w_085_4566, w_085_4567, w_085_4569, w_085_4570, w_085_4571, w_085_4572, w_085_4575, w_085_4579, w_085_4582, w_085_4586, w_085_4588, w_085_4589, w_085_4590, w_085_4591, w_085_4592, w_085_4595, w_085_4596, w_085_4599, w_085_4602, w_085_4606, w_085_4610, w_085_4614, w_085_4615, w_085_4616, w_085_4618, w_085_4619, w_085_4623, w_085_4628, w_085_4630, w_085_4632, w_085_4634, w_085_4636, w_085_4639, w_085_4641, w_085_4643, w_085_4645, w_085_4653, w_085_4654, w_085_4656, w_085_4658, w_085_4659, w_085_4663, w_085_4664, w_085_4665, w_085_4666, w_085_4668, w_085_4676, w_085_4677, w_085_4678, w_085_4680, w_085_4681, w_085_4685, w_085_4695, w_085_4696, w_085_4701, w_085_4704, w_085_4708, w_085_4712, w_085_4720, w_085_4722, w_085_4724, w_085_4738, w_085_4739, w_085_4744, w_085_4746, w_085_4760, w_085_4763, w_085_4768, w_085_4769, w_085_4782, w_085_4783, w_085_4787, w_085_4788, w_085_4789, w_085_4790, w_085_4792, w_085_4798, w_085_4800, w_085_4805, w_085_4809, w_085_4811, w_085_4813, w_085_4817, w_085_4818, w_085_4819, w_085_4825, w_085_4826, w_085_4828, w_085_4830, w_085_4833, w_085_4837, w_085_4847, w_085_4849, w_085_4855, w_085_4857, w_085_4865, w_085_4868, w_085_4869, w_085_4871, w_085_4872, w_085_4876, w_085_4878, w_085_4881, w_085_4889, w_085_4892, w_085_4893, w_085_4898, w_085_4900, w_085_4901, w_085_4906, w_085_4912, w_085_4918, w_085_4920, w_085_4922, w_085_4926, w_085_4927, w_085_4933, w_085_4934, w_085_4935, w_085_4936, w_085_4939, w_085_4944, w_085_4947, w_085_4948, w_085_4960, w_085_4970, w_085_4972, w_085_4973, w_085_4975, w_085_4976, w_085_4988, w_085_4989, w_085_4990, w_085_4993, w_085_4994, w_085_4999, w_085_5005, w_085_5006, w_085_5010, w_085_5020, w_085_5021, w_085_5026, w_085_5031, w_085_5033, w_085_5038, w_085_5039, w_085_5044, w_085_5046, w_085_5047, w_085_5051, w_085_5052, w_085_5054, w_085_5055, w_085_5058, w_085_5064, w_085_5065, w_085_5070, w_085_5076, w_085_5082, w_085_5086, w_085_5089, w_085_5093, w_085_5096, w_085_5098, w_085_5104, w_085_5107, w_085_5121, w_085_5128, w_085_5131, w_085_5132, w_085_5133, w_085_5137, w_085_5141, w_085_5143, w_085_5146, w_085_5149, w_085_5152, w_085_5153, w_085_5156, w_085_5181, w_085_5182, w_085_5185, w_085_5187, w_085_5188, w_085_5192, w_085_5197, w_085_5200, w_085_5206, w_085_5207, w_085_5208, w_085_5212, w_085_5216, w_085_5225, w_085_5231, w_085_5234, w_085_5240, w_085_5243, w_085_5247, w_085_5257, w_085_5260, w_085_5263, w_085_5265, w_085_5267, w_085_5269, w_085_5272, w_085_5278, w_085_5285, w_085_5286, w_085_5291, w_085_5303, w_085_5313;
  wire w_086_000, w_086_004, w_086_005, w_086_006, w_086_007, w_086_009, w_086_010, w_086_012, w_086_013, w_086_014, w_086_018, w_086_020, w_086_021, w_086_023, w_086_025, w_086_026, w_086_027, w_086_028, w_086_031, w_086_032, w_086_033, w_086_034, w_086_036, w_086_039, w_086_042, w_086_043, w_086_044, w_086_045, w_086_046, w_086_047, w_086_050, w_086_061, w_086_063, w_086_064, w_086_065, w_086_068, w_086_069, w_086_074, w_086_076, w_086_078, w_086_081, w_086_082, w_086_084, w_086_085, w_086_087, w_086_089, w_086_091, w_086_092, w_086_094, w_086_095, w_086_096, w_086_097, w_086_098, w_086_100, w_086_102, w_086_104, w_086_107, w_086_109, w_086_112, w_086_113, w_086_114, w_086_116, w_086_118, w_086_119, w_086_121, w_086_123, w_086_125, w_086_126, w_086_127, w_086_129, w_086_131, w_086_132, w_086_133, w_086_134, w_086_139, w_086_141, w_086_142, w_086_146, w_086_147, w_086_149, w_086_150, w_086_154, w_086_157, w_086_159, w_086_169, w_086_170, w_086_172, w_086_174, w_086_175, w_086_177, w_086_179, w_086_183, w_086_184, w_086_185, w_086_187, w_086_190, w_086_191, w_086_193, w_086_195, w_086_197, w_086_199, w_086_202, w_086_205, w_086_206, w_086_208, w_086_209, w_086_215, w_086_216, w_086_217, w_086_219, w_086_220, w_086_221, w_086_224, w_086_234, w_086_240, w_086_241, w_086_245, w_086_249, w_086_251, w_086_252, w_086_253, w_086_255, w_086_257, w_086_258, w_086_263, w_086_264, w_086_265, w_086_270, w_086_271, w_086_278, w_086_279, w_086_281, w_086_284, w_086_286, w_086_289, w_086_296, w_086_297, w_086_303, w_086_304, w_086_305, w_086_306, w_086_311, w_086_314, w_086_315, w_086_316, w_086_318, w_086_323, w_086_328, w_086_330, w_086_331, w_086_333, w_086_340, w_086_341, w_086_343, w_086_349, w_086_351, w_086_352, w_086_353, w_086_357, w_086_359, w_086_362, w_086_365, w_086_367, w_086_373, w_086_374, w_086_375, w_086_376, w_086_377, w_086_378, w_086_379, w_086_380, w_086_382, w_086_384, w_086_385, w_086_389, w_086_391, w_086_392, w_086_395, w_086_397, w_086_400, w_086_405, w_086_406, w_086_410, w_086_411, w_086_416, w_086_417, w_086_421, w_086_423, w_086_424, w_086_426, w_086_427, w_086_428, w_086_430, w_086_431, w_086_432, w_086_433, w_086_436, w_086_437, w_086_438, w_086_439, w_086_444, w_086_451, w_086_452, w_086_454, w_086_459, w_086_461, w_086_466, w_086_468, w_086_469, w_086_470, w_086_471, w_086_472, w_086_473, w_086_475, w_086_481, w_086_482, w_086_488, w_086_489, w_086_490, w_086_494, w_086_495, w_086_500, w_086_502, w_086_504, w_086_505, w_086_506, w_086_512, w_086_514, w_086_515, w_086_526, w_086_527, w_086_528, w_086_529, w_086_532, w_086_533, w_086_534, w_086_536, w_086_537, w_086_538, w_086_539, w_086_544, w_086_545, w_086_546, w_086_547, w_086_551, w_086_554, w_086_555, w_086_557, w_086_558, w_086_560, w_086_561, w_086_563, w_086_564, w_086_565, w_086_569, w_086_570, w_086_571, w_086_572, w_086_578, w_086_579, w_086_581, w_086_583, w_086_585, w_086_590, w_086_592, w_086_593, w_086_594, w_086_598, w_086_603, w_086_605, w_086_606, w_086_609, w_086_613, w_086_614, w_086_615, w_086_616, w_086_617, w_086_619, w_086_621, w_086_622, w_086_624, w_086_625, w_086_628, w_086_629, w_086_630, w_086_631, w_086_633, w_086_636, w_086_637, w_086_638, w_086_644, w_086_646, w_086_647, w_086_649, w_086_650, w_086_652, w_086_655, w_086_660, w_086_665, w_086_666, w_086_667, w_086_668, w_086_669, w_086_672, w_086_676, w_086_678, w_086_679, w_086_680, w_086_690, w_086_692, w_086_694, w_086_699, w_086_703, w_086_704, w_086_705, w_086_706, w_086_707, w_086_708, w_086_710, w_086_711, w_086_713, w_086_718, w_086_719, w_086_720, w_086_724, w_086_728, w_086_729, w_086_734, w_086_735, w_086_736, w_086_740, w_086_742, w_086_743, w_086_747, w_086_749, w_086_751, w_086_752, w_086_754, w_086_756, w_086_757, w_086_759, w_086_762, w_086_764, w_086_770, w_086_771, w_086_772, w_086_773, w_086_776, w_086_777, w_086_779, w_086_781, w_086_782, w_086_783, w_086_784, w_086_785, w_086_791, w_086_792, w_086_793, w_086_794, w_086_796, w_086_798, w_086_799, w_086_801, w_086_802, w_086_808, w_086_809, w_086_812, w_086_814, w_086_815, w_086_816, w_086_818, w_086_819, w_086_820, w_086_822, w_086_825, w_086_827, w_086_828, w_086_832, w_086_835, w_086_836, w_086_838, w_086_839, w_086_841, w_086_842, w_086_845, w_086_848, w_086_850, w_086_851, w_086_854, w_086_855, w_086_856, w_086_859, w_086_861, w_086_862, w_086_863, w_086_864, w_086_869, w_086_876, w_086_883, w_086_884, w_086_885, w_086_888, w_086_894, w_086_897, w_086_898, w_086_899, w_086_906, w_086_907, w_086_910, w_086_912, w_086_914, w_086_915, w_086_918, w_086_920, w_086_922, w_086_924, w_086_930, w_086_933, w_086_934, w_086_939, w_086_941, w_086_944, w_086_947, w_086_949, w_086_951, w_086_952, w_086_954, w_086_960, w_086_961, w_086_963, w_086_966, w_086_973, w_086_975, w_086_977, w_086_978, w_086_979, w_086_982, w_086_983, w_086_987, w_086_990, w_086_993, w_086_996, w_086_997, w_086_1001, w_086_1002, w_086_1003, w_086_1004, w_086_1007, w_086_1008, w_086_1014, w_086_1019, w_086_1020, w_086_1023, w_086_1024, w_086_1025, w_086_1028, w_086_1031, w_086_1036, w_086_1038, w_086_1040, w_086_1042, w_086_1045, w_086_1051, w_086_1052, w_086_1054, w_086_1059, w_086_1060, w_086_1064, w_086_1067, w_086_1069, w_086_1070, w_086_1071, w_086_1073, w_086_1074, w_086_1078, w_086_1079, w_086_1080, w_086_1081, w_086_1084, w_086_1086, w_086_1089, w_086_1095, w_086_1098, w_086_1102, w_086_1104, w_086_1106, w_086_1109, w_086_1110, w_086_1111, w_086_1115, w_086_1118, w_086_1119, w_086_1123, w_086_1125, w_086_1126, w_086_1128, w_086_1129, w_086_1131, w_086_1135, w_086_1136, w_086_1137, w_086_1139, w_086_1140, w_086_1141, w_086_1143, w_086_1146, w_086_1149, w_086_1150, w_086_1153, w_086_1154, w_086_1155, w_086_1158, w_086_1159, w_086_1160, w_086_1164, w_086_1167, w_086_1168, w_086_1170, w_086_1175, w_086_1177, w_086_1179, w_086_1183, w_086_1184, w_086_1185, w_086_1186, w_086_1187, w_086_1188, w_086_1190, w_086_1194, w_086_1195, w_086_1196, w_086_1199, w_086_1201, w_086_1203, w_086_1204, w_086_1206, w_086_1208, w_086_1214, w_086_1215, w_086_1217, w_086_1218, w_086_1220, w_086_1221, w_086_1222, w_086_1225, w_086_1226, w_086_1228, w_086_1229, w_086_1231, w_086_1233, w_086_1234, w_086_1238, w_086_1241, w_086_1243, w_086_1244, w_086_1248, w_086_1251, w_086_1256, w_086_1260, w_086_1261, w_086_1262, w_086_1263, w_086_1264, w_086_1265, w_086_1266, w_086_1267, w_086_1268, w_086_1272, w_086_1273, w_086_1275, w_086_1277, w_086_1280, w_086_1281, w_086_1283, w_086_1285, w_086_1293, w_086_1294, w_086_1295, w_086_1298, w_086_1300, w_086_1304, w_086_1306, w_086_1309, w_086_1312, w_086_1316, w_086_1317, w_086_1319, w_086_1322, w_086_1323, w_086_1329, w_086_1338, w_086_1339, w_086_1342, w_086_1345, w_086_1347, w_086_1348, w_086_1349, w_086_1350, w_086_1352, w_086_1353, w_086_1354, w_086_1362, w_086_1365, w_086_1368, w_086_1370, w_086_1371, w_086_1373, w_086_1378, w_086_1380, w_086_1383, w_086_1384, w_086_1385, w_086_1386, w_086_1387, w_086_1388, w_086_1390, w_086_1392, w_086_1393, w_086_1395, w_086_1397, w_086_1399, w_086_1400, w_086_1401, w_086_1402, w_086_1404, w_086_1406, w_086_1408, w_086_1409, w_086_1412, w_086_1413, w_086_1414, w_086_1415, w_086_1418, w_086_1419, w_086_1420, w_086_1421, w_086_1431, w_086_1434, w_086_1437, w_086_1438, w_086_1441, w_086_1443, w_086_1444, w_086_1449, w_086_1452, w_086_1453, w_086_1459, w_086_1462, w_086_1464, w_086_1465, w_086_1466, w_086_1467, w_086_1468, w_086_1470, w_086_1474, w_086_1475, w_086_1477, w_086_1479, w_086_1480, w_086_1481, w_086_1482, w_086_1484, w_086_1487, w_086_1489, w_086_1491, w_086_1494, w_086_1495, w_086_1496, w_086_1498, w_086_1500, w_086_1502, w_086_1503, w_086_1504, w_086_1505, w_086_1507, w_086_1511, w_086_1513, w_086_1514, w_086_1515, w_086_1516, w_086_1518, w_086_1523, w_086_1527, w_086_1528, w_086_1529, w_086_1534, w_086_1535, w_086_1538, w_086_1540, w_086_1541, w_086_1542, w_086_1543, w_086_1548, w_086_1551, w_086_1557, w_086_1558, w_086_1559, w_086_1562, w_086_1563, w_086_1567, w_086_1570, w_086_1571, w_086_1573, w_086_1574, w_086_1575, w_086_1576, w_086_1578, w_086_1579, w_086_1580, w_086_1581, w_086_1586, w_086_1588, w_086_1590, w_086_1591, w_086_1592, w_086_1595, w_086_1597, w_086_1598, w_086_1601, w_086_1602, w_086_1604, w_086_1606, w_086_1607, w_086_1609, w_086_1610, w_086_1612, w_086_1613, w_086_1622, w_086_1623, w_086_1625, w_086_1626, w_086_1630, w_086_1636, w_086_1638, w_086_1639, w_086_1640, w_086_1641, w_086_1643, w_086_1649, w_086_1651, w_086_1652, w_086_1654, w_086_1656, w_086_1659, w_086_1660, w_086_1663, w_086_1664, w_086_1671, w_086_1672, w_086_1673, w_086_1674, w_086_1676, w_086_1679, w_086_1682, w_086_1685, w_086_1686, w_086_1687, w_086_1688, w_086_1689, w_086_1690, w_086_1693, w_086_1694, w_086_1696, w_086_1699, w_086_1705, w_086_1706, w_086_1707, w_086_1711, w_086_1712, w_086_1715, w_086_1716, w_086_1718, w_086_1721, w_086_1722, w_086_1724, w_086_1728, w_086_1733, w_086_1734, w_086_1738, w_086_1739, w_086_1740, w_086_1741, w_086_1743, w_086_1744, w_086_1745, w_086_1746, w_086_1751, w_086_1752, w_086_1754, w_086_1755, w_086_1757, w_086_1758, w_086_1759, w_086_1760, w_086_1763, w_086_1764, w_086_1766, w_086_1767, w_086_1771, w_086_1772, w_086_1774, w_086_1775, w_086_1776, w_086_1778, w_086_1779, w_086_1780, w_086_1781, w_086_1783, w_086_1785, w_086_1790, w_086_1791, w_086_1794, w_086_1795, w_086_1797, w_086_1799, w_086_1800, w_086_1801, w_086_1802, w_086_1804, w_086_1809, w_086_1814, w_086_1816, w_086_1818, w_086_1824, w_086_1825, w_086_1827, w_086_1833, w_086_1834, w_086_1835, w_086_1836, w_086_1837, w_086_1838, w_086_1840, w_086_1843, w_086_1845, w_086_1846, w_086_1852, w_086_1853, w_086_1855, w_086_1856, w_086_1858, w_086_1859, w_086_1861, w_086_1863, w_086_1864, w_086_1868, w_086_1869, w_086_1872, w_086_1877, w_086_1878, w_086_1882, w_086_1884, w_086_1886, w_086_1887, w_086_1888, w_086_1891, w_086_1893, w_086_1895, w_086_1897, w_086_1898, w_086_1899, w_086_1903, w_086_1905, w_086_1906, w_086_1908, w_086_1912, w_086_1913, w_086_1914, w_086_1917, w_086_1919, w_086_1922, w_086_1924, w_086_1925, w_086_1928, w_086_1929, w_086_1932, w_086_1934, w_086_1938, w_086_1940, w_086_1943, w_086_1945, w_086_1948, w_086_1951, w_086_1952, w_086_1956, w_086_1957, w_086_1959, w_086_1960, w_086_1961, w_086_1970, w_086_1972, w_086_1974, w_086_1975, w_086_1979, w_086_1981, w_086_1982, w_086_1983, w_086_1984, w_086_1986, w_086_1987, w_086_1992, w_086_1993, w_086_1995, w_086_2001, w_086_2002, w_086_2006, w_086_2011, w_086_2012, w_086_2014, w_086_2017, w_086_2020, w_086_2021, w_086_2024, w_086_2027, w_086_2029, w_086_2031, w_086_2034, w_086_2035, w_086_2037, w_086_2043, w_086_2047, w_086_2048, w_086_2049, w_086_2051, w_086_2052, w_086_2053, w_086_2055, w_086_2058, w_086_2060, w_086_2063, w_086_2065, w_086_2067, w_086_2069, w_086_2071, w_086_2074, w_086_2076, w_086_2077, w_086_2082, w_086_2085, w_086_2087, w_086_2088, w_086_2091, w_086_2092, w_086_2093, w_086_2094, w_086_2096, w_086_2098, w_086_2099, w_086_2100, w_086_2102, w_086_2106, w_086_2109, w_086_2113, w_086_2116, w_086_2117, w_086_2120, w_086_2121, w_086_2122, w_086_2123, w_086_2124, w_086_2128, w_086_2130, w_086_2131, w_086_2136, w_086_2137, w_086_2139, w_086_2140, w_086_2143, w_086_2144, w_086_2147, w_086_2148, w_086_2149, w_086_2154, w_086_2157, w_086_2158, w_086_2159, w_086_2162, w_086_2163, w_086_2168, w_086_2170, w_086_2171, w_086_2174, w_086_2175, w_086_2178, w_086_2180, w_086_2181, w_086_2189, w_086_2195, w_086_2196, w_086_2197, w_086_2198, w_086_2199, w_086_2202, w_086_2204, w_086_2205, w_086_2206, w_086_2207, w_086_2208, w_086_2210, w_086_2213, w_086_2214, w_086_2215, w_086_2217, w_086_2224, w_086_2227, w_086_2228, w_086_2231, w_086_2232, w_086_2233, w_086_2236, w_086_2237, w_086_2246, w_086_2249, w_086_2251, w_086_2252, w_086_2253, w_086_2257, w_086_2260, w_086_2269, w_086_2270, w_086_2272, w_086_2273, w_086_2276, w_086_2281, w_086_2283, w_086_2287, w_086_2289, w_086_2290, w_086_2291, w_086_2292, w_086_2293, w_086_2295, w_086_2297, w_086_2304, w_086_2305, w_086_2307, w_086_2308, w_086_2310, w_086_2314, w_086_2318, w_086_2319, w_086_2320, w_086_2321, w_086_2323, w_086_2324, w_086_2325, w_086_2326, w_086_2327, w_086_2329, w_086_2330, w_086_2332, w_086_2334, w_086_2336, w_086_2337, w_086_2338, w_086_2339, w_086_2340, w_086_2341, w_086_2342, w_086_2343, w_086_2344, w_086_2346, w_086_2348, w_086_2351, w_086_2352, w_086_2355, w_086_2356, w_086_2358, w_086_2359, w_086_2362, w_086_2364, w_086_2365, w_086_2370, w_086_2373, w_086_2374, w_086_2375, w_086_2381, w_086_2382, w_086_2385, w_086_2392, w_086_2393, w_086_2397, w_086_2398, w_086_2399, w_086_2400, w_086_2401, w_086_2403, w_086_2404, w_086_2406, w_086_2410, w_086_2411, w_086_2412, w_086_2418, w_086_2423, w_086_2424, w_086_2428, w_086_2430, w_086_2431, w_086_2432, w_086_2433, w_086_2435, w_086_2438, w_086_2441, w_086_2444, w_086_2446, w_086_2447, w_086_2448, w_086_2449, w_086_2450, w_086_2451, w_086_2452, w_086_2454, w_086_2459, w_086_2464, w_086_2467, w_086_2468, w_086_2469, w_086_2472, w_086_2474, w_086_2475, w_086_2479, w_086_2480, w_086_2481, w_086_2485, w_086_2486, w_086_2487, w_086_2492, w_086_2493, w_086_2495, w_086_2497, w_086_2500, w_086_2506, w_086_2509, w_086_2511, w_086_2512, w_086_2514, w_086_2515, w_086_2516, w_086_2518, w_086_2520, w_086_2524, w_086_2528, w_086_2529, w_086_2530, w_086_2531, w_086_2533, w_086_2538, w_086_2539, w_086_2541, w_086_2542, w_086_2543, w_086_2544, w_086_2549, w_086_2550, w_086_2552, w_086_2553, w_086_2562, w_086_2564, w_086_2566, w_086_2567, w_086_2570, w_086_2573, w_086_2575, w_086_2577, w_086_2584, w_086_2585, w_086_2586, w_086_2588, w_086_2590, w_086_2591, w_086_2595, w_086_2596, w_086_2597, w_086_2598, w_086_2601, w_086_2602, w_086_2605, w_086_2607, w_086_2608, w_086_2609, w_086_2614, w_086_2616, w_086_2618, w_086_2619, w_086_2620, w_086_2621, w_086_2624, w_086_2625, w_086_2627, w_086_2629, w_086_2630, w_086_2633, w_086_2638, w_086_2639, w_086_2643, w_086_2644, w_086_2648, w_086_2651, w_086_2652, w_086_2655, w_086_2656, w_086_2657, w_086_2658, w_086_2659, w_086_2662, w_086_2668, w_086_2669, w_086_2670, w_086_2671, w_086_2672, w_086_2679, w_086_2680, w_086_2681, w_086_2682, w_086_2683, w_086_2687, w_086_2690, w_086_2693, w_086_2696, w_086_2698, w_086_2701, w_086_2702, w_086_2704, w_086_2705, w_086_2708, w_086_2713, w_086_2714, w_086_2718, w_086_2719, w_086_2722, w_086_2723, w_086_2724, w_086_2726, w_086_2729, w_086_2731, w_086_2732, w_086_2733, w_086_2734, w_086_2736, w_086_2742, w_086_2744, w_086_2745, w_086_2746, w_086_2749, w_086_2751, w_086_2754, w_086_2757, w_086_2761, w_086_2762, w_086_2765, w_086_2766, w_086_2767, w_086_2770, w_086_2772, w_086_2782, w_086_2784, w_086_2785, w_086_2788, w_086_2791, w_086_2792, w_086_2797, w_086_2798, w_086_2799, w_086_2801, w_086_2802, w_086_2803, w_086_2805, w_086_2806, w_086_2807, w_086_2808, w_086_2812, w_086_2813, w_086_2815, w_086_2817, w_086_2818, w_086_2821, w_086_2829, w_086_2835, w_086_2836, w_086_2837, w_086_2838, w_086_2842, w_086_2846, w_086_2847, w_086_2848, w_086_2851, w_086_2853, w_086_2854, w_086_2859, w_086_2862, w_086_2864, w_086_2869, w_086_2870, w_086_2876, w_086_2877, w_086_2883, w_086_2885, w_086_2886, w_086_2887, w_086_2888, w_086_2890, w_086_2891, w_086_2898, w_086_2899, w_086_2903, w_086_2904, w_086_2905, w_086_2906, w_086_2908, w_086_2920, w_086_2924, w_086_2925, w_086_2926, w_086_2928, w_086_2931, w_086_2936, w_086_2937, w_086_2938, w_086_2939, w_086_2941, w_086_2943, w_086_2945, w_086_2949, w_086_2952, w_086_2953, w_086_2956, w_086_2958, w_086_2961, w_086_2966, w_086_2969, w_086_2974, w_086_2977, w_086_2983, w_086_2988, w_086_2989, w_086_2991, w_086_2994, w_086_2995, w_086_2996, w_086_2998, w_086_3001, w_086_3003, w_086_3004, w_086_3017, w_086_3027, w_086_3029, w_086_3035, w_086_3040, w_086_3049, w_086_3055, w_086_3059, w_086_3060, w_086_3061, w_086_3062, w_086_3063, w_086_3064, w_086_3067, w_086_3070, w_086_3073, w_086_3076, w_086_3078, w_086_3084, w_086_3085, w_086_3086, w_086_3092, w_086_3094, w_086_3100, w_086_3104, w_086_3106, w_086_3109, w_086_3112, w_086_3120, w_086_3127, w_086_3129, w_086_3133, w_086_3137, w_086_3138, w_086_3139, w_086_3140, w_086_3145, w_086_3147, w_086_3148, w_086_3151, w_086_3152, w_086_3153, w_086_3159, w_086_3161, w_086_3164, w_086_3166, w_086_3167, w_086_3181, w_086_3186, w_086_3199, w_086_3200, w_086_3203, w_086_3205, w_086_3207, w_086_3208, w_086_3213, w_086_3221, w_086_3234, w_086_3236, w_086_3238, w_086_3259, w_086_3264, w_086_3266, w_086_3273, w_086_3274, w_086_3281, w_086_3285, w_086_3288, w_086_3299, w_086_3301, w_086_3311, w_086_3313, w_086_3315, w_086_3319, w_086_3321, w_086_3323, w_086_3324, w_086_3331, w_086_3333, w_086_3334, w_086_3343, w_086_3348, w_086_3349, w_086_3350, w_086_3358, w_086_3359, w_086_3360, w_086_3367, w_086_3370, w_086_3382, w_086_3390, w_086_3391, w_086_3393, w_086_3395, w_086_3405, w_086_3408, w_086_3409, w_086_3414, w_086_3426, w_086_3436, w_086_3439, w_086_3440, w_086_3442, w_086_3444, w_086_3446, w_086_3447, w_086_3450, w_086_3454, w_086_3457, w_086_3465, w_086_3466, w_086_3468, w_086_3479, w_086_3481, w_086_3502, w_086_3504, w_086_3510, w_086_3513, w_086_3516, w_086_3519, w_086_3520, w_086_3521, w_086_3527, w_086_3528, w_086_3530, w_086_3533, w_086_3535, w_086_3539, w_086_3542, w_086_3544, w_086_3545, w_086_3548, w_086_3549, w_086_3556, w_086_3558, w_086_3567, w_086_3576, w_086_3587, w_086_3588, w_086_3591, w_086_3597, w_086_3599, w_086_3601, w_086_3603, w_086_3607, w_086_3612, w_086_3617, w_086_3618, w_086_3626, w_086_3637, w_086_3638, w_086_3640, w_086_3643, w_086_3646, w_086_3648, w_086_3653, w_086_3661, w_086_3668, w_086_3670, w_086_3673, w_086_3677, w_086_3679, w_086_3680, w_086_3682, w_086_3683, w_086_3690, w_086_3693, w_086_3696, w_086_3698, w_086_3700, w_086_3707, w_086_3715, w_086_3716, w_086_3719, w_086_3721, w_086_3726, w_086_3729, w_086_3735, w_086_3736, w_086_3742, w_086_3743, w_086_3748, w_086_3755, w_086_3756, w_086_3757, w_086_3763, w_086_3764, w_086_3767, w_086_3769, w_086_3770, w_086_3772, w_086_3774, w_086_3776, w_086_3777, w_086_3782, w_086_3789, w_086_3794, w_086_3799, w_086_3802, w_086_3809, w_086_3812, w_086_3815, w_086_3823, w_086_3827, w_086_3833, w_086_3836, w_086_3839, w_086_3848, w_086_3851, w_086_3854, w_086_3856, w_086_3857, w_086_3859, w_086_3862, w_086_3880, w_086_3888, w_086_3889, w_086_3892, w_086_3896, w_086_3903, w_086_3906, w_086_3909, w_086_3910, w_086_3917, w_086_3922, w_086_3923, w_086_3926, w_086_3931, w_086_3933, w_086_3936, w_086_3942, w_086_3946, w_086_3947, w_086_3949, w_086_3954, w_086_3957, w_086_3962, w_086_3963, w_086_3966, w_086_3971, w_086_3973, w_086_3978, w_086_3980, w_086_3983, w_086_3985, w_086_3986, w_086_3987, w_086_3990, w_086_3994, w_086_3997, w_086_4010, w_086_4013, w_086_4022, w_086_4024, w_086_4031, w_086_4032, w_086_4035, w_086_4039, w_086_4042, w_086_4044, w_086_4047, w_086_4049, w_086_4050, w_086_4051, w_086_4062, w_086_4063, w_086_4064, w_086_4069, w_086_4070, w_086_4072, w_086_4089, w_086_4090, w_086_4093, w_086_4102, w_086_4105, w_086_4106, w_086_4107, w_086_4108, w_086_4115, w_086_4131, w_086_4133, w_086_4134, w_086_4146, w_086_4148, w_086_4151, w_086_4153, w_086_4161, w_086_4165, w_086_4188, w_086_4194, w_086_4198, w_086_4206, w_086_4214, w_086_4218, w_086_4224, w_086_4229, w_086_4231, w_086_4238, w_086_4240, w_086_4242, w_086_4244, w_086_4245, w_086_4247, w_086_4250, w_086_4253, w_086_4254, w_086_4255, w_086_4264, w_086_4265, w_086_4269, w_086_4272, w_086_4276, w_086_4305, w_086_4309, w_086_4313, w_086_4316, w_086_4331, w_086_4333, w_086_4337, w_086_4342, w_086_4346, w_086_4348, w_086_4353, w_086_4359, w_086_4362, w_086_4365, w_086_4366, w_086_4373, w_086_4375, w_086_4377, w_086_4381, w_086_4383, w_086_4384, w_086_4385, w_086_4390, w_086_4394, w_086_4397, w_086_4403, w_086_4407, w_086_4411, w_086_4415, w_086_4421, w_086_4425, w_086_4433, w_086_4438, w_086_4440, w_086_4441, w_086_4443, w_086_4445, w_086_4446, w_086_4450, w_086_4451, w_086_4453, w_086_4457, w_086_4463, w_086_4469, w_086_4474, w_086_4479, w_086_4482, w_086_4484, w_086_4485, w_086_4488, w_086_4493, w_086_4496, w_086_4503, w_086_4506, w_086_4508, w_086_4515, w_086_4517, w_086_4521, w_086_4527, w_086_4529, w_086_4530, w_086_4531, w_086_4534, w_086_4536, w_086_4555, w_086_4560, w_086_4561, w_086_4562, w_086_4572, w_086_4575, w_086_4577, w_086_4578, w_086_4587, w_086_4590, w_086_4591, w_086_4592, w_086_4594, w_086_4596, w_086_4598, w_086_4602, w_086_4604, w_086_4606, w_086_4609, w_086_4618, w_086_4620, w_086_4621, w_086_4623, w_086_4632, w_086_4637, w_086_4640, w_086_4642, w_086_4645, w_086_4647, w_086_4650, w_086_4651, w_086_4652, w_086_4654, w_086_4655, w_086_4662, w_086_4666, w_086_4669, w_086_4670, w_086_4680, w_086_4692, w_086_4697, w_086_4699, w_086_4700, w_086_4709, w_086_4711, w_086_4713, w_086_4714, w_086_4715, w_086_4721, w_086_4732, w_086_4737, w_086_4745, w_086_4746, w_086_4749, w_086_4752, w_086_4754, w_086_4759, w_086_4760, w_086_4765, w_086_4768, w_086_4769, w_086_4773, w_086_4778, w_086_4785, w_086_4798, w_086_4802, w_086_4804, w_086_4807, w_086_4815, w_086_4819, w_086_4823, w_086_4835, w_086_4841, w_086_4843, w_086_4844, w_086_4847, w_086_4855, w_086_4864, w_086_4873, w_086_4877, w_086_4891, w_086_4892, w_086_4893, w_086_4897, w_086_4899, w_086_4900, w_086_4905, w_086_4909, w_086_4914, w_086_4916, w_086_4918, w_086_4926, w_086_4932, w_086_4941, w_086_4947, w_086_4952, w_086_4955, w_086_4956, w_086_4957, w_086_4960, w_086_4970, w_086_4973, w_086_4981, w_086_4988, w_086_5008, w_086_5012, w_086_5013, w_086_5014, w_086_5017, w_086_5020, w_086_5026, w_086_5029, w_086_5037, w_086_5038, w_086_5039, w_086_5041, w_086_5046, w_086_5049, w_086_5050, w_086_5054, w_086_5057, w_086_5059, w_086_5064, w_086_5065, w_086_5066, w_086_5067, w_086_5072, w_086_5073, w_086_5080, w_086_5082, w_086_5090, w_086_5094, w_086_5096, w_086_5100, w_086_5108, w_086_5113, w_086_5115, w_086_5118, w_086_5126, w_086_5130, w_086_5135, w_086_5144, w_086_5146, w_086_5148, w_086_5151, w_086_5158, w_086_5162, w_086_5170, w_086_5173, w_086_5176, w_086_5177, w_086_5181, w_086_5185, w_086_5187, w_086_5188, w_086_5191, w_086_5192, w_086_5193, w_086_5196, w_086_5199, w_086_5201, w_086_5205, w_086_5206, w_086_5207, w_086_5210, w_086_5213, w_086_5218, w_086_5220, w_086_5222, w_086_5225, w_086_5228, w_086_5244, w_086_5251, w_086_5256, w_086_5261, w_086_5265, w_086_5267, w_086_5269, w_086_5271, w_086_5272, w_086_5274, w_086_5275, w_086_5281, w_086_5285, w_086_5289, w_086_5290, w_086_5292, w_086_5297, w_086_5301, w_086_5302, w_086_5305, w_086_5306, w_086_5307, w_086_5315, w_086_5329, w_086_5331, w_086_5333, w_086_5337, w_086_5338, w_086_5340, w_086_5345, w_086_5347, w_086_5348, w_086_5351, w_086_5352, w_086_5354, w_086_5356, w_086_5360, w_086_5362, w_086_5367, w_086_5370, w_086_5371, w_086_5377, w_086_5378, w_086_5386, w_086_5389, w_086_5390, w_086_5393, w_086_5398, w_086_5399, w_086_5400, w_086_5404, w_086_5415, w_086_5419, w_086_5421, w_086_5423, w_086_5427, w_086_5429, w_086_5430, w_086_5435, w_086_5436, w_086_5441, w_086_5442, w_086_5446, w_086_5447, w_086_5451, w_086_5457, w_086_5460, w_086_5469, w_086_5472, w_086_5480, w_086_5488, w_086_5490, w_086_5493, w_086_5498, w_086_5499, w_086_5500, w_086_5502, w_086_5503, w_086_5504, w_086_5507, w_086_5516, w_086_5517, w_086_5519, w_086_5520, w_086_5526, w_086_5527, w_086_5528, w_086_5533, w_086_5537, w_086_5538, w_086_5539, w_086_5540, w_086_5542, w_086_5544, w_086_5545, w_086_5555, w_086_5556, w_086_5559, w_086_5560, w_086_5564, w_086_5567, w_086_5574, w_086_5575, w_086_5578, w_086_5586, w_086_5589, w_086_5592, w_086_5596, w_086_5597, w_086_5611, w_086_5615, w_086_5616, w_086_5618, w_086_5624, w_086_5632, w_086_5639, w_086_5640, w_086_5647, w_086_5648, w_086_5652, w_086_5654, w_086_5656, w_086_5663, w_086_5678, w_086_5680, w_086_5681, w_086_5682, w_086_5685, w_086_5689, w_086_5694, w_086_5696, w_086_5699, w_086_5701, w_086_5705, w_086_5706, w_086_5709, w_086_5716, w_086_5718, w_086_5723, w_086_5733, w_086_5745, w_086_5749, w_086_5752, w_086_5755, w_086_5756, w_086_5757, w_086_5758, w_086_5760, w_086_5763, w_086_5765, w_086_5766, w_086_5768, w_086_5786, w_086_5791, w_086_5795, w_086_5799, w_086_5805, w_086_5807, w_086_5809, w_086_5812, w_086_5815, w_086_5818, w_086_5821, w_086_5825, w_086_5827, w_086_5828, w_086_5836, w_086_5838, w_086_5840, w_086_5841, w_086_5842, w_086_5843, w_086_5849, w_086_5850, w_086_5853, w_086_5856, w_086_5857, w_086_5860, w_086_5862, w_086_5863, w_086_5879, w_086_5884, w_086_5888, w_086_5896, w_086_5899, w_086_5904, w_086_5905, w_086_5909, w_086_5913, w_086_5915, w_086_5916, w_086_5917, w_086_5919, w_086_5920, w_086_5922, w_086_5925, w_086_5926, w_086_5928, w_086_5932, w_086_5935, w_086_5937, w_086_5939, w_086_5944, w_086_5946, w_086_5949, w_086_5951, w_086_5952, w_086_5958, w_086_5961, w_086_5962, w_086_5975, w_086_5978, w_086_5982, w_086_5993, w_086_5999, w_086_6000, w_086_6004, w_086_6006, w_086_6008, w_086_6013, w_086_6014, w_086_6019, w_086_6022, w_086_6023, w_086_6024, w_086_6025, w_086_6026, w_086_6036, w_086_6039, w_086_6044, w_086_6046, w_086_6051, w_086_6052, w_086_6053, w_086_6056, w_086_6059, w_086_6063, w_086_6066, w_086_6071, w_086_6072, w_086_6081, w_086_6082, w_086_6090, w_086_6094, w_086_6095, w_086_6099, w_086_6101, w_086_6103, w_086_6106, w_086_6107, w_086_6111, w_086_6117, w_086_6119, w_086_6121, w_086_6122, w_086_6129, w_086_6139, w_086_6143, w_086_6144, w_086_6146, w_086_6149, w_086_6152, w_086_6153, w_086_6155, w_086_6156, w_086_6157, w_086_6158, w_086_6163, w_086_6164, w_086_6167, w_086_6168, w_086_6170, w_086_6176, w_086_6178, w_086_6182, w_086_6184, w_086_6192, w_086_6196, w_086_6197, w_086_6199, w_086_6201, w_086_6207, w_086_6208, w_086_6210, w_086_6212, w_086_6214, w_086_6216, w_086_6223, w_086_6227, w_086_6229, w_086_6235, w_086_6237, w_086_6241, w_086_6242, w_086_6245, w_086_6247, w_086_6248, w_086_6256, w_086_6259, w_086_6261, w_086_6267, w_086_6272, w_086_6273, w_086_6274, w_086_6275, w_086_6284, w_086_6287, w_086_6297, w_086_6308, w_086_6313, w_086_6314, w_086_6316, w_086_6317, w_086_6319, w_086_6321, w_086_6323, w_086_6324, w_086_6334, w_086_6335, w_086_6339, w_086_6342, w_086_6343, w_086_6344, w_086_6347, w_086_6350, w_086_6351, w_086_6356, w_086_6362, w_086_6363, w_086_6386, w_086_6387, w_086_6389, w_086_6390, w_086_6393, w_086_6404, w_086_6417, w_086_6419, w_086_6422, w_086_6424, w_086_6426, w_086_6427, w_086_6434, w_086_6436, w_086_6441, w_086_6443, w_086_6448, w_086_6453, w_086_6455, w_086_6457, w_086_6459, w_086_6461, w_086_6466, w_086_6473, w_086_6477, w_086_6478, w_086_6483, w_086_6485, w_086_6493, w_086_6496, w_086_6499, w_086_6504, w_086_6511, w_086_6512, w_086_6514, w_086_6517, w_086_6520, w_086_6521, w_086_6525, w_086_6526, w_086_6534, w_086_6538, w_086_6539, w_086_6541, w_086_6542, w_086_6543, w_086_6549, w_086_6558, w_086_6568, w_086_6569, w_086_6574, w_086_6575, w_086_6580, w_086_6582, w_086_6587, w_086_6589, w_086_6591, w_086_6592, w_086_6594, w_086_6602, w_086_6616, w_086_6624, w_086_6628, w_086_6629, w_086_6631, w_086_6640, w_086_6646, w_086_6648, w_086_6652, w_086_6656, w_086_6663, w_086_6664, w_086_6669, w_086_6673, w_086_6676, w_086_6685, w_086_6697, w_086_6703, w_086_6705, w_086_6708, w_086_6711, w_086_6713, w_086_6717, w_086_6718, w_086_6724, w_086_6727, w_086_6729, w_086_6730, w_086_6733, w_086_6744, w_086_6749, w_086_6751, w_086_6754, w_086_6757, w_086_6764, w_086_6768, w_086_6771, w_086_6774, w_086_6780, w_086_6782, w_086_6784, w_086_6785, w_086_6789, w_086_6792, w_086_6806, w_086_6808, w_086_6814, w_086_6817, w_086_6821, w_086_6825, w_086_6830, w_086_6835, w_086_6846, w_086_6848, w_086_6850, w_086_6866, w_086_6867, w_086_6872, w_086_6874, w_086_6880, w_086_6881, w_086_6882, w_086_6883, w_086_6884, w_086_6888, w_086_6889, w_086_6892, w_086_6903, w_086_6914, w_086_6923, w_086_6930, w_086_6935, w_086_6936, w_086_6938, w_086_6940, w_086_6944, w_086_6945, w_086_6948, w_086_6951, w_086_6952, w_086_6953, w_086_6957, w_086_6959, w_086_6963, w_086_6970, w_086_6973, w_086_6976, w_086_6978, w_086_6980, w_086_6982, w_086_6990, w_086_6996, w_086_6999, w_086_7002;
  wire w_087_004, w_087_005, w_087_008, w_087_009, w_087_011, w_087_012, w_087_013, w_087_016, w_087_017, w_087_018, w_087_020, w_087_021, w_087_024, w_087_029, w_087_031, w_087_036, w_087_037, w_087_042, w_087_043, w_087_044, w_087_045, w_087_046, w_087_049, w_087_050, w_087_051, w_087_052, w_087_053, w_087_055, w_087_061, w_087_066, w_087_067, w_087_070, w_087_073, w_087_074, w_087_075, w_087_079, w_087_081, w_087_082, w_087_084, w_087_085, w_087_086, w_087_087, w_087_089, w_087_090, w_087_092, w_087_096, w_087_098, w_087_099, w_087_101, w_087_103, w_087_106, w_087_107, w_087_108, w_087_110, w_087_112, w_087_113, w_087_114, w_087_117, w_087_118, w_087_119, w_087_121, w_087_122, w_087_123, w_087_124, w_087_125, w_087_126, w_087_127, w_087_129, w_087_132, w_087_134, w_087_136, w_087_137, w_087_139, w_087_140, w_087_141, w_087_142, w_087_143, w_087_145, w_087_146, w_087_149, w_087_151, w_087_153, w_087_156, w_087_160, w_087_161, w_087_162, w_087_163, w_087_166, w_087_169, w_087_171, w_087_172, w_087_173, w_087_176, w_087_177, w_087_179, w_087_185, w_087_187, w_087_188, w_087_191, w_087_192, w_087_193, w_087_194, w_087_195, w_087_201, w_087_202, w_087_205, w_087_206, w_087_207, w_087_209, w_087_218, w_087_220, w_087_222, w_087_226, w_087_227, w_087_228, w_087_229, w_087_230, w_087_231, w_087_232, w_087_233, w_087_235, w_087_236, w_087_237, w_087_245, w_087_246, w_087_247, w_087_249, w_087_251, w_087_252, w_087_258, w_087_259, w_087_260, w_087_264, w_087_267, w_087_268, w_087_269, w_087_270, w_087_271, w_087_272, w_087_275, w_087_276, w_087_277, w_087_278, w_087_279, w_087_283, w_087_286, w_087_289, w_087_290, w_087_292, w_087_296, w_087_297, w_087_298, w_087_299, w_087_301, w_087_305, w_087_306, w_087_307, w_087_308, w_087_309, w_087_310, w_087_311, w_087_312, w_087_314, w_087_317, w_087_319, w_087_324, w_087_325, w_087_326, w_087_328, w_087_329, w_087_332, w_087_333, w_087_339, w_087_340, w_087_346, w_087_350, w_087_352, w_087_355, w_087_358, w_087_359, w_087_362, w_087_366, w_087_367, w_087_369, w_087_370, w_087_373, w_087_374, w_087_376, w_087_378, w_087_382, w_087_388, w_087_391, w_087_392, w_087_401, w_087_403, w_087_406, w_087_411, w_087_412, w_087_413, w_087_417, w_087_420, w_087_422, w_087_424, w_087_429, w_087_430, w_087_432, w_087_433, w_087_437, w_087_438, w_087_439, w_087_440, w_087_443, w_087_444, w_087_445, w_087_447, w_087_449, w_087_450, w_087_452, w_087_454, w_087_457, w_087_458, w_087_460, w_087_463, w_087_466, w_087_467, w_087_468, w_087_469, w_087_470, w_087_472, w_087_473, w_087_474, w_087_476, w_087_478, w_087_482, w_087_487, w_087_488, w_087_489, w_087_490, w_087_492, w_087_495, w_087_497, w_087_502, w_087_503, w_087_504, w_087_505, w_087_507, w_087_508, w_087_509, w_087_510, w_087_512, w_087_515, w_087_516, w_087_517, w_087_518, w_087_521, w_087_523, w_087_525, w_087_526, w_087_528, w_087_535, w_087_536, w_087_540, w_087_541, w_087_542, w_087_545, w_087_546, w_087_547, w_087_548, w_087_550, w_087_552, w_087_556, w_087_558, w_087_562, w_087_563, w_087_566, w_087_568, w_087_569, w_087_570, w_087_575, w_087_576, w_087_577, w_087_580, w_087_581, w_087_586, w_087_587, w_087_589, w_087_593, w_087_594, w_087_597, w_087_598, w_087_601, w_087_605, w_087_606, w_087_608, w_087_609, w_087_611, w_087_614, w_087_616, w_087_618, w_087_619, w_087_621, w_087_624, w_087_626, w_087_627, w_087_628, w_087_629, w_087_631, w_087_634, w_087_635, w_087_637, w_087_639, w_087_641, w_087_644, w_087_646, w_087_648, w_087_649, w_087_650, w_087_653, w_087_654, w_087_658, w_087_659, w_087_661, w_087_662, w_087_665, w_087_666, w_087_667, w_087_671, w_087_674, w_087_677, w_087_678, w_087_680, w_087_681, w_087_685, w_087_688, w_087_689, w_087_691, w_087_695, w_087_696, w_087_697, w_087_698, w_087_699, w_087_700, w_087_704, w_087_705, w_087_707, w_087_708, w_087_709, w_087_711, w_087_716, w_087_717, w_087_719, w_087_721, w_087_723, w_087_724, w_087_726, w_087_727, w_087_729, w_087_737, w_087_738, w_087_743, w_087_744, w_087_745, w_087_752, w_087_754, w_087_759, w_087_760, w_087_761, w_087_762, w_087_763, w_087_765, w_087_768, w_087_769, w_087_771, w_087_774, w_087_775, w_087_778, w_087_781, w_087_782, w_087_783, w_087_785, w_087_787, w_087_788, w_087_789, w_087_790, w_087_793, w_087_795, w_087_797, w_087_804, w_087_807, w_087_812, w_087_815, w_087_820, w_087_822, w_087_824, w_087_825, w_087_826, w_087_827, w_087_829, w_087_832, w_087_834, w_087_835, w_087_839, w_087_841, w_087_842, w_087_845, w_087_846, w_087_848, w_087_849, w_087_854, w_087_859, w_087_861, w_087_863, w_087_864, w_087_868, w_087_870, w_087_873, w_087_875, w_087_876, w_087_881, w_087_884, w_087_887, w_087_891, w_087_892, w_087_893, w_087_896, w_087_901, w_087_908, w_087_911, w_087_912, w_087_913, w_087_915, w_087_917, w_087_918, w_087_920, w_087_921, w_087_924, w_087_926, w_087_929, w_087_932, w_087_935, w_087_939, w_087_941, w_087_946, w_087_949, w_087_950, w_087_955, w_087_960, w_087_962, w_087_969, w_087_970, w_087_972, w_087_973, w_087_974, w_087_980, w_087_983, w_087_986, w_087_991, w_087_994, w_087_996, w_087_997, w_087_1003, w_087_1007, w_087_1009, w_087_1010, w_087_1013, w_087_1015, w_087_1017, w_087_1018, w_087_1020, w_087_1023, w_087_1029, w_087_1030, w_087_1033, w_087_1034, w_087_1035, w_087_1036, w_087_1039, w_087_1040, w_087_1043, w_087_1044, w_087_1045, w_087_1048, w_087_1049, w_087_1050, w_087_1053, w_087_1056, w_087_1057, w_087_1058, w_087_1060, w_087_1061, w_087_1063, w_087_1064, w_087_1065, w_087_1066, w_087_1069, w_087_1070, w_087_1071, w_087_1074, w_087_1077, w_087_1078, w_087_1080, w_087_1081, w_087_1083, w_087_1087, w_087_1089, w_087_1090, w_087_1091, w_087_1093, w_087_1097, w_087_1098, w_087_1099, w_087_1107, w_087_1116, w_087_1117, w_087_1123, w_087_1124, w_087_1126, w_087_1127, w_087_1130, w_087_1132, w_087_1134, w_087_1136, w_087_1139, w_087_1141, w_087_1142, w_087_1143, w_087_1145, w_087_1146, w_087_1150, w_087_1154, w_087_1157, w_087_1159, w_087_1160, w_087_1161, w_087_1164, w_087_1165, w_087_1168, w_087_1170, w_087_1171, w_087_1172, w_087_1174, w_087_1178, w_087_1181, w_087_1186, w_087_1187, w_087_1188, w_087_1189, w_087_1191, w_087_1193, w_087_1195, w_087_1197, w_087_1198, w_087_1200, w_087_1207, w_087_1209, w_087_1210, w_087_1211, w_087_1217, w_087_1223, w_087_1226, w_087_1230, w_087_1232, w_087_1233, w_087_1234, w_087_1236, w_087_1238, w_087_1239, w_087_1243, w_087_1251, w_087_1252, w_087_1254, w_087_1256, w_087_1257, w_087_1261, w_087_1262, w_087_1263, w_087_1264, w_087_1265, w_087_1267, w_087_1269, w_087_1270, w_087_1271, w_087_1272, w_087_1279, w_087_1280, w_087_1286, w_087_1293, w_087_1295, w_087_1296, w_087_1298, w_087_1302, w_087_1303, w_087_1307, w_087_1308, w_087_1316, w_087_1320, w_087_1321, w_087_1322, w_087_1323, w_087_1327, w_087_1335, w_087_1336, w_087_1339, w_087_1341, w_087_1343, w_087_1346, w_087_1347, w_087_1349, w_087_1351, w_087_1356, w_087_1357, w_087_1358, w_087_1361, w_087_1363, w_087_1366, w_087_1370, w_087_1371, w_087_1373, w_087_1378, w_087_1379, w_087_1380, w_087_1381, w_087_1382, w_087_1384, w_087_1385, w_087_1390, w_087_1394, w_087_1400, w_087_1402, w_087_1403, w_087_1405, w_087_1407, w_087_1408, w_087_1412, w_087_1413, w_087_1416, w_087_1417, w_087_1418, w_087_1419, w_087_1421, w_087_1428, w_087_1431, w_087_1433, w_087_1434, w_087_1435, w_087_1436, w_087_1437, w_087_1441, w_087_1442, w_087_1443, w_087_1444, w_087_1447, w_087_1448, w_087_1454, w_087_1455, w_087_1458, w_087_1459, w_087_1460, w_087_1461, w_087_1464, w_087_1465, w_087_1466, w_087_1467, w_087_1469, w_087_1470, w_087_1474, w_087_1477, w_087_1482, w_087_1484, w_087_1485, w_087_1488, w_087_1490, w_087_1491, w_087_1494, w_087_1503, w_087_1505, w_087_1511, w_087_1512, w_087_1519, w_087_1522, w_087_1524, w_087_1526, w_087_1528, w_087_1529, w_087_1531, w_087_1532, w_087_1534, w_087_1535, w_087_1536, w_087_1537, w_087_1538, w_087_1541, w_087_1544, w_087_1547, w_087_1550, w_087_1551, w_087_1552, w_087_1553, w_087_1557, w_087_1558, w_087_1559, w_087_1561, w_087_1569, w_087_1571, w_087_1572, w_087_1573, w_087_1577, w_087_1578, w_087_1579, w_087_1582, w_087_1583, w_087_1584, w_087_1586, w_087_1588, w_087_1590, w_087_1591, w_087_1593, w_087_1594, w_087_1600, w_087_1605, w_087_1606, w_087_1609, w_087_1612, w_087_1616, w_087_1617, w_087_1619, w_087_1621, w_087_1624, w_087_1625, w_087_1630, w_087_1631, w_087_1632, w_087_1638, w_087_1639, w_087_1642, w_087_1645, w_087_1646, w_087_1648, w_087_1651, w_087_1653, w_087_1654, w_087_1656, w_087_1658, w_087_1659, w_087_1662, w_087_1663, w_087_1664, w_087_1668, w_087_1672, w_087_1675, w_087_1677, w_087_1679, w_087_1681, w_087_1682, w_087_1685, w_087_1687, w_087_1688, w_087_1690, w_087_1694, w_087_1695, w_087_1696, w_087_1697, w_087_1698, w_087_1702, w_087_1709, w_087_1710, w_087_1714, w_087_1716, w_087_1717, w_087_1718, w_087_1719, w_087_1720, w_087_1722, w_087_1723, w_087_1725, w_087_1728, w_087_1730, w_087_1731, w_087_1734, w_087_1736, w_087_1737, w_087_1739, w_087_1742, w_087_1743, w_087_1745, w_087_1750, w_087_1752, w_087_1755, w_087_1756, w_087_1760, w_087_1762, w_087_1763, w_087_1764, w_087_1765, w_087_1766, w_087_1768, w_087_1769, w_087_1771, w_087_1772, w_087_1773, w_087_1774, w_087_1775, w_087_1778, w_087_1780, w_087_1781, w_087_1785, w_087_1790, w_087_1792, w_087_1794, w_087_1795, w_087_1804, w_087_1807, w_087_1808, w_087_1810, w_087_1811, w_087_1812, w_087_1813, w_087_1814, w_087_1815, w_087_1816, w_087_1819, w_087_1820, w_087_1822, w_087_1824, w_087_1827, w_087_1829, w_087_1832, w_087_1833, w_087_1834, w_087_1835, w_087_1837, w_087_1841, w_087_1843, w_087_1846, w_087_1852, w_087_1853, w_087_1854, w_087_1856, w_087_1857, w_087_1861, w_087_1862, w_087_1865, w_087_1866, w_087_1867, w_087_1871, w_087_1872, w_087_1873, w_087_1879, w_087_1881, w_087_1884, w_087_1885, w_087_1886, w_087_1888, w_087_1891, w_087_1892, w_087_1898, w_087_1900, w_087_1901, w_087_1904, w_087_1906, w_087_1913, w_087_1915, w_087_1917, w_087_1921, w_087_1923, w_087_1924, w_087_1925, w_087_1927, w_087_1928, w_087_1937, w_087_1942, w_087_1943, w_087_1944, w_087_1949, w_087_1951, w_087_1952, w_087_1955, w_087_1956, w_087_1957, w_087_1959, w_087_1961, w_087_1966, w_087_1967, w_087_1968, w_087_1969, w_087_1971, w_087_1972, w_087_1977, w_087_1984, w_087_1985, w_087_1988, w_087_1990, w_087_1995, w_087_1996, w_087_1998, w_087_1999, w_087_2002, w_087_2003, w_087_2005, w_087_2006, w_087_2008, w_087_2009, w_087_2011, w_087_2012, w_087_2013, w_087_2015, w_087_2016, w_087_2017, w_087_2018, w_087_2023, w_087_2025, w_087_2028, w_087_2031, w_087_2032, w_087_2037, w_087_2038, w_087_2041, w_087_2042, w_087_2043, w_087_2051, w_087_2055, w_087_2059, w_087_2067, w_087_2068, w_087_2069, w_087_2070, w_087_2071, w_087_2073, w_087_2080, w_087_2085, w_087_2086, w_087_2087, w_087_2090, w_087_2092, w_087_2093, w_087_2094, w_087_2099, w_087_2100, w_087_2101, w_087_2102, w_087_2105, w_087_2108, w_087_2112, w_087_2113, w_087_2114, w_087_2116, w_087_2118, w_087_2119, w_087_2120, w_087_2122, w_087_2123, w_087_2126, w_087_2127, w_087_2128, w_087_2130, w_087_2131, w_087_2133, w_087_2135, w_087_2136, w_087_2137, w_087_2142, w_087_2145, w_087_2146, w_087_2147, w_087_2150, w_087_2151, w_087_2152, w_087_2159, w_087_2160, w_087_2163, w_087_2164, w_087_2165, w_087_2167, w_087_2178, w_087_2180, w_087_2181, w_087_2185, w_087_2186, w_087_2193, w_087_2202, w_087_2204, w_087_2206, w_087_2207, w_087_2209, w_087_2212, w_087_2213, w_087_2215, w_087_2216, w_087_2217, w_087_2218, w_087_2219, w_087_2222, w_087_2223, w_087_2226, w_087_2231, w_087_2233, w_087_2237, w_087_2238, w_087_2239, w_087_2240, w_087_2244, w_087_2245, w_087_2247, w_087_2251, w_087_2252, w_087_2253, w_087_2255, w_087_2257, w_087_2258, w_087_2260, w_087_2261, w_087_2262, w_087_2265, w_087_2267, w_087_2269, w_087_2270, w_087_2272, w_087_2273, w_087_2279, w_087_2281, w_087_2282, w_087_2284, w_087_2285, w_087_2286, w_087_2288, w_087_2290, w_087_2294, w_087_2300, w_087_2302, w_087_2303, w_087_2304, w_087_2307, w_087_2308, w_087_2309, w_087_2311, w_087_2313, w_087_2316, w_087_2317, w_087_2318, w_087_2319, w_087_2320, w_087_2321, w_087_2323, w_087_2325, w_087_2326, w_087_2327, w_087_2330, w_087_2331, w_087_2332, w_087_2333, w_087_2339, w_087_2346, w_087_2347, w_087_2349, w_087_2351, w_087_2353, w_087_2354, w_087_2356, w_087_2357, w_087_2358, w_087_2359, w_087_2360, w_087_2362, w_087_2364, w_087_2366, w_087_2367, w_087_2368, w_087_2370, w_087_2371, w_087_2373, w_087_2376, w_087_2379, w_087_2380, w_087_2381, w_087_2384, w_087_2386, w_087_2389, w_087_2390, w_087_2391, w_087_2392, w_087_2396, w_087_2400, w_087_2402, w_087_2404, w_087_2406, w_087_2407, w_087_2408, w_087_2412, w_087_2418, w_087_2420, w_087_2424, w_087_2428, w_087_2429, w_087_2433, w_087_2434, w_087_2435, w_087_2436, w_087_2437, w_087_2438, w_087_2439, w_087_2445, w_087_2446, w_087_2451, w_087_2453, w_087_2454, w_087_2455, w_087_2456, w_087_2458, w_087_2461, w_087_2464, w_087_2468, w_087_2469, w_087_2473, w_087_2475, w_087_2477, w_087_2480, w_087_2481, w_087_2482, w_087_2483, w_087_2484, w_087_2485, w_087_2487, w_087_2495, w_087_2502, w_087_2503, w_087_2505, w_087_2506, w_087_2508, w_087_2512, w_087_2513, w_087_2516, w_087_2518, w_087_2519, w_087_2520, w_087_2521, w_087_2522, w_087_2523, w_087_2524, w_087_2527, w_087_2528, w_087_2530, w_087_2531, w_087_2532, w_087_2533, w_087_2537, w_087_2538, w_087_2541, w_087_2543, w_087_2544, w_087_2545, w_087_2547, w_087_2548, w_087_2550, w_087_2552, w_087_2553, w_087_2559, w_087_2560, w_087_2561, w_087_2563, w_087_2567, w_087_2571, w_087_2573, w_087_2574, w_087_2576, w_087_2578, w_087_2579, w_087_2586, w_087_2588, w_087_2589, w_087_2590, w_087_2593, w_087_2595, w_087_2596, w_087_2598, w_087_2600, w_087_2601, w_087_2602, w_087_2603, w_087_2604, w_087_2605, w_087_2608, w_087_2609, w_087_2610, w_087_2612, w_087_2614, w_087_2619, w_087_2623, w_087_2625, w_087_2626, w_087_2639, w_087_2640, w_087_2641, w_087_2642, w_087_2644, w_087_2648, w_087_2650, w_087_2653, w_087_2659, w_087_2662, w_087_2665, w_087_2666, w_087_2668, w_087_2670, w_087_2671, w_087_2673, w_087_2675, w_087_2679, w_087_2680, w_087_2684, w_087_2686, w_087_2688, w_087_2689, w_087_2691, w_087_2695, w_087_2696, w_087_2700, w_087_2701, w_087_2705, w_087_2706, w_087_2710, w_087_2713, w_087_2714, w_087_2718, w_087_2722, w_087_2723, w_087_2726, w_087_2730, w_087_2736, w_087_2737, w_087_2746, w_087_2747, w_087_2748, w_087_2751, w_087_2752, w_087_2757, w_087_2758, w_087_2759, w_087_2760, w_087_2763, w_087_2769, w_087_2770, w_087_2775, w_087_2780, w_087_2783, w_087_2784, w_087_2785, w_087_2786, w_087_2789, w_087_2793, w_087_2794, w_087_2795, w_087_2797, w_087_2803, w_087_2809, w_087_2811, w_087_2818, w_087_2821, w_087_2824, w_087_2825, w_087_2827, w_087_2828, w_087_2830, w_087_2835, w_087_2836, w_087_2843, w_087_2845, w_087_2846, w_087_2848, w_087_2849, w_087_2851, w_087_2853, w_087_2854, w_087_2855, w_087_2856, w_087_2857, w_087_2860, w_087_2862, w_087_2863, w_087_2864, w_087_2865, w_087_2869, w_087_2870, w_087_2872, w_087_2875, w_087_2877, w_087_2881, w_087_2883, w_087_2884, w_087_2885, w_087_2886, w_087_2892, w_087_2893, w_087_2895, w_087_2896, w_087_2897, w_087_2898, w_087_2900, w_087_2903, w_087_2908, w_087_2912, w_087_2914, w_087_2917, w_087_2920, w_087_2921, w_087_2923, w_087_2924, w_087_2925, w_087_2928, w_087_2929, w_087_2931, w_087_2932, w_087_2933, w_087_2935, w_087_2936, w_087_2938, w_087_2941, w_087_2942, w_087_2943, w_087_2944, w_087_2945, w_087_2946, w_087_2949, w_087_2950, w_087_2951, w_087_2952, w_087_2953, w_087_2955, w_087_2957, w_087_2960, w_087_2961, w_087_2965, w_087_2967, w_087_2968, w_087_2969, w_087_2976, w_087_2978, w_087_2979, w_087_2980, w_087_2981, w_087_2982, w_087_2985, w_087_2986, w_087_2988, w_087_2989, w_087_2990, w_087_2991, w_087_2992, w_087_2993, w_087_2997, w_087_3000, w_087_3002, w_087_3003, w_087_3004, w_087_3008, w_087_3009, w_087_3012, w_087_3021, w_087_3023, w_087_3028, w_087_3030, w_087_3031, w_087_3032, w_087_3033, w_087_3035, w_087_3038, w_087_3042, w_087_3045, w_087_3048, w_087_3049, w_087_3052, w_087_3053, w_087_3054, w_087_3056, w_087_3059, w_087_3060, w_087_3063, w_087_3065, w_087_3069, w_087_3072, w_087_3074, w_087_3078, w_087_3079, w_087_3081, w_087_3085, w_087_3087, w_087_3091, w_087_3093, w_087_3097, w_087_3098, w_087_3099, w_087_3102, w_087_3104, w_087_3105, w_087_3109, w_087_3111, w_087_3113, w_087_3117, w_087_3119, w_087_3121, w_087_3123, w_087_3124, w_087_3128, w_087_3129, w_087_3131, w_087_3136, w_087_3137, w_087_3138, w_087_3140, w_087_3141, w_087_3144, w_087_3148, w_087_3152, w_087_3157, w_087_3158, w_087_3163, w_087_3164, w_087_3165, w_087_3166, w_087_3170, w_087_3172, w_087_3175, w_087_3177, w_087_3178, w_087_3180, w_087_3181, w_087_3182, w_087_3183, w_087_3184, w_087_3186, w_087_3187, w_087_3188, w_087_3189, w_087_3193, w_087_3197, w_087_3198, w_087_3199, w_087_3200, w_087_3201, w_087_3205, w_087_3206, w_087_3208, w_087_3210, w_087_3213, w_087_3214, w_087_3216, w_087_3219, w_087_3221, w_087_3224, w_087_3228, w_087_3229, w_087_3230, w_087_3231, w_087_3233, w_087_3234, w_087_3236, w_087_3242, w_087_3244, w_087_3247, w_087_3248, w_087_3250, w_087_3251, w_087_3254, w_087_3256, w_087_3257, w_087_3260, w_087_3261, w_087_3265, w_087_3272, w_087_3273, w_087_3275, w_087_3276, w_087_3277, w_087_3278, w_087_3280, w_087_3281, w_087_3285, w_087_3286, w_087_3289, w_087_3291, w_087_3293, w_087_3295, w_087_3297, w_087_3301, w_087_3302, w_087_3303, w_087_3304, w_087_3305, w_087_3313, w_087_3314, w_087_3315, w_087_3316, w_087_3317, w_087_3322, w_087_3323, w_087_3326, w_087_3330, w_087_3334, w_087_3335, w_087_3337, w_087_3341, w_087_3347, w_087_3349, w_087_3351, w_087_3352, w_087_3355, w_087_3356, w_087_3357, w_087_3361, w_087_3366, w_087_3367, w_087_3368, w_087_3373, w_087_3374, w_087_3377, w_087_3385, w_087_3386, w_087_3390, w_087_3392, w_087_3393, w_087_3394, w_087_3397, w_087_3398, w_087_3400, w_087_3401, w_087_3402, w_087_3406, w_087_3407, w_087_3409, w_087_3410, w_087_3413, w_087_3417, w_087_3418, w_087_3419, w_087_3420, w_087_3422, w_087_3423, w_087_3425, w_087_3428, w_087_3429, w_087_3430, w_087_3431, w_087_3434, w_087_3435, w_087_3436, w_087_3441, w_087_3442, w_087_3444, w_087_3446, w_087_3449, w_087_3451, w_087_3452, w_087_3453, w_087_3454, w_087_3457, w_087_3460, w_087_3467, w_087_3469, w_087_3471, w_087_3473, w_087_3475, w_087_3477, w_087_3479, w_087_3480, w_087_3481, w_087_3487, w_087_3492, w_087_3493, w_087_3498, w_087_3500, w_087_3501, w_087_3502, w_087_3505, w_087_3509, w_087_3511, w_087_3512, w_087_3513, w_087_3516, w_087_3517, w_087_3518, w_087_3520, w_087_3525, w_087_3526, w_087_3533, w_087_3534, w_087_3536, w_087_3538, w_087_3541, w_087_3544, w_087_3545, w_087_3546, w_087_3547, w_087_3548, w_087_3551, w_087_3552, w_087_3556, w_087_3557, w_087_3561, w_087_3562, w_087_3564, w_087_3566, w_087_3568, w_087_3572, w_087_3573, w_087_3574, w_087_3578, w_087_3579, w_087_3582, w_087_3583, w_087_3584, w_087_3587, w_087_3593, w_087_3595, w_087_3597, w_087_3601, w_087_3602, w_087_3603, w_087_3606, w_087_3611, w_087_3614, w_087_3615, w_087_3616, w_087_3619, w_087_3625, w_087_3626, w_087_3628, w_087_3631, w_087_3634, w_087_3637, w_087_3639, w_087_3640, w_087_3642, w_087_3643, w_087_3644, w_087_3647, w_087_3648, w_087_3649, w_087_3650, w_087_3651, w_087_3656, w_087_3657, w_087_3660, w_087_3664, w_087_3665, w_087_3666, w_087_3667, w_087_3669, w_087_3672, w_087_3673, w_087_3674, w_087_3675, w_087_3677, w_087_3679, w_087_3687, w_087_3691, w_087_3692, w_087_3697, w_087_3698, w_087_3700, w_087_3702, w_087_3706, w_087_3711, w_087_3712, w_087_3713, w_087_3718, w_087_3728, w_087_3734, w_087_3735, w_087_3737, w_087_3744, w_087_3745, w_087_3747, w_087_3763, w_087_3769, w_087_3780, w_087_3782, w_087_3796, w_087_3803, w_087_3808, w_087_3811, w_087_3813, w_087_3815, w_087_3816, w_087_3828, w_087_3831, w_087_3834, w_087_3841, w_087_3843, w_087_3854, w_087_3859, w_087_3860, w_087_3861, w_087_3866, w_087_3885, w_087_3886, w_087_3889, w_087_3890, w_087_3895, w_087_3897, w_087_3899, w_087_3900, w_087_3909, w_087_3915, w_087_3921, w_087_3923, w_087_3924, w_087_3926, w_087_3929, w_087_3932, w_087_3941, w_087_3948, w_087_3952, w_087_3953, w_087_3954, w_087_3965, w_087_3967, w_087_3968, w_087_3973, w_087_3975, w_087_3977, w_087_3979, w_087_3984, w_087_3985, w_087_3988, w_087_3993, w_087_3994, w_087_3996, w_087_3999, w_087_4005, w_087_4011, w_087_4015, w_087_4016, w_087_4018, w_087_4020, w_087_4026, w_087_4027, w_087_4033, w_087_4039, w_087_4043, w_087_4047, w_087_4056, w_087_4063, w_087_4068, w_087_4072, w_087_4081, w_087_4084, w_087_4097, w_087_4102, w_087_4104, w_087_4107, w_087_4112, w_087_4118, w_087_4123, w_087_4124, w_087_4133, w_087_4142, w_087_4149, w_087_4150, w_087_4152, w_087_4155, w_087_4156, w_087_4162, w_087_4163, w_087_4165, w_087_4167, w_087_4170, w_087_4174, w_087_4175, w_087_4176, w_087_4177, w_087_4182, w_087_4190, w_087_4192, w_087_4194, w_087_4203, w_087_4208, w_087_4212, w_087_4221, w_087_4225, w_087_4226, w_087_4235, w_087_4238, w_087_4239, w_087_4245, w_087_4246, w_087_4247, w_087_4251, w_087_4260, w_087_4264, w_087_4268, w_087_4274, w_087_4281, w_087_4294, w_087_4296, w_087_4297, w_087_4303, w_087_4308, w_087_4311, w_087_4314, w_087_4321, w_087_4322, w_087_4323, w_087_4324, w_087_4329, w_087_4330, w_087_4335, w_087_4344, w_087_4346, w_087_4348, w_087_4354, w_087_4359, w_087_4361, w_087_4362, w_087_4365, w_087_4367, w_087_4369, w_087_4371, w_087_4374, w_087_4377, w_087_4383, w_087_4384, w_087_4389, w_087_4390, w_087_4395, w_087_4410, w_087_4411, w_087_4412, w_087_4415, w_087_4430, w_087_4431, w_087_4433, w_087_4439, w_087_4448, w_087_4451, w_087_4454, w_087_4455, w_087_4456, w_087_4457, w_087_4458, w_087_4460, w_087_4464, w_087_4466, w_087_4467, w_087_4475, w_087_4477, w_087_4479, w_087_4481, w_087_4485, w_087_4486, w_087_4491, w_087_4493, w_087_4494, w_087_4495, w_087_4496, w_087_4500, w_087_4501, w_087_4507, w_087_4508, w_087_4509, w_087_4512, w_087_4515, w_087_4533, w_087_4539, w_087_4540, w_087_4542, w_087_4543, w_087_4544, w_087_4545, w_087_4549, w_087_4551, w_087_4553, w_087_4554, w_087_4558, w_087_4561, w_087_4562, w_087_4564, w_087_4568, w_087_4571, w_087_4572, w_087_4573, w_087_4574, w_087_4576, w_087_4578, w_087_4582, w_087_4584, w_087_4594, w_087_4599, w_087_4603, w_087_4608, w_087_4615, w_087_4625, w_087_4628, w_087_4629, w_087_4631, w_087_4636, w_087_4640, w_087_4642, w_087_4647, w_087_4655, w_087_4657, w_087_4658, w_087_4660, w_087_4661, w_087_4667, w_087_4669, w_087_4673, w_087_4690, w_087_4696, w_087_4701, w_087_4705, w_087_4710, w_087_4712, w_087_4716, w_087_4719, w_087_4721, w_087_4727, w_087_4730, w_087_4734, w_087_4735, w_087_4740, w_087_4742, w_087_4743, w_087_4746, w_087_4752, w_087_4753, w_087_4757, w_087_4762, w_087_4764, w_087_4765, w_087_4769, w_087_4770, w_087_4772, w_087_4774, w_087_4776, w_087_4777, w_087_4802, w_087_4803, w_087_4805, w_087_4810, w_087_4813, w_087_4815, w_087_4816, w_087_4817, w_087_4819, w_087_4821, w_087_4825, w_087_4829, w_087_4831, w_087_4835, w_087_4836, w_087_4837, w_087_4843, w_087_4847, w_087_4848, w_087_4862, w_087_4868, w_087_4870, w_087_4871, w_087_4878, w_087_4883, w_087_4888, w_087_4893, w_087_4897, w_087_4922, w_087_4924, w_087_4925, w_087_4926, w_087_4929, w_087_4938, w_087_4942, w_087_4943, w_087_4947, w_087_4960, w_087_4963, w_087_4971, w_087_4977, w_087_4978, w_087_4982, w_087_4983, w_087_4989, w_087_4990, w_087_4993, w_087_5007, w_087_5012, w_087_5013, w_087_5027, w_087_5030, w_087_5031, w_087_5035, w_087_5037, w_087_5045, w_087_5048, w_087_5052, w_087_5053, w_087_5057, w_087_5059, w_087_5064, w_087_5065, w_087_5068, w_087_5072, w_087_5074, w_087_5076, w_087_5077, w_087_5078, w_087_5086, w_087_5090, w_087_5092, w_087_5111, w_087_5114, w_087_5119, w_087_5120, w_087_5128, w_087_5130, w_087_5132, w_087_5135, w_087_5149, w_087_5152, w_087_5154, w_087_5158, w_087_5159, w_087_5164, w_087_5165, w_087_5167, w_087_5174, w_087_5175, w_087_5177, w_087_5191, w_087_5200, w_087_5203, w_087_5211, w_087_5218, w_087_5222, w_087_5224, w_087_5235, w_087_5238, w_087_5245, w_087_5247, w_087_5249, w_087_5257, w_087_5258, w_087_5260, w_087_5263, w_087_5267, w_087_5271, w_087_5273, w_087_5274, w_087_5275, w_087_5283, w_087_5285, w_087_5286, w_087_5294, w_087_5295, w_087_5296, w_087_5301, w_087_5302, w_087_5303, w_087_5304, w_087_5305, w_087_5310, w_087_5311, w_087_5312, w_087_5313, w_087_5319, w_087_5321, w_087_5322, w_087_5332, w_087_5335, w_087_5337, w_087_5344, w_087_5345, w_087_5350, w_087_5352, w_087_5357, w_087_5359, w_087_5362, w_087_5389, w_087_5390, w_087_5391, w_087_5393, w_087_5395, w_087_5400, w_087_5401, w_087_5407, w_087_5409, w_087_5411, w_087_5412, w_087_5413, w_087_5418, w_087_5421, w_087_5422, w_087_5424, w_087_5425, w_087_5430, w_087_5437, w_087_5446, w_087_5449, w_087_5450, w_087_5453, w_087_5457, w_087_5458, w_087_5463, w_087_5472, w_087_5477, w_087_5478, w_087_5482, w_087_5488, w_087_5494, w_087_5496, w_087_5508, w_087_5509, w_087_5510, w_087_5511, w_087_5514, w_087_5516, w_087_5527, w_087_5528, w_087_5529, w_087_5540, w_087_5543, w_087_5544, w_087_5547, w_087_5548, w_087_5557, w_087_5558, w_087_5562, w_087_5579, w_087_5580, w_087_5582, w_087_5586, w_087_5589, w_087_5595, w_087_5597, w_087_5598, w_087_5601, w_087_5603, w_087_5606, w_087_5608, w_087_5609, w_087_5611, w_087_5613, w_087_5617, w_087_5631, w_087_5632, w_087_5633, w_087_5636, w_087_5638, w_087_5642, w_087_5645, w_087_5649, w_087_5651, w_087_5673, w_087_5675, w_087_5682, w_087_5683, w_087_5685, w_087_5687, w_087_5690, w_087_5692, w_087_5701, w_087_5702, w_087_5707, w_087_5718, w_087_5720, w_087_5727, w_087_5728, w_087_5732, w_087_5733, w_087_5735, w_087_5737, w_087_5739, w_087_5741, w_087_5746, w_087_5747, w_087_5748, w_087_5749, w_087_5750, w_087_5751, w_087_5752, w_087_5754, w_087_5755, w_087_5762, w_087_5763, w_087_5766, w_087_5769, w_087_5777, w_087_5778, w_087_5784, w_087_5787, w_087_5792, w_087_5796, w_087_5798, w_087_5799, w_087_5800, w_087_5801, w_087_5806, w_087_5813, w_087_5820, w_087_5826, w_087_5827, w_087_5828, w_087_5830, w_087_5839, w_087_5844, w_087_5847, w_087_5853, w_087_5857, w_087_5866, w_087_5867, w_087_5885, w_087_5890, w_087_5899, w_087_5900, w_087_5901, w_087_5909, w_087_5911, w_087_5916, w_087_5920, w_087_5925, w_087_5927, w_087_5928, w_087_5929, w_087_5931, w_087_5933, w_087_5934, w_087_5935, w_087_5938, w_087_5944, w_087_5945, w_087_5959, w_087_5963, w_087_5970, w_087_5973, w_087_5979, w_087_5981, w_087_5983, w_087_5986, w_087_5990, w_087_5994, w_087_5995, w_087_6002, w_087_6005, w_087_6007, w_087_6010, w_087_6021, w_087_6024, w_087_6025, w_087_6030, w_087_6031, w_087_6032, w_087_6033, w_087_6034, w_087_6041, w_087_6053, w_087_6055, w_087_6059, w_087_6060, w_087_6062, w_087_6067, w_087_6068, w_087_6069, w_087_6070, w_087_6073, w_087_6079, w_087_6081, w_087_6082, w_087_6087, w_087_6090, w_087_6095, w_087_6096, w_087_6100, w_087_6104, w_087_6105, w_087_6110, w_087_6111, w_087_6113, w_087_6118, w_087_6124, w_087_6127, w_087_6139, w_087_6157, w_087_6158, w_087_6161, w_087_6163, w_087_6165, w_087_6166, w_087_6169, w_087_6171, w_087_6175, w_087_6176, w_087_6177, w_087_6180, w_087_6191, w_087_6196, w_087_6202, w_087_6203, w_087_6208, w_087_6213, w_087_6222, w_087_6227, w_087_6231, w_087_6238, w_087_6244, w_087_6245, w_087_6249, w_087_6250, w_087_6251, w_087_6252, w_087_6268, w_087_6269, w_087_6270, w_087_6273, w_087_6274, w_087_6280, w_087_6286, w_087_6288, w_087_6291;
  wire w_088_001, w_088_008, w_088_009, w_088_010, w_088_013, w_088_017, w_088_019, w_088_020, w_088_025, w_088_028, w_088_029, w_088_030, w_088_034, w_088_037, w_088_038, w_088_039, w_088_044, w_088_045, w_088_049, w_088_052, w_088_055, w_088_056, w_088_058, w_088_060, w_088_061, w_088_062, w_088_063, w_088_067, w_088_070, w_088_073, w_088_074, w_088_075, w_088_077, w_088_080, w_088_083, w_088_084, w_088_085, w_088_092, w_088_094, w_088_096, w_088_097, w_088_098, w_088_101, w_088_103, w_088_105, w_088_115, w_088_118, w_088_120, w_088_123, w_088_125, w_088_129, w_088_130, w_088_132, w_088_135, w_088_139, w_088_140, w_088_141, w_088_144, w_088_151, w_088_155, w_088_158, w_088_159, w_088_160, w_088_164, w_088_165, w_088_166, w_088_173, w_088_174, w_088_179, w_088_181, w_088_182, w_088_183, w_088_188, w_088_189, w_088_190, w_088_191, w_088_192, w_088_193, w_088_195, w_088_196, w_088_198, w_088_199, w_088_201, w_088_203, w_088_207, w_088_208, w_088_211, w_088_215, w_088_216, w_088_220, w_088_222, w_088_225, w_088_228, w_088_231, w_088_234, w_088_235, w_088_237, w_088_240, w_088_241, w_088_242, w_088_244, w_088_247, w_088_248, w_088_249, w_088_250, w_088_251, w_088_253, w_088_261, w_088_262, w_088_263, w_088_265, w_088_268, w_088_271, w_088_273, w_088_274, w_088_275, w_088_278, w_088_279, w_088_280, w_088_281, w_088_282, w_088_284, w_088_286, w_088_289, w_088_295, w_088_296, w_088_298, w_088_299, w_088_300, w_088_301, w_088_305, w_088_306, w_088_309, w_088_311, w_088_313, w_088_314, w_088_315, w_088_318, w_088_320, w_088_322, w_088_326, w_088_327, w_088_328, w_088_329, w_088_330, w_088_331, w_088_332, w_088_334, w_088_335, w_088_336, w_088_337, w_088_341, w_088_343, w_088_344, w_088_346, w_088_347, w_088_350, w_088_354, w_088_355, w_088_356, w_088_357, w_088_358, w_088_360, w_088_363, w_088_365, w_088_366, w_088_367, w_088_368, w_088_369, w_088_370, w_088_371, w_088_373, w_088_374, w_088_375, w_088_376, w_088_379, w_088_380, w_088_383, w_088_384, w_088_385, w_088_387, w_088_389, w_088_392, w_088_396, w_088_398, w_088_403, w_088_404, w_088_405, w_088_408, w_088_409, w_088_410, w_088_411, w_088_412, w_088_414, w_088_415, w_088_416, w_088_417, w_088_420, w_088_425, w_088_426, w_088_443, w_088_446, w_088_448, w_088_449, w_088_455, w_088_461, w_088_462, w_088_468, w_088_469, w_088_471, w_088_473, w_088_474, w_088_475, w_088_477, w_088_479, w_088_482, w_088_484, w_088_485, w_088_486, w_088_489, w_088_490, w_088_495, w_088_498, w_088_502, w_088_503, w_088_505, w_088_508, w_088_509, w_088_510, w_088_511, w_088_513, w_088_517, w_088_520, w_088_521, w_088_522, w_088_524, w_088_528, w_088_529, w_088_531, w_088_534, w_088_536, w_088_540, w_088_542, w_088_544, w_088_545, w_088_549, w_088_553, w_088_554, w_088_555, w_088_556, w_088_561, w_088_562, w_088_563, w_088_564, w_088_566, w_088_567, w_088_568, w_088_570, w_088_572, w_088_574, w_088_576, w_088_577, w_088_578, w_088_579, w_088_580, w_088_584, w_088_586, w_088_589, w_088_590, w_088_593, w_088_594, w_088_598, w_088_600, w_088_603, w_088_612, w_088_617, w_088_621, w_088_624, w_088_630, w_088_633, w_088_634, w_088_637, w_088_639, w_088_640, w_088_642, w_088_643, w_088_644, w_088_646, w_088_648, w_088_649, w_088_654, w_088_656, w_088_658, w_088_660, w_088_663, w_088_671, w_088_672, w_088_675, w_088_676, w_088_677, w_088_678, w_088_681, w_088_684, w_088_689, w_088_690, w_088_691, w_088_692, w_088_693, w_088_695, w_088_696, w_088_697, w_088_699, w_088_700, w_088_704, w_088_705, w_088_706, w_088_707, w_088_708, w_088_709, w_088_710, w_088_712, w_088_715, w_088_717, w_088_718, w_088_720, w_088_728, w_088_729, w_088_731, w_088_732, w_088_736, w_088_739, w_088_742, w_088_743, w_088_744, w_088_746, w_088_750, w_088_751, w_088_753, w_088_755, w_088_758, w_088_759, w_088_762, w_088_763, w_088_770, w_088_771, w_088_772, w_088_774, w_088_777, w_088_780, w_088_787, w_088_789, w_088_791, w_088_794, w_088_795, w_088_798, w_088_801, w_088_803, w_088_804, w_088_805, w_088_806, w_088_807, w_088_808, w_088_811, w_088_813, w_088_814, w_088_815, w_088_816, w_088_817, w_088_823, w_088_824, w_088_826, w_088_827, w_088_829, w_088_831, w_088_836, w_088_845, w_088_849, w_088_850, w_088_851, w_088_854, w_088_856, w_088_857, w_088_860, w_088_866, w_088_871, w_088_876, w_088_877, w_088_878, w_088_880, w_088_881, w_088_882, w_088_883, w_088_887, w_088_893, w_088_894, w_088_895, w_088_897, w_088_898, w_088_899, w_088_900, w_088_907, w_088_909, w_088_912, w_088_916, w_088_917, w_088_919, w_088_920, w_088_921, w_088_925, w_088_926, w_088_930, w_088_931, w_088_932, w_088_936, w_088_937, w_088_940, w_088_942, w_088_943, w_088_944, w_088_946, w_088_947, w_088_951, w_088_957, w_088_958, w_088_962, w_088_964, w_088_965, w_088_968, w_088_974, w_088_975, w_088_977, w_088_980, w_088_981, w_088_985, w_088_989, w_088_992, w_088_998, w_088_1003, w_088_1006, w_088_1008, w_088_1009, w_088_1011, w_088_1012, w_088_1014, w_088_1015, w_088_1016, w_088_1018, w_088_1020, w_088_1022, w_088_1023, w_088_1024, w_088_1025, w_088_1026, w_088_1029, w_088_1030, w_088_1035, w_088_1037, w_088_1038, w_088_1039, w_088_1040, w_088_1042, w_088_1047, w_088_1049, w_088_1052, w_088_1053, w_088_1058, w_088_1059, w_088_1061, w_088_1062, w_088_1068, w_088_1071, w_088_1073, w_088_1074, w_088_1076, w_088_1078, w_088_1083, w_088_1084, w_088_1085, w_088_1087, w_088_1088, w_088_1090, w_088_1092, w_088_1093, w_088_1094, w_088_1098, w_088_1100, w_088_1102, w_088_1103, w_088_1104, w_088_1116, w_088_1118, w_088_1122, w_088_1123, w_088_1124, w_088_1125, w_088_1129, w_088_1130, w_088_1131, w_088_1134, w_088_1138, w_088_1141, w_088_1144, w_088_1146, w_088_1147, w_088_1148, w_088_1149, w_088_1151, w_088_1153, w_088_1155, w_088_1156, w_088_1158, w_088_1160, w_088_1161, w_088_1162, w_088_1163, w_088_1164, w_088_1165, w_088_1166, w_088_1168, w_088_1169, w_088_1170, w_088_1173, w_088_1175, w_088_1176, w_088_1182, w_088_1185, w_088_1186, w_088_1189, w_088_1190, w_088_1192, w_088_1193, w_088_1198, w_088_1199, w_088_1200, w_088_1201, w_088_1203, w_088_1204, w_088_1205, w_088_1209, w_088_1210, w_088_1217, w_088_1218, w_088_1221, w_088_1222, w_088_1225, w_088_1226, w_088_1229, w_088_1231, w_088_1236, w_088_1238, w_088_1240, w_088_1248, w_088_1250, w_088_1252, w_088_1254, w_088_1256, w_088_1258, w_088_1259, w_088_1260, w_088_1264, w_088_1267, w_088_1271, w_088_1274, w_088_1276, w_088_1279, w_088_1280, w_088_1281, w_088_1282, w_088_1287, w_088_1289, w_088_1291, w_088_1292, w_088_1293, w_088_1294, w_088_1295, w_088_1298, w_088_1299, w_088_1300, w_088_1302, w_088_1305, w_088_1306, w_088_1307, w_088_1309, w_088_1310, w_088_1315, w_088_1322, w_088_1323, w_088_1324, w_088_1326, w_088_1328, w_088_1329, w_088_1332, w_088_1334, w_088_1336, w_088_1341, w_088_1344, w_088_1346, w_088_1350, w_088_1354, w_088_1356, w_088_1357, w_088_1361, w_088_1365, w_088_1368, w_088_1370, w_088_1373, w_088_1374, w_088_1376, w_088_1378, w_088_1383, w_088_1384, w_088_1385, w_088_1386, w_088_1388, w_088_1390, w_088_1391, w_088_1397, w_088_1401, w_088_1402, w_088_1403, w_088_1404, w_088_1407, w_088_1410, w_088_1411, w_088_1412, w_088_1414, w_088_1415, w_088_1418, w_088_1423, w_088_1432, w_088_1433, w_088_1434, w_088_1436, w_088_1437, w_088_1438, w_088_1440, w_088_1442, w_088_1443, w_088_1447, w_088_1452, w_088_1453, w_088_1454, w_088_1457, w_088_1458, w_088_1463, w_088_1464, w_088_1467, w_088_1469, w_088_1471, w_088_1472, w_088_1473, w_088_1474, w_088_1475, w_088_1477, w_088_1480, w_088_1481, w_088_1483, w_088_1486, w_088_1487, w_088_1488, w_088_1490, w_088_1492, w_088_1497, w_088_1498, w_088_1501, w_088_1502, w_088_1503, w_088_1505, w_088_1508, w_088_1512, w_088_1513, w_088_1514, w_088_1515, w_088_1518, w_088_1520, w_088_1521, w_088_1525, w_088_1527, w_088_1529, w_088_1530, w_088_1531, w_088_1535, w_088_1536, w_088_1537, w_088_1538, w_088_1540, w_088_1541, w_088_1543, w_088_1546, w_088_1549, w_088_1552, w_088_1553, w_088_1555, w_088_1556, w_088_1560, w_088_1562, w_088_1563, w_088_1565, w_088_1567, w_088_1570, w_088_1571, w_088_1572, w_088_1573, w_088_1577, w_088_1581, w_088_1582, w_088_1584, w_088_1586, w_088_1588, w_088_1591, w_088_1592, w_088_1593, w_088_1594, w_088_1600, w_088_1601, w_088_1602, w_088_1605, w_088_1606, w_088_1607, w_088_1608, w_088_1612, w_088_1613, w_088_1614, w_088_1616, w_088_1618, w_088_1622, w_088_1624, w_088_1625, w_088_1628, w_088_1629, w_088_1630, w_088_1632, w_088_1633, w_088_1635, w_088_1640, w_088_1644, w_088_1645, w_088_1646, w_088_1648, w_088_1650, w_088_1653, w_088_1656, w_088_1659, w_088_1660, w_088_1662, w_088_1664, w_088_1667, w_088_1668, w_088_1669, w_088_1670, w_088_1672, w_088_1673, w_088_1680, w_088_1690, w_088_1691, w_088_1692, w_088_1698, w_088_1700, w_088_1701, w_088_1705, w_088_1707, w_088_1714, w_088_1715, w_088_1716, w_088_1722, w_088_1723, w_088_1725, w_088_1727, w_088_1731, w_088_1732, w_088_1733, w_088_1738, w_088_1744, w_088_1745, w_088_1747, w_088_1749, w_088_1751, w_088_1752, w_088_1755, w_088_1759, w_088_1760, w_088_1761, w_088_1771, w_088_1778, w_088_1781, w_088_1787, w_088_1790, w_088_1791, w_088_1798, w_088_1803, w_088_1805, w_088_1806, w_088_1809, w_088_1818, w_088_1820, w_088_1823, w_088_1824, w_088_1825, w_088_1828, w_088_1829, w_088_1830, w_088_1841, w_088_1845, w_088_1846, w_088_1847, w_088_1850, w_088_1851, w_088_1856, w_088_1858, w_088_1865, w_088_1871, w_088_1872, w_088_1879, w_088_1880, w_088_1881, w_088_1883, w_088_1884, w_088_1887, w_088_1889, w_088_1891, w_088_1895, w_088_1896, w_088_1901, w_088_1908, w_088_1918, w_088_1920, w_088_1926, w_088_1931, w_088_1932, w_088_1935, w_088_1939, w_088_1940, w_088_1942, w_088_1944, w_088_1963, w_088_1964, w_088_1967, w_088_1969, w_088_1970, w_088_1972, w_088_1977, w_088_1981, w_088_1985, w_088_1991, w_088_1993, w_088_1994, w_088_1996, w_088_2007, w_088_2009, w_088_2015, w_088_2019, w_088_2020, w_088_2023, w_088_2027, w_088_2028, w_088_2033, w_088_2039, w_088_2044, w_088_2048, w_088_2050, w_088_2070, w_088_2073, w_088_2074, w_088_2082, w_088_2086, w_088_2092, w_088_2093, w_088_2096, w_088_2104, w_088_2108, w_088_2120, w_088_2126, w_088_2129, w_088_2132, w_088_2135, w_088_2139, w_088_2141, w_088_2143, w_088_2148, w_088_2149, w_088_2153, w_088_2155, w_088_2159, w_088_2167, w_088_2171, w_088_2177, w_088_2179, w_088_2183, w_088_2188, w_088_2189, w_088_2191, w_088_2200, w_088_2201, w_088_2205, w_088_2209, w_088_2213, w_088_2216, w_088_2228, w_088_2232, w_088_2235, w_088_2236, w_088_2243, w_088_2244, w_088_2250, w_088_2252, w_088_2253, w_088_2254, w_088_2257, w_088_2262, w_088_2270, w_088_2271, w_088_2272, w_088_2274, w_088_2275, w_088_2276, w_088_2281, w_088_2283, w_088_2289, w_088_2290, w_088_2293, w_088_2294, w_088_2295, w_088_2297, w_088_2298, w_088_2299, w_088_2300, w_088_2301, w_088_2302, w_088_2303, w_088_2309, w_088_2311, w_088_2314, w_088_2317, w_088_2319, w_088_2320, w_088_2325, w_088_2332, w_088_2335, w_088_2339, w_088_2341, w_088_2343, w_088_2345, w_088_2349, w_088_2364, w_088_2367, w_088_2370, w_088_2371, w_088_2373, w_088_2376, w_088_2382, w_088_2383, w_088_2398, w_088_2401, w_088_2404, w_088_2407, w_088_2408, w_088_2413, w_088_2416, w_088_2420, w_088_2423, w_088_2428, w_088_2430, w_088_2431, w_088_2433, w_088_2437, w_088_2438, w_088_2444, w_088_2455, w_088_2463, w_088_2467, w_088_2468, w_088_2472, w_088_2478, w_088_2481, w_088_2483, w_088_2485, w_088_2491, w_088_2492, w_088_2497, w_088_2498, w_088_2502, w_088_2508, w_088_2514, w_088_2515, w_088_2516, w_088_2519, w_088_2522, w_088_2523, w_088_2526, w_088_2533, w_088_2536, w_088_2541, w_088_2548, w_088_2553, w_088_2560, w_088_2565, w_088_2567, w_088_2577, w_088_2580, w_088_2583, w_088_2586, w_088_2587, w_088_2588, w_088_2610, w_088_2616, w_088_2620, w_088_2623, w_088_2624, w_088_2626, w_088_2632, w_088_2633, w_088_2635, w_088_2644, w_088_2647, w_088_2648, w_088_2651, w_088_2653, w_088_2662, w_088_2668, w_088_2671, w_088_2675, w_088_2676, w_088_2680, w_088_2687, w_088_2700, w_088_2702, w_088_2705, w_088_2706, w_088_2708, w_088_2716, w_088_2727, w_088_2728, w_088_2731, w_088_2734, w_088_2737, w_088_2745, w_088_2746, w_088_2747, w_088_2752, w_088_2756, w_088_2765, w_088_2774, w_088_2778, w_088_2786, w_088_2789, w_088_2790, w_088_2792, w_088_2793, w_088_2796, w_088_2797, w_088_2810, w_088_2816, w_088_2822, w_088_2829, w_088_2832, w_088_2837, w_088_2840, w_088_2844, w_088_2847, w_088_2849, w_088_2862, w_088_2866, w_088_2870, w_088_2874, w_088_2876, w_088_2878, w_088_2885, w_088_2886, w_088_2898, w_088_2902, w_088_2910, w_088_2914, w_088_2916, w_088_2920, w_088_2921, w_088_2926, w_088_2928, w_088_2935, w_088_2938, w_088_2939, w_088_2941, w_088_2944, w_088_2945, w_088_2955, w_088_2957, w_088_2959, w_088_2960, w_088_2969, w_088_2972, w_088_2977, w_088_2996, w_088_2999, w_088_3001, w_088_3003, w_088_3008, w_088_3015, w_088_3018, w_088_3019, w_088_3025, w_088_3029, w_088_3030, w_088_3040, w_088_3046, w_088_3048, w_088_3053, w_088_3055, w_088_3056, w_088_3057, w_088_3058, w_088_3062, w_088_3076, w_088_3077, w_088_3080, w_088_3086, w_088_3087, w_088_3089, w_088_3090, w_088_3095, w_088_3096, w_088_3102, w_088_3112, w_088_3115, w_088_3121, w_088_3122, w_088_3125, w_088_3126, w_088_3131, w_088_3132, w_088_3134, w_088_3136, w_088_3143, w_088_3144, w_088_3145, w_088_3146, w_088_3148, w_088_3150, w_088_3153, w_088_3156, w_088_3159, w_088_3162, w_088_3176, w_088_3178, w_088_3182, w_088_3183, w_088_3188, w_088_3189, w_088_3191, w_088_3192, w_088_3198, w_088_3200, w_088_3210, w_088_3217, w_088_3219, w_088_3221, w_088_3222, w_088_3223, w_088_3232, w_088_3233, w_088_3235, w_088_3238, w_088_3240, w_088_3242, w_088_3243, w_088_3244, w_088_3246, w_088_3254, w_088_3258, w_088_3259, w_088_3260, w_088_3263, w_088_3264, w_088_3265, w_088_3270, w_088_3273, w_088_3279, w_088_3284, w_088_3288, w_088_3292, w_088_3295, w_088_3296, w_088_3298, w_088_3299, w_088_3300, w_088_3302, w_088_3312, w_088_3321, w_088_3322, w_088_3325, w_088_3327, w_088_3330, w_088_3333, w_088_3334, w_088_3337, w_088_3340, w_088_3341, w_088_3345, w_088_3346, w_088_3349, w_088_3353, w_088_3356, w_088_3359, w_088_3360, w_088_3366, w_088_3368, w_088_3372, w_088_3377, w_088_3382, w_088_3386, w_088_3388, w_088_3393, w_088_3394, w_088_3397, w_088_3400, w_088_3401, w_088_3404, w_088_3411, w_088_3414, w_088_3422, w_088_3425, w_088_3427, w_088_3429, w_088_3432, w_088_3433, w_088_3434, w_088_3436, w_088_3439, w_088_3440, w_088_3442, w_088_3444, w_088_3446, w_088_3457, w_088_3465, w_088_3470, w_088_3472, w_088_3474, w_088_3476, w_088_3479, w_088_3483, w_088_3484, w_088_3485, w_088_3487, w_088_3490, w_088_3499, w_088_3512, w_088_3515, w_088_3519, w_088_3520, w_088_3525, w_088_3529, w_088_3536, w_088_3539, w_088_3540, w_088_3545, w_088_3547, w_088_3548, w_088_3554, w_088_3555, w_088_3556, w_088_3557, w_088_3558, w_088_3560, w_088_3566, w_088_3570, w_088_3573, w_088_3576, w_088_3579, w_088_3583, w_088_3586, w_088_3588, w_088_3593, w_088_3597, w_088_3605, w_088_3608, w_088_3610, w_088_3613, w_088_3619, w_088_3626, w_088_3628, w_088_3630, w_088_3631, w_088_3632, w_088_3634, w_088_3642, w_088_3652, w_088_3656, w_088_3662, w_088_3663, w_088_3673, w_088_3674, w_088_3675, w_088_3680, w_088_3681, w_088_3683, w_088_3687, w_088_3688, w_088_3694, w_088_3695, w_088_3696, w_088_3700, w_088_3703, w_088_3704, w_088_3705, w_088_3707, w_088_3710, w_088_3712, w_088_3723, w_088_3724, w_088_3740, w_088_3745, w_088_3751, w_088_3755, w_088_3760, w_088_3761, w_088_3762, w_088_3764, w_088_3778, w_088_3779, w_088_3783, w_088_3784, w_088_3789, w_088_3796, w_088_3801, w_088_3803, w_088_3809, w_088_3819, w_088_3823, w_088_3824, w_088_3825, w_088_3828, w_088_3834, w_088_3835, w_088_3841, w_088_3845, w_088_3846, w_088_3848, w_088_3849, w_088_3853, w_088_3858, w_088_3865, w_088_3870, w_088_3872, w_088_3880, w_088_3881, w_088_3888, w_088_3891, w_088_3894, w_088_3899, w_088_3902, w_088_3903, w_088_3904, w_088_3908, w_088_3911, w_088_3915, w_088_3916, w_088_3919, w_088_3920, w_088_3921, w_088_3925, w_088_3927, w_088_3932, w_088_3934, w_088_3936, w_088_3942, w_088_3943, w_088_3948, w_088_3952, w_088_3953, w_088_3959, w_088_3962, w_088_3966, w_088_3971, w_088_3972, w_088_3975, w_088_3977, w_088_3982, w_088_3984, w_088_3986, w_088_3988, w_088_3997, w_088_3999, w_088_4003, w_088_4006, w_088_4019, w_088_4020, w_088_4022, w_088_4023, w_088_4026, w_088_4036, w_088_4037, w_088_4038, w_088_4046, w_088_4049, w_088_4051, w_088_4056, w_088_4059, w_088_4060, w_088_4062, w_088_4065, w_088_4066, w_088_4067, w_088_4068, w_088_4071, w_088_4073, w_088_4085, w_088_4090, w_088_4092, w_088_4094, w_088_4096, w_088_4097, w_088_4098, w_088_4102, w_088_4110, w_088_4115, w_088_4117, w_088_4118, w_088_4122, w_088_4126, w_088_4127, w_088_4128, w_088_4132, w_088_4134, w_088_4140, w_088_4144, w_088_4151, w_088_4153, w_088_4154, w_088_4158, w_088_4159, w_088_4161, w_088_4163, w_088_4167, w_088_4168, w_088_4172, w_088_4174, w_088_4178, w_088_4181, w_088_4182, w_088_4185, w_088_4188, w_088_4194, w_088_4198, w_088_4202, w_088_4205, w_088_4218, w_088_4222, w_088_4228, w_088_4231, w_088_4235, w_088_4237, w_088_4241, w_088_4244, w_088_4246, w_088_4254, w_088_4256, w_088_4258, w_088_4267, w_088_4269, w_088_4272, w_088_4278, w_088_4280, w_088_4282, w_088_4283, w_088_4300, w_088_4307, w_088_4314, w_088_4320, w_088_4321, w_088_4324, w_088_4326, w_088_4331, w_088_4341, w_088_4343, w_088_4346, w_088_4347, w_088_4351, w_088_4353, w_088_4355, w_088_4362, w_088_4365, w_088_4371, w_088_4378, w_088_4380, w_088_4391, w_088_4392, w_088_4399, w_088_4401, w_088_4406, w_088_4410, w_088_4414, w_088_4415, w_088_4416, w_088_4422, w_088_4425, w_088_4426, w_088_4428, w_088_4435, w_088_4442, w_088_4445, w_088_4453, w_088_4458, w_088_4460, w_088_4461, w_088_4462, w_088_4463, w_088_4464, w_088_4465, w_088_4471, w_088_4477, w_088_4493, w_088_4494, w_088_4497, w_088_4498, w_088_4500, w_088_4506, w_088_4508, w_088_4514, w_088_4519, w_088_4526, w_088_4527, w_088_4533, w_088_4535, w_088_4541, w_088_4549, w_088_4554, w_088_4555, w_088_4578, w_088_4588, w_088_4590, w_088_4592, w_088_4596, w_088_4606, w_088_4612, w_088_4616, w_088_4617, w_088_4624, w_088_4627, w_088_4628, w_088_4632, w_088_4638, w_088_4640, w_088_4645, w_088_4649, w_088_4652, w_088_4657, w_088_4660, w_088_4663, w_088_4665, w_088_4667, w_088_4676, w_088_4686, w_088_4692, w_088_4693, w_088_4694, w_088_4699, w_088_4700, w_088_4702, w_088_4704, w_088_4707, w_088_4715, w_088_4717, w_088_4718, w_088_4719, w_088_4721, w_088_4724, w_088_4727, w_088_4728, w_088_4735, w_088_4737, w_088_4742, w_088_4744, w_088_4747, w_088_4754, w_088_4757, w_088_4762, w_088_4763, w_088_4766, w_088_4767, w_088_4768, w_088_4773, w_088_4774, w_088_4782, w_088_4785, w_088_4787, w_088_4792, w_088_4799, w_088_4803, w_088_4805, w_088_4813, w_088_4815, w_088_4817, w_088_4820, w_088_4822, w_088_4823, w_088_4825, w_088_4830, w_088_4831, w_088_4835, w_088_4841, w_088_4842, w_088_4844, w_088_4848, w_088_4853, w_088_4883, w_088_4887, w_088_4891, w_088_4899, w_088_4903, w_088_4905, w_088_4906, w_088_4907, w_088_4921, w_088_4932, w_088_4940, w_088_4941, w_088_4943, w_088_4948, w_088_4950, w_088_4951, w_088_4957, w_088_4960, w_088_4965, w_088_4968, w_088_4970, w_088_4974, w_088_4975, w_088_4980, w_088_4985, w_088_4987, w_088_4989, w_088_5001, w_088_5004, w_088_5005, w_088_5006, w_088_5007, w_088_5014, w_088_5023, w_088_5025, w_088_5027, w_088_5038, w_088_5042, w_088_5045, w_088_5048, w_088_5049, w_088_5051, w_088_5052, w_088_5053, w_088_5055, w_088_5056, w_088_5061, w_088_5064, w_088_5065, w_088_5067, w_088_5068, w_088_5074, w_088_5079, w_088_5083, w_088_5090, w_088_5094, w_088_5095, w_088_5096, w_088_5112, w_088_5127, w_088_5128, w_088_5129, w_088_5135, w_088_5137, w_088_5138, w_088_5141, w_088_5143, w_088_5147, w_088_5169, w_088_5171, w_088_5178, w_088_5184, w_088_5186, w_088_5188, w_088_5190, w_088_5199, w_088_5201, w_088_5203, w_088_5210, w_088_5218, w_088_5219, w_088_5226, w_088_5231, w_088_5232, w_088_5234, w_088_5237, w_088_5240, w_088_5244, w_088_5247, w_088_5250, w_088_5252, w_088_5253, w_088_5256, w_088_5261, w_088_5270, w_088_5272, w_088_5273, w_088_5275, w_088_5279, w_088_5281, w_088_5282, w_088_5285, w_088_5287, w_088_5288, w_088_5291, w_088_5296, w_088_5298, w_088_5304, w_088_5305, w_088_5309, w_088_5313, w_088_5317, w_088_5321, w_088_5323, w_088_5326, w_088_5329, w_088_5332, w_088_5334, w_088_5337, w_088_5338, w_088_5339, w_088_5343, w_088_5347, w_088_5349, w_088_5350, w_088_5355, w_088_5356, w_088_5358, w_088_5365, w_088_5368, w_088_5369, w_088_5374, w_088_5377, w_088_5383, w_088_5387, w_088_5391, w_088_5393, w_088_5394, w_088_5395, w_088_5399, w_088_5405, w_088_5412, w_088_5414, w_088_5415, w_088_5419, w_088_5420, w_088_5423, w_088_5434, w_088_5437, w_088_5441, w_088_5443, w_088_5444, w_088_5450, w_088_5451, w_088_5452, w_088_5453, w_088_5454, w_088_5455, w_088_5456, w_088_5457, w_088_5461, w_088_5462, w_088_5465, w_088_5466, w_088_5467, w_088_5475, w_088_5476, w_088_5479, w_088_5481, w_088_5484, w_088_5488, w_088_5490, w_088_5491, w_088_5493, w_088_5494, w_088_5496, w_088_5497, w_088_5502, w_088_5503, w_088_5510, w_088_5520, w_088_5522, w_088_5525, w_088_5529, w_088_5533, w_088_5539, w_088_5560, w_088_5565, w_088_5572, w_088_5582, w_088_5584, w_088_5587, w_088_5589, w_088_5594, w_088_5598, w_088_5602, w_088_5605, w_088_5607, w_088_5610, w_088_5611, w_088_5613, w_088_5622, w_088_5624, w_088_5625, w_088_5627, w_088_5629, w_088_5631, w_088_5646, w_088_5657, w_088_5658, w_088_5659, w_088_5663, w_088_5674, w_088_5675, w_088_5684, w_088_5686, w_088_5690, w_088_5705, w_088_5717, w_088_5718, w_088_5720, w_088_5722, w_088_5723, w_088_5727, w_088_5738, w_088_5740, w_088_5755, w_088_5757, w_088_5758, w_088_5768, w_088_5774, w_088_5776, w_088_5785, w_088_5786, w_088_5787, w_088_5803, w_088_5808, w_088_5809, w_088_5824, w_088_5825, w_088_5827, w_088_5832, w_088_5836, w_088_5842, w_088_5844, w_088_5845, w_088_5849, w_088_5852, w_088_5859, w_088_5876, w_088_5879, w_088_5886, w_088_5889, w_088_5892, w_088_5895, w_088_5901, w_088_5905, w_088_5922, w_088_5929, w_088_5932, w_088_5934, w_088_5935, w_088_5941, w_088_5942, w_088_5944, w_088_5947, w_088_5949, w_088_5952, w_088_5960, w_088_5961, w_088_5968, w_088_5972, w_088_5975, w_088_5982, w_088_5984, w_088_5988, w_088_5991, w_088_5996, w_088_6001, w_088_6006, w_088_6011, w_088_6017, w_088_6019, w_088_6020, w_088_6021, w_088_6027, w_088_6031, w_088_6036, w_088_6037, w_088_6038, w_088_6040, w_088_6046, w_088_6049, w_088_6052, w_088_6054, w_088_6055, w_088_6056, w_088_6058, w_088_6059, w_088_6060, w_088_6070, w_088_6072, w_088_6073, w_088_6077, w_088_6079, w_088_6086, w_088_6089, w_088_6090, w_088_6097, w_088_6098, w_088_6101, w_088_6107, w_088_6115, w_088_6118, w_088_6125, w_088_6133, w_088_6135, w_088_6136, w_088_6141, w_088_6142, w_088_6146, w_088_6149, w_088_6151, w_088_6152, w_088_6157, w_088_6158, w_088_6159, w_088_6160, w_088_6161, w_088_6162, w_088_6165, w_088_6168, w_088_6190, w_088_6198, w_088_6202, w_088_6209, w_088_6213, w_088_6215, w_088_6217, w_088_6222, w_088_6224, w_088_6225, w_088_6228, w_088_6230, w_088_6243, w_088_6247, w_088_6250, w_088_6253, w_088_6259, w_088_6271, w_088_6273, w_088_6276, w_088_6277, w_088_6289, w_088_6296, w_088_6298, w_088_6300, w_088_6313, w_088_6319, w_088_6322, w_088_6329, w_088_6334, w_088_6337, w_088_6340, w_088_6347, w_088_6349, w_088_6350, w_088_6358, w_088_6360, w_088_6361, w_088_6377, w_088_6378, w_088_6384, w_088_6385, w_088_6392, w_088_6397, w_088_6399, w_088_6405, w_088_6407, w_088_6409, w_088_6415, w_088_6417, w_088_6422, w_088_6424, w_088_6426, w_088_6430, w_088_6434, w_088_6438, w_088_6439, w_088_6441, w_088_6442, w_088_6452, w_088_6453, w_088_6454, w_088_6461, w_088_6464, w_088_6466, w_088_6477, w_088_6487, w_088_6490, w_088_6495, w_088_6496, w_088_6499, w_088_6504, w_088_6505, w_088_6508, w_088_6518, w_088_6528, w_088_6533, w_088_6535, w_088_6536, w_088_6537, w_088_6545, w_088_6547, w_088_6548, w_088_6549, w_088_6556, w_088_6557, w_088_6569, w_088_6571, w_088_6574, w_088_6575, w_088_6578, w_088_6580, w_088_6592, w_088_6596, w_088_6598, w_088_6605, w_088_6613, w_088_6614, w_088_6621, w_088_6631, w_088_6633, w_088_6634, w_088_6636, w_088_6639, w_088_6642, w_088_6644, w_088_6646, w_088_6650, w_088_6651, w_088_6657, w_088_6658, w_088_6661, w_088_6662, w_088_6663, w_088_6672, w_088_6681, w_088_6686, w_088_6687, w_088_6690, w_088_6696, w_088_6697, w_088_6704, w_088_6705, w_088_6708, w_088_6711, w_088_6723, w_088_6726, w_088_6728, w_088_6735, w_088_6743, w_088_6744, w_088_6757, w_088_6759, w_088_6763, w_088_6766, w_088_6771, w_088_6775, w_088_6779, w_088_6786, w_088_6788, w_088_6792, w_088_6797, w_088_6801, w_088_6814, w_088_6817, w_088_6820, w_088_6825, w_088_6826, w_088_6829, w_088_6833, w_088_6835, w_088_6837, w_088_6838, w_088_6839, w_088_6849, w_088_6852, w_088_6862, w_088_6866, w_088_6871, w_088_6874, w_088_6876, w_088_6881, w_088_6884, w_088_6891, w_088_6897, w_088_6899, w_088_6905, w_088_6912, w_088_6913, w_088_6914, w_088_6915, w_088_6931, w_088_6940, w_088_6946, w_088_6952, w_088_6954, w_088_6955, w_088_6958, w_088_6964, w_088_6968, w_088_6975, w_088_6979, w_088_6981, w_088_6983, w_088_6984, w_088_6986, w_088_6988, w_088_6994, w_088_6999, w_088_7004, w_088_7008, w_088_7010, w_088_7012, w_088_7023, w_088_7024, w_088_7027, w_088_7034, w_088_7036, w_088_7039, w_088_7040, w_088_7042, w_088_7043, w_088_7046, w_088_7050, w_088_7057, w_088_7059, w_088_7066, w_088_7068, w_088_7078, w_088_7083, w_088_7086, w_088_7092, w_088_7093, w_088_7096, w_088_7098, w_088_7099, w_088_7107, w_088_7113, w_088_7119, w_088_7132, w_088_7135, w_088_7137, w_088_7141, w_088_7143, w_088_7146, w_088_7154, w_088_7159, w_088_7160, w_088_7161, w_088_7168, w_088_7176, w_088_7179, w_088_7182, w_088_7188, w_088_7194, w_088_7208, w_088_7210, w_088_7211, w_088_7213, w_088_7218, w_088_7219, w_088_7224, w_088_7230, w_088_7242, w_088_7243, w_088_7248, w_088_7249, w_088_7252, w_088_7253, w_088_7256, w_088_7259, w_088_7260, w_088_7266, w_088_7271, w_088_7273, w_088_7278, w_088_7279, w_088_7281, w_088_7283, w_088_7288, w_088_7289, w_088_7308, w_088_7310, w_088_7312, w_088_7319, w_088_7323, w_088_7324, w_088_7329, w_088_7337, w_088_7338, w_088_7343, w_088_7344, w_088_7352, w_088_7353, w_088_7355, w_088_7362, w_088_7363, w_088_7364, w_088_7366, w_088_7372, w_088_7373, w_088_7377, w_088_7379, w_088_7383, w_088_7389, w_088_7393, w_088_7394, w_088_7397, w_088_7399, w_088_7400, w_088_7404, w_088_7408, w_088_7411, w_088_7412, w_088_7413, w_088_7417, w_088_7419, w_088_7429, w_088_7431, w_088_7434, w_088_7435, w_088_7438, w_088_7442, w_088_7443, w_088_7444, w_088_7447, w_088_7452, w_088_7460, w_088_7466, w_088_7471, w_088_7474, w_088_7476, w_088_7481, w_088_7482, w_088_7483, w_088_7486, w_088_7487, w_088_7491, w_088_7495, w_088_7498, w_088_7500, w_088_7502, w_088_7505, w_088_7508, w_088_7510, w_088_7511, w_088_7513, w_088_7521, w_088_7522, w_088_7524, w_088_7527, w_088_7530, w_088_7532, w_088_7543, w_088_7545, w_088_7546, w_088_7552, w_088_7553, w_088_7556, w_088_7558, w_088_7560, w_088_7563, w_088_7584, w_088_7585, w_088_7588, w_088_7589, w_088_7590, w_088_7606, w_088_7609, w_088_7612, w_088_7613, w_088_7619, w_088_7620, w_088_7622, w_088_7624, w_088_7629, w_088_7633, w_088_7639, w_088_7652, w_088_7661, w_088_7666, w_088_7667, w_088_7677, w_088_7680, w_088_7681, w_088_7682, w_088_7687, w_088_7692, w_088_7703, w_088_7705, w_088_7712, w_088_7716, w_088_7724, w_088_7727, w_088_7731, w_088_7732, w_088_7735, w_088_7738, w_088_7743, w_088_7745, w_088_7747, w_088_7748, w_088_7750, w_088_7751, w_088_7752, w_088_7759, w_088_7760, w_088_7761, w_088_7765, w_088_7767, w_088_7770, w_088_7771, w_088_7772, w_088_7773, w_088_7775, w_088_7776, w_088_7777, w_088_7781, w_088_7782, w_088_7783, w_088_7788, w_088_7793, w_088_7794, w_088_7796, w_088_7797, w_088_7810, w_088_7814, w_088_7817, w_088_7822, w_088_7823, w_088_7824, w_088_7828, w_088_7831, w_088_7850, w_088_7853, w_088_7854, w_088_7862, w_088_7863, w_088_7869, w_088_7872, w_088_7873, w_088_7883, w_088_7888, w_088_7890, w_088_7892, w_088_7893, w_088_7896, w_088_7901, w_088_7902, w_088_7915, w_088_7921, w_088_7923, w_088_7925, w_088_7929, w_088_7940, w_088_7946, w_088_7948, w_088_7954, w_088_7955, w_088_7956, w_088_7957, w_088_7958, w_088_7959, w_088_7962, w_088_7965, w_088_7970, w_088_7971, w_088_7978, w_088_7983, w_088_7985, w_088_7987, w_088_7991, w_088_8000, w_088_8006, w_088_8010, w_088_8018, w_088_8022, w_088_8025, w_088_8026, w_088_8031, w_088_8037, w_088_8039, w_088_8049, w_088_8050, w_088_8059, w_088_8061, w_088_8064, w_088_8065, w_088_8067, w_088_8068, w_088_8070, w_088_8086, w_088_8087, w_088_8093, w_088_8094, w_088_8095, w_088_8113, w_088_8114, w_088_8118, w_088_8120, w_088_8125, w_088_8126, w_088_8128, w_088_8130, w_088_8136, w_088_8146, w_088_8151, w_088_8154, w_088_8164, w_088_8169, w_088_8170, w_088_8182, w_088_8183, w_088_8184, w_088_8185, w_088_8194, w_088_8195, w_088_8197, w_088_8198, w_088_8204, w_088_8210, w_088_8213, w_088_8217, w_088_8220;
  wire w_089_000, w_089_001, w_089_002, w_089_003, w_089_004, w_089_006, w_089_008, w_089_009, w_089_011, w_089_013, w_089_014, w_089_015, w_089_016, w_089_017, w_089_018, w_089_020, w_089_021, w_089_022, w_089_023, w_089_026, w_089_027, w_089_028, w_089_029, w_089_030, w_089_031, w_089_032, w_089_033, w_089_034, w_089_035, w_089_036, w_089_037, w_089_038, w_089_039, w_089_040, w_089_042, w_089_043, w_089_046, w_089_048, w_089_049, w_089_052, w_089_054, w_089_056, w_089_057, w_089_058, w_089_059, w_089_060, w_089_061, w_089_063, w_089_064, w_089_066, w_089_067, w_089_068, w_089_069, w_089_071, w_089_072, w_089_073, w_089_074, w_089_076, w_089_077, w_089_082, w_089_083, w_089_087, w_089_090, w_089_091, w_089_092, w_089_093, w_089_094, w_089_095, w_089_096, w_089_098, w_089_101, w_089_102, w_089_104, w_089_105, w_089_106, w_089_107, w_089_108, w_089_109, w_089_110, w_089_111, w_089_112, w_089_113, w_089_116, w_089_117, w_089_118, w_089_119, w_089_120, w_089_121, w_089_122, w_089_123, w_089_125, w_089_126, w_089_127, w_089_128, w_089_129, w_089_130, w_089_131, w_089_132, w_089_133, w_089_134, w_089_135, w_089_136, w_089_137, w_089_138, w_089_139, w_089_141, w_089_142, w_089_143, w_089_144, w_089_145, w_089_146, w_089_147, w_089_148, w_089_149, w_089_150, w_089_151, w_089_154, w_089_155, w_089_156, w_089_157, w_089_158, w_089_159, w_089_163, w_089_166, w_089_167, w_089_168, w_089_170, w_089_171, w_089_172, w_089_173, w_089_175, w_089_176, w_089_177, w_089_178, w_089_179, w_089_180, w_089_181, w_089_182, w_089_183, w_089_185, w_089_186, w_089_187, w_089_188, w_089_189, w_089_190, w_089_191, w_089_193, w_089_194, w_089_195, w_089_196, w_089_197, w_089_198, w_089_199, w_089_200, w_089_201, w_089_203, w_089_205, w_089_206, w_089_207, w_089_208, w_089_209, w_089_210, w_089_212, w_089_213, w_089_215, w_089_217, w_089_218, w_089_220, w_089_223, w_089_224, w_089_225, w_089_226, w_089_227, w_089_228, w_089_229, w_089_230, w_089_231, w_089_232, w_089_234, w_089_235, w_089_239, w_089_240, w_089_242, w_089_245, w_089_246, w_089_247, w_089_249, w_089_250, w_089_251, w_089_252, w_089_253, w_089_255, w_089_256, w_089_257, w_089_258, w_089_259, w_089_263, w_089_264, w_089_265, w_089_267, w_089_268, w_089_269, w_089_270, w_089_271, w_089_272, w_089_275, w_089_276, w_089_278, w_089_279, w_089_280, w_089_281, w_089_282, w_089_286, w_089_287, w_089_288, w_089_290, w_089_291, w_089_292, w_089_293, w_089_294, w_089_295, w_089_296, w_089_297, w_089_298, w_089_299, w_089_300, w_089_301, w_089_302, w_089_304, w_089_306, w_089_307, w_089_308, w_089_310, w_089_311, w_089_312, w_089_313, w_089_314, w_089_315, w_089_317, w_089_318, w_089_320, w_089_321, w_089_323, w_089_324, w_089_325, w_089_326, w_089_327, w_089_329, w_089_330, w_089_331, w_089_333, w_089_334, w_089_335, w_089_336, w_089_337, w_089_338, w_089_340, w_089_342, w_089_344, w_089_345, w_089_347, w_089_348, w_089_349, w_089_350, w_089_352, w_089_353, w_089_354, w_089_355, w_089_357, w_089_358, w_089_360, w_089_361, w_089_363, w_089_364, w_089_366, w_089_367, w_089_370, w_089_373, w_089_375, w_089_376, w_089_377, w_089_378, w_089_379, w_089_380, w_089_381, w_089_382, w_089_383, w_089_384, w_089_385, w_089_386, w_089_387, w_089_389, w_089_390, w_089_392, w_089_393, w_089_394, w_089_395, w_089_396, w_089_398, w_089_399, w_089_401, w_089_402, w_089_403, w_089_404, w_089_405, w_089_406, w_089_408, w_089_410, w_089_411, w_089_412, w_089_413, w_089_416, w_089_418, w_089_421, w_089_422, w_089_423, w_089_424, w_089_425, w_089_426, w_089_427, w_089_429, w_089_430, w_089_432, w_089_433, w_089_434, w_089_435, w_089_436, w_089_437, w_089_438, w_089_439, w_089_440, w_089_441, w_089_442, w_089_443, w_089_446, w_089_447, w_089_448, w_089_449, w_089_452, w_089_453, w_089_454, w_089_455, w_089_458, w_089_459, w_089_460, w_089_461, w_089_462, w_089_463, w_089_465, w_089_466, w_089_467, w_089_468, w_089_469, w_089_470, w_089_471, w_089_472, w_089_473, w_089_476, w_089_479, w_089_480, w_089_481, w_089_482, w_089_484, w_089_485, w_089_486, w_089_487, w_089_488, w_089_490, w_089_492, w_089_493, w_089_494, w_089_495, w_089_496, w_089_497, w_089_499, w_089_500, w_089_502, w_089_503, w_089_504, w_089_505, w_089_508, w_089_509, w_089_510, w_089_512, w_089_514, w_089_515, w_089_517, w_089_518, w_089_519, w_089_520, w_089_521, w_089_522, w_089_523, w_089_525, w_089_526, w_089_527, w_089_528, w_089_530, w_089_531, w_089_532, w_089_533, w_089_534, w_089_535, w_089_536, w_089_537, w_089_538, w_089_542, w_089_543, w_089_544, w_089_545, w_089_546, w_089_547, w_089_548, w_089_549, w_089_550, w_089_551, w_089_552, w_089_554, w_089_555, w_089_556, w_089_557, w_089_559, w_089_560, w_089_561, w_089_562, w_089_563, w_089_565, w_089_566, w_089_567, w_089_568, w_089_570, w_089_571, w_089_572, w_089_573, w_089_575, w_089_576, w_089_578, w_089_579, w_089_580, w_089_581, w_089_582, w_089_583, w_089_585, w_089_586, w_089_589, w_089_590, w_089_591, w_089_592, w_089_596, w_089_597, w_089_598, w_089_600, w_089_601, w_089_602, w_089_605, w_089_606, w_089_607, w_089_608, w_089_609, w_089_611, w_089_612, w_089_613, w_089_617, w_089_619, w_089_621, w_089_623, w_089_624, w_089_628, w_089_629, w_089_630, w_089_632, w_089_634, w_089_635, w_089_637, w_089_639, w_089_642, w_089_645, w_089_647, w_089_648, w_089_649, w_089_650, w_089_651, w_089_652, w_089_653, w_089_654, w_089_655, w_089_656, w_089_657, w_089_658, w_089_659, w_089_660, w_089_662, w_089_666, w_089_667, w_089_669, w_089_670, w_089_671, w_089_672, w_089_674, w_089_677, w_089_678, w_089_680, w_089_681, w_089_682, w_089_684, w_089_685, w_089_686, w_089_689, w_089_690, w_089_691, w_089_694, w_089_695, w_089_696, w_089_697, w_089_698, w_089_699, w_089_701, w_089_702, w_089_703, w_089_704, w_089_705, w_089_706, w_089_707, w_089_708, w_089_709, w_089_710, w_089_711, w_089_713, w_089_714, w_089_715, w_089_716, w_089_717, w_089_718, w_089_719, w_089_721, w_089_722, w_089_723, w_089_724, w_089_725, w_089_727, w_089_728, w_089_729, w_089_730, w_089_733, w_089_734, w_089_735, w_089_736, w_089_737, w_089_738, w_089_739, w_089_740, w_089_741, w_089_744, w_089_745, w_089_746, w_089_748, w_089_749, w_089_750, w_089_751, w_089_752, w_089_753, w_089_754, w_089_755, w_089_756, w_089_757, w_089_758, w_089_759, w_089_760, w_089_761, w_089_762, w_089_763, w_089_764, w_089_765, w_089_766, w_089_767, w_089_770, w_089_772, w_089_773, w_089_774, w_089_775, w_089_776, w_089_777, w_089_778, w_089_779, w_089_780, w_089_781, w_089_782, w_089_783, w_089_784, w_089_785, w_089_786, w_089_787, w_089_788, w_089_789, w_089_790, w_089_791, w_089_793, w_089_794, w_089_795, w_089_796, w_089_797, w_089_798, w_089_799, w_089_802, w_089_803, w_089_804, w_089_805, w_089_806, w_089_807, w_089_808, w_089_809, w_089_810, w_089_811, w_089_813, w_089_815, w_089_816, w_089_818, w_089_820, w_089_821, w_089_822, w_089_823, w_089_824, w_089_825, w_089_828, w_089_829, w_089_831, w_089_832, w_089_833, w_089_834, w_089_837, w_089_838, w_089_839, w_089_840, w_089_841, w_089_842, w_089_843, w_089_844, w_089_845, w_089_846, w_089_847, w_089_849, w_089_850, w_089_851, w_089_852, w_089_854, w_089_855, w_089_856, w_089_858, w_089_859, w_089_861, w_089_862, w_089_865, w_089_866, w_089_867, w_089_868, w_089_869, w_089_871, w_089_872, w_089_873, w_089_874, w_089_876, w_089_877, w_089_878, w_089_880, w_089_881, w_089_882, w_089_883, w_089_884, w_089_885, w_089_886, w_089_887, w_089_889, w_089_890, w_089_891, w_089_892, w_089_893, w_089_895, w_089_897, w_089_898, w_089_899, w_089_902, w_089_903, w_089_904, w_089_906, w_089_907, w_089_908, w_089_910, w_089_912, w_089_914, w_089_915, w_089_916, w_089_917, w_089_918, w_089_919, w_089_920, w_089_921, w_089_922, w_089_923, w_089_924, w_089_927, w_089_929, w_089_930, w_089_932, w_089_935, w_089_936, w_089_937, w_089_938, w_089_939, w_089_940, w_089_941, w_089_942, w_089_945, w_089_946, w_089_947, w_089_948, w_089_949, w_089_950, w_089_951, w_089_954, w_089_955, w_089_957, w_089_958, w_089_959, w_089_960, w_089_962, w_089_963, w_089_964, w_089_965, w_089_967, w_089_968, w_089_970, w_089_971, w_089_972, w_089_973, w_089_974, w_089_976, w_089_977, w_089_979, w_089_980, w_089_981, w_089_984, w_089_986, w_089_987, w_089_988, w_089_990, w_089_992, w_089_993, w_089_994, w_089_995, w_089_996, w_089_997, w_089_999, w_089_1000, w_089_1001, w_089_1003, w_089_1004, w_089_1006, w_089_1009, w_089_1011, w_089_1012, w_089_1013, w_089_1014, w_089_1015, w_089_1016, w_089_1017, w_089_1018, w_089_1019, w_089_1020, w_089_1021, w_089_1022, w_089_1023, w_089_1024, w_089_1026, w_089_1027, w_089_1028, w_089_1030, w_089_1031, w_089_1033, w_089_1035, w_089_1036, w_089_1037, w_089_1038, w_089_1039, w_089_1042, w_089_1043, w_089_1044, w_089_1047, w_089_1048, w_089_1049, w_089_1050, w_089_1051, w_089_1052, w_089_1053, w_089_1055, w_089_1056, w_089_1058, w_089_1059, w_089_1060, w_089_1062, w_089_1063, w_089_1064, w_089_1065, w_089_1066, w_089_1067, w_089_1068, w_089_1069, w_089_1070, w_089_1071, w_089_1072, w_089_1075, w_089_1076, w_089_1077, w_089_1079, w_089_1080, w_089_1081, w_089_1082, w_089_1086, w_089_1087, w_089_1090, w_089_1092, w_089_1095, w_089_1096, w_089_1097, w_089_1098, w_089_1099, w_089_1101, w_089_1102, w_089_1104, w_089_1105, w_089_1106, w_089_1109, w_089_1110, w_089_1111, w_089_1112, w_089_1113, w_089_1114, w_089_1117, w_089_1118, w_089_1120, w_089_1122, w_089_1123, w_089_1124, w_089_1125, w_089_1127, w_089_1128, w_089_1129, w_089_1130, w_089_1131, w_089_1132, w_089_1133, w_089_1135, w_089_1136, w_089_1137, w_089_1138, w_089_1139, w_089_1142, w_089_1147, w_089_1149, w_089_1150, w_089_1153, w_089_1155, w_089_1159, w_089_1160, w_089_1162, w_089_1163, w_089_1164, w_089_1165, w_089_1166, w_089_1169, w_089_1171, w_089_1173, w_089_1174, w_089_1175, w_089_1176, w_089_1178, w_089_1179, w_089_1180, w_089_1181, w_089_1183, w_089_1184, w_089_1186, w_089_1187, w_089_1188, w_089_1189, w_089_1191, w_089_1192, w_089_1193, w_089_1194, w_089_1197, w_089_1198, w_089_1199, w_089_1201, w_089_1203, w_089_1204, w_089_1205, w_089_1206, w_089_1207, w_089_1208, w_089_1210, w_089_1211, w_089_1212, w_089_1214, w_089_1215, w_089_1216, w_089_1217, w_089_1218, w_089_1219, w_089_1222, w_089_1224, w_089_1225, w_089_1226, w_089_1228, w_089_1229, w_089_1231, w_089_1232, w_089_1233, w_089_1234, w_089_1235, w_089_1236, w_089_1237, w_089_1238, w_089_1240, w_089_1241, w_089_1242, w_089_1243, w_089_1244, w_089_1245, w_089_1249, w_089_1250, w_089_1251, w_089_1252, w_089_1253, w_089_1254, w_089_1255, w_089_1256, w_089_1258, w_089_1259, w_089_1260, w_089_1263, w_089_1267, w_089_1269, w_089_1271, w_089_1273, w_089_1274, w_089_1275, w_089_1276, w_089_1277, w_089_1279, w_089_1282, w_089_1283, w_089_1284, w_089_1285, w_089_1287, w_089_1288, w_089_1293, w_089_1294, w_089_1295, w_089_1297, w_089_1300, w_089_1302, w_089_1303, w_089_1307, w_089_1308, w_089_1309, w_089_1310, w_089_1311, w_089_1312, w_089_1313, w_089_1314, w_089_1315, w_089_1316, w_089_1318, w_089_1319, w_089_1320, w_089_1321, w_089_1323, w_089_1326, w_089_1327, w_089_1328, w_089_1329, w_089_1331, w_089_1332, w_089_1333, w_089_1335, w_089_1336, w_089_1337, w_089_1338, w_089_1339, w_089_1340, w_089_1342, w_089_1343, w_089_1347, w_089_1348, w_089_1350, w_089_1352, w_089_1353, w_089_1354, w_089_1355, w_089_1356, w_089_1357, w_089_1361, w_089_1362, w_089_1363, w_089_1364, w_089_1365, w_089_1366, w_089_1368, w_089_1370, w_089_1372, w_089_1374, w_089_1377, w_089_1380, w_089_1381, w_089_1382, w_089_1383, w_089_1385, w_089_1388, w_089_1391, w_089_1392, w_089_1394, w_089_1395, w_089_1397, w_089_1398, w_089_1399, w_089_1402, w_089_1403, w_089_1404, w_089_1405, w_089_1406, w_089_1411, w_089_1412, w_089_1414, w_089_1415, w_089_1416, w_089_1417, w_089_1418, w_089_1420, w_089_1422, w_089_1423, w_089_1424, w_089_1425, w_089_1427, w_089_1428, w_089_1430, w_089_1432, w_089_1433, w_089_1434, w_089_1435, w_089_1436, w_089_1437, w_089_1439, w_089_1440, w_089_1441, w_089_1444, w_089_1445, w_089_1446, w_089_1447, w_089_1448, w_089_1450, w_089_1451, w_089_1452, w_089_1453, w_089_1454, w_089_1455, w_089_1457, w_089_1458, w_089_1459, w_089_1461, w_089_1462, w_089_1463, w_089_1465, w_089_1466, w_089_1468, w_089_1469, w_089_1470, w_089_1473, w_089_1474, w_089_1475, w_089_1477, w_089_1478, w_089_1479, w_089_1481, w_089_1482, w_089_1483, w_089_1484, w_089_1485, w_089_1486, w_089_1489, w_089_1491, w_089_1492, w_089_1493, w_089_1496, w_089_1497, w_089_1498, w_089_1500, w_089_1503, w_089_1504, w_089_1505, w_089_1506, w_089_1507, w_089_1508, w_089_1509, w_089_1510, w_089_1512, w_089_1513, w_089_1514, w_089_1515, w_089_1517, w_089_1519, w_089_1521, w_089_1524, w_089_1525, w_089_1527, w_089_1528, w_089_1529, w_089_1530, w_089_1531, w_089_1532, w_089_1535, w_089_1536, w_089_1537, w_089_1538, w_089_1540, w_089_1542, w_089_1543, w_089_1545, w_089_1546, w_089_1547, w_089_1548, w_089_1549, w_089_1550, w_089_1553, w_089_1555, w_089_1556, w_089_1558, w_089_1560, w_089_1561, w_089_1562, w_089_1564, w_089_1565, w_089_1566, w_089_1568, w_089_1571, w_089_1572, w_089_1573, w_089_1577, w_089_1580, w_089_1582, w_089_1583, w_089_1585, w_089_1586, w_089_1587, w_089_1588, w_089_1589, w_089_1591, w_089_1592, w_089_1593, w_089_1594, w_089_1597, w_089_1598, w_089_1599, w_089_1600, w_089_1601, w_089_1602, w_089_1603, w_089_1604, w_089_1605, w_089_1606, w_089_1608, w_089_1610, w_089_1613, w_089_1614, w_089_1615, w_089_1616, w_089_1617, w_089_1618, w_089_1619, w_089_1620, w_089_1622, w_089_1624, w_089_1626, w_089_1628, w_089_1629, w_089_1630, w_089_1631, w_089_1632, w_089_1634, w_089_1635, w_089_1637, w_089_1638, w_089_1640, w_089_1641, w_089_1642, w_089_1643, w_089_1644, w_089_1645, w_089_1646, w_089_1647, w_089_1649, w_089_1650, w_089_1651, w_089_1652, w_089_1653, w_089_1655, w_089_1659, w_089_1660, w_089_1662, w_089_1663, w_089_1666, w_089_1667, w_089_1668, w_089_1669, w_089_1670, w_089_1671, w_089_1672, w_089_1675, w_089_1676, w_089_1677, w_089_1678, w_089_1680, w_089_1681, w_089_1682, w_089_1684, w_089_1685, w_089_1686, w_089_1687, w_089_1688, w_089_1689, w_089_1692, w_089_1693, w_089_1695, w_089_1696, w_089_1697, w_089_1698, w_089_1699, w_089_1700, w_089_1703, w_089_1705, w_089_1706, w_089_1707, w_089_1709, w_089_1710, w_089_1711, w_089_1714, w_089_1719, w_089_1720, w_089_1721, w_089_1722, w_089_1723, w_089_1724, w_089_1728, w_089_1729, w_089_1730, w_089_1731, w_089_1733, w_089_1734, w_089_1735, w_089_1736, w_089_1737, w_089_1740, w_089_1741, w_089_1743, w_089_1744, w_089_1745, w_089_1746, w_089_1747, w_089_1748, w_089_1750, w_089_1751, w_089_1752, w_089_1753, w_089_1755, w_089_1756, w_089_1757, w_089_1758, w_089_1759, w_089_1761, w_089_1762, w_089_1763, w_089_1767, w_089_1768, w_089_1769, w_089_1771, w_089_1772, w_089_1773, w_089_1774, w_089_1778, w_089_1779, w_089_1780, w_089_1782, w_089_1783, w_089_1785, w_089_1786, w_089_1788, w_089_1789, w_089_1790, w_089_1791, w_089_1792, w_089_1793, w_089_1794, w_089_1795, w_089_1798, w_089_1803, w_089_1804, w_089_1805, w_089_1807, w_089_1810, w_089_1811, w_089_1812, w_089_1813, w_089_1816, w_089_1817, w_089_1818, w_089_1819, w_089_1820, w_089_1821, w_089_1823, w_089_1824, w_089_1826, w_089_1828, w_089_1829, w_089_1830, w_089_1831, w_089_1832, w_089_1833, w_089_1836, w_089_1838, w_089_1839, w_089_1840, w_089_1842, w_089_1843, w_089_1844, w_089_1845, w_089_1847, w_089_1848, w_089_1849, w_089_1850, w_089_1851, w_089_1852, w_089_1853, w_089_1854, w_089_1855, w_089_1856, w_089_1857, w_089_1860, w_089_1861, w_089_1862, w_089_1864, w_089_1866, w_089_1869, w_089_1870, w_089_1871, w_089_1872, w_089_1873, w_089_1874, w_089_1876, w_089_1877, w_089_1878, w_089_1880, w_089_1883, w_089_1884, w_089_1885, w_089_1887, w_089_1889, w_089_1890, w_089_1892, w_089_1893, w_089_1894, w_089_1895, w_089_1896, w_089_1899, w_089_1900, w_089_1901, w_089_1903, w_089_1904, w_089_1906, w_089_1907, w_089_1910, w_089_1911, w_089_1912, w_089_1913, w_089_1914, w_089_1915, w_089_1916, w_089_1917, w_089_1918, w_089_1919, w_089_1920, w_089_1921, w_089_1923, w_089_1925, w_089_1928, w_089_1929, w_089_1930, w_089_1931, w_089_1932, w_089_1934, w_089_1935, w_089_1937, w_089_1939, w_089_1940, w_089_1941, w_089_1942, w_089_1943, w_089_1944, w_089_1945, w_089_1946, w_089_1947, w_089_1948, w_089_1953, w_089_1955, w_089_1957, w_089_1958, w_089_1959, w_089_1960, w_089_1961, w_089_1963, w_089_1964, w_089_1965, w_089_1967, w_089_1968, w_089_1969, w_089_1970, w_089_1971, w_089_1973, w_089_1975, w_089_1977, w_089_1978, w_089_1979, w_089_1981, w_089_1985, w_089_1988, w_089_1989, w_089_1990, w_089_1991, w_089_1992, w_089_1993, w_089_1994, w_089_1995, w_089_1997, w_089_1999, w_089_2000, w_089_2001, w_089_2002, w_089_2004, w_089_2006, w_089_2009, w_089_2012, w_089_2015, w_089_2018, w_089_2019, w_089_2020, w_089_2021, w_089_2022, w_089_2023, w_089_2025, w_089_2026, w_089_2029, w_089_2030, w_089_2031, w_089_2032, w_089_2033, w_089_2034, w_089_2036, w_089_2037, w_089_2039, w_089_2040, w_089_2043, w_089_2044, w_089_2046, w_089_2047, w_089_2048, w_089_2049, w_089_2050, w_089_2051, w_089_2052, w_089_2053, w_089_2054, w_089_2055, w_089_2056, w_089_2057, w_089_2058, w_089_2059, w_089_2060, w_089_2061, w_089_2062, w_089_2063, w_089_2065, w_089_2066, w_089_2067, w_089_2069, w_089_2071, w_089_2072, w_089_2074, w_089_2075, w_089_2077, w_089_2078, w_089_2079, w_089_2080, w_089_2082, w_089_2083, w_089_2084, w_089_2085, w_089_2086, w_089_2087, w_089_2088, w_089_2090, w_089_2092, w_089_2093, w_089_2096, w_089_2097, w_089_2098, w_089_2100, w_089_2101, w_089_2102, w_089_2103, w_089_2105, w_089_2106, w_089_2107, w_089_2108, w_089_2109, w_089_2110, w_089_2111, w_089_2114, w_089_2115, w_089_2117, w_089_2119, w_089_2121, w_089_2122, w_089_2124, w_089_2125, w_089_2126, w_089_2128, w_089_2129, w_089_2130, w_089_2131, w_089_2132, w_089_2134, w_089_2135, w_089_2136, w_089_2137, w_089_2138, w_089_2139, w_089_2140, w_089_2142, w_089_2143, w_089_2146, w_089_2147, w_089_2148, w_089_2149, w_089_2151, w_089_2152, w_089_2153, w_089_2157, w_089_2158, w_089_2159, w_089_2161, w_089_2162, w_089_2163, w_089_2164, w_089_2167, w_089_2168, w_089_2169, w_089_2170, w_089_2171, w_089_2172, w_089_2175, w_089_2176, w_089_2178, w_089_2179, w_089_2180, w_089_2181, w_089_2183, w_089_2186, w_089_2187, w_089_2188, w_089_2189, w_089_2190, w_089_2193, w_089_2194, w_089_2195, w_089_2197, w_089_2198, w_089_2199, w_089_2200, w_089_2202, w_089_2205, w_089_2207, w_089_2210, w_089_2211, w_089_2212, w_089_2213, w_089_2214, w_089_2215, w_089_2216, w_089_2217, w_089_2218, w_089_2219, w_089_2220, w_089_2222, w_089_2223, w_089_2224, w_089_2226, w_089_2227, w_089_2230, w_089_2231, w_089_2232, w_089_2233, w_089_2234, w_089_2236, w_089_2237, w_089_2239, w_089_2240, w_089_2241, w_089_2242, w_089_2243, w_089_2245, w_089_2248, w_089_2251, w_089_2252, w_089_2253, w_089_2257, w_089_2259, w_089_2261, w_089_2266;
  wire w_090_001, w_090_003, w_090_004, w_090_005, w_090_006, w_090_007, w_090_008, w_090_010, w_090_012, w_090_015, w_090_020, w_090_021, w_090_022, w_090_023, w_090_024, w_090_026, w_090_030, w_090_032, w_090_033, w_090_034, w_090_035, w_090_036, w_090_038, w_090_040, w_090_043, w_090_044, w_090_045, w_090_046, w_090_047, w_090_048, w_090_049, w_090_050, w_090_051, w_090_052, w_090_053, w_090_054, w_090_056, w_090_057, w_090_059, w_090_060, w_090_061, w_090_063, w_090_064, w_090_065, w_090_066, w_090_074, w_090_075, w_090_076, w_090_077, w_090_078, w_090_079, w_090_080, w_090_081, w_090_082, w_090_083, w_090_084, w_090_086, w_090_087, w_090_088, w_090_090, w_090_092, w_090_093, w_090_094, w_090_096, w_090_097, w_090_099, w_090_101, w_090_103, w_090_107, w_090_108, w_090_110, w_090_111, w_090_112, w_090_114, w_090_115, w_090_117, w_090_125, w_090_128, w_090_129, w_090_130, w_090_132, w_090_134, w_090_136, w_090_138, w_090_139, w_090_140, w_090_144, w_090_145, w_090_148, w_090_149, w_090_150, w_090_151, w_090_153, w_090_157, w_090_158, w_090_160, w_090_161, w_090_164, w_090_165, w_090_167, w_090_168, w_090_170, w_090_172, w_090_174, w_090_177, w_090_179, w_090_182, w_090_183, w_090_184, w_090_187, w_090_193, w_090_195, w_090_196, w_090_200, w_090_201, w_090_205, w_090_206, w_090_207, w_090_209, w_090_214, w_090_215, w_090_218, w_090_219, w_090_220, w_090_224, w_090_225, w_090_227, w_090_228, w_090_230, w_090_231, w_090_232, w_090_233, w_090_238, w_090_239, w_090_242, w_090_244, w_090_246, w_090_247, w_090_248, w_090_249, w_090_250, w_090_252, w_090_253, w_090_254, w_090_257, w_090_258, w_090_259, w_090_262, w_090_263, w_090_265, w_090_267, w_090_268, w_090_271, w_090_272, w_090_273, w_090_274, w_090_275, w_090_276, w_090_279, w_090_280, w_090_281, w_090_282, w_090_283, w_090_284, w_090_285, w_090_287, w_090_288, w_090_290, w_090_291, w_090_292, w_090_293, w_090_295, w_090_296, w_090_298, w_090_299, w_090_300, w_090_301, w_090_302, w_090_303, w_090_304, w_090_306, w_090_307, w_090_309, w_090_311, w_090_315, w_090_316, w_090_318, w_090_321, w_090_325, w_090_326, w_090_327, w_090_328, w_090_329, w_090_330, w_090_331, w_090_332, w_090_334, w_090_336, w_090_337, w_090_338, w_090_339, w_090_343, w_090_344, w_090_346, w_090_348, w_090_351, w_090_352, w_090_353, w_090_354, w_090_358, w_090_363, w_090_365, w_090_367, w_090_368, w_090_370, w_090_371, w_090_373, w_090_374, w_090_375, w_090_376, w_090_377, w_090_378, w_090_380, w_090_382, w_090_383, w_090_386, w_090_387, w_090_389, w_090_392, w_090_396, w_090_398, w_090_400, w_090_401, w_090_405, w_090_407, w_090_409, w_090_411, w_090_412, w_090_415, w_090_416, w_090_419, w_090_420, w_090_421, w_090_424, w_090_425, w_090_426, w_090_427, w_090_428, w_090_429, w_090_432, w_090_433, w_090_434, w_090_436, w_090_438, w_090_439, w_090_441, w_090_442, w_090_445, w_090_447, w_090_448, w_090_450, w_090_451, w_090_452, w_090_453, w_090_454, w_090_455, w_090_460, w_090_461, w_090_462, w_090_464, w_090_465, w_090_466, w_090_467, w_090_468, w_090_469, w_090_471, w_090_474, w_090_475, w_090_476, w_090_478, w_090_479, w_090_480, w_090_482, w_090_484, w_090_485, w_090_486, w_090_487, w_090_488, w_090_489, w_090_490, w_090_491, w_090_493, w_090_495, w_090_496, w_090_499, w_090_500, w_090_501, w_090_502, w_090_503, w_090_504, w_090_505, w_090_506, w_090_507, w_090_508, w_090_509, w_090_510, w_090_511, w_090_513, w_090_517, w_090_519, w_090_520, w_090_522, w_090_524, w_090_525, w_090_528, w_090_529, w_090_531, w_090_532, w_090_533, w_090_534, w_090_537, w_090_538, w_090_539, w_090_542, w_090_544, w_090_545, w_090_547, w_090_548, w_090_549, w_090_551, w_090_556, w_090_557, w_090_558, w_090_559, w_090_562, w_090_564, w_090_565, w_090_566, w_090_569, w_090_571, w_090_572, w_090_573, w_090_574, w_090_575, w_090_577, w_090_578, w_090_579, w_090_580, w_090_581, w_090_583, w_090_585, w_090_586, w_090_587, w_090_588, w_090_589, w_090_590, w_090_591, w_090_592, w_090_594, w_090_596, w_090_597, w_090_599, w_090_600, w_090_601, w_090_602, w_090_604, w_090_605, w_090_607, w_090_608, w_090_610, w_090_613, w_090_617, w_090_620, w_090_625, w_090_626, w_090_627, w_090_628, w_090_629, w_090_630, w_090_631, w_090_633, w_090_636, w_090_637, w_090_638, w_090_639, w_090_641, w_090_643, w_090_645, w_090_647, w_090_649, w_090_655, w_090_656, w_090_659, w_090_660, w_090_662, w_090_665, w_090_667, w_090_668, w_090_670, w_090_671, w_090_672, w_090_674, w_090_675, w_090_676, w_090_677, w_090_679, w_090_680, w_090_682, w_090_683, w_090_684, w_090_687, w_090_688, w_090_692, w_090_696, w_090_697, w_090_699, w_090_705, w_090_710, w_090_711, w_090_712, w_090_713, w_090_715, w_090_716, w_090_717, w_090_720, w_090_721, w_090_724, w_090_725, w_090_728, w_090_732, w_090_734, w_090_735, w_090_739, w_090_740, w_090_742, w_090_744, w_090_746, w_090_748, w_090_749, w_090_750, w_090_751, w_090_752, w_090_753, w_090_756, w_090_758, w_090_759, w_090_761, w_090_762, w_090_763, w_090_764, w_090_768, w_090_770, w_090_771, w_090_775, w_090_778, w_090_781, w_090_782, w_090_785, w_090_786, w_090_787, w_090_790, w_090_791, w_090_792, w_090_793, w_090_794, w_090_795, w_090_798, w_090_799, w_090_801, w_090_805, w_090_806, w_090_807, w_090_808, w_090_811, w_090_813, w_090_816, w_090_817, w_090_818, w_090_819, w_090_822, w_090_824, w_090_825, w_090_827, w_090_828, w_090_829, w_090_830, w_090_831, w_090_833, w_090_834, w_090_835, w_090_836, w_090_839, w_090_841, w_090_842, w_090_844, w_090_847, w_090_850, w_090_852, w_090_855, w_090_856, w_090_857, w_090_859, w_090_860, w_090_861, w_090_864, w_090_866, w_090_867, w_090_868, w_090_869, w_090_871, w_090_872, w_090_875, w_090_877, w_090_878, w_090_880, w_090_881, w_090_884, w_090_886, w_090_887, w_090_888, w_090_890, w_090_894, w_090_895, w_090_897, w_090_899, w_090_901, w_090_902, w_090_903, w_090_904, w_090_906, w_090_907, w_090_908, w_090_909, w_090_911, w_090_912, w_090_913, w_090_914, w_090_915, w_090_916, w_090_917, w_090_920, w_090_922, w_090_923, w_090_924, w_090_927, w_090_928, w_090_929, w_090_930, w_090_931, w_090_933, w_090_934, w_090_935, w_090_937, w_090_939, w_090_942, w_090_944, w_090_945, w_090_946, w_090_948, w_090_949, w_090_950, w_090_953, w_090_955, w_090_957, w_090_958, w_090_959, w_090_961, w_090_965, w_090_966, w_090_967, w_090_968, w_090_970, w_090_973, w_090_976, w_090_980, w_090_982, w_090_984, w_090_986, w_090_987, w_090_988, w_090_992, w_090_993, w_090_995, w_090_998, w_090_999, w_090_1002, w_090_1003, w_090_1005, w_090_1006, w_090_1007, w_090_1010, w_090_1011, w_090_1014, w_090_1015, w_090_1016, w_090_1019, w_090_1020, w_090_1021, w_090_1023, w_090_1024, w_090_1026, w_090_1027, w_090_1028, w_090_1029, w_090_1031, w_090_1032, w_090_1033, w_090_1034, w_090_1035, w_090_1038, w_090_1039, w_090_1040, w_090_1041, w_090_1043, w_090_1045, w_090_1046, w_090_1048, w_090_1050, w_090_1051, w_090_1052, w_090_1054, w_090_1056, w_090_1057, w_090_1058, w_090_1059, w_090_1062, w_090_1066, w_090_1069, w_090_1070, w_090_1071, w_090_1072, w_090_1073, w_090_1074, w_090_1076, w_090_1078, w_090_1080, w_090_1082, w_090_1084, w_090_1086, w_090_1088, w_090_1090, w_090_1092, w_090_1093, w_090_1095, w_090_1096, w_090_1097, w_090_1099, w_090_1100, w_090_1102, w_090_1105, w_090_1106, w_090_1107, w_090_1108, w_090_1112, w_090_1114, w_090_1116, w_090_1117, w_090_1118, w_090_1119, w_090_1120, w_090_1121, w_090_1123, w_090_1124, w_090_1126, w_090_1127, w_090_1130, w_090_1133, w_090_1134, w_090_1136, w_090_1137, w_090_1140, w_090_1142, w_090_1143, w_090_1147, w_090_1149, w_090_1150, w_090_1151, w_090_1152, w_090_1153, w_090_1155, w_090_1157, w_090_1160, w_090_1162, w_090_1165, w_090_1166, w_090_1168, w_090_1170, w_090_1173, w_090_1174, w_090_1176, w_090_1178, w_090_1180, w_090_1183, w_090_1186, w_090_1187, w_090_1188, w_090_1190, w_090_1191, w_090_1192, w_090_1194, w_090_1195, w_090_1198, w_090_1199, w_090_1200, w_090_1201, w_090_1203, w_090_1207, w_090_1212, w_090_1213, w_090_1214, w_090_1216, w_090_1217, w_090_1219, w_090_1220, w_090_1223, w_090_1226, w_090_1229, w_090_1230, w_090_1231, w_090_1232, w_090_1234, w_090_1240, w_090_1244, w_090_1246, w_090_1248, w_090_1249, w_090_1251, w_090_1253, w_090_1259, w_090_1260, w_090_1262, w_090_1264, w_090_1267, w_090_1270, w_090_1271, w_090_1275, w_090_1277, w_090_1278, w_090_1283, w_090_1284, w_090_1285, w_090_1286, w_090_1289, w_090_1290, w_090_1292, w_090_1293, w_090_1294, w_090_1295, w_090_1296, w_090_1297, w_090_1299, w_090_1300, w_090_1303, w_090_1305, w_090_1306, w_090_1308, w_090_1309, w_090_1312, w_090_1313, w_090_1315, w_090_1318, w_090_1319, w_090_1325, w_090_1326, w_090_1327, w_090_1329, w_090_1330, w_090_1331, w_090_1332, w_090_1333, w_090_1335, w_090_1336, w_090_1338, w_090_1339, w_090_1340, w_090_1342, w_090_1344, w_090_1346, w_090_1347, w_090_1350, w_090_1351, w_090_1354, w_090_1356, w_090_1357, w_090_1359, w_090_1361, w_090_1362, w_090_1368, w_090_1369, w_090_1370, w_090_1372, w_090_1373, w_090_1375, w_090_1376, w_090_1378, w_090_1380, w_090_1381, w_090_1384, w_090_1386, w_090_1387, w_090_1389, w_090_1390, w_090_1391, w_090_1392, w_090_1393, w_090_1394, w_090_1395, w_090_1398, w_090_1399, w_090_1401, w_090_1403, w_090_1407, w_090_1408, w_090_1411, w_090_1414, w_090_1417, w_090_1420, w_090_1423, w_090_1424, w_090_1426, w_090_1427, w_090_1429, w_090_1430, w_090_1431, w_090_1434, w_090_1438, w_090_1439, w_090_1440, w_090_1441, w_090_1442, w_090_1447, w_090_1449, w_090_1450, w_090_1451, w_090_1452, w_090_1453, w_090_1454, w_090_1456, w_090_1458, w_090_1459, w_090_1460, w_090_1462, w_090_1465, w_090_1466, w_090_1467, w_090_1468, w_090_1469, w_090_1470, w_090_1471, w_090_1472, w_090_1473, w_090_1476, w_090_1478, w_090_1480, w_090_1481, w_090_1482, w_090_1484, w_090_1485, w_090_1486, w_090_1490, w_090_1491, w_090_1493, w_090_1494, w_090_1498, w_090_1500, w_090_1501, w_090_1505, w_090_1506, w_090_1508, w_090_1509, w_090_1512, w_090_1513, w_090_1514, w_090_1516, w_090_1519, w_090_1520, w_090_1521, w_090_1522, w_090_1523, w_090_1525, w_090_1526, w_090_1529, w_090_1530, w_090_1532, w_090_1533, w_090_1538, w_090_1539, w_090_1540, w_090_1542, w_090_1543, w_090_1544, w_090_1546, w_090_1548, w_090_1549, w_090_1550, w_090_1552, w_090_1554, w_090_1555, w_090_1556, w_090_1557, w_090_1558, w_090_1559, w_090_1560, w_090_1561, w_090_1562, w_090_1563, w_090_1564, w_090_1566, w_090_1567, w_090_1568, w_090_1572, w_090_1573, w_090_1575, w_090_1578, w_090_1584, w_090_1587, w_090_1589, w_090_1590, w_090_1591, w_090_1592, w_090_1593, w_090_1596, w_090_1598, w_090_1601, w_090_1602, w_090_1603, w_090_1604, w_090_1605, w_090_1607, w_090_1609, w_090_1610, w_090_1612, w_090_1614, w_090_1618, w_090_1621, w_090_1624, w_090_1626, w_090_1627, w_090_1628, w_090_1629, w_090_1631, w_090_1634, w_090_1635, w_090_1637, w_090_1638, w_090_1639, w_090_1640, w_090_1641, w_090_1642, w_090_1643, w_090_1644, w_090_1645, w_090_1646, w_090_1652, w_090_1653, w_090_1654, w_090_1657, w_090_1659, w_090_1661, w_090_1666, w_090_1668, w_090_1671, w_090_1675, w_090_1677, w_090_1678, w_090_1682, w_090_1683, w_090_1684, w_090_1685, w_090_1687, w_090_1690, w_090_1691, w_090_1692, w_090_1694, w_090_1696, w_090_1697, w_090_1698, w_090_1701, w_090_1702, w_090_1703, w_090_1704, w_090_1706, w_090_1707, w_090_1710, w_090_1712, w_090_1714, w_090_1715, w_090_1716, w_090_1719, w_090_1721, w_090_1722, w_090_1724, w_090_1725, w_090_1726, w_090_1728, w_090_1729, w_090_1730, w_090_1731, w_090_1732, w_090_1735, w_090_1737, w_090_1738, w_090_1740, w_090_1741, w_090_1742, w_090_1743, w_090_1747, w_090_1750, w_090_1752, w_090_1753, w_090_1754, w_090_1755, w_090_1756, w_090_1757, w_090_1758, w_090_1761, w_090_1762, w_090_1763, w_090_1764, w_090_1767, w_090_1769, w_090_1770, w_090_1771, w_090_1772, w_090_1773, w_090_1774, w_090_1775, w_090_1778, w_090_1779, w_090_1780, w_090_1782, w_090_1783, w_090_1784, w_090_1786, w_090_1787, w_090_1788, w_090_1790, w_090_1791, w_090_1793, w_090_1794, w_090_1796, w_090_1797, w_090_1798, w_090_1799, w_090_1800, w_090_1802, w_090_1803, w_090_1807, w_090_1808, w_090_1809, w_090_1810, w_090_1812, w_090_1814, w_090_1817, w_090_1818, w_090_1823, w_090_1824, w_090_1825, w_090_1827, w_090_1831, w_090_1833, w_090_1836, w_090_1837, w_090_1841, w_090_1842, w_090_1844, w_090_1847, w_090_1848, w_090_1849, w_090_1851, w_090_1852, w_090_1853, w_090_1854, w_090_1859, w_090_1862, w_090_1864, w_090_1865, w_090_1866, w_090_1868, w_090_1869, w_090_1870, w_090_1871, w_090_1876, w_090_1878, w_090_1879, w_090_1886, w_090_1887, w_090_1890, w_090_1892, w_090_1893, w_090_1894, w_090_1896, w_090_1897, w_090_1898, w_090_1899, w_090_1900, w_090_1901, w_090_1903, w_090_1906, w_090_1907, w_090_1908, w_090_1909, w_090_1910, w_090_1911, w_090_1912, w_090_1913, w_090_1916, w_090_1917, w_090_1918, w_090_1920, w_090_1921, w_090_1922, w_090_1923, w_090_1924, w_090_1925, w_090_1927, w_090_1928, w_090_1929, w_090_1930, w_090_1931, w_090_1932, w_090_1933, w_090_1935, w_090_1937, w_090_1939, w_090_1941, w_090_1944, w_090_1947, w_090_1948, w_090_1949, w_090_1951, w_090_1952, w_090_1957, w_090_1960, w_090_1964, w_090_1965, w_090_1969, w_090_1970, w_090_1973, w_090_1974, w_090_1975, w_090_1979, w_090_1981, w_090_1983, w_090_1987, w_090_1989, w_090_1990, w_090_1992, w_090_1993, w_090_1995, w_090_1996, w_090_2000, w_090_2001, w_090_2002, w_090_2005, w_090_2007, w_090_2013, w_090_2015, w_090_2018, w_090_2019, w_090_2020, w_090_2022, w_090_2023, w_090_2025, w_090_2026, w_090_2027, w_090_2028, w_090_2029, w_090_2033, w_090_2035, w_090_2038, w_090_2039, w_090_2040, w_090_2041, w_090_2042, w_090_2044, w_090_2045, w_090_2047, w_090_2049, w_090_2050, w_090_2052, w_090_2053, w_090_2054, w_090_2055, w_090_2058, w_090_2060, w_090_2061, w_090_2063, w_090_2065, w_090_2067, w_090_2068, w_090_2070, w_090_2071, w_090_2075, w_090_2076, w_090_2077, w_090_2078, w_090_2080, w_090_2082, w_090_2084, w_090_2087, w_090_2089, w_090_2090, w_090_2091, w_090_2094, w_090_2095, w_090_2096, w_090_2099, w_090_2100, w_090_2102, w_090_2103, w_090_2106, w_090_2107, w_090_2109, w_090_2110, w_090_2111, w_090_2113, w_090_2114, w_090_2118, w_090_2119, w_090_2121, w_090_2122, w_090_2124, w_090_2126, w_090_2130, w_090_2132, w_090_2134, w_090_2135, w_090_2137, w_090_2138, w_090_2140, w_090_2142, w_090_2144, w_090_2147, w_090_2148, w_090_2150, w_090_2151, w_090_2152, w_090_2157, w_090_2158, w_090_2160, w_090_2162, w_090_2165, w_090_2172, w_090_2173, w_090_2174, w_090_2175, w_090_2179, w_090_2180, w_090_2183, w_090_2184, w_090_2185, w_090_2186, w_090_2190, w_090_2191, w_090_2192, w_090_2194, w_090_2195, w_090_2196, w_090_2197, w_090_2199, w_090_2200, w_090_2201, w_090_2202, w_090_2204, w_090_2207, w_090_2208, w_090_2211, w_090_2212, w_090_2214, w_090_2215, w_090_2216, w_090_2217, w_090_2218, w_090_2221, w_090_2222, w_090_2223, w_090_2225, w_090_2229, w_090_2230, w_090_2231, w_090_2232, w_090_2237, w_090_2239, w_090_2245, w_090_2246, w_090_2250, w_090_2251, w_090_2252, w_090_2254, w_090_2255, w_090_2256, w_090_2257, w_090_2258, w_090_2260, w_090_2261, w_090_2263, w_090_2268, w_090_2269, w_090_2275, w_090_2276, w_090_2277, w_090_2282, w_090_2283, w_090_2285, w_090_2289, w_090_2292, w_090_2293, w_090_2294, w_090_2295, w_090_2296, w_090_2297, w_090_2299, w_090_2301, w_090_2303, w_090_2304, w_090_2308, w_090_2309, w_090_2311, w_090_2312, w_090_2317, w_090_2318, w_090_2321, w_090_2324, w_090_2325, w_090_2327, w_090_2329, w_090_2330, w_090_2331, w_090_2333, w_090_2334, w_090_2335, w_090_2336, w_090_2337, w_090_2339, w_090_2340, w_090_2344, w_090_2347, w_090_2348, w_090_2350, w_090_2352, w_090_2355, w_090_2356, w_090_2357, w_090_2358, w_090_2359, w_090_2360, w_090_2362, w_090_2364, w_090_2365, w_090_2367, w_090_2368, w_090_2371, w_090_2373, w_090_2375, w_090_2376, w_090_2379, w_090_2382, w_090_2385, w_090_2387, w_090_2389, w_090_2392, w_090_2395, w_090_2400, w_090_2401, w_090_2403, w_090_2406, w_090_2410, w_090_2415, w_090_2416, w_090_2420, w_090_2421, w_090_2422, w_090_2423, w_090_2425, w_090_2426, w_090_2427, w_090_2428, w_090_2429, w_090_2430, w_090_2431, w_090_2432, w_090_2433, w_090_2435, w_090_2438, w_090_2439, w_090_2440, w_090_2441, w_090_2442, w_090_2443, w_090_2446, w_090_2449, w_090_2450, w_090_2453, w_090_2455, w_090_2456, w_090_2457, w_090_2459, w_090_2460, w_090_2461, w_090_2465, w_090_2468, w_090_2469, w_090_2471, w_090_2473, w_090_2474, w_090_2475, w_090_2476, w_090_2478, w_090_2479, w_090_2480, w_090_2482, w_090_2484, w_090_2485, w_090_2489, w_090_2491, w_090_2492, w_090_2493, w_090_2496, w_090_2498, w_090_2500, w_090_2501, w_090_2504, w_090_2505, w_090_2506, w_090_2508, w_090_2510, w_090_2514, w_090_2516, w_090_2517, w_090_2518, w_090_2519, w_090_2520, w_090_2522, w_090_2525, w_090_2526, w_090_2527, w_090_2528, w_090_2529, w_090_2530, w_090_2535, w_090_2536, w_090_2539, w_090_2540, w_090_2541, w_090_2542, w_090_2544, w_090_2548, w_090_2550, w_090_2554, w_090_2555, w_090_2559, w_090_2560, w_090_2561, w_090_2563, w_090_2566, w_090_2567, w_090_2570, w_090_2571, w_090_2573, w_090_2577, w_090_2580, w_090_2583, w_090_2584, w_090_2586, w_090_2589, w_090_2590, w_090_2593, w_090_2599, w_090_2600, w_090_2601, w_090_2602, w_090_2604, w_090_2607, w_090_2608, w_090_2609, w_090_2612, w_090_2614, w_090_2615, w_090_2616, w_090_2619, w_090_2620, w_090_2621, w_090_2622, w_090_2624, w_090_2625, w_090_2630, w_090_2632, w_090_2633, w_090_2634, w_090_2635, w_090_2640, w_090_2642, w_090_2644, w_090_2646, w_090_2647, w_090_2648, w_090_2649, w_090_2653, w_090_2654, w_090_2660, w_090_2662, w_090_2666, w_090_2669, w_090_2671, w_090_2672, w_090_2674, w_090_2676, w_090_2678, w_090_2679, w_090_2680, w_090_2681, w_090_2682, w_090_2683, w_090_2684, w_090_2685, w_090_2688, w_090_2690, w_090_2691, w_090_2693, w_090_2695, w_090_2697, w_090_2698, w_090_2699, w_090_2700, w_090_2703, w_090_2704, w_090_2709, w_090_2710, w_090_2711, w_090_2713, w_090_2714, w_090_2715, w_090_2717, w_090_2720, w_090_2722, w_090_2723, w_090_2727, w_090_2728, w_090_2730, w_090_2734, w_090_2736, w_090_2738, w_090_2739, w_090_2740, w_090_2741, w_090_2744, w_090_2745, w_090_2746, w_090_2747, w_090_2748, w_090_2749, w_090_2750, w_090_2752, w_090_2754, w_090_2755, w_090_2756, w_090_2757, w_090_2758, w_090_2760, w_090_2761, w_090_2762, w_090_2763, w_090_2764, w_090_2765, w_090_2767, w_090_2769, w_090_2770, w_090_2771, w_090_2773, w_090_2774, w_090_2775, w_090_2776, w_090_2777, w_090_2778, w_090_2783, w_090_2784, w_090_2786, w_090_2788, w_090_2789, w_090_2792, w_090_2794, w_090_2796, w_090_2798, w_090_2799, w_090_2801, w_090_2802, w_090_2804, w_090_2805, w_090_2807, w_090_2808, w_090_2813, w_090_2817, w_090_2819, w_090_2820, w_090_2822, w_090_2823, w_090_2824, w_090_2827, w_090_2828, w_090_2829, w_090_2832, w_090_2834, w_090_2835, w_090_2836, w_090_2838, w_090_2840, w_090_2842, w_090_2843, w_090_2844, w_090_2845, w_090_2846, w_090_2847, w_090_2848, w_090_2849, w_090_2851, w_090_2852, w_090_2853, w_090_2854, w_090_2855, w_090_2856, w_090_2857, w_090_2858, w_090_2860, w_090_2867, w_090_2868, w_090_2869, w_090_2870, w_090_2871, w_090_2877, w_090_2878, w_090_2879, w_090_2882, w_090_2883, w_090_2884, w_090_2885, w_090_2891, w_090_2893, w_090_2894, w_090_2895, w_090_2897, w_090_2898, w_090_2899, w_090_2900, w_090_2901, w_090_2902, w_090_2904, w_090_2906, w_090_2908, w_090_2909, w_090_2914, w_090_2915, w_090_2917, w_090_2918, w_090_2919, w_090_2920, w_090_2921, w_090_2922, w_090_2923, w_090_2924, w_090_2925, w_090_2927, w_090_2928, w_090_2930, w_090_2932, w_090_2933, w_090_2935, w_090_2936, w_090_2941, w_090_2943, w_090_2944, w_090_2945, w_090_2946, w_090_2947, w_090_2948, w_090_2949, w_090_2950, w_090_2951, w_090_2953, w_090_2954, w_090_2955, w_090_2956, w_090_2957, w_090_2959, w_090_2963, w_090_2967, w_090_2969, w_090_2970, w_090_2976, w_090_2977, w_090_2979, w_090_2980, w_090_2983, w_090_2984, w_090_2985, w_090_2988, w_090_2992, w_090_2995, w_090_2996, w_090_2997, w_090_2999, w_090_3001, w_090_3004, w_090_3007, w_090_3008, w_090_3009, w_090_3011, w_090_3013, w_090_3014, w_090_3015, w_090_3016, w_090_3017, w_090_3019, w_090_3020, w_090_3022, w_090_3025, w_090_3026, w_090_3029, w_090_3034, w_090_3035, w_090_3039, w_090_3040, w_090_3041, w_090_3042, w_090_3043, w_090_3045, w_090_3046, w_090_3047, w_090_3049, w_090_3050, w_090_3051, w_090_3053, w_090_3054, w_090_3055, w_090_3056, w_090_3057, w_090_3060, w_090_3062, w_090_3064, w_090_3065, w_090_3067, w_090_3071, w_090_3072, w_090_3073, w_090_3075, w_090_3076, w_090_3077, w_090_3079, w_090_3081, w_090_3082, w_090_3084, w_090_3085, w_090_3087, w_090_3088, w_090_3090, w_090_3091, w_090_3092, w_090_3094, w_090_3096, w_090_3097, w_090_3100, w_090_3102, w_090_3103, w_090_3105, w_090_3106, w_090_3108, w_090_3109, w_090_3110, w_090_3112, w_090_3114, w_090_3115, w_090_3117, w_090_3118, w_090_3119, w_090_3121, w_090_3122, w_090_3125, w_090_3126, w_090_3128, w_090_3130, w_090_3131, w_090_3132, w_090_3134, w_090_3135, w_090_3138, w_090_3140, w_090_3141, w_090_3143, w_090_3144, w_090_3145, w_090_3146, w_090_3148, w_090_3149, w_090_3152, w_090_3154, w_090_3156, w_090_3157, w_090_3158, w_090_3159, w_090_3160, w_090_3162, w_090_3164, w_090_3165, w_090_3167, w_090_3168, w_090_3169, w_090_3170, w_090_3172, w_090_3174, w_090_3175, w_090_3176, w_090_3178, w_090_3179, w_090_3180, w_090_3181, w_090_3182, w_090_3186, w_090_3188, w_090_3189, w_090_3192, w_090_3195, w_090_3196, w_090_3197, w_090_3198, w_090_3199, w_090_3202, w_090_3205, w_090_3206, w_090_3208, w_090_3211, w_090_3212, w_090_3213, w_090_3215, w_090_3216, w_090_3217, w_090_3218, w_090_3220, w_090_3221, w_090_3222, w_090_3223, w_090_3225, w_090_3226, w_090_3227, w_090_3228, w_090_3229, w_090_3230, w_090_3233, w_090_3236, w_090_3240, w_090_3241, w_090_3243, w_090_3244, w_090_3246, w_090_3248, w_090_3249, w_090_3254, w_090_3256, w_090_3258, w_090_3263, w_090_3265, w_090_3266, w_090_3270, w_090_3271, w_090_3274, w_090_3276, w_090_3279, w_090_3280, w_090_3281, w_090_3282, w_090_3283, w_090_3284, w_090_3285, w_090_3286, w_090_3288, w_090_3289, w_090_3290, w_090_3293, w_090_3297, w_090_3298, w_090_3299, w_090_3300, w_090_3302, w_090_3303, w_090_3304, w_090_3305, w_090_3306, w_090_3308, w_090_3309, w_090_3312, w_090_3314, w_090_3315, w_090_3316, w_090_3317, w_090_3321, w_090_3322, w_090_3323, w_090_3326, w_090_3327, w_090_3328, w_090_3329, w_090_3334, w_090_3335, w_090_3336, w_090_3339, w_090_3342;
  wire w_091_000, w_091_009, w_091_012, w_091_014, w_091_016, w_091_017, w_091_018, w_091_022, w_091_023, w_091_028, w_091_031, w_091_032, w_091_034, w_091_036, w_091_037, w_091_038, w_091_039, w_091_040, w_091_041, w_091_045, w_091_049, w_091_050, w_091_052, w_091_055, w_091_057, w_091_059, w_091_060, w_091_062, w_091_066, w_091_067, w_091_070, w_091_075, w_091_076, w_091_077, w_091_078, w_091_079, w_091_080, w_091_081, w_091_084, w_091_085, w_091_086, w_091_087, w_091_092, w_091_097, w_091_098, w_091_100, w_091_101, w_091_102, w_091_104, w_091_106, w_091_108, w_091_109, w_091_110, w_091_111, w_091_114, w_091_124, w_091_125, w_091_126, w_091_127, w_091_132, w_091_133, w_091_136, w_091_138, w_091_142, w_091_143, w_091_146, w_091_150, w_091_155, w_091_161, w_091_163, w_091_166, w_091_169, w_091_173, w_091_174, w_091_180, w_091_181, w_091_186, w_091_187, w_091_188, w_091_189, w_091_190, w_091_194, w_091_196, w_091_197, w_091_198, w_091_201, w_091_203, w_091_204, w_091_206, w_091_207, w_091_212, w_091_213, w_091_214, w_091_215, w_091_219, w_091_222, w_091_224, w_091_234, w_091_237, w_091_240, w_091_241, w_091_242, w_091_243, w_091_244, w_091_245, w_091_248, w_091_249, w_091_250, w_091_253, w_091_254, w_091_260, w_091_261, w_091_263, w_091_265, w_091_267, w_091_268, w_091_270, w_091_271, w_091_272, w_091_273, w_091_277, w_091_278, w_091_280, w_091_285, w_091_286, w_091_287, w_091_288, w_091_291, w_091_292, w_091_293, w_091_296, w_091_298, w_091_300, w_091_304, w_091_305, w_091_307, w_091_309, w_091_312, w_091_313, w_091_314, w_091_316, w_091_319, w_091_320, w_091_321, w_091_322, w_091_325, w_091_327, w_091_328, w_091_330, w_091_331, w_091_334, w_091_341, w_091_343, w_091_346, w_091_348, w_091_350, w_091_351, w_091_352, w_091_354, w_091_355, w_091_359, w_091_361, w_091_367, w_091_369, w_091_371, w_091_372, w_091_375, w_091_377, w_091_378, w_091_379, w_091_384, w_091_386, w_091_387, w_091_390, w_091_393, w_091_394, w_091_397, w_091_398, w_091_400, w_091_402, w_091_403, w_091_405, w_091_408, w_091_411, w_091_416, w_091_418, w_091_424, w_091_427, w_091_428, w_091_433, w_091_436, w_091_439, w_091_440, w_091_441, w_091_442, w_091_443, w_091_445, w_091_447, w_091_449, w_091_453, w_091_455, w_091_456, w_091_457, w_091_458, w_091_461, w_091_465, w_091_467, w_091_468, w_091_472, w_091_482, w_091_483, w_091_484, w_091_485, w_091_486, w_091_487, w_091_489, w_091_492, w_091_494, w_091_496, w_091_498, w_091_500, w_091_501, w_091_502, w_091_503, w_091_505, w_091_507, w_091_508, w_091_511, w_091_512, w_091_516, w_091_517, w_091_518, w_091_520, w_091_522, w_091_529, w_091_530, w_091_535, w_091_541, w_091_542, w_091_545, w_091_547, w_091_552, w_091_558, w_091_561, w_091_562, w_091_564, w_091_565, w_091_568, w_091_569, w_091_571, w_091_572, w_091_574, w_091_575, w_091_576, w_091_577, w_091_578, w_091_579, w_091_580, w_091_581, w_091_582, w_091_589, w_091_590, w_091_596, w_091_598, w_091_599, w_091_601, w_091_603, w_091_605, w_091_607, w_091_608, w_091_611, w_091_613, w_091_615, w_091_621, w_091_622, w_091_624, w_091_627, w_091_628, w_091_630, w_091_634, w_091_639, w_091_641, w_091_642, w_091_644, w_091_651, w_091_655, w_091_658, w_091_659, w_091_660, w_091_661, w_091_662, w_091_665, w_091_675, w_091_677, w_091_679, w_091_681, w_091_683, w_091_688, w_091_692, w_091_695, w_091_696, w_091_697, w_091_698, w_091_699, w_091_704, w_091_710, w_091_711, w_091_712, w_091_715, w_091_723, w_091_724, w_091_730, w_091_734, w_091_735, w_091_738, w_091_739, w_091_740, w_091_742, w_091_743, w_091_745, w_091_747, w_091_756, w_091_757, w_091_760, w_091_761, w_091_762, w_091_763, w_091_764, w_091_767, w_091_768, w_091_769, w_091_772, w_091_776, w_091_777, w_091_779, w_091_780, w_091_784, w_091_785, w_091_786, w_091_789, w_091_791, w_091_792, w_091_794, w_091_798, w_091_800, w_091_801, w_091_802, w_091_803, w_091_804, w_091_807, w_091_808, w_091_817, w_091_819, w_091_821, w_091_822, w_091_824, w_091_827, w_091_829, w_091_831, w_091_835, w_091_837, w_091_840, w_091_843, w_091_844, w_091_850, w_091_855, w_091_858, w_091_860, w_091_861, w_091_863, w_091_864, w_091_865, w_091_871, w_091_876, w_091_878, w_091_881, w_091_892, w_091_894, w_091_895, w_091_900, w_091_901, w_091_903, w_091_904, w_091_905, w_091_907, w_091_908, w_091_913, w_091_917, w_091_919, w_091_920, w_091_921, w_091_922, w_091_923, w_091_925, w_091_927, w_091_928, w_091_931, w_091_932, w_091_933, w_091_934, w_091_936, w_091_938, w_091_940, w_091_941, w_091_944, w_091_946, w_091_947, w_091_948, w_091_951, w_091_952, w_091_953, w_091_954, w_091_955, w_091_960, w_091_961, w_091_962, w_091_963, w_091_966, w_091_967, w_091_968, w_091_969, w_091_971, w_091_973, w_091_974, w_091_976, w_091_980, w_091_982, w_091_983, w_091_985, w_091_987, w_091_990, w_091_992, w_091_993, w_091_995, w_091_998, w_091_1000, w_091_1001, w_091_1002, w_091_1006, w_091_1007, w_091_1017, w_091_1018, w_091_1022, w_091_1025, w_091_1026, w_091_1028, w_091_1030, w_091_1033, w_091_1035, w_091_1036, w_091_1038, w_091_1040, w_091_1042, w_091_1043, w_091_1044, w_091_1047, w_091_1048, w_091_1053, w_091_1057, w_091_1059, w_091_1061, w_091_1062, w_091_1068, w_091_1070, w_091_1071, w_091_1078, w_091_1080, w_091_1083, w_091_1085, w_091_1086, w_091_1089, w_091_1092, w_091_1097, w_091_1102, w_091_1103, w_091_1104, w_091_1105, w_091_1106, w_091_1108, w_091_1110, w_091_1111, w_091_1112, w_091_1114, w_091_1118, w_091_1119, w_091_1122, w_091_1126, w_091_1129, w_091_1134, w_091_1135, w_091_1136, w_091_1138, w_091_1139, w_091_1141, w_091_1146, w_091_1149, w_091_1150, w_091_1151, w_091_1154, w_091_1156, w_091_1159, w_091_1160, w_091_1161, w_091_1162, w_091_1165, w_091_1167, w_091_1171, w_091_1172, w_091_1173, w_091_1175, w_091_1179, w_091_1182, w_091_1185, w_091_1187, w_091_1189, w_091_1190, w_091_1194, w_091_1197, w_091_1201, w_091_1208, w_091_1214, w_091_1217, w_091_1218, w_091_1220, w_091_1228, w_091_1231, w_091_1233, w_091_1235, w_091_1238, w_091_1239, w_091_1241, w_091_1243, w_091_1250, w_091_1255, w_091_1257, w_091_1258, w_091_1260, w_091_1263, w_091_1264, w_091_1267, w_091_1269, w_091_1272, w_091_1275, w_091_1276, w_091_1279, w_091_1280, w_091_1282, w_091_1283, w_091_1284, w_091_1292, w_091_1295, w_091_1298, w_091_1304, w_091_1306, w_091_1309, w_091_1311, w_091_1313, w_091_1314, w_091_1317, w_091_1318, w_091_1323, w_091_1326, w_091_1333, w_091_1337, w_091_1338, w_091_1341, w_091_1344, w_091_1345, w_091_1350, w_091_1351, w_091_1352, w_091_1354, w_091_1358, w_091_1360, w_091_1362, w_091_1365, w_091_1370, w_091_1371, w_091_1377, w_091_1379, w_091_1380, w_091_1381, w_091_1382, w_091_1383, w_091_1384, w_091_1385, w_091_1387, w_091_1393, w_091_1394, w_091_1396, w_091_1397, w_091_1398, w_091_1402, w_091_1404, w_091_1405, w_091_1406, w_091_1410, w_091_1416, w_091_1418, w_091_1420, w_091_1421, w_091_1424, w_091_1429, w_091_1430, w_091_1432, w_091_1435, w_091_1437, w_091_1438, w_091_1439, w_091_1440, w_091_1442, w_091_1446, w_091_1448, w_091_1449, w_091_1451, w_091_1456, w_091_1458, w_091_1460, w_091_1465, w_091_1466, w_091_1468, w_091_1469, w_091_1470, w_091_1472, w_091_1473, w_091_1476, w_091_1478, w_091_1479, w_091_1482, w_091_1484, w_091_1486, w_091_1488, w_091_1491, w_091_1494, w_091_1497, w_091_1501, w_091_1503, w_091_1506, w_091_1507, w_091_1508, w_091_1509, w_091_1510, w_091_1514, w_091_1515, w_091_1518, w_091_1519, w_091_1522, w_091_1527, w_091_1528, w_091_1535, w_091_1536, w_091_1541, w_091_1542, w_091_1543, w_091_1544, w_091_1545, w_091_1546, w_091_1547, w_091_1549, w_091_1550, w_091_1551, w_091_1552, w_091_1553, w_091_1556, w_091_1557, w_091_1559, w_091_1560, w_091_1562, w_091_1564, w_091_1574, w_091_1575, w_091_1578, w_091_1579, w_091_1580, w_091_1584, w_091_1586, w_091_1587, w_091_1588, w_091_1589, w_091_1590, w_091_1594, w_091_1595, w_091_1600, w_091_1602, w_091_1604, w_091_1605, w_091_1612, w_091_1613, w_091_1616, w_091_1617, w_091_1618, w_091_1619, w_091_1620, w_091_1622, w_091_1625, w_091_1626, w_091_1629, w_091_1631, w_091_1633, w_091_1635, w_091_1638, w_091_1639, w_091_1647, w_091_1648, w_091_1654, w_091_1658, w_091_1661, w_091_1664, w_091_1665, w_091_1666, w_091_1672, w_091_1674, w_091_1677, w_091_1680, w_091_1684, w_091_1687, w_091_1689, w_091_1695, w_091_1698, w_091_1700, w_091_1705, w_091_1716, w_091_1717, w_091_1720, w_091_1721, w_091_1722, w_091_1723, w_091_1725, w_091_1726, w_091_1727, w_091_1736, w_091_1738, w_091_1739, w_091_1748, w_091_1749, w_091_1750, w_091_1752, w_091_1753, w_091_1754, w_091_1756, w_091_1763, w_091_1765, w_091_1766, w_091_1768, w_091_1770, w_091_1771, w_091_1772, w_091_1773, w_091_1778, w_091_1779, w_091_1783, w_091_1784, w_091_1786, w_091_1787, w_091_1788, w_091_1789, w_091_1791, w_091_1792, w_091_1795, w_091_1796, w_091_1797, w_091_1798, w_091_1802, w_091_1804, w_091_1809, w_091_1813, w_091_1817, w_091_1819, w_091_1821, w_091_1822, w_091_1828, w_091_1831, w_091_1838, w_091_1842, w_091_1844, w_091_1845, w_091_1846, w_091_1847, w_091_1848, w_091_1853, w_091_1856, w_091_1859, w_091_1862, w_091_1865, w_091_1867, w_091_1868, w_091_1871, w_091_1873, w_091_1877, w_091_1888, w_091_1893, w_091_1895, w_091_1896, w_091_1898, w_091_1900, w_091_1903, w_091_1905, w_091_1906, w_091_1914, w_091_1916, w_091_1918, w_091_1922, w_091_1927, w_091_1928, w_091_1929, w_091_1930, w_091_1934, w_091_1936, w_091_1938, w_091_1940, w_091_1941, w_091_1944, w_091_1947, w_091_1948, w_091_1953, w_091_1958, w_091_1960, w_091_1963, w_091_1965, w_091_1967, w_091_1968, w_091_1969, w_091_1973, w_091_1974, w_091_1975, w_091_1976, w_091_1977, w_091_1981, w_091_1985, w_091_1987, w_091_1989, w_091_1990, w_091_1991, w_091_1992, w_091_1994, w_091_1998, w_091_1999, w_091_2003, w_091_2004, w_091_2009, w_091_2012, w_091_2015, w_091_2016, w_091_2020, w_091_2022, w_091_2024, w_091_2025, w_091_2029, w_091_2030, w_091_2032, w_091_2033, w_091_2034, w_091_2035, w_091_2039, w_091_2044, w_091_2046, w_091_2051, w_091_2054, w_091_2055, w_091_2056, w_091_2058, w_091_2059, w_091_2067, w_091_2069, w_091_2074, w_091_2078, w_091_2081, w_091_2082, w_091_2086, w_091_2087, w_091_2088, w_091_2092, w_091_2094, w_091_2096, w_091_2098, w_091_2099, w_091_2100, w_091_2103, w_091_2104, w_091_2105, w_091_2108, w_091_2109, w_091_2111, w_091_2115, w_091_2116, w_091_2123, w_091_2124, w_091_2125, w_091_2126, w_091_2128, w_091_2129, w_091_2137, w_091_2142, w_091_2145, w_091_2146, w_091_2148, w_091_2149, w_091_2150, w_091_2151, w_091_2154, w_091_2157, w_091_2159, w_091_2161, w_091_2166, w_091_2169, w_091_2171, w_091_2173, w_091_2175, w_091_2176, w_091_2179, w_091_2180, w_091_2184, w_091_2189, w_091_2192, w_091_2193, w_091_2195, w_091_2196, w_091_2197, w_091_2198, w_091_2200, w_091_2201, w_091_2205, w_091_2210, w_091_2212, w_091_2213, w_091_2217, w_091_2221, w_091_2222, w_091_2223, w_091_2225, w_091_2226, w_091_2232, w_091_2233, w_091_2235, w_091_2238, w_091_2239, w_091_2245, w_091_2246, w_091_2248, w_091_2250, w_091_2251, w_091_2255, w_091_2257, w_091_2258, w_091_2261, w_091_2265, w_091_2266, w_091_2268, w_091_2269, w_091_2273, w_091_2276, w_091_2277, w_091_2279, w_091_2282, w_091_2289, w_091_2293, w_091_2295, w_091_2296, w_091_2298, w_091_2299, w_091_2305, w_091_2308, w_091_2309, w_091_2314, w_091_2315, w_091_2320, w_091_2321, w_091_2324, w_091_2327, w_091_2333, w_091_2334, w_091_2335, w_091_2336, w_091_2338, w_091_2340, w_091_2341, w_091_2343, w_091_2344, w_091_2349, w_091_2352, w_091_2353, w_091_2356, w_091_2357, w_091_2358, w_091_2359, w_091_2361, w_091_2362, w_091_2367, w_091_2370, w_091_2373, w_091_2374, w_091_2375, w_091_2376, w_091_2378, w_091_2379, w_091_2380, w_091_2381, w_091_2383, w_091_2386, w_091_2388, w_091_2389, w_091_2392, w_091_2393, w_091_2394, w_091_2395, w_091_2397, w_091_2399, w_091_2400, w_091_2402, w_091_2403, w_091_2404, w_091_2405, w_091_2406, w_091_2407, w_091_2408, w_091_2410, w_091_2414, w_091_2415, w_091_2419, w_091_2434, w_091_2442, w_091_2443, w_091_2448, w_091_2449, w_091_2450, w_091_2455, w_091_2458, w_091_2466, w_091_2468, w_091_2470, w_091_2475, w_091_2482, w_091_2494, w_091_2496, w_091_2504, w_091_2507, w_091_2508, w_091_2520, w_091_2522, w_091_2526, w_091_2529, w_091_2530, w_091_2531, w_091_2541, w_091_2547, w_091_2549, w_091_2563, w_091_2570, w_091_2571, w_091_2574, w_091_2583, w_091_2598, w_091_2599, w_091_2612, w_091_2616, w_091_2617, w_091_2619, w_091_2621, w_091_2624, w_091_2631, w_091_2638, w_091_2639, w_091_2641, w_091_2643, w_091_2645, w_091_2652, w_091_2655, w_091_2657, w_091_2660, w_091_2663, w_091_2667, w_091_2674, w_091_2679, w_091_2681, w_091_2686, w_091_2687, w_091_2689, w_091_2690, w_091_2694, w_091_2700, w_091_2704, w_091_2718, w_091_2722, w_091_2735, w_091_2736, w_091_2740, w_091_2744, w_091_2746, w_091_2747, w_091_2748, w_091_2750, w_091_2756, w_091_2757, w_091_2761, w_091_2765, w_091_2766, w_091_2775, w_091_2786, w_091_2792, w_091_2794, w_091_2806, w_091_2808, w_091_2811, w_091_2815, w_091_2816, w_091_2826, w_091_2828, w_091_2835, w_091_2836, w_091_2838, w_091_2839, w_091_2840, w_091_2848, w_091_2849, w_091_2850, w_091_2853, w_091_2854, w_091_2857, w_091_2869, w_091_2872, w_091_2877, w_091_2882, w_091_2884, w_091_2889, w_091_2891, w_091_2894, w_091_2896, w_091_2907, w_091_2914, w_091_2921, w_091_2922, w_091_2930, w_091_2931, w_091_2936, w_091_2947, w_091_2951, w_091_2954, w_091_2955, w_091_2962, w_091_2963, w_091_2967, w_091_2971, w_091_2972, w_091_2981, w_091_2988, w_091_2990, w_091_2991, w_091_2994, w_091_2996, w_091_2997, w_091_3004, w_091_3006, w_091_3012, w_091_3014, w_091_3019, w_091_3023, w_091_3024, w_091_3025, w_091_3026, w_091_3029, w_091_3032, w_091_3033, w_091_3036, w_091_3039, w_091_3042, w_091_3057, w_091_3061, w_091_3070, w_091_3074, w_091_3078, w_091_3081, w_091_3085, w_091_3086, w_091_3091, w_091_3093, w_091_3100, w_091_3103, w_091_3105, w_091_3109, w_091_3111, w_091_3114, w_091_3115, w_091_3116, w_091_3118, w_091_3122, w_091_3123, w_091_3128, w_091_3132, w_091_3133, w_091_3135, w_091_3137, w_091_3139, w_091_3143, w_091_3145, w_091_3153, w_091_3157, w_091_3159, w_091_3162, w_091_3165, w_091_3167, w_091_3182, w_091_3189, w_091_3197, w_091_3204, w_091_3207, w_091_3217, w_091_3219, w_091_3223, w_091_3227, w_091_3228, w_091_3229, w_091_3231, w_091_3232, w_091_3234, w_091_3242, w_091_3244, w_091_3258, w_091_3260, w_091_3263, w_091_3266, w_091_3270, w_091_3271, w_091_3272, w_091_3278, w_091_3279, w_091_3283, w_091_3286, w_091_3287, w_091_3289, w_091_3290, w_091_3291, w_091_3306, w_091_3307, w_091_3308, w_091_3310, w_091_3314, w_091_3317, w_091_3320, w_091_3321, w_091_3326, w_091_3331, w_091_3337, w_091_3341, w_091_3346, w_091_3347, w_091_3353, w_091_3358, w_091_3363, w_091_3365, w_091_3367, w_091_3369, w_091_3370, w_091_3374, w_091_3381, w_091_3386, w_091_3393, w_091_3398, w_091_3402, w_091_3411, w_091_3414, w_091_3429, w_091_3433, w_091_3435, w_091_3436, w_091_3439, w_091_3440, w_091_3445, w_091_3446, w_091_3447, w_091_3454, w_091_3466, w_091_3468, w_091_3469, w_091_3474, w_091_3477, w_091_3487, w_091_3489, w_091_3501, w_091_3507, w_091_3510, w_091_3513, w_091_3522, w_091_3530, w_091_3531, w_091_3534, w_091_3539, w_091_3548, w_091_3552, w_091_3553, w_091_3554, w_091_3558, w_091_3565, w_091_3567, w_091_3569, w_091_3570, w_091_3573, w_091_3577, w_091_3580, w_091_3581, w_091_3586, w_091_3599, w_091_3601, w_091_3602, w_091_3605, w_091_3607, w_091_3609, w_091_3620, w_091_3621, w_091_3622, w_091_3624, w_091_3626, w_091_3632, w_091_3636, w_091_3637, w_091_3639, w_091_3643, w_091_3645, w_091_3646, w_091_3651, w_091_3658, w_091_3659, w_091_3665, w_091_3666, w_091_3673, w_091_3678, w_091_3685, w_091_3689, w_091_3691, w_091_3695, w_091_3697, w_091_3705, w_091_3706, w_091_3714, w_091_3735, w_091_3743, w_091_3747, w_091_3748, w_091_3754, w_091_3761, w_091_3763, w_091_3766, w_091_3772, w_091_3773, w_091_3776, w_091_3778, w_091_3784, w_091_3785, w_091_3788, w_091_3790, w_091_3791, w_091_3796, w_091_3802, w_091_3803, w_091_3810, w_091_3811, w_091_3828, w_091_3832, w_091_3836, w_091_3838, w_091_3844, w_091_3848, w_091_3851, w_091_3853, w_091_3856, w_091_3861, w_091_3863, w_091_3865, w_091_3868, w_091_3874, w_091_3876, w_091_3885, w_091_3886, w_091_3887, w_091_3893, w_091_3895, w_091_3899, w_091_3901, w_091_3903, w_091_3907, w_091_3909, w_091_3911, w_091_3917, w_091_3922, w_091_3926, w_091_3930, w_091_3932, w_091_3933, w_091_3942, w_091_3943, w_091_3947, w_091_3949, w_091_3956, w_091_3959, w_091_3962, w_091_3964, w_091_3965, w_091_3970, w_091_3971, w_091_3980, w_091_3988, w_091_3990, w_091_3991, w_091_3993, w_091_3996, w_091_3997, w_091_3999, w_091_4008, w_091_4010, w_091_4012, w_091_4013, w_091_4014, w_091_4015, w_091_4018, w_091_4028, w_091_4030, w_091_4032, w_091_4035, w_091_4037, w_091_4038, w_091_4040, w_091_4041, w_091_4048, w_091_4052, w_091_4053, w_091_4064, w_091_4065, w_091_4066, w_091_4069, w_091_4073, w_091_4083, w_091_4085, w_091_4094, w_091_4105, w_091_4106, w_091_4110, w_091_4113, w_091_4114, w_091_4115, w_091_4120, w_091_4121, w_091_4125, w_091_4127, w_091_4128, w_091_4132, w_091_4134, w_091_4140, w_091_4143, w_091_4145, w_091_4147, w_091_4149, w_091_4153, w_091_4157, w_091_4159, w_091_4165, w_091_4169, w_091_4170, w_091_4171, w_091_4172, w_091_4177, w_091_4183, w_091_4188, w_091_4191, w_091_4193, w_091_4194, w_091_4202, w_091_4203, w_091_4208, w_091_4209, w_091_4211, w_091_4219, w_091_4220, w_091_4225, w_091_4228, w_091_4230, w_091_4231, w_091_4233, w_091_4235, w_091_4236, w_091_4241, w_091_4242, w_091_4243, w_091_4245, w_091_4255, w_091_4260, w_091_4261, w_091_4263, w_091_4265, w_091_4267, w_091_4271, w_091_4281, w_091_4284, w_091_4285, w_091_4286, w_091_4287, w_091_4295, w_091_4303, w_091_4304, w_091_4305, w_091_4307, w_091_4313, w_091_4317, w_091_4320, w_091_4321, w_091_4326, w_091_4332, w_091_4345, w_091_4351, w_091_4352, w_091_4361, w_091_4362, w_091_4365, w_091_4366, w_091_4375, w_091_4376, w_091_4382, w_091_4387, w_091_4388, w_091_4391, w_091_4392, w_091_4399, w_091_4409, w_091_4412, w_091_4419, w_091_4425, w_091_4433, w_091_4436, w_091_4439, w_091_4442, w_091_4453, w_091_4457, w_091_4459, w_091_4464, w_091_4468, w_091_4479, w_091_4480, w_091_4481, w_091_4482, w_091_4483, w_091_4485, w_091_4486, w_091_4487, w_091_4488, w_091_4492, w_091_4496, w_091_4501, w_091_4504, w_091_4505, w_091_4507, w_091_4508, w_091_4509, w_091_4513, w_091_4516, w_091_4520, w_091_4522, w_091_4527, w_091_4528, w_091_4529, w_091_4539, w_091_4541, w_091_4544, w_091_4546, w_091_4548, w_091_4555, w_091_4560, w_091_4562, w_091_4563, w_091_4569, w_091_4571, w_091_4576, w_091_4578, w_091_4582, w_091_4584, w_091_4587, w_091_4596, w_091_4597, w_091_4598, w_091_4604, w_091_4610, w_091_4623, w_091_4626, w_091_4630, w_091_4636, w_091_4641, w_091_4643, w_091_4644, w_091_4645, w_091_4648, w_091_4668, w_091_4671, w_091_4673, w_091_4676, w_091_4678, w_091_4680, w_091_4682, w_091_4690, w_091_4699, w_091_4700, w_091_4701, w_091_4704, w_091_4708, w_091_4714, w_091_4728, w_091_4731, w_091_4734, w_091_4737, w_091_4739, w_091_4740, w_091_4742, w_091_4747, w_091_4758, w_091_4760, w_091_4767, w_091_4772, w_091_4773, w_091_4774, w_091_4778, w_091_4779, w_091_4783, w_091_4785, w_091_4788, w_091_4807, w_091_4812, w_091_4815, w_091_4818, w_091_4819, w_091_4820, w_091_4825, w_091_4838, w_091_4843, w_091_4859, w_091_4860, w_091_4863, w_091_4870, w_091_4880, w_091_4881, w_091_4882, w_091_4883, w_091_4886, w_091_4892, w_091_4894, w_091_4901, w_091_4908, w_091_4923, w_091_4935, w_091_4943, w_091_4944, w_091_4948, w_091_4949, w_091_4956, w_091_4963, w_091_4966, w_091_4967, w_091_4969, w_091_4976, w_091_4977, w_091_4981, w_091_4982, w_091_4985, w_091_4987, w_091_4991, w_091_4995, w_091_5004, w_091_5008, w_091_5010, w_091_5015, w_091_5018, w_091_5023, w_091_5026, w_091_5027, w_091_5040, w_091_5049, w_091_5050, w_091_5051, w_091_5052, w_091_5065, w_091_5067, w_091_5073, w_091_5074, w_091_5075, w_091_5082, w_091_5092, w_091_5095, w_091_5100, w_091_5113, w_091_5121, w_091_5125, w_091_5127, w_091_5128, w_091_5135, w_091_5139, w_091_5140, w_091_5144, w_091_5152, w_091_5153, w_091_5173, w_091_5175, w_091_5177, w_091_5181, w_091_5185, w_091_5195, w_091_5197, w_091_5198, w_091_5200, w_091_5211, w_091_5213, w_091_5217, w_091_5218, w_091_5219, w_091_5220, w_091_5230, w_091_5235, w_091_5236, w_091_5239, w_091_5244, w_091_5249, w_091_5251, w_091_5259, w_091_5269, w_091_5277, w_091_5285, w_091_5287, w_091_5288, w_091_5293, w_091_5301, w_091_5306, w_091_5307, w_091_5309, w_091_5316, w_091_5323, w_091_5326, w_091_5330, w_091_5331, w_091_5333, w_091_5336, w_091_5338, w_091_5347, w_091_5349, w_091_5355, w_091_5356, w_091_5362, w_091_5363, w_091_5364, w_091_5367, w_091_5369, w_091_5370, w_091_5372, w_091_5373, w_091_5386, w_091_5389, w_091_5391, w_091_5392, w_091_5395, w_091_5403, w_091_5409, w_091_5416, w_091_5423, w_091_5428, w_091_5429, w_091_5431, w_091_5441, w_091_5443, w_091_5444, w_091_5448, w_091_5450, w_091_5457, w_091_5458, w_091_5460, w_091_5461, w_091_5463, w_091_5472, w_091_5478, w_091_5480, w_091_5484, w_091_5486, w_091_5487, w_091_5488, w_091_5491, w_091_5496, w_091_5500, w_091_5501, w_091_5502, w_091_5506, w_091_5512, w_091_5513, w_091_5516, w_091_5517, w_091_5521, w_091_5522, w_091_5531, w_091_5535, w_091_5540, w_091_5541, w_091_5546, w_091_5549, w_091_5557, w_091_5560, w_091_5562, w_091_5565, w_091_5567, w_091_5570, w_091_5578, w_091_5596, w_091_5620, w_091_5621, w_091_5627, w_091_5628, w_091_5633, w_091_5648, w_091_5649, w_091_5650, w_091_5654, w_091_5659, w_091_5660, w_091_5666, w_091_5668, w_091_5673, w_091_5674, w_091_5677, w_091_5679, w_091_5680, w_091_5682, w_091_5684, w_091_5685, w_091_5687, w_091_5692, w_091_5699, w_091_5701, w_091_5709, w_091_5711, w_091_5714, w_091_5717, w_091_5722, w_091_5729, w_091_5731, w_091_5735, w_091_5746, w_091_5748, w_091_5749, w_091_5753, w_091_5760, w_091_5762, w_091_5765, w_091_5768, w_091_5769, w_091_5770, w_091_5771, w_091_5772, w_091_5780, w_091_5783, w_091_5786, w_091_5789, w_091_5797, w_091_5801, w_091_5808, w_091_5814, w_091_5826, w_091_5828, w_091_5836, w_091_5838, w_091_5840, w_091_5844, w_091_5846, w_091_5851, w_091_5853, w_091_5857, w_091_5863, w_091_5866, w_091_5876, w_091_5881, w_091_5883, w_091_5885, w_091_5890, w_091_5891, w_091_5904, w_091_5905, w_091_5908, w_091_5914, w_091_5915, w_091_5916, w_091_5920, w_091_5924, w_091_5926, w_091_5927, w_091_5928, w_091_5955, w_091_5957, w_091_5965, w_091_5973, w_091_5977, w_091_5978, w_091_5979, w_091_5982, w_091_5984, w_091_5985, w_091_5988, w_091_5990, w_091_5991, w_091_6000, w_091_6004, w_091_6006, w_091_6007, w_091_6011, w_091_6012, w_091_6014, w_091_6015, w_091_6026, w_091_6027, w_091_6031, w_091_6040, w_091_6044, w_091_6055, w_091_6057, w_091_6062, w_091_6064, w_091_6066, w_091_6072, w_091_6073, w_091_6076, w_091_6077, w_091_6083, w_091_6090, w_091_6098, w_091_6104, w_091_6108, w_091_6110, w_091_6111, w_091_6113, w_091_6119, w_091_6123, w_091_6128, w_091_6131, w_091_6132, w_091_6134, w_091_6136, w_091_6137, w_091_6139, w_091_6141, w_091_6143, w_091_6145, w_091_6151, w_091_6153, w_091_6164, w_091_6178, w_091_6189, w_091_6193, w_091_6206, w_091_6210, w_091_6215, w_091_6228, w_091_6236, w_091_6238, w_091_6246, w_091_6258, w_091_6274, w_091_6277, w_091_6278, w_091_6283, w_091_6286, w_091_6290, w_091_6291, w_091_6294, w_091_6299, w_091_6300, w_091_6301, w_091_6306, w_091_6310, w_091_6311, w_091_6316, w_091_6318, w_091_6319, w_091_6326, w_091_6329, w_091_6334, w_091_6340, w_091_6348, w_091_6351, w_091_6352, w_091_6356, w_091_6361, w_091_6363, w_091_6365, w_091_6369, w_091_6370, w_091_6372, w_091_6374, w_091_6376, w_091_6377, w_091_6387, w_091_6389, w_091_6392, w_091_6396, w_091_6398, w_091_6403, w_091_6405, w_091_6409, w_091_6411, w_091_6412, w_091_6415, w_091_6420, w_091_6429, w_091_6437, w_091_6441, w_091_6442, w_091_6444, w_091_6447, w_091_6451, w_091_6453, w_091_6457, w_091_6458, w_091_6459, w_091_6461, w_091_6466, w_091_6476, w_091_6477, w_091_6479, w_091_6481, w_091_6486, w_091_6489, w_091_6490, w_091_6493, w_091_6494, w_091_6499, w_091_6503, w_091_6504, w_091_6509, w_091_6510, w_091_6513, w_091_6523, w_091_6524, w_091_6528, w_091_6529, w_091_6532, w_091_6534, w_091_6537, w_091_6538, w_091_6540, w_091_6542, w_091_6547, w_091_6550, w_091_6551, w_091_6553, w_091_6554, w_091_6563, w_091_6566, w_091_6570, w_091_6582, w_091_6586, w_091_6587, w_091_6592, w_091_6605, w_091_6606, w_091_6607, w_091_6608, w_091_6610, w_091_6614, w_091_6615, w_091_6617, w_091_6624, w_091_6625, w_091_6627, w_091_6628, w_091_6630, w_091_6634, w_091_6642, w_091_6643, w_091_6646, w_091_6649, w_091_6652, w_091_6659, w_091_6661, w_091_6662, w_091_6665, w_091_6669, w_091_6670, w_091_6675, w_091_6676, w_091_6678, w_091_6679, w_091_6683, w_091_6685, w_091_6694, w_091_6695, w_091_6696, w_091_6697, w_091_6698, w_091_6700, w_091_6701, w_091_6704, w_091_6728, w_091_6729, w_091_6730, w_091_6732, w_091_6738, w_091_6740, w_091_6751, w_091_6752, w_091_6754, w_091_6759, w_091_6762, w_091_6772, w_091_6773, w_091_6774, w_091_6775, w_091_6777, w_091_6785, w_091_6788, w_091_6790, w_091_6793, w_091_6796, w_091_6797, w_091_6804, w_091_6807, w_091_6809, w_091_6817, w_091_6820, w_091_6830, w_091_6834, w_091_6835, w_091_6845, w_091_6847, w_091_6848, w_091_6849, w_091_6850, w_091_6852, w_091_6863, w_091_6869, w_091_6870, w_091_6873, w_091_6876, w_091_6883, w_091_6889, w_091_6892, w_091_6893, w_091_6899, w_091_6900, w_091_6902, w_091_6904, w_091_6908, w_091_6911, w_091_6914, w_091_6922, w_091_6927, w_091_6929, w_091_6933, w_091_6934, w_091_6954, w_091_6963, w_091_6967, w_091_6970, w_091_6971, w_091_6975, w_091_6978, w_091_6992, w_091_6996, w_091_7003, w_091_7012, w_091_7015, w_091_7023, w_091_7024, w_091_7027, w_091_7033, w_091_7041, w_091_7043, w_091_7044, w_091_7047, w_091_7048, w_091_7058, w_091_7060, w_091_7066, w_091_7076, w_091_7078, w_091_7079, w_091_7086, w_091_7087, w_091_7089, w_091_7093, w_091_7094, w_091_7101, w_091_7104, w_091_7105, w_091_7111, w_091_7123, w_091_7124, w_091_7128, w_091_7129, w_091_7135, w_091_7139, w_091_7141, w_091_7146, w_091_7150, w_091_7154, w_091_7159, w_091_7161, w_091_7162, w_091_7163, w_091_7168, w_091_7169, w_091_7173, w_091_7180, w_091_7182, w_091_7183, w_091_7188, w_091_7190, w_091_7192, w_091_7193, w_091_7196, w_091_7198, w_091_7200, w_091_7203, w_091_7208, w_091_7210, w_091_7212, w_091_7214, w_091_7216, w_091_7219, w_091_7222, w_091_7228, w_091_7232, w_091_7240, w_091_7243, w_091_7245, w_091_7247, w_091_7248, w_091_7251, w_091_7253, w_091_7257, w_091_7262, w_091_7269, w_091_7271, w_091_7275, w_091_7276, w_091_7283, w_091_7287, w_091_7290, w_091_7291, w_091_7296, w_091_7298, w_091_7299, w_091_7301, w_091_7305, w_091_7306, w_091_7308, w_091_7319, w_091_7326, w_091_7329, w_091_7330, w_091_7331, w_091_7335, w_091_7336, w_091_7337, w_091_7339, w_091_7340, w_091_7348, w_091_7350, w_091_7358, w_091_7359, w_091_7365, w_091_7376, w_091_7388, w_091_7393, w_091_7400, w_091_7404, w_091_7410, w_091_7412, w_091_7414, w_091_7420, w_091_7425, w_091_7431, w_091_7433, w_091_7436, w_091_7438, w_091_7439, w_091_7447, w_091_7461, w_091_7464, w_091_7465, w_091_7467, w_091_7468, w_091_7478, w_091_7480, w_091_7481, w_091_7483, w_091_7485, w_091_7490, w_091_7494, w_091_7501, w_091_7505, w_091_7506, w_091_7507, w_091_7511, w_091_7513, w_091_7519, w_091_7523, w_091_7524, w_091_7537, w_091_7539, w_091_7541, w_091_7543, w_091_7546, w_091_7550, w_091_7551, w_091_7552, w_091_7560, w_091_7562, w_091_7564, w_091_7565, w_091_7566;
  wire w_092_003, w_092_004, w_092_006, w_092_014, w_092_015, w_092_016, w_092_018, w_092_021, w_092_022, w_092_024, w_092_025, w_092_026, w_092_028, w_092_034, w_092_035, w_092_036, w_092_037, w_092_038, w_092_039, w_092_040, w_092_044, w_092_045, w_092_048, w_092_049, w_092_057, w_092_058, w_092_063, w_092_064, w_092_065, w_092_067, w_092_068, w_092_071, w_092_072, w_092_078, w_092_080, w_092_083, w_092_085, w_092_087, w_092_088, w_092_092, w_092_093, w_092_096, w_092_099, w_092_100, w_092_101, w_092_107, w_092_108, w_092_111, w_092_116, w_092_117, w_092_118, w_092_119, w_092_120, w_092_121, w_092_122, w_092_124, w_092_134, w_092_136, w_092_139, w_092_143, w_092_150, w_092_152, w_092_154, w_092_155, w_092_157, w_092_158, w_092_161, w_092_165, w_092_169, w_092_170, w_092_171, w_092_172, w_092_174, w_092_176, w_092_177, w_092_179, w_092_183, w_092_184, w_092_187, w_092_191, w_092_192, w_092_194, w_092_197, w_092_198, w_092_199, w_092_204, w_092_206, w_092_207, w_092_209, w_092_210, w_092_213, w_092_214, w_092_216, w_092_218, w_092_220, w_092_225, w_092_226, w_092_227, w_092_231, w_092_234, w_092_238, w_092_242, w_092_243, w_092_245, w_092_248, w_092_249, w_092_251, w_092_253, w_092_254, w_092_257, w_092_260, w_092_261, w_092_271, w_092_273, w_092_277, w_092_278, w_092_285, w_092_288, w_092_289, w_092_290, w_092_293, w_092_294, w_092_295, w_092_296, w_092_297, w_092_298, w_092_299, w_092_301, w_092_302, w_092_305, w_092_308, w_092_309, w_092_313, w_092_314, w_092_316, w_092_319, w_092_325, w_092_326, w_092_327, w_092_329, w_092_330, w_092_331, w_092_333, w_092_335, w_092_336, w_092_337, w_092_338, w_092_339, w_092_343, w_092_344, w_092_345, w_092_346, w_092_347, w_092_351, w_092_355, w_092_359, w_092_364, w_092_369, w_092_370, w_092_374, w_092_375, w_092_377, w_092_379, w_092_381, w_092_382, w_092_383, w_092_387, w_092_391, w_092_393, w_092_402, w_092_411, w_092_413, w_092_415, w_092_417, w_092_422, w_092_424, w_092_425, w_092_428, w_092_430, w_092_433, w_092_434, w_092_435, w_092_438, w_092_448, w_092_451, w_092_458, w_092_459, w_092_460, w_092_461, w_092_462, w_092_464, w_092_466, w_092_468, w_092_472, w_092_474, w_092_477, w_092_485, w_092_487, w_092_488, w_092_490, w_092_491, w_092_492, w_092_493, w_092_496, w_092_497, w_092_498, w_092_500, w_092_502, w_092_503, w_092_504, w_092_507, w_092_510, w_092_514, w_092_515, w_092_516, w_092_519, w_092_522, w_092_523, w_092_524, w_092_526, w_092_528, w_092_529, w_092_531, w_092_532, w_092_534, w_092_537, w_092_540, w_092_543, w_092_545, w_092_546, w_092_547, w_092_548, w_092_554, w_092_555, w_092_560, w_092_562, w_092_564, w_092_567, w_092_570, w_092_572, w_092_574, w_092_581, w_092_582, w_092_584, w_092_585, w_092_586, w_092_589, w_092_590, w_092_592, w_092_595, w_092_596, w_092_598, w_092_600, w_092_604, w_092_605, w_092_606, w_092_609, w_092_613, w_092_615, w_092_621, w_092_622, w_092_625, w_092_629, w_092_633, w_092_634, w_092_640, w_092_644, w_092_646, w_092_647, w_092_648, w_092_650, w_092_654, w_092_655, w_092_656, w_092_657, w_092_659, w_092_661, w_092_663, w_092_665, w_092_666, w_092_667, w_092_669, w_092_675, w_092_680, w_092_683, w_092_689, w_092_691, w_092_692, w_092_696, w_092_697, w_092_699, w_092_701, w_092_707, w_092_708, w_092_711, w_092_712, w_092_714, w_092_716, w_092_717, w_092_718, w_092_720, w_092_721, w_092_722, w_092_723, w_092_727, w_092_728, w_092_732, w_092_733, w_092_738, w_092_740, w_092_741, w_092_743, w_092_748, w_092_749, w_092_753, w_092_754, w_092_766, w_092_772, w_092_773, w_092_774, w_092_776, w_092_777, w_092_778, w_092_782, w_092_783, w_092_784, w_092_785, w_092_787, w_092_788, w_092_790, w_092_791, w_092_793, w_092_795, w_092_798, w_092_801, w_092_802, w_092_803, w_092_806, w_092_807, w_092_811, w_092_813, w_092_816, w_092_817, w_092_818, w_092_821, w_092_822, w_092_823, w_092_825, w_092_827, w_092_829, w_092_831, w_092_832, w_092_836, w_092_837, w_092_838, w_092_839, w_092_841, w_092_842, w_092_844, w_092_846, w_092_851, w_092_853, w_092_858, w_092_859, w_092_860, w_092_861, w_092_862, w_092_863, w_092_866, w_092_868, w_092_872, w_092_875, w_092_876, w_092_883, w_092_889, w_092_890, w_092_894, w_092_900, w_092_901, w_092_903, w_092_909, w_092_912, w_092_914, w_092_916, w_092_919, w_092_920, w_092_921, w_092_924, w_092_926, w_092_930, w_092_935, w_092_937, w_092_940, w_092_941, w_092_943, w_092_946, w_092_947, w_092_949, w_092_950, w_092_951, w_092_954, w_092_955, w_092_957, w_092_959, w_092_960, w_092_967, w_092_969, w_092_971, w_092_973, w_092_974, w_092_975, w_092_980, w_092_981, w_092_990, w_092_991, w_092_993, w_092_994, w_092_998, w_092_1001, w_092_1008, w_092_1011, w_092_1012, w_092_1013, w_092_1014, w_092_1017, w_092_1019, w_092_1024, w_092_1025, w_092_1027, w_092_1034, w_092_1035, w_092_1036, w_092_1037, w_092_1044, w_092_1050, w_092_1058, w_092_1063, w_092_1069, w_092_1070, w_092_1071, w_092_1074, w_092_1080, w_092_1081, w_092_1083, w_092_1084, w_092_1085, w_092_1087, w_092_1091, w_092_1092, w_092_1094, w_092_1099, w_092_1101, w_092_1102, w_092_1106, w_092_1116, w_092_1117, w_092_1127, w_092_1131, w_092_1132, w_092_1134, w_092_1137, w_092_1140, w_092_1147, w_092_1148, w_092_1161, w_092_1163, w_092_1172, w_092_1174, w_092_1175, w_092_1182, w_092_1190, w_092_1207, w_092_1215, w_092_1220, w_092_1234, w_092_1237, w_092_1238, w_092_1239, w_092_1240, w_092_1242, w_092_1243, w_092_1247, w_092_1248, w_092_1257, w_092_1268, w_092_1278, w_092_1279, w_092_1286, w_092_1290, w_092_1293, w_092_1297, w_092_1309, w_092_1312, w_092_1314, w_092_1316, w_092_1320, w_092_1326, w_092_1331, w_092_1337, w_092_1340, w_092_1344, w_092_1352, w_092_1356, w_092_1359, w_092_1362, w_092_1364, w_092_1365, w_092_1369, w_092_1372, w_092_1373, w_092_1384, w_092_1387, w_092_1392, w_092_1396, w_092_1400, w_092_1402, w_092_1412, w_092_1414, w_092_1417, w_092_1418, w_092_1421, w_092_1424, w_092_1431, w_092_1434, w_092_1435, w_092_1438, w_092_1445, w_092_1450, w_092_1453, w_092_1454, w_092_1455, w_092_1459, w_092_1465, w_092_1473, w_092_1478, w_092_1483, w_092_1484, w_092_1485, w_092_1486, w_092_1489, w_092_1491, w_092_1492, w_092_1496, w_092_1498, w_092_1501, w_092_1505, w_092_1509, w_092_1515, w_092_1517, w_092_1518, w_092_1521, w_092_1523, w_092_1532, w_092_1534, w_092_1538, w_092_1540, w_092_1543, w_092_1551, w_092_1553, w_092_1572, w_092_1580, w_092_1589, w_092_1592, w_092_1593, w_092_1600, w_092_1608, w_092_1612, w_092_1614, w_092_1621, w_092_1624, w_092_1633, w_092_1634, w_092_1635, w_092_1638, w_092_1643, w_092_1645, w_092_1646, w_092_1659, w_092_1660, w_092_1661, w_092_1668, w_092_1671, w_092_1672, w_092_1673, w_092_1675, w_092_1683, w_092_1684, w_092_1685, w_092_1694, w_092_1700, w_092_1705, w_092_1716, w_092_1719, w_092_1726, w_092_1727, w_092_1739, w_092_1741, w_092_1747, w_092_1752, w_092_1755, w_092_1759, w_092_1763, w_092_1767, w_092_1771, w_092_1776, w_092_1779, w_092_1785, w_092_1786, w_092_1787, w_092_1790, w_092_1797, w_092_1800, w_092_1806, w_092_1817, w_092_1820, w_092_1822, w_092_1825, w_092_1832, w_092_1834, w_092_1840, w_092_1842, w_092_1860, w_092_1864, w_092_1868, w_092_1870, w_092_1871, w_092_1875, w_092_1881, w_092_1883, w_092_1888, w_092_1895, w_092_1897, w_092_1909, w_092_1915, w_092_1921, w_092_1922, w_092_1927, w_092_1930, w_092_1934, w_092_1938, w_092_1939, w_092_1941, w_092_1949, w_092_1952, w_092_1955, w_092_1956, w_092_1959, w_092_1961, w_092_1964, w_092_1965, w_092_1970, w_092_1976, w_092_1996, w_092_1997, w_092_1999, w_092_2000, w_092_2002, w_092_2011, w_092_2012, w_092_2016, w_092_2017, w_092_2018, w_092_2020, w_092_2022, w_092_2027, w_092_2028, w_092_2038, w_092_2039, w_092_2053, w_092_2054, w_092_2062, w_092_2066, w_092_2075, w_092_2084, w_092_2086, w_092_2097, w_092_2102, w_092_2108, w_092_2113, w_092_2116, w_092_2119, w_092_2120, w_092_2121, w_092_2122, w_092_2124, w_092_2125, w_092_2126, w_092_2128, w_092_2130, w_092_2131, w_092_2143, w_092_2149, w_092_2152, w_092_2153, w_092_2155, w_092_2159, w_092_2160, w_092_2162, w_092_2164, w_092_2165, w_092_2171, w_092_2184, w_092_2185, w_092_2188, w_092_2190, w_092_2193, w_092_2195, w_092_2197, w_092_2199, w_092_2201, w_092_2203, w_092_2205, w_092_2207, w_092_2209, w_092_2210, w_092_2222, w_092_2224, w_092_2227, w_092_2232, w_092_2233, w_092_2238, w_092_2239, w_092_2241, w_092_2242, w_092_2251, w_092_2253, w_092_2254, w_092_2255, w_092_2262, w_092_2264, w_092_2270, w_092_2273, w_092_2281, w_092_2282, w_092_2283, w_092_2286, w_092_2288, w_092_2294, w_092_2297, w_092_2299, w_092_2304, w_092_2305, w_092_2306, w_092_2314, w_092_2316, w_092_2322, w_092_2336, w_092_2338, w_092_2339, w_092_2343, w_092_2346, w_092_2350, w_092_2351, w_092_2362, w_092_2363, w_092_2367, w_092_2368, w_092_2375, w_092_2376, w_092_2381, w_092_2385, w_092_2388, w_092_2394, w_092_2400, w_092_2401, w_092_2403, w_092_2404, w_092_2405, w_092_2409, w_092_2412, w_092_2427, w_092_2428, w_092_2431, w_092_2433, w_092_2442, w_092_2443, w_092_2446, w_092_2447, w_092_2460, w_092_2465, w_092_2470, w_092_2483, w_092_2492, w_092_2508, w_092_2509, w_092_2510, w_092_2518, w_092_2526, w_092_2531, w_092_2532, w_092_2533, w_092_2534, w_092_2543, w_092_2544, w_092_2549, w_092_2550, w_092_2566, w_092_2567, w_092_2570, w_092_2572, w_092_2582, w_092_2586, w_092_2591, w_092_2601, w_092_2606, w_092_2613, w_092_2614, w_092_2615, w_092_2619, w_092_2620, w_092_2621, w_092_2626, w_092_2628, w_092_2635, w_092_2637, w_092_2646, w_092_2649, w_092_2651, w_092_2652, w_092_2657, w_092_2665, w_092_2667, w_092_2669, w_092_2671, w_092_2672, w_092_2674, w_092_2676, w_092_2678, w_092_2679, w_092_2680, w_092_2682, w_092_2684, w_092_2685, w_092_2686, w_092_2690, w_092_2693, w_092_2696, w_092_2701, w_092_2708, w_092_2715, w_092_2719, w_092_2721, w_092_2740, w_092_2743, w_092_2749, w_092_2753, w_092_2757, w_092_2761, w_092_2763, w_092_2775, w_092_2776, w_092_2792, w_092_2795, w_092_2800, w_092_2801, w_092_2802, w_092_2803, w_092_2807, w_092_2808, w_092_2809, w_092_2811, w_092_2817, w_092_2828, w_092_2830, w_092_2831, w_092_2832, w_092_2835, w_092_2844, w_092_2848, w_092_2849, w_092_2857, w_092_2859, w_092_2861, w_092_2863, w_092_2868, w_092_2878, w_092_2880, w_092_2881, w_092_2891, w_092_2899, w_092_2904, w_092_2913, w_092_2917, w_092_2918, w_092_2930, w_092_2932, w_092_2935, w_092_2940, w_092_2941, w_092_2948, w_092_2953, w_092_2960, w_092_2962, w_092_2971, w_092_2972, w_092_2976, w_092_2982, w_092_2990, w_092_2991, w_092_2993, w_092_2995, w_092_3002, w_092_3012, w_092_3019, w_092_3020, w_092_3023, w_092_3026, w_092_3028, w_092_3032, w_092_3036, w_092_3038, w_092_3040, w_092_3041, w_092_3052, w_092_3053, w_092_3055, w_092_3062, w_092_3063, w_092_3072, w_092_3075, w_092_3084, w_092_3085, w_092_3088, w_092_3089, w_092_3092, w_092_3105, w_092_3108, w_092_3115, w_092_3121, w_092_3123, w_092_3124, w_092_3126, w_092_3128, w_092_3132, w_092_3143, w_092_3146, w_092_3147, w_092_3148, w_092_3158, w_092_3163, w_092_3169, w_092_3175, w_092_3179, w_092_3183, w_092_3185, w_092_3191, w_092_3201, w_092_3207, w_092_3209, w_092_3211, w_092_3214, w_092_3222, w_092_3231, w_092_3238, w_092_3239, w_092_3244, w_092_3245, w_092_3247, w_092_3249, w_092_3251, w_092_3254, w_092_3265, w_092_3268, w_092_3269, w_092_3272, w_092_3281, w_092_3282, w_092_3284, w_092_3285, w_092_3287, w_092_3298, w_092_3304, w_092_3305, w_092_3306, w_092_3311, w_092_3313, w_092_3315, w_092_3320, w_092_3323, w_092_3324, w_092_3326, w_092_3333, w_092_3335, w_092_3338, w_092_3340, w_092_3341, w_092_3351, w_092_3352, w_092_3365, w_092_3369, w_092_3380, w_092_3389, w_092_3390, w_092_3392, w_092_3393, w_092_3394, w_092_3406, w_092_3409, w_092_3410, w_092_3424, w_092_3439, w_092_3448, w_092_3451, w_092_3452, w_092_3458, w_092_3459, w_092_3477, w_092_3478, w_092_3481, w_092_3487, w_092_3488, w_092_3491, w_092_3499, w_092_3504, w_092_3513, w_092_3514, w_092_3519, w_092_3524, w_092_3525, w_092_3526, w_092_3529, w_092_3534, w_092_3537, w_092_3543, w_092_3545, w_092_3547, w_092_3556, w_092_3559, w_092_3562, w_092_3565, w_092_3573, w_092_3581, w_092_3584, w_092_3588, w_092_3597, w_092_3604, w_092_3610, w_092_3618, w_092_3623, w_092_3625, w_092_3640, w_092_3641, w_092_3646, w_092_3652, w_092_3654, w_092_3657, w_092_3675, w_092_3677, w_092_3680, w_092_3695, w_092_3701, w_092_3703, w_092_3707, w_092_3708, w_092_3709, w_092_3722, w_092_3731, w_092_3733, w_092_3734, w_092_3735, w_092_3736, w_092_3740, w_092_3745, w_092_3750, w_092_3751, w_092_3753, w_092_3755, w_092_3756, w_092_3764, w_092_3774, w_092_3776, w_092_3778, w_092_3779, w_092_3781, w_092_3782, w_092_3788, w_092_3792, w_092_3796, w_092_3798, w_092_3809, w_092_3817, w_092_3821, w_092_3823, w_092_3824, w_092_3828, w_092_3831, w_092_3835, w_092_3836, w_092_3837, w_092_3842, w_092_3843, w_092_3844, w_092_3847, w_092_3853, w_092_3859, w_092_3864, w_092_3867, w_092_3869, w_092_3871, w_092_3873, w_092_3879, w_092_3880, w_092_3888, w_092_3889, w_092_3890, w_092_3892, w_092_3896, w_092_3901, w_092_3906, w_092_3907, w_092_3910, w_092_3912, w_092_3914, w_092_3916, w_092_3918, w_092_3923, w_092_3927, w_092_3937, w_092_3944, w_092_3945, w_092_3946, w_092_3951, w_092_3952, w_092_3958, w_092_3959, w_092_3964, w_092_3971, w_092_3973, w_092_3976, w_092_3977, w_092_3978, w_092_3979, w_092_3984, w_092_3985, w_092_3987, w_092_3989, w_092_3995, w_092_3997, w_092_4017, w_092_4019, w_092_4023, w_092_4024, w_092_4027, w_092_4029, w_092_4033, w_092_4037, w_092_4038, w_092_4041, w_092_4042, w_092_4047, w_092_4053, w_092_4059, w_092_4064, w_092_4068, w_092_4078, w_092_4079, w_092_4083, w_092_4084, w_092_4086, w_092_4091, w_092_4094, w_092_4101, w_092_4102, w_092_4104, w_092_4107, w_092_4108, w_092_4113, w_092_4116, w_092_4117, w_092_4118, w_092_4121, w_092_4128, w_092_4139, w_092_4145, w_092_4147, w_092_4150, w_092_4151, w_092_4162, w_092_4176, w_092_4186, w_092_4187, w_092_4188, w_092_4193, w_092_4197, w_092_4204, w_092_4210, w_092_4217, w_092_4228, w_092_4232, w_092_4239, w_092_4242, w_092_4244, w_092_4251, w_092_4253, w_092_4257, w_092_4258, w_092_4259, w_092_4280, w_092_4283, w_092_4286, w_092_4299, w_092_4311, w_092_4320, w_092_4322, w_092_4329, w_092_4345, w_092_4357, w_092_4363, w_092_4371, w_092_4372, w_092_4376, w_092_4377, w_092_4388, w_092_4390, w_092_4391, w_092_4397, w_092_4401, w_092_4407, w_092_4412, w_092_4414, w_092_4415, w_092_4416, w_092_4419, w_092_4425, w_092_4432, w_092_4433, w_092_4450, w_092_4453, w_092_4456, w_092_4462, w_092_4464, w_092_4470, w_092_4478, w_092_4481, w_092_4483, w_092_4488, w_092_4492, w_092_4493, w_092_4500, w_092_4506, w_092_4508, w_092_4518, w_092_4520, w_092_4527, w_092_4531, w_092_4568, w_092_4573, w_092_4577, w_092_4580, w_092_4581, w_092_4589, w_092_4594, w_092_4595, w_092_4598, w_092_4601, w_092_4606, w_092_4611, w_092_4612, w_092_4613, w_092_4616, w_092_4621, w_092_4624, w_092_4626, w_092_4627, w_092_4635, w_092_4644, w_092_4648, w_092_4649, w_092_4652, w_092_4658, w_092_4661, w_092_4662, w_092_4665, w_092_4667, w_092_4671, w_092_4681, w_092_4684, w_092_4693, w_092_4695, w_092_4698, w_092_4701, w_092_4702, w_092_4711, w_092_4715, w_092_4725, w_092_4731, w_092_4732, w_092_4734, w_092_4735, w_092_4737, w_092_4738, w_092_4740, w_092_4744, w_092_4745, w_092_4748, w_092_4754, w_092_4755, w_092_4761, w_092_4766, w_092_4776, w_092_4779, w_092_4783, w_092_4791, w_092_4792, w_092_4799, w_092_4800, w_092_4804, w_092_4806, w_092_4807, w_092_4814, w_092_4819, w_092_4843, w_092_4859, w_092_4864, w_092_4865, w_092_4866, w_092_4870, w_092_4880, w_092_4884, w_092_4886, w_092_4887, w_092_4895, w_092_4899, w_092_4902, w_092_4905, w_092_4906, w_092_4907, w_092_4909, w_092_4922, w_092_4926, w_092_4928, w_092_4930, w_092_4935, w_092_4939, w_092_4941, w_092_4942, w_092_4943, w_092_4944, w_092_4945, w_092_4946, w_092_4950, w_092_4951, w_092_4954, w_092_4956, w_092_4958, w_092_4965, w_092_4969, w_092_4972, w_092_4975, w_092_4976, w_092_4978, w_092_5008, w_092_5009, w_092_5012, w_092_5014, w_092_5016, w_092_5035, w_092_5040, w_092_5041, w_092_5042, w_092_5046, w_092_5049, w_092_5050, w_092_5056, w_092_5061, w_092_5065, w_092_5071, w_092_5076, w_092_5077, w_092_5078, w_092_5079, w_092_5082, w_092_5090, w_092_5092, w_092_5106, w_092_5110, w_092_5115, w_092_5119, w_092_5121, w_092_5129, w_092_5131, w_092_5135, w_092_5139, w_092_5143, w_092_5147, w_092_5148, w_092_5149, w_092_5151, w_092_5153, w_092_5154, w_092_5155, w_092_5157, w_092_5158, w_092_5159, w_092_5163, w_092_5165, w_092_5168, w_092_5193, w_092_5197, w_092_5211, w_092_5216, w_092_5220, w_092_5223, w_092_5224, w_092_5234, w_092_5246, w_092_5248, w_092_5255, w_092_5256, w_092_5257, w_092_5259, w_092_5260, w_092_5261, w_092_5262, w_092_5264, w_092_5277, w_092_5279, w_092_5285, w_092_5288, w_092_5291, w_092_5296, w_092_5298, w_092_5302, w_092_5305, w_092_5307, w_092_5312, w_092_5317, w_092_5318, w_092_5321, w_092_5322, w_092_5325, w_092_5333, w_092_5337, w_092_5346, w_092_5349, w_092_5350, w_092_5351, w_092_5354, w_092_5355, w_092_5361, w_092_5365, w_092_5370, w_092_5371, w_092_5372, w_092_5381, w_092_5384, w_092_5388, w_092_5389, w_092_5394, w_092_5402, w_092_5405, w_092_5414, w_092_5415, w_092_5423, w_092_5428, w_092_5432, w_092_5445, w_092_5451, w_092_5454, w_092_5464, w_092_5476, w_092_5483, w_092_5487, w_092_5500, w_092_5503, w_092_5507, w_092_5512, w_092_5513, w_092_5517, w_092_5519, w_092_5523, w_092_5527, w_092_5531, w_092_5538, w_092_5552, w_092_5553, w_092_5557, w_092_5559, w_092_5574, w_092_5581, w_092_5583, w_092_5586, w_092_5587, w_092_5588, w_092_5593, w_092_5596, w_092_5603, w_092_5606, w_092_5611, w_092_5612, w_092_5615, w_092_5616, w_092_5621, w_092_5623, w_092_5628, w_092_5638, w_092_5640, w_092_5644, w_092_5649, w_092_5650, w_092_5658, w_092_5664, w_092_5670, w_092_5671, w_092_5672, w_092_5674, w_092_5677, w_092_5684, w_092_5688, w_092_5696, w_092_5697, w_092_5699, w_092_5701, w_092_5710, w_092_5715, w_092_5718, w_092_5720, w_092_5728, w_092_5743, w_092_5744, w_092_5749, w_092_5753, w_092_5754, w_092_5759, w_092_5767, w_092_5770, w_092_5771, w_092_5773, w_092_5775, w_092_5778, w_092_5785, w_092_5786, w_092_5788, w_092_5789, w_092_5794, w_092_5799, w_092_5800, w_092_5803, w_092_5808, w_092_5809, w_092_5812, w_092_5823, w_092_5827, w_092_5829, w_092_5832, w_092_5840, w_092_5843, w_092_5848, w_092_5850, w_092_5852, w_092_5859, w_092_5860, w_092_5863, w_092_5864, w_092_5866, w_092_5868, w_092_5872, w_092_5873, w_092_5879, w_092_5880, w_092_5885, w_092_5886, w_092_5890, w_092_5892, w_092_5894, w_092_5895, w_092_5896, w_092_5897, w_092_5906, w_092_5908, w_092_5916, w_092_5919, w_092_5930, w_092_5932, w_092_5939, w_092_5940, w_092_5941, w_092_5944, w_092_5949, w_092_5950, w_092_5955, w_092_5961, w_092_5964, w_092_5965, w_092_5974, w_092_5979, w_092_5984, w_092_5989, w_092_5993, w_092_5996, w_092_5998, w_092_6000, w_092_6007, w_092_6008, w_092_6014, w_092_6015, w_092_6016, w_092_6018, w_092_6022, w_092_6023, w_092_6025, w_092_6035, w_092_6036, w_092_6037, w_092_6040, w_092_6054, w_092_6055, w_092_6058, w_092_6072, w_092_6087, w_092_6096, w_092_6097, w_092_6102, w_092_6103, w_092_6104, w_092_6108, w_092_6109, w_092_6110, w_092_6114, w_092_6119, w_092_6127, w_092_6129, w_092_6137, w_092_6144, w_092_6146, w_092_6149, w_092_6150, w_092_6151, w_092_6155, w_092_6158, w_092_6161, w_092_6179, w_092_6180, w_092_6187, w_092_6190, w_092_6191, w_092_6192, w_092_6196, w_092_6198, w_092_6199, w_092_6200, w_092_6212, w_092_6222, w_092_6227, w_092_6229, w_092_6230, w_092_6231, w_092_6232, w_092_6240, w_092_6245, w_092_6253, w_092_6257, w_092_6264, w_092_6265, w_092_6266, w_092_6269, w_092_6270, w_092_6275, w_092_6278, w_092_6298, w_092_6305, w_092_6306, w_092_6307, w_092_6311, w_092_6315, w_092_6316, w_092_6322, w_092_6323, w_092_6324, w_092_6328, w_092_6330, w_092_6337, w_092_6340, w_092_6347, w_092_6348, w_092_6351, w_092_6353, w_092_6356, w_092_6360, w_092_6368, w_092_6376, w_092_6378, w_092_6379, w_092_6380, w_092_6385, w_092_6394, w_092_6402, w_092_6404, w_092_6406, w_092_6411, w_092_6416, w_092_6418, w_092_6419, w_092_6420, w_092_6426, w_092_6433, w_092_6440, w_092_6441, w_092_6443, w_092_6448, w_092_6451, w_092_6460, w_092_6466, w_092_6471, w_092_6478, w_092_6482, w_092_6485, w_092_6486, w_092_6488, w_092_6492, w_092_6494, w_092_6507, w_092_6508, w_092_6515, w_092_6517, w_092_6520, w_092_6522, w_092_6525, w_092_6530, w_092_6537, w_092_6539, w_092_6541, w_092_6551, w_092_6553, w_092_6556, w_092_6558, w_092_6562, w_092_6564, w_092_6567, w_092_6570, w_092_6580, w_092_6582, w_092_6584, w_092_6586, w_092_6587, w_092_6596, w_092_6598, w_092_6601, w_092_6605, w_092_6606, w_092_6607, w_092_6612, w_092_6618, w_092_6622, w_092_6626, w_092_6635, w_092_6637, w_092_6638, w_092_6640, w_092_6641, w_092_6643, w_092_6652, w_092_6655, w_092_6662, w_092_6665, w_092_6666, w_092_6674, w_092_6681, w_092_6686, w_092_6687, w_092_6697, w_092_6700, w_092_6702, w_092_6708, w_092_6709, w_092_6716, w_092_6718, w_092_6732, w_092_6734, w_092_6739, w_092_6741, w_092_6747, w_092_6752, w_092_6753, w_092_6759, w_092_6776, w_092_6779, w_092_6792, w_092_6801, w_092_6805, w_092_6807, w_092_6809, w_092_6810, w_092_6813, w_092_6816, w_092_6824, w_092_6827, w_092_6829, w_092_6830, w_092_6833, w_092_6834, w_092_6846, w_092_6851, w_092_6861, w_092_6864, w_092_6866, w_092_6869, w_092_6872, w_092_6876, w_092_6877, w_092_6878, w_092_6883, w_092_6887, w_092_6893, w_092_6894, w_092_6896, w_092_6899, w_092_6900, w_092_6906, w_092_6911, w_092_6913, w_092_6925, w_092_6928, w_092_6934, w_092_6936, w_092_6938, w_092_6942, w_092_6943, w_092_6948, w_092_6949, w_092_6950, w_092_6951, w_092_6952, w_092_6956, w_092_6961, w_092_6963, w_092_6966, w_092_6976, w_092_6979, w_092_6997, w_092_6998, w_092_6999, w_092_7001, w_092_7003, w_092_7009, w_092_7011, w_092_7013, w_092_7021, w_092_7027, w_092_7028, w_092_7031, w_092_7036, w_092_7041, w_092_7044, w_092_7051, w_092_7053, w_092_7061, w_092_7070, w_092_7079, w_092_7080, w_092_7085, w_092_7086, w_092_7087, w_092_7096, w_092_7099, w_092_7102, w_092_7113, w_092_7118, w_092_7122, w_092_7132, w_092_7134, w_092_7135, w_092_7140, w_092_7141, w_092_7148, w_092_7152, w_092_7154, w_092_7155, w_092_7161, w_092_7167, w_092_7173, w_092_7174, w_092_7178, w_092_7179, w_092_7182, w_092_7184, w_092_7187, w_092_7192, w_092_7196, w_092_7198, w_092_7203, w_092_7204, w_092_7213, w_092_7216, w_092_7218, w_092_7221, w_092_7224, w_092_7227, w_092_7230, w_092_7231, w_092_7233, w_092_7235, w_092_7237, w_092_7242, w_092_7246, w_092_7255, w_092_7257, w_092_7258, w_092_7262, w_092_7263, w_092_7269, w_092_7270, w_092_7293, w_092_7305, w_092_7306, w_092_7307, w_092_7311, w_092_7313, w_092_7314, w_092_7324, w_092_7331, w_092_7334, w_092_7335, w_092_7338, w_092_7341, w_092_7342, w_092_7346, w_092_7355, w_092_7359, w_092_7360, w_092_7368, w_092_7387, w_092_7392, w_092_7395, w_092_7396, w_092_7397, w_092_7401, w_092_7402, w_092_7405, w_092_7409, w_092_7412, w_092_7415, w_092_7418, w_092_7422, w_092_7425, w_092_7428, w_092_7432, w_092_7434, w_092_7435, w_092_7439, w_092_7442, w_092_7443, w_092_7446, w_092_7452, w_092_7469, w_092_7475, w_092_7492, w_092_7500, w_092_7505, w_092_7506, w_092_7519, w_092_7520, w_092_7525, w_092_7529, w_092_7532, w_092_7533, w_092_7534, w_092_7535, w_092_7540, w_092_7543, w_092_7544, w_092_7545, w_092_7548, w_092_7549, w_092_7551, w_092_7554, w_092_7561, w_092_7562, w_092_7571, w_092_7578, w_092_7580, w_092_7583, w_092_7587, w_092_7588, w_092_7592, w_092_7598, w_092_7600, w_092_7603, w_092_7610, w_092_7613, w_092_7618, w_092_7619, w_092_7625, w_092_7635, w_092_7638, w_092_7639, w_092_7644, w_092_7646, w_092_7649, w_092_7650, w_092_7653, w_092_7662, w_092_7663, w_092_7664, w_092_7668, w_092_7670, w_092_7672, w_092_7674, w_092_7677, w_092_7683, w_092_7684, w_092_7687, w_092_7691, w_092_7694, w_092_7701, w_092_7702, w_092_7712, w_092_7718, w_092_7720, w_092_7721, w_092_7722, w_092_7724, w_092_7726, w_092_7732, w_092_7734, w_092_7739, w_092_7746, w_092_7750, w_092_7758, w_092_7763, w_092_7764, w_092_7766, w_092_7770, w_092_7771, w_092_7773, w_092_7778, w_092_7780, w_092_7783, w_092_7787, w_092_7791, w_092_7793, w_092_7796, w_092_7800, w_092_7803, w_092_7818, w_092_7822, w_092_7828, w_092_7832, w_092_7835, w_092_7843, w_092_7845, w_092_7849, w_092_7852, w_092_7856, w_092_7859, w_092_7860, w_092_7861, w_092_7863, w_092_7865, w_092_7871, w_092_7875, w_092_7879, w_092_7880, w_092_7884, w_092_7885, w_092_7888, w_092_7889, w_092_7892, w_092_7896, w_092_7905, w_092_7907, w_092_7911, w_092_7915, w_092_7928, w_092_7929, w_092_7933, w_092_7937, w_092_7939, w_092_7940, w_092_7947, w_092_7949, w_092_7951, w_092_7953, w_092_7957, w_092_7959, w_092_7970, w_092_7982, w_092_7983, w_092_7986, w_092_7988, w_092_7992, w_092_8000, w_092_8005, w_092_8008, w_092_8010, w_092_8014, w_092_8019, w_092_8021, w_092_8026, w_092_8028, w_092_8035, w_092_8040, w_092_8045, w_092_8047, w_092_8051, w_092_8053, w_092_8055, w_092_8062, w_092_8064, w_092_8067, w_092_8084, w_092_8085, w_092_8086, w_092_8097, w_092_8098, w_092_8101, w_092_8106, w_092_8114, w_092_8115, w_092_8120, w_092_8121, w_092_8124, w_092_8125, w_092_8126, w_092_8133, w_092_8136, w_092_8137, w_092_8139, w_092_8147, w_092_8148, w_092_8150, w_092_8156, w_092_8157, w_092_8164, w_092_8169, w_092_8173, w_092_8177, w_092_8184, w_092_8193, w_092_8206, w_092_8209, w_092_8217, w_092_8227, w_092_8234, w_092_8236, w_092_8251, w_092_8253, w_092_8254, w_092_8258, w_092_8264, w_092_8265, w_092_8268, w_092_8270, w_092_8272, w_092_8275, w_092_8278, w_092_8279, w_092_8285, w_092_8286, w_092_8288, w_092_8296, w_092_8298, w_092_8302, w_092_8303, w_092_8310, w_092_8313, w_092_8317, w_092_8319, w_092_8320, w_092_8324, w_092_8326, w_092_8328, w_092_8329, w_092_8336, w_092_8343, w_092_8354, w_092_8358, w_092_8374, w_092_8382, w_092_8388, w_092_8390, w_092_8391, w_092_8395, w_092_8397, w_092_8402, w_092_8406, w_092_8417, w_092_8422, w_092_8423, w_092_8426, w_092_8427, w_092_8431, w_092_8433, w_092_8441, w_092_8443, w_092_8444, w_092_8457, w_092_8459, w_092_8462, w_092_8463, w_092_8464, w_092_8465, w_092_8469, w_092_8474, w_092_8477, w_092_8478, w_092_8479, w_092_8484, w_092_8488, w_092_8498, w_092_8500, w_092_8503, w_092_8504, w_092_8505, w_092_8514, w_092_8516, w_092_8526, w_092_8534, w_092_8535, w_092_8536, w_092_8545, w_092_8552, w_092_8561, w_092_8562, w_092_8571, w_092_8572, w_092_8576, w_092_8578, w_092_8588, w_092_8591, w_092_8592, w_092_8597, w_092_8603, w_092_8604, w_092_8606, w_092_8614, w_092_8620, w_092_8632, w_092_8635, w_092_8639, w_092_8641, w_092_8647, w_092_8648, w_092_8649, w_092_8650, w_092_8659, w_092_8663, w_092_8665, w_092_8667, w_092_8672, w_092_8679, w_092_8685, w_092_8687, w_092_8689, w_092_8690, w_092_8691, w_092_8692, w_092_8694, w_092_8695, w_092_8697, w_092_8705, w_092_8706, w_092_8707, w_092_8708, w_092_8711, w_092_8714, w_092_8715, w_092_8717, w_092_8724, w_092_8726, w_092_8743, w_092_8748, w_092_8751, w_092_8753, w_092_8757, w_092_8761, w_092_8764, w_092_8765, w_092_8766, w_092_8771, w_092_8773, w_092_8774, w_092_8776, w_092_8783, w_092_8789, w_092_8790, w_092_8797, w_092_8802, w_092_8813, w_092_8816, w_092_8825, w_092_8827, w_092_8833, w_092_8836, w_092_8848, w_092_8852, w_092_8859, w_092_8861, w_092_8863, w_092_8866, w_092_8871, w_092_8874, w_092_8879, w_092_8881, w_092_8882, w_092_8885, w_092_8893, w_092_8894, w_092_8895, w_092_8899, w_092_8902;
  wire w_093_000, w_093_002, w_093_004, w_093_010, w_093_011, w_093_016, w_093_017, w_093_022, w_093_023, w_093_027, w_093_028, w_093_029, w_093_030, w_093_032, w_093_034, w_093_036, w_093_037, w_093_038, w_093_041, w_093_042, w_093_043, w_093_044, w_093_053, w_093_055, w_093_057, w_093_059, w_093_062, w_093_063, w_093_064, w_093_066, w_093_067, w_093_069, w_093_072, w_093_075, w_093_080, w_093_083, w_093_086, w_093_089, w_093_092, w_093_096, w_093_099, w_093_103, w_093_104, w_093_105, w_093_106, w_093_107, w_093_110, w_093_112, w_093_114, w_093_117, w_093_122, w_093_124, w_093_127, w_093_129, w_093_133, w_093_141, w_093_143, w_093_147, w_093_148, w_093_150, w_093_152, w_093_157, w_093_159, w_093_162, w_093_164, w_093_165, w_093_170, w_093_172, w_093_174, w_093_175, w_093_176, w_093_177, w_093_182, w_093_183, w_093_186, w_093_190, w_093_191, w_093_193, w_093_194, w_093_195, w_093_198, w_093_200, w_093_201, w_093_204, w_093_206, w_093_207, w_093_208, w_093_210, w_093_212, w_093_215, w_093_217, w_093_221, w_093_223, w_093_224, w_093_225, w_093_226, w_093_227, w_093_229, w_093_232, w_093_234, w_093_236, w_093_238, w_093_239, w_093_240, w_093_242, w_093_245, w_093_246, w_093_249, w_093_251, w_093_252, w_093_253, w_093_254, w_093_256, w_093_257, w_093_259, w_093_260, w_093_262, w_093_266, w_093_271, w_093_275, w_093_278, w_093_279, w_093_280, w_093_281, w_093_284, w_093_286, w_093_289, w_093_291, w_093_293, w_093_294, w_093_295, w_093_296, w_093_300, w_093_303, w_093_305, w_093_308, w_093_310, w_093_314, w_093_315, w_093_318, w_093_320, w_093_323, w_093_327, w_093_330, w_093_332, w_093_333, w_093_335, w_093_336, w_093_342, w_093_348, w_093_349, w_093_352, w_093_353, w_093_356, w_093_357, w_093_363, w_093_368, w_093_371, w_093_373, w_093_374, w_093_376, w_093_377, w_093_378, w_093_379, w_093_384, w_093_385, w_093_389, w_093_391, w_093_393, w_093_397, w_093_399, w_093_401, w_093_405, w_093_406, w_093_407, w_093_408, w_093_409, w_093_413, w_093_414, w_093_415, w_093_416, w_093_417, w_093_421, w_093_423, w_093_424, w_093_429, w_093_430, w_093_437, w_093_439, w_093_442, w_093_444, w_093_447, w_093_449, w_093_450, w_093_451, w_093_454, w_093_455, w_093_458, w_093_459, w_093_460, w_093_461, w_093_464, w_093_465, w_093_466, w_093_468, w_093_470, w_093_472, w_093_473, w_093_480, w_093_484, w_093_486, w_093_489, w_093_492, w_093_493, w_093_494, w_093_495, w_093_496, w_093_497, w_093_500, w_093_503, w_093_504, w_093_506, w_093_507, w_093_509, w_093_510, w_093_514, w_093_516, w_093_517, w_093_519, w_093_522, w_093_526, w_093_529, w_093_530, w_093_531, w_093_535, w_093_539, w_093_540, w_093_542, w_093_543, w_093_544, w_093_546, w_093_551, w_093_554, w_093_556, w_093_557, w_093_558, w_093_564, w_093_565, w_093_566, w_093_569, w_093_573, w_093_574, w_093_575, w_093_577, w_093_588, w_093_589, w_093_593, w_093_596, w_093_598, w_093_603, w_093_605, w_093_612, w_093_614, w_093_616, w_093_621, w_093_622, w_093_623, w_093_625, w_093_627, w_093_628, w_093_630, w_093_631, w_093_632, w_093_634, w_093_635, w_093_637, w_093_643, w_093_645, w_093_646, w_093_649, w_093_650, w_093_651, w_093_653, w_093_655, w_093_657, w_093_658, w_093_659, w_093_661, w_093_663, w_093_665, w_093_668, w_093_669, w_093_672, w_093_678, w_093_681, w_093_682, w_093_683, w_093_687, w_093_689, w_093_694, w_093_701, w_093_702, w_093_703, w_093_707, w_093_709, w_093_710, w_093_711, w_093_712, w_093_713, w_093_717, w_093_719, w_093_721, w_093_723, w_093_727, w_093_729, w_093_731, w_093_732, w_093_735, w_093_737, w_093_738, w_093_740, w_093_741, w_093_742, w_093_745, w_093_747, w_093_751, w_093_753, w_093_755, w_093_757, w_093_758, w_093_759, w_093_760, w_093_761, w_093_767, w_093_768, w_093_771, w_093_775, w_093_779, w_093_780, w_093_781, w_093_782, w_093_783, w_093_789, w_093_791, w_093_793, w_093_795, w_093_796, w_093_801, w_093_805, w_093_807, w_093_808, w_093_809, w_093_811, w_093_813, w_093_814, w_093_817, w_093_826, w_093_828, w_093_829, w_093_833, w_093_834, w_093_837, w_093_845, w_093_847, w_093_848, w_093_849, w_093_852, w_093_856, w_093_857, w_093_858, w_093_859, w_093_865, w_093_866, w_093_870, w_093_871, w_093_873, w_093_875, w_093_876, w_093_877, w_093_878, w_093_885, w_093_889, w_093_892, w_093_901, w_093_903, w_093_910, w_093_911, w_093_912, w_093_915, w_093_916, w_093_917, w_093_921, w_093_926, w_093_927, w_093_929, w_093_930, w_093_935, w_093_938, w_093_943, w_093_944, w_093_950, w_093_952, w_093_955, w_093_956, w_093_959, w_093_960, w_093_964, w_093_966, w_093_967, w_093_974, w_093_981, w_093_986, w_093_987, w_093_989, w_093_990, w_093_992, w_093_994, w_093_995, w_093_997, w_093_998, w_093_1002, w_093_1007, w_093_1008, w_093_1009, w_093_1012, w_093_1013, w_093_1016, w_093_1018, w_093_1020, w_093_1029, w_093_1030, w_093_1032, w_093_1036, w_093_1037, w_093_1039, w_093_1040, w_093_1044, w_093_1046, w_093_1047, w_093_1049, w_093_1050, w_093_1052, w_093_1053, w_093_1056, w_093_1057, w_093_1060, w_093_1062, w_093_1064, w_093_1065, w_093_1067, w_093_1069, w_093_1072, w_093_1077, w_093_1078, w_093_1081, w_093_1084, w_093_1085, w_093_1086, w_093_1089, w_093_1091, w_093_1092, w_093_1093, w_093_1094, w_093_1097, w_093_1098, w_093_1103, w_093_1104, w_093_1105, w_093_1106, w_093_1107, w_093_1111, w_093_1117, w_093_1118, w_093_1123, w_093_1127, w_093_1128, w_093_1132, w_093_1133, w_093_1134, w_093_1139, w_093_1143, w_093_1144, w_093_1145, w_093_1146, w_093_1152, w_093_1157, w_093_1158, w_093_1159, w_093_1160, w_093_1167, w_093_1171, w_093_1180, w_093_1184, w_093_1185, w_093_1187, w_093_1188, w_093_1189, w_093_1190, w_093_1192, w_093_1193, w_093_1195, w_093_1196, w_093_1198, w_093_1205, w_093_1207, w_093_1208, w_093_1209, w_093_1210, w_093_1212, w_093_1216, w_093_1217, w_093_1221, w_093_1224, w_093_1228, w_093_1230, w_093_1232, w_093_1233, w_093_1234, w_093_1237, w_093_1241, w_093_1242, w_093_1245, w_093_1248, w_093_1249, w_093_1256, w_093_1258, w_093_1260, w_093_1261, w_093_1262, w_093_1267, w_093_1270, w_093_1271, w_093_1272, w_093_1274, w_093_1277, w_093_1278, w_093_1279, w_093_1283, w_093_1288, w_093_1291, w_093_1295, w_093_1299, w_093_1300, w_093_1301, w_093_1302, w_093_1305, w_093_1317, w_093_1318, w_093_1319, w_093_1321, w_093_1326, w_093_1329, w_093_1330, w_093_1332, w_093_1339, w_093_1342, w_093_1343, w_093_1344, w_093_1345, w_093_1346, w_093_1347, w_093_1348, w_093_1354, w_093_1355, w_093_1356, w_093_1358, w_093_1359, w_093_1362, w_093_1364, w_093_1365, w_093_1368, w_093_1369, w_093_1373, w_093_1376, w_093_1377, w_093_1380, w_093_1382, w_093_1383, w_093_1386, w_093_1388, w_093_1390, w_093_1391, w_093_1392, w_093_1394, w_093_1396, w_093_1399, w_093_1404, w_093_1411, w_093_1412, w_093_1419, w_093_1420, w_093_1431, w_093_1433, w_093_1440, w_093_1441, w_093_1443, w_093_1449, w_093_1450, w_093_1451, w_093_1452, w_093_1454, w_093_1456, w_093_1457, w_093_1459, w_093_1461, w_093_1464, w_093_1466, w_093_1468, w_093_1470, w_093_1471, w_093_1473, w_093_1474, w_093_1475, w_093_1485, w_093_1487, w_093_1491, w_093_1496, w_093_1506, w_093_1507, w_093_1517, w_093_1521, w_093_1522, w_093_1523, w_093_1525, w_093_1526, w_093_1530, w_093_1531, w_093_1534, w_093_1535, w_093_1536, w_093_1538, w_093_1542, w_093_1543, w_093_1549, w_093_1553, w_093_1556, w_093_1557, w_093_1561, w_093_1563, w_093_1565, w_093_1567, w_093_1568, w_093_1570, w_093_1571, w_093_1573, w_093_1575, w_093_1576, w_093_1577, w_093_1579, w_093_1582, w_093_1583, w_093_1584, w_093_1586, w_093_1588, w_093_1591, w_093_1593, w_093_1597, w_093_1598, w_093_1599, w_093_1603, w_093_1604, w_093_1605, w_093_1606, w_093_1607, w_093_1609, w_093_1615, w_093_1617, w_093_1620, w_093_1621, w_093_1623, w_093_1624, w_093_1627, w_093_1628, w_093_1629, w_093_1630, w_093_1637, w_093_1640, w_093_1642, w_093_1643, w_093_1644, w_093_1650, w_093_1651, w_093_1655, w_093_1658, w_093_1660, w_093_1662, w_093_1663, w_093_1670, w_093_1674, w_093_1675, w_093_1677, w_093_1678, w_093_1679, w_093_1684, w_093_1685, w_093_1688, w_093_1692, w_093_1695, w_093_1696, w_093_1699, w_093_1703, w_093_1705, w_093_1706, w_093_1711, w_093_1713, w_093_1715, w_093_1720, w_093_1722, w_093_1723, w_093_1726, w_093_1728, w_093_1729, w_093_1730, w_093_1731, w_093_1733, w_093_1735, w_093_1736, w_093_1738, w_093_1739, w_093_1744, w_093_1746, w_093_1754, w_093_1756, w_093_1761, w_093_1764, w_093_1774, w_093_1776, w_093_1777, w_093_1778, w_093_1780, w_093_1784, w_093_1785, w_093_1787, w_093_1790, w_093_1793, w_093_1794, w_093_1795, w_093_1796, w_093_1797, w_093_1798, w_093_1800, w_093_1803, w_093_1804, w_093_1809, w_093_1810, w_093_1811, w_093_1813, w_093_1816, w_093_1821, w_093_1823, w_093_1824, w_093_1826, w_093_1827, w_093_1831, w_093_1833, w_093_1836, w_093_1837, w_093_1838, w_093_1840, w_093_1845, w_093_1847, w_093_1849, w_093_1860, w_093_1862, w_093_1865, w_093_1868, w_093_1869, w_093_1870, w_093_1875, w_093_1877, w_093_1879, w_093_1881, w_093_1882, w_093_1883, w_093_1887, w_093_1888, w_093_1889, w_093_1890, w_093_1894, w_093_1896, w_093_1897, w_093_1900, w_093_1905, w_093_1906, w_093_1910, w_093_1914, w_093_1917, w_093_1918, w_093_1919, w_093_1923, w_093_1925, w_093_1926, w_093_1927, w_093_1929, w_093_1930, w_093_1932, w_093_1933, w_093_1935, w_093_1936, w_093_1937, w_093_1939, w_093_1941, w_093_1944, w_093_1945, w_093_1950, w_093_1955, w_093_1957, w_093_1959, w_093_1961, w_093_1962, w_093_1963, w_093_1966, w_093_1968, w_093_1972, w_093_1973, w_093_1975, w_093_1978, w_093_1981, w_093_1983, w_093_1985, w_093_1987, w_093_1988, w_093_1989, w_093_1991, w_093_1992, w_093_1993, w_093_1995, w_093_1996, w_093_1997, w_093_2000, w_093_2001, w_093_2003, w_093_2010, w_093_2012, w_093_2017, w_093_2021, w_093_2024, w_093_2025, w_093_2028, w_093_2033, w_093_2034, w_093_2036, w_093_2037, w_093_2040, w_093_2041, w_093_2042, w_093_2046, w_093_2051, w_093_2052, w_093_2054, w_093_2055, w_093_2056, w_093_2057, w_093_2059, w_093_2067, w_093_2068, w_093_2069, w_093_2073, w_093_2074, w_093_2078, w_093_2083, w_093_2086, w_093_2088, w_093_2089, w_093_2092, w_093_2093, w_093_2096, w_093_2099, w_093_2100, w_093_2107, w_093_2109, w_093_2110, w_093_2116, w_093_2118, w_093_2120, w_093_2121, w_093_2123, w_093_2135, w_093_2143, w_093_2145, w_093_2146, w_093_2152, w_093_2153, w_093_2155, w_093_2156, w_093_2161, w_093_2165, w_093_2166, w_093_2167, w_093_2169, w_093_2171, w_093_2172, w_093_2176, w_093_2177, w_093_2179, w_093_2183, w_093_2184, w_093_2185, w_093_2188, w_093_2190, w_093_2191, w_093_2192, w_093_2197, w_093_2204, w_093_2207, w_093_2210, w_093_2213, w_093_2215, w_093_2219, w_093_2220, w_093_2225, w_093_2226, w_093_2227, w_093_2228, w_093_2229, w_093_2231, w_093_2234, w_093_2238, w_093_2240, w_093_2241, w_093_2242, w_093_2245, w_093_2253, w_093_2256, w_093_2257, w_093_2258, w_093_2261, w_093_2262, w_093_2267, w_093_2268, w_093_2270, w_093_2272, w_093_2273, w_093_2278, w_093_2280, w_093_2283, w_093_2284, w_093_2285, w_093_2289, w_093_2290, w_093_2295, w_093_2298, w_093_2300, w_093_2303, w_093_2304, w_093_2305, w_093_2306, w_093_2309, w_093_2312, w_093_2313, w_093_2314, w_093_2316, w_093_2320, w_093_2323, w_093_2324, w_093_2327, w_093_2328, w_093_2329, w_093_2331, w_093_2332, w_093_2335, w_093_2337, w_093_2340, w_093_2341, w_093_2345, w_093_2346, w_093_2348, w_093_2349, w_093_2350, w_093_2351, w_093_2353, w_093_2357, w_093_2359, w_093_2360, w_093_2362, w_093_2366, w_093_2367, w_093_2368, w_093_2369, w_093_2370, w_093_2372, w_093_2375, w_093_2376, w_093_2384, w_093_2386, w_093_2387, w_093_2388, w_093_2390, w_093_2393, w_093_2404, w_093_2406, w_093_2407, w_093_2411, w_093_2412, w_093_2415, w_093_2417, w_093_2420, w_093_2421, w_093_2423, w_093_2425, w_093_2426, w_093_2433, w_093_2434, w_093_2435, w_093_2437, w_093_2439, w_093_2442, w_093_2461, w_093_2467, w_093_2474, w_093_2478, w_093_2485, w_093_2487, w_093_2492, w_093_2501, w_093_2512, w_093_2515, w_093_2520, w_093_2524, w_093_2543, w_093_2548, w_093_2550, w_093_2556, w_093_2558, w_093_2562, w_093_2563, w_093_2564, w_093_2565, w_093_2572, w_093_2573, w_093_2578, w_093_2580, w_093_2581, w_093_2584, w_093_2588, w_093_2598, w_093_2603, w_093_2604, w_093_2614, w_093_2618, w_093_2636, w_093_2638, w_093_2639, w_093_2641, w_093_2647, w_093_2649, w_093_2655, w_093_2657, w_093_2658, w_093_2663, w_093_2664, w_093_2667, w_093_2670, w_093_2672, w_093_2673, w_093_2676, w_093_2678, w_093_2687, w_093_2688, w_093_2689, w_093_2692, w_093_2695, w_093_2698, w_093_2704, w_093_2705, w_093_2709, w_093_2710, w_093_2712, w_093_2713, w_093_2720, w_093_2725, w_093_2728, w_093_2733, w_093_2735, w_093_2736, w_093_2740, w_093_2742, w_093_2748, w_093_2750, w_093_2751, w_093_2758, w_093_2771, w_093_2778, w_093_2781, w_093_2783, w_093_2788, w_093_2789, w_093_2790, w_093_2797, w_093_2798, w_093_2803, w_093_2808, w_093_2816, w_093_2818, w_093_2820, w_093_2824, w_093_2826, w_093_2828, w_093_2832, w_093_2833, w_093_2839, w_093_2841, w_093_2844, w_093_2845, w_093_2846, w_093_2848, w_093_2849, w_093_2850, w_093_2851, w_093_2855, w_093_2860, w_093_2867, w_093_2872, w_093_2874, w_093_2881, w_093_2882, w_093_2888, w_093_2889, w_093_2896, w_093_2904, w_093_2915, w_093_2921, w_093_2924, w_093_2930, w_093_2937, w_093_2939, w_093_2942, w_093_2943, w_093_2945, w_093_2949, w_093_2952, w_093_2955, w_093_2957, w_093_2959, w_093_2962, w_093_2963, w_093_2964, w_093_2967, w_093_2968, w_093_2973, w_093_2978, w_093_2979, w_093_2981, w_093_2983, w_093_2985, w_093_2986, w_093_2995, w_093_3002, w_093_3003, w_093_3004, w_093_3005, w_093_3010, w_093_3015, w_093_3018, w_093_3032, w_093_3038, w_093_3039, w_093_3043, w_093_3059, w_093_3061, w_093_3070, w_093_3074, w_093_3076, w_093_3082, w_093_3083, w_093_3085, w_093_3087, w_093_3088, w_093_3092, w_093_3094, w_093_3095, w_093_3101, w_093_3103, w_093_3111, w_093_3113, w_093_3122, w_093_3130, w_093_3138, w_093_3142, w_093_3146, w_093_3147, w_093_3155, w_093_3159, w_093_3172, w_093_3175, w_093_3177, w_093_3183, w_093_3188, w_093_3190, w_093_3194, w_093_3206, w_093_3210, w_093_3217, w_093_3224, w_093_3225, w_093_3226, w_093_3228, w_093_3241, w_093_3246, w_093_3251, w_093_3260, w_093_3263, w_093_3271, w_093_3272, w_093_3279, w_093_3280, w_093_3281, w_093_3283, w_093_3286, w_093_3288, w_093_3294, w_093_3295, w_093_3296, w_093_3301, w_093_3308, w_093_3319, w_093_3323, w_093_3327, w_093_3332, w_093_3338, w_093_3341, w_093_3342, w_093_3344, w_093_3348, w_093_3349, w_093_3353, w_093_3358, w_093_3362, w_093_3363, w_093_3364, w_093_3365, w_093_3372, w_093_3374, w_093_3376, w_093_3378, w_093_3384, w_093_3385, w_093_3387, w_093_3388, w_093_3389, w_093_3393, w_093_3394, w_093_3395, w_093_3403, w_093_3404, w_093_3405, w_093_3418, w_093_3420, w_093_3422, w_093_3427, w_093_3434, w_093_3440, w_093_3443, w_093_3444, w_093_3445, w_093_3446, w_093_3447, w_093_3448, w_093_3450, w_093_3454, w_093_3460, w_093_3463, w_093_3465, w_093_3472, w_093_3474, w_093_3477, w_093_3485, w_093_3486, w_093_3487, w_093_3488, w_093_3491, w_093_3499, w_093_3506, w_093_3512, w_093_3517, w_093_3523, w_093_3524, w_093_3528, w_093_3531, w_093_3536, w_093_3541, w_093_3544, w_093_3548, w_093_3549, w_093_3553, w_093_3557, w_093_3564, w_093_3566, w_093_3568, w_093_3572, w_093_3577, w_093_3578, w_093_3583, w_093_3587, w_093_3591, w_093_3597, w_093_3600, w_093_3601, w_093_3608, w_093_3611, w_093_3615, w_093_3617, w_093_3632, w_093_3638, w_093_3639, w_093_3640, w_093_3641, w_093_3644, w_093_3647, w_093_3652, w_093_3654, w_093_3655, w_093_3656, w_093_3663, w_093_3665, w_093_3669, w_093_3675, w_093_3680, w_093_3681, w_093_3682, w_093_3690, w_093_3697, w_093_3700, w_093_3708, w_093_3710, w_093_3719, w_093_3722, w_093_3725, w_093_3732, w_093_3734, w_093_3736, w_093_3751, w_093_3752, w_093_3779, w_093_3783, w_093_3787, w_093_3788, w_093_3791, w_093_3792, w_093_3794, w_093_3798, w_093_3799, w_093_3809, w_093_3810, w_093_3817, w_093_3821, w_093_3823, w_093_3824, w_093_3827, w_093_3829, w_093_3831, w_093_3847, w_093_3848, w_093_3860, w_093_3865, w_093_3869, w_093_3870, w_093_3871, w_093_3879, w_093_3883, w_093_3886, w_093_3888, w_093_3892, w_093_3895, w_093_3899, w_093_3915, w_093_3919, w_093_3922, w_093_3928, w_093_3931, w_093_3932, w_093_3935, w_093_3938, w_093_3939, w_093_3952, w_093_3958, w_093_3959, w_093_3963, w_093_3974, w_093_3986, w_093_3988, w_093_3993, w_093_4003, w_093_4005, w_093_4006, w_093_4027, w_093_4037, w_093_4038, w_093_4039, w_093_4040, w_093_4041, w_093_4043, w_093_4051, w_093_4064, w_093_4068, w_093_4071, w_093_4078, w_093_4079, w_093_4082, w_093_4087, w_093_4088, w_093_4090, w_093_4101, w_093_4103, w_093_4106, w_093_4115, w_093_4119, w_093_4127, w_093_4130, w_093_4139, w_093_4140, w_093_4144, w_093_4148, w_093_4149, w_093_4154, w_093_4158, w_093_4165, w_093_4171, w_093_4173, w_093_4174, w_093_4175, w_093_4183, w_093_4192, w_093_4196, w_093_4206, w_093_4207, w_093_4211, w_093_4212, w_093_4214, w_093_4218, w_093_4226, w_093_4230, w_093_4231, w_093_4232, w_093_4236, w_093_4238, w_093_4241, w_093_4244, w_093_4245, w_093_4247, w_093_4250, w_093_4256, w_093_4258, w_093_4264, w_093_4277, w_093_4284, w_093_4289, w_093_4298, w_093_4302, w_093_4305, w_093_4310, w_093_4318, w_093_4321, w_093_4323, w_093_4325, w_093_4341, w_093_4343, w_093_4344, w_093_4348, w_093_4352, w_093_4361, w_093_4362, w_093_4367, w_093_4373, w_093_4376, w_093_4382, w_093_4384, w_093_4385, w_093_4398, w_093_4412, w_093_4422, w_093_4428, w_093_4437, w_093_4438, w_093_4448, w_093_4449, w_093_4453, w_093_4455, w_093_4470, w_093_4476, w_093_4481, w_093_4483, w_093_4487, w_093_4489, w_093_4490, w_093_4491, w_093_4497, w_093_4498, w_093_4503, w_093_4505, w_093_4513, w_093_4517, w_093_4520, w_093_4521, w_093_4528, w_093_4533, w_093_4534, w_093_4539, w_093_4548, w_093_4553, w_093_4554, w_093_4557, w_093_4558, w_093_4566, w_093_4571, w_093_4582, w_093_4587, w_093_4600, w_093_4609, w_093_4610, w_093_4613, w_093_4614, w_093_4619, w_093_4625, w_093_4631, w_093_4634, w_093_4635, w_093_4645, w_093_4648, w_093_4656, w_093_4657, w_093_4659, w_093_4660, w_093_4671, w_093_4673, w_093_4674, w_093_4676, w_093_4686, w_093_4700, w_093_4703, w_093_4704, w_093_4706, w_093_4711, w_093_4713, w_093_4714, w_093_4719, w_093_4722, w_093_4725, w_093_4729, w_093_4736, w_093_4738, w_093_4742, w_093_4745, w_093_4749, w_093_4751, w_093_4756, w_093_4757, w_093_4758, w_093_4764, w_093_4768, w_093_4769, w_093_4774, w_093_4777, w_093_4778, w_093_4786, w_093_4789, w_093_4795, w_093_4802, w_093_4807, w_093_4815, w_093_4816, w_093_4824, w_093_4830, w_093_4831, w_093_4836, w_093_4841, w_093_4845, w_093_4846, w_093_4847, w_093_4857, w_093_4858, w_093_4859, w_093_4872, w_093_4879, w_093_4884, w_093_4887, w_093_4888, w_093_4889, w_093_4893, w_093_4897, w_093_4898, w_093_4900, w_093_4902, w_093_4903, w_093_4910, w_093_4919, w_093_4920, w_093_4924, w_093_4931, w_093_4936, w_093_4937, w_093_4942, w_093_4948, w_093_4951, w_093_4953, w_093_4954, w_093_4956, w_093_4958, w_093_4960, w_093_4966, w_093_4969, w_093_4981, w_093_4985, w_093_4992, w_093_5000, w_093_5006, w_093_5007, w_093_5009, w_093_5021, w_093_5026, w_093_5027, w_093_5031, w_093_5035, w_093_5039, w_093_5047, w_093_5050, w_093_5056, w_093_5060, w_093_5061, w_093_5070, w_093_5071, w_093_5078, w_093_5080, w_093_5082, w_093_5087, w_093_5088, w_093_5095, w_093_5096, w_093_5106, w_093_5111, w_093_5114, w_093_5122, w_093_5123, w_093_5126, w_093_5139, w_093_5141, w_093_5145, w_093_5148, w_093_5154, w_093_5159, w_093_5160, w_093_5161, w_093_5164, w_093_5169, w_093_5170, w_093_5171, w_093_5174, w_093_5176, w_093_5180, w_093_5188, w_093_5194, w_093_5196, w_093_5199, w_093_5204, w_093_5207, w_093_5208, w_093_5210, w_093_5213, w_093_5214, w_093_5216, w_093_5220, w_093_5223, w_093_5226, w_093_5228, w_093_5231, w_093_5233, w_093_5236, w_093_5240, w_093_5243, w_093_5247, w_093_5248, w_093_5249, w_093_5252, w_093_5265, w_093_5267, w_093_5268, w_093_5274, w_093_5279, w_093_5282, w_093_5284, w_093_5286, w_093_5289, w_093_5290, w_093_5300, w_093_5301, w_093_5306, w_093_5308, w_093_5318, w_093_5331, w_093_5333, w_093_5338, w_093_5339, w_093_5342, w_093_5354, w_093_5359, w_093_5364, w_093_5366, w_093_5370, w_093_5377, w_093_5380, w_093_5385, w_093_5390, w_093_5411, w_093_5412, w_093_5413, w_093_5421, w_093_5429, w_093_5430, w_093_5431, w_093_5432, w_093_5434, w_093_5435, w_093_5440, w_093_5441, w_093_5442, w_093_5444, w_093_5450, w_093_5451, w_093_5456, w_093_5461, w_093_5463, w_093_5470, w_093_5471, w_093_5472, w_093_5478, w_093_5483, w_093_5489, w_093_5494, w_093_5498, w_093_5499, w_093_5510, w_093_5511, w_093_5512, w_093_5521, w_093_5524, w_093_5530, w_093_5532, w_093_5536, w_093_5547, w_093_5549, w_093_5557, w_093_5569, w_093_5570, w_093_5572, w_093_5575, w_093_5579, w_093_5585, w_093_5589, w_093_5590, w_093_5592, w_093_5593, w_093_5596, w_093_5597, w_093_5610, w_093_5617, w_093_5618, w_093_5624, w_093_5629, w_093_5641, w_093_5642, w_093_5647, w_093_5649, w_093_5650, w_093_5656, w_093_5665, w_093_5668, w_093_5674, w_093_5678, w_093_5682, w_093_5683, w_093_5684, w_093_5691, w_093_5692, w_093_5695, w_093_5702, w_093_5707, w_093_5711, w_093_5712, w_093_5714, w_093_5721, w_093_5725, w_093_5729, w_093_5730, w_093_5742, w_093_5743, w_093_5744, w_093_5747, w_093_5755, w_093_5757, w_093_5777, w_093_5786, w_093_5789, w_093_5799, w_093_5808, w_093_5819, w_093_5825, w_093_5826, w_093_5830, w_093_5834, w_093_5841, w_093_5845, w_093_5846, w_093_5847, w_093_5849, w_093_5851, w_093_5852, w_093_5853, w_093_5863, w_093_5872, w_093_5877, w_093_5890, w_093_5892, w_093_5893, w_093_5896, w_093_5900, w_093_5901, w_093_5902, w_093_5903, w_093_5905, w_093_5912, w_093_5913, w_093_5914, w_093_5916, w_093_5917, w_093_5919, w_093_5920, w_093_5921, w_093_5926, w_093_5931, w_093_5936, w_093_5937, w_093_5945, w_093_5946, w_093_5949, w_093_5951, w_093_5954, w_093_5959, w_093_5966, w_093_5968, w_093_5969, w_093_5980, w_093_5985, w_093_5987, w_093_5989, w_093_5990, w_093_5991, w_093_5996, w_093_5999, w_093_6004, w_093_6007, w_093_6009, w_093_6016, w_093_6017, w_093_6022, w_093_6025, w_093_6030, w_093_6031, w_093_6039, w_093_6050, w_093_6051, w_093_6056, w_093_6060, w_093_6066, w_093_6069, w_093_6080, w_093_6084, w_093_6085, w_093_6087, w_093_6094, w_093_6101, w_093_6102, w_093_6113, w_093_6114, w_093_6119, w_093_6125, w_093_6127, w_093_6138, w_093_6139, w_093_6143, w_093_6148, w_093_6149, w_093_6153, w_093_6155, w_093_6157, w_093_6159, w_093_6164, w_093_6166, w_093_6169, w_093_6172, w_093_6174, w_093_6183, w_093_6186, w_093_6189, w_093_6197, w_093_6225, w_093_6226, w_093_6233, w_093_6235, w_093_6237, w_093_6245, w_093_6246, w_093_6247, w_093_6248, w_093_6249, w_093_6259, w_093_6261, w_093_6263, w_093_6264, w_093_6265, w_093_6267, w_093_6271, w_093_6272, w_093_6278, w_093_6280, w_093_6285, w_093_6291, w_093_6300, w_093_6309, w_093_6315, w_093_6324, w_093_6325, w_093_6338, w_093_6340, w_093_6348, w_093_6349, w_093_6350, w_093_6355, w_093_6356, w_093_6359, w_093_6361, w_093_6364, w_093_6366, w_093_6367, w_093_6375, w_093_6384, w_093_6392, w_093_6393, w_093_6397, w_093_6398, w_093_6399, w_093_6403, w_093_6405, w_093_6413, w_093_6421, w_093_6425, w_093_6432, w_093_6433, w_093_6438, w_093_6439, w_093_6445, w_093_6451, w_093_6454, w_093_6455, w_093_6456, w_093_6464, w_093_6469, w_093_6473, w_093_6476, w_093_6480, w_093_6485, w_093_6493, w_093_6497, w_093_6504, w_093_6505, w_093_6506, w_093_6507, w_093_6522, w_093_6528, w_093_6533, w_093_6535, w_093_6537, w_093_6539, w_093_6541, w_093_6544, w_093_6549, w_093_6552, w_093_6555, w_093_6564, w_093_6575, w_093_6578, w_093_6579, w_093_6582, w_093_6583, w_093_6586, w_093_6590, w_093_6595, w_093_6600, w_093_6623, w_093_6624, w_093_6626, w_093_6627, w_093_6647, w_093_6656, w_093_6670, w_093_6673, w_093_6675, w_093_6677, w_093_6679, w_093_6680, w_093_6682, w_093_6684, w_093_6687, w_093_6689, w_093_6692, w_093_6694, w_093_6713, w_093_6724, w_093_6725, w_093_6728, w_093_6734, w_093_6737, w_093_6739, w_093_6740, w_093_6746, w_093_6751, w_093_6766, w_093_6771, w_093_6778, w_093_6786, w_093_6792, w_093_6801, w_093_6808, w_093_6816, w_093_6817, w_093_6820, w_093_6821, w_093_6823, w_093_6831, w_093_6833, w_093_6834, w_093_6835, w_093_6837, w_093_6839, w_093_6844, w_093_6847, w_093_6852, w_093_6854, w_093_6856, w_093_6858, w_093_6868, w_093_6871, w_093_6873, w_093_6875, w_093_6876, w_093_6880, w_093_6887, w_093_6888, w_093_6893, w_093_6899, w_093_6903, w_093_6906, w_093_6907, w_093_6909, w_093_6910, w_093_6911, w_093_6912, w_093_6916, w_093_6917, w_093_6920, w_093_6921, w_093_6925, w_093_6926, w_093_6930, w_093_6932, w_093_6941, w_093_6945, w_093_6947, w_093_6952, w_093_6967, w_093_6973, w_093_6974, w_093_6977, w_093_6980, w_093_6983, w_093_6991, w_093_6992, w_093_6993, w_093_6994, w_093_7011, w_093_7013, w_093_7016, w_093_7019, w_093_7023, w_093_7024, w_093_7026, w_093_7035, w_093_7039, w_093_7041, w_093_7054, w_093_7055, w_093_7056, w_093_7069, w_093_7073, w_093_7077, w_093_7084, w_093_7089, w_093_7091, w_093_7094, w_093_7095, w_093_7098, w_093_7106, w_093_7113, w_093_7117, w_093_7118, w_093_7121, w_093_7123, w_093_7128, w_093_7129, w_093_7135, w_093_7136, w_093_7137, w_093_7139, w_093_7140, w_093_7141, w_093_7146, w_093_7156, w_093_7165, w_093_7167, w_093_7179, w_093_7181, w_093_7189, w_093_7190, w_093_7191, w_093_7192, w_093_7202, w_093_7203, w_093_7208, w_093_7212, w_093_7231, w_093_7241, w_093_7242, w_093_7252, w_093_7253, w_093_7259, w_093_7269, w_093_7279, w_093_7286, w_093_7287, w_093_7289, w_093_7291, w_093_7292, w_093_7301, w_093_7302, w_093_7305, w_093_7309, w_093_7310, w_093_7320, w_093_7321, w_093_7333, w_093_7338, w_093_7346, w_093_7349, w_093_7359, w_093_7360, w_093_7368, w_093_7369, w_093_7372, w_093_7377, w_093_7381, w_093_7386, w_093_7399, w_093_7403, w_093_7405, w_093_7406, w_093_7409, w_093_7412, w_093_7413, w_093_7417, w_093_7425, w_093_7426, w_093_7434, w_093_7441, w_093_7451, w_093_7461, w_093_7463, w_093_7464, w_093_7466, w_093_7467, w_093_7468, w_093_7470, w_093_7475, w_093_7478, w_093_7480, w_093_7481, w_093_7492, w_093_7493, w_093_7495, w_093_7498, w_093_7499, w_093_7503, w_093_7522, w_093_7525, w_093_7527, w_093_7529, w_093_7532, w_093_7534, w_093_7535, w_093_7537, w_093_7539;
  wire w_094_001, w_094_002, w_094_003, w_094_004, w_094_008, w_094_009, w_094_011, w_094_012, w_094_016, w_094_017, w_094_018, w_094_020, w_094_021, w_094_022, w_094_023, w_094_024, w_094_026, w_094_027, w_094_028, w_094_029, w_094_030, w_094_032, w_094_034, w_094_035, w_094_036, w_094_038, w_094_039, w_094_041, w_094_042, w_094_045, w_094_047, w_094_050, w_094_051, w_094_052, w_094_054, w_094_055, w_094_056, w_094_059, w_094_061, w_094_064, w_094_067, w_094_068, w_094_069, w_094_071, w_094_074, w_094_075, w_094_076, w_094_077, w_094_078, w_094_079, w_094_080, w_094_082, w_094_086, w_094_088, w_094_089, w_094_090, w_094_091, w_094_092, w_094_096, w_094_097, w_094_098, w_094_099, w_094_100, w_094_101, w_094_102, w_094_103, w_094_105, w_094_107, w_094_108, w_094_109, w_094_110, w_094_116, w_094_117, w_094_118, w_094_120, w_094_122, w_094_123, w_094_127, w_094_128, w_094_130, w_094_134, w_094_135, w_094_136, w_094_137, w_094_138, w_094_139, w_094_140, w_094_144, w_094_145, w_094_149, w_094_150, w_094_152, w_094_153, w_094_154, w_094_155, w_094_156, w_094_157, w_094_159, w_094_161, w_094_162, w_094_166, w_094_167, w_094_169, w_094_170, w_094_174, w_094_175, w_094_176, w_094_178, w_094_179, w_094_180, w_094_181, w_094_182, w_094_183, w_094_184, w_094_188, w_094_191, w_094_193, w_094_195, w_094_196, w_094_199, w_094_201, w_094_203, w_094_205, w_094_206, w_094_207, w_094_208, w_094_209, w_094_210, w_094_211, w_094_212, w_094_213, w_094_215, w_094_217, w_094_221, w_094_223, w_094_225, w_094_230, w_094_231, w_094_232, w_094_235, w_094_237, w_094_238, w_094_239, w_094_240, w_094_241, w_094_242, w_094_244, w_094_245, w_094_246, w_094_249, w_094_251, w_094_253, w_094_256, w_094_259, w_094_260, w_094_261, w_094_262, w_094_264, w_094_265, w_094_266, w_094_267, w_094_269, w_094_270, w_094_271, w_094_275, w_094_276, w_094_277, w_094_278, w_094_279, w_094_280, w_094_281, w_094_282, w_094_283, w_094_284, w_094_285, w_094_286, w_094_287, w_094_288, w_094_291, w_094_295, w_094_297, w_094_298, w_094_299, w_094_301, w_094_302, w_094_304, w_094_305, w_094_306, w_094_308, w_094_309, w_094_311, w_094_312, w_094_313, w_094_314, w_094_315, w_094_317, w_094_318, w_094_319, w_094_323, w_094_325, w_094_327, w_094_329, w_094_330, w_094_331, w_094_332, w_094_334, w_094_336, w_094_337, w_094_338, w_094_340, w_094_341, w_094_343, w_094_345, w_094_346, w_094_347, w_094_348, w_094_352, w_094_354, w_094_355, w_094_356, w_094_359, w_094_360, w_094_362, w_094_363, w_094_364, w_094_365, w_094_366, w_094_369, w_094_371, w_094_373, w_094_374, w_094_375, w_094_376, w_094_377, w_094_379, w_094_381, w_094_384, w_094_385, w_094_387, w_094_388, w_094_390, w_094_391, w_094_393, w_094_394, w_094_395, w_094_397, w_094_398, w_094_400, w_094_401, w_094_402, w_094_403, w_094_404, w_094_405, w_094_407, w_094_408, w_094_409, w_094_411, w_094_412, w_094_413, w_094_414, w_094_415, w_094_416, w_094_417, w_094_418, w_094_419, w_094_420, w_094_421, w_094_423, w_094_427, w_094_428, w_094_429, w_094_431, w_094_434, w_094_436, w_094_437, w_094_438, w_094_439, w_094_440, w_094_442, w_094_443, w_094_444, w_094_446, w_094_452, w_094_455, w_094_457, w_094_458, w_094_460, w_094_461, w_094_462, w_094_465, w_094_468, w_094_469, w_094_472, w_094_473, w_094_474, w_094_475, w_094_476, w_094_478, w_094_479, w_094_480, w_094_481, w_094_482, w_094_483, w_094_486, w_094_487, w_094_489, w_094_492, w_094_493, w_094_495, w_094_496, w_094_498, w_094_500, w_094_501, w_094_502, w_094_504, w_094_506, w_094_507, w_094_508, w_094_510, w_094_513, w_094_514, w_094_516, w_094_517, w_094_520, w_094_522, w_094_523, w_094_524, w_094_525, w_094_527, w_094_528, w_094_529, w_094_530, w_094_532, w_094_533, w_094_536, w_094_538, w_094_540, w_094_541, w_094_542, w_094_543, w_094_545, w_094_548, w_094_550, w_094_551, w_094_552, w_094_553, w_094_554, w_094_556, w_094_557, w_094_560, w_094_561, w_094_562, w_094_563, w_094_564, w_094_565, w_094_566, w_094_568, w_094_571, w_094_572, w_094_573, w_094_574, w_094_575, w_094_576, w_094_577, w_094_579, w_094_580, w_094_581, w_094_583, w_094_585, w_094_587, w_094_588, w_094_590, w_094_591, w_094_592, w_094_593, w_094_594, w_094_595, w_094_596, w_094_598, w_094_599, w_094_600, w_094_601, w_094_602, w_094_603, w_094_605, w_094_606, w_094_608, w_094_611, w_094_612, w_094_613, w_094_616, w_094_619, w_094_620, w_094_623, w_094_625, w_094_626, w_094_627, w_094_628, w_094_631, w_094_632, w_094_634, w_094_636, w_094_637, w_094_638, w_094_639, w_094_640, w_094_643, w_094_644, w_094_645, w_094_646, w_094_647, w_094_650, w_094_652, w_094_657, w_094_659, w_094_661, w_094_662, w_094_663, w_094_665, w_094_667, w_094_669, w_094_670, w_094_671, w_094_673, w_094_674, w_094_675, w_094_676, w_094_678, w_094_680, w_094_682, w_094_684, w_094_686, w_094_687, w_094_688, w_094_690, w_094_691, w_094_692, w_094_693, w_094_694, w_094_695, w_094_696, w_094_699, w_094_700, w_094_703, w_094_704, w_094_705, w_094_708, w_094_710, w_094_711, w_094_712, w_094_713, w_094_715, w_094_716, w_094_718, w_094_719, w_094_720, w_094_721, w_094_722, w_094_723, w_094_727, w_094_728, w_094_731, w_094_733, w_094_734, w_094_737, w_094_742, w_094_743, w_094_744, w_094_745, w_094_746, w_094_749, w_094_750, w_094_753, w_094_754, w_094_756, w_094_757, w_094_758, w_094_759, w_094_761, w_094_762, w_094_763, w_094_765, w_094_766, w_094_768, w_094_770, w_094_775, w_094_776, w_094_777, w_094_778, w_094_780, w_094_781, w_094_782, w_094_783, w_094_784, w_094_786, w_094_787, w_094_788, w_094_789, w_094_790, w_094_792, w_094_793, w_094_794, w_094_795, w_094_796, w_094_797, w_094_798, w_094_799, w_094_800, w_094_802, w_094_803, w_094_805, w_094_806, w_094_807, w_094_808, w_094_809, w_094_810, w_094_811, w_094_812, w_094_815, w_094_817, w_094_818, w_094_819, w_094_820, w_094_822, w_094_823, w_094_826, w_094_827, w_094_828, w_094_829, w_094_830, w_094_831, w_094_832, w_094_833, w_094_838, w_094_839, w_094_842, w_094_845, w_094_846, w_094_847, w_094_848, w_094_849, w_094_851, w_094_852, w_094_853, w_094_854, w_094_855, w_094_857, w_094_858, w_094_859, w_094_860, w_094_863, w_094_865, w_094_868, w_094_869, w_094_870, w_094_871, w_094_873, w_094_875, w_094_876, w_094_879, w_094_880, w_094_882, w_094_884, w_094_885, w_094_887, w_094_890, w_094_891, w_094_892, w_094_893, w_094_894, w_094_895, w_094_898, w_094_899, w_094_900, w_094_901, w_094_902, w_094_903, w_094_904, w_094_905, w_094_906, w_094_908, w_094_909, w_094_911, w_094_912, w_094_913, w_094_915, w_094_916, w_094_917, w_094_920, w_094_921, w_094_923, w_094_924, w_094_925, w_094_926, w_094_927, w_094_928, w_094_929, w_094_930, w_094_932, w_094_933, w_094_934, w_094_935, w_094_936, w_094_937, w_094_938, w_094_939, w_094_940, w_094_942, w_094_944, w_094_947, w_094_948, w_094_949, w_094_950, w_094_951, w_094_954, w_094_956, w_094_958, w_094_959, w_094_960, w_094_963, w_094_964, w_094_966, w_094_967, w_094_968, w_094_969, w_094_970, w_094_972, w_094_974, w_094_975, w_094_976, w_094_977, w_094_980, w_094_982, w_094_983, w_094_984, w_094_985, w_094_987, w_094_988, w_094_989, w_094_991, w_094_992, w_094_993, w_094_994, w_094_996, w_094_997, w_094_999, w_094_1000, w_094_1002, w_094_1004, w_094_1005, w_094_1007, w_094_1008, w_094_1009, w_094_1010, w_094_1011, w_094_1012, w_094_1013, w_094_1015, w_094_1018, w_094_1019, w_094_1024, w_094_1025, w_094_1027, w_094_1028, w_094_1029, w_094_1032, w_094_1033, w_094_1036, w_094_1041, w_094_1042, w_094_1044, w_094_1045, w_094_1047, w_094_1048, w_094_1050, w_094_1052, w_094_1053, w_094_1054, w_094_1057, w_094_1061, w_094_1063, w_094_1064, w_094_1067, w_094_1068, w_094_1069, w_094_1070, w_094_1071, w_094_1072, w_094_1073, w_094_1074, w_094_1077, w_094_1078, w_094_1080, w_094_1081, w_094_1084, w_094_1085, w_094_1086, w_094_1088, w_094_1089, w_094_1090, w_094_1091, w_094_1093, w_094_1095, w_094_1096, w_094_1097, w_094_1098, w_094_1100, w_094_1102, w_094_1105, w_094_1106, w_094_1108, w_094_1109, w_094_1110, w_094_1113, w_094_1114, w_094_1116, w_094_1119, w_094_1121, w_094_1122, w_094_1123, w_094_1124, w_094_1125, w_094_1126, w_094_1127, w_094_1128, w_094_1129, w_094_1130, w_094_1131, w_094_1132, w_094_1139, w_094_1140, w_094_1143, w_094_1144, w_094_1145, w_094_1146, w_094_1147, w_094_1148, w_094_1149, w_094_1150, w_094_1151, w_094_1152, w_094_1153, w_094_1154, w_094_1155, w_094_1157, w_094_1158, w_094_1159, w_094_1162, w_094_1164, w_094_1165, w_094_1166, w_094_1167, w_094_1168, w_094_1170, w_094_1171, w_094_1172, w_094_1173, w_094_1176, w_094_1177, w_094_1179, w_094_1180, w_094_1181, w_094_1184, w_094_1185, w_094_1187, w_094_1188, w_094_1189, w_094_1190, w_094_1191, w_094_1192, w_094_1193, w_094_1198, w_094_1199, w_094_1202, w_094_1203, w_094_1204, w_094_1205, w_094_1207, w_094_1208, w_094_1209, w_094_1210, w_094_1212, w_094_1213, w_094_1215, w_094_1216, w_094_1217, w_094_1219, w_094_1220, w_094_1221, w_094_1222, w_094_1223, w_094_1225, w_094_1226, w_094_1227, w_094_1228, w_094_1229, w_094_1231, w_094_1232, w_094_1234, w_094_1236, w_094_1237, w_094_1238, w_094_1239, w_094_1240, w_094_1242, w_094_1245, w_094_1248, w_094_1249, w_094_1250, w_094_1251, w_094_1252, w_094_1253, w_094_1254, w_094_1255, w_094_1257, w_094_1258, w_094_1260, w_094_1262, w_094_1264, w_094_1269, w_094_1271, w_094_1272, w_094_1274, w_094_1275, w_094_1276, w_094_1278, w_094_1279, w_094_1280, w_094_1282, w_094_1284, w_094_1285, w_094_1286, w_094_1287, w_094_1290, w_094_1293, w_094_1294, w_094_1295, w_094_1296, w_094_1297, w_094_1299, w_094_1301, w_094_1302, w_094_1317, w_094_1319, w_094_1320, w_094_1321, w_094_1323, w_094_1324, w_094_1325, w_094_1326, w_094_1327, w_094_1328, w_094_1331, w_094_1332, w_094_1333, w_094_1336, w_094_1338, w_094_1339, w_094_1340, w_094_1342, w_094_1343, w_094_1344, w_094_1345, w_094_1346, w_094_1347, w_094_1349, w_094_1350, w_094_1351, w_094_1355, w_094_1356, w_094_1357, w_094_1359, w_094_1361, w_094_1362, w_094_1364, w_094_1365, w_094_1368, w_094_1369, w_094_1370, w_094_1372, w_094_1373, w_094_1374, w_094_1375, w_094_1376, w_094_1378, w_094_1379, w_094_1383, w_094_1384, w_094_1385, w_094_1386, w_094_1388, w_094_1391, w_094_1392, w_094_1395, w_094_1398, w_094_1399, w_094_1401, w_094_1404, w_094_1405, w_094_1406, w_094_1407, w_094_1408, w_094_1409, w_094_1413, w_094_1415, w_094_1417, w_094_1421, w_094_1422, w_094_1423, w_094_1424, w_094_1426, w_094_1427, w_094_1432, w_094_1434, w_094_1435, w_094_1439, w_094_1440, w_094_1441, w_094_1443, w_094_1444, w_094_1447, w_094_1449, w_094_1450, w_094_1451, w_094_1454, w_094_1455, w_094_1457, w_094_1458, w_094_1459, w_094_1461, w_094_1463, w_094_1464, w_094_1465, w_094_1466, w_094_1467, w_094_1468, w_094_1471, w_094_1472, w_094_1474, w_094_1479, w_094_1480, w_094_1484, w_094_1490, w_094_1492, w_094_1493, w_094_1495, w_094_1496, w_094_1497, w_094_1499, w_094_1501, w_094_1502, w_094_1503, w_094_1505, w_094_1506, w_094_1509, w_094_1510, w_094_1512, w_094_1514, w_094_1515, w_094_1516, w_094_1518, w_094_1521, w_094_1523, w_094_1525, w_094_1526, w_094_1527, w_094_1528, w_094_1531, w_094_1533, w_094_1535, w_094_1536, w_094_1537, w_094_1540, w_094_1541, w_094_1542, w_094_1543, w_094_1544, w_094_1546, w_094_1548, w_094_1550, w_094_1551, w_094_1555, w_094_1556, w_094_1558, w_094_1563, w_094_1564, w_094_1565, w_094_1566, w_094_1568, w_094_1570, w_094_1572, w_094_1573, w_094_1574, w_094_1575, w_094_1580, w_094_1582, w_094_1585, w_094_1586, w_094_1593, w_094_1595, w_094_1599, w_094_1602, w_094_1603, w_094_1604, w_094_1607, w_094_1611, w_094_1612, w_094_1613, w_094_1614, w_094_1615, w_094_1617, w_094_1619, w_094_1620, w_094_1621, w_094_1624, w_094_1625, w_094_1626, w_094_1627, w_094_1629, w_094_1633, w_094_1634, w_094_1639, w_094_1640, w_094_1643, w_094_1644, w_094_1645, w_094_1648, w_094_1650, w_094_1652, w_094_1653, w_094_1654, w_094_1655, w_094_1656, w_094_1657, w_094_1658, w_094_1660, w_094_1662, w_094_1664, w_094_1665, w_094_1666, w_094_1667, w_094_1673, w_094_1675, w_094_1676, w_094_1681, w_094_1683, w_094_1689, w_094_1690, w_094_1691, w_094_1692, w_094_1694, w_094_1698, w_094_1699, w_094_1700, w_094_1701, w_094_1705, w_094_1706, w_094_1707, w_094_1709, w_094_1711, w_094_1714, w_094_1716, w_094_1717, w_094_1720, w_094_1721, w_094_1722, w_094_1723, w_094_1725, w_094_1727, w_094_1731, w_094_1734, w_094_1735, w_094_1736, w_094_1737, w_094_1738, w_094_1742, w_094_1745, w_094_1746, w_094_1747, w_094_1751, w_094_1752, w_094_1754, w_094_1757, w_094_1759, w_094_1761, w_094_1762, w_094_1764, w_094_1765, w_094_1766, w_094_1767, w_094_1768, w_094_1769, w_094_1770, w_094_1771, w_094_1780, w_094_1781, w_094_1783, w_094_1785, w_094_1786, w_094_1788, w_094_1790, w_094_1791, w_094_1792, w_094_1795, w_094_1796, w_094_1797, w_094_1799, w_094_1801, w_094_1802, w_094_1804, w_094_1805, w_094_1807, w_094_1808, w_094_1809, w_094_1811, w_094_1812, w_094_1813, w_094_1814, w_094_1815, w_094_1816, w_094_1820, w_094_1821, w_094_1822, w_094_1823, w_094_1825, w_094_1826, w_094_1829, w_094_1830, w_094_1832, w_094_1834, w_094_1835, w_094_1836, w_094_1837, w_094_1838, w_094_1839, w_094_1840, w_094_1841, w_094_1843, w_094_1844, w_094_1845, w_094_1847, w_094_1848, w_094_1851, w_094_1853, w_094_1854, w_094_1856, w_094_1858, w_094_1859, w_094_1860, w_094_1861, w_094_1862, w_094_1864, w_094_1865, w_094_1868, w_094_1869, w_094_1870, w_094_1872, w_094_1874, w_094_1875, w_094_1877, w_094_1878, w_094_1879, w_094_1882, w_094_1883, w_094_1884, w_094_1885, w_094_1887, w_094_1888, w_094_1889, w_094_1890, w_094_1891, w_094_1892, w_094_1896, w_094_1898, w_094_1899, w_094_1900, w_094_1901, w_094_1902, w_094_1903, w_094_1905, w_094_1906, w_094_1907, w_094_1908, w_094_1909, w_094_1910, w_094_1912, w_094_1913, w_094_1914, w_094_1917, w_094_1918, w_094_1921, w_094_1922, w_094_1923, w_094_1925, w_094_1927, w_094_1928, w_094_1931, w_094_1932, w_094_1934, w_094_1936, w_094_1938, w_094_1939, w_094_1940, w_094_1942, w_094_1943, w_094_1947, w_094_1948, w_094_1949, w_094_1950, w_094_1956, w_094_1959, w_094_1961, w_094_1963, w_094_1964, w_094_1965, w_094_1968, w_094_1969, w_094_1973, w_094_1975, w_094_1977, w_094_1982, w_094_1983, w_094_1984, w_094_1987, w_094_1988, w_094_1989, w_094_1990, w_094_1991, w_094_1993, w_094_1994, w_094_1996, w_094_1998, w_094_1999, w_094_2001, w_094_2002, w_094_2003, w_094_2004, w_094_2005, w_094_2010, w_094_2012, w_094_2014, w_094_2016, w_094_2019, w_094_2021, w_094_2022, w_094_2024, w_094_2025, w_094_2027, w_094_2029, w_094_2030, w_094_2033, w_094_2034, w_094_2035, w_094_2036, w_094_2037, w_094_2040, w_094_2041, w_094_2043, w_094_2045, w_094_2047, w_094_2048, w_094_2052, w_094_2056, w_094_2058, w_094_2059, w_094_2062, w_094_2063, w_094_2066, w_094_2067, w_094_2068, w_094_2071, w_094_2072, w_094_2074, w_094_2076, w_094_2083, w_094_2087, w_094_2088, w_094_2091, w_094_2093, w_094_2095, w_094_2098, w_094_2099, w_094_2100, w_094_2101, w_094_2102, w_094_2103, w_094_2104, w_094_2105, w_094_2106, w_094_2108, w_094_2110, w_094_2111, w_094_2114, w_094_2115, w_094_2117, w_094_2118, w_094_2119, w_094_2121, w_094_2122, w_094_2126, w_094_2127, w_094_2128, w_094_2130, w_094_2131, w_094_2134, w_094_2135, w_094_2137, w_094_2138, w_094_2139, w_094_2141, w_094_2145, w_094_2148, w_094_2150, w_094_2151, w_094_2152, w_094_2154, w_094_2156, w_094_2160, w_094_2162, w_094_2163, w_094_2165, w_094_2167, w_094_2168, w_094_2169, w_094_2170, w_094_2171, w_094_2173, w_094_2174, w_094_2177, w_094_2178, w_094_2179, w_094_2180, w_094_2182, w_094_2183, w_094_2184, w_094_2186, w_094_2188, w_094_2189, w_094_2190, w_094_2191, w_094_2192, w_094_2193, w_094_2194, w_094_2197, w_094_2199, w_094_2202, w_094_2203, w_094_2205, w_094_2206, w_094_2208, w_094_2209, w_094_2212, w_094_2214, w_094_2215, w_094_2218, w_094_2219, w_094_2221, w_094_2222, w_094_2223, w_094_2225, w_094_2227, w_094_2230, w_094_2231, w_094_2233, w_094_2234, w_094_2236, w_094_2238, w_094_2242, w_094_2246, w_094_2247, w_094_2249, w_094_2250, w_094_2251, w_094_2254, w_094_2257, w_094_2258, w_094_2259, w_094_2261, w_094_2263, w_094_2267, w_094_2270, w_094_2273, w_094_2274, w_094_2277, w_094_2281, w_094_2282, w_094_2283, w_094_2284, w_094_2285, w_094_2287, w_094_2289, w_094_2290, w_094_2291, w_094_2292, w_094_2293, w_094_2296, w_094_2298, w_094_2299, w_094_2302, w_094_2304, w_094_2307, w_094_2310, w_094_2311, w_094_2313, w_094_2315, w_094_2316, w_094_2318, w_094_2319, w_094_2320, w_094_2321, w_094_2323, w_094_2325, w_094_2327, w_094_2329, w_094_2330, w_094_2333, w_094_2335, w_094_2336, w_094_2337, w_094_2338, w_094_2339, w_094_2343, w_094_2350, w_094_2357, w_094_2360, w_094_2362, w_094_2363, w_094_2364, w_094_2368, w_094_2370, w_094_2371, w_094_2372, w_094_2374, w_094_2376, w_094_2377, w_094_2379, w_094_2380, w_094_2381, w_094_2382, w_094_2384, w_094_2385, w_094_2389, w_094_2390, w_094_2391, w_094_2393, w_094_2397, w_094_2399, w_094_2401, w_094_2402, w_094_2403, w_094_2406, w_094_2408, w_094_2411, w_094_2413, w_094_2414, w_094_2415, w_094_2418, w_094_2419, w_094_2421, w_094_2422, w_094_2424, w_094_2426, w_094_2428, w_094_2433, w_094_2434, w_094_2436, w_094_2437, w_094_2438, w_094_2439, w_094_2442, w_094_2444, w_094_2445, w_094_2448, w_094_2449, w_094_2450, w_094_2452, w_094_2454, w_094_2455, w_094_2456, w_094_2457, w_094_2458, w_094_2461, w_094_2463, w_094_2468, w_094_2469, w_094_2470, w_094_2471, w_094_2479, w_094_2482, w_094_2485, w_094_2486, w_094_2488, w_094_2489, w_094_2492, w_094_2493, w_094_2496, w_094_2497, w_094_2498, w_094_2503, w_094_2505, w_094_2507, w_094_2508, w_094_2510, w_094_2512, w_094_2513, w_094_2514, w_094_2515, w_094_2517, w_094_2518, w_094_2519, w_094_2520, w_094_2526, w_094_2527, w_094_2528, w_094_2529, w_094_2533, w_094_2534, w_094_2535, w_094_2536, w_094_2538, w_094_2539, w_094_2541, w_094_2542, w_094_2545, w_094_2550, w_094_2551, w_094_2552, w_094_2556, w_094_2558, w_094_2559, w_094_2564, w_094_2566, w_094_2568, w_094_2569, w_094_2570, w_094_2571, w_094_2576, w_094_2577, w_094_2579, w_094_2580, w_094_2584, w_094_2585, w_094_2586, w_094_2587, w_094_2589, w_094_2592, w_094_2593, w_094_2595, w_094_2598, w_094_2599, w_094_2600, w_094_2602, w_094_2604, w_094_2605, w_094_2606, w_094_2607, w_094_2613, w_094_2616, w_094_2617, w_094_2621, w_094_2622, w_094_2625, w_094_2627, w_094_2628, w_094_2630, w_094_2631, w_094_2632, w_094_2637, w_094_2639, w_094_2640, w_094_2641, w_094_2643, w_094_2646, w_094_2647, w_094_2648, w_094_2649, w_094_2650, w_094_2654, w_094_2655, w_094_2656, w_094_2660, w_094_2661, w_094_2664, w_094_2665, w_094_2667, w_094_2668, w_094_2669, w_094_2670, w_094_2671, w_094_2674, w_094_2675, w_094_2676, w_094_2678, w_094_2679, w_094_2680, w_094_2681, w_094_2682, w_094_2683, w_094_2687, w_094_2690, w_094_2691, w_094_2692, w_094_2694, w_094_2695, w_094_2696, w_094_2697, w_094_2699, w_094_2703, w_094_2705, w_094_2706, w_094_2708, w_094_2709, w_094_2711, w_094_2712, w_094_2715, w_094_2718, w_094_2719, w_094_2720, w_094_2721, w_094_2722, w_094_2726, w_094_2727, w_094_2728, w_094_2730, w_094_2731, w_094_2734, w_094_2738, w_094_2740, w_094_2741, w_094_2742, w_094_2744, w_094_2745, w_094_2746, w_094_2748, w_094_2749, w_094_2750, w_094_2757, w_094_2758, w_094_2761, w_094_2763, w_094_2767, w_094_2768, w_094_2769, w_094_2770, w_094_2771, w_094_2772, w_094_2773, w_094_2776, w_094_2777, w_094_2779, w_094_2781, w_094_2782, w_094_2783, w_094_2787, w_094_2791, w_094_2793, w_094_2794, w_094_2797, w_094_2799, w_094_2800, w_094_2802, w_094_2804, w_094_2806, w_094_2809, w_094_2810, w_094_2811, w_094_2813, w_094_2814, w_094_2818, w_094_2820, w_094_2821, w_094_2822, w_094_2824, w_094_2826, w_094_2828, w_094_2834, w_094_2835, w_094_2836, w_094_2837, w_094_2838, w_094_2839, w_094_2840, w_094_2843, w_094_2845, w_094_2847, w_094_2849, w_094_2850, w_094_2852, w_094_2855, w_094_2856, w_094_2857, w_094_2858, w_094_2860, w_094_2861, w_094_2862, w_094_2865;
  wire w_095_001, w_095_003, w_095_004, w_095_005, w_095_006, w_095_009, w_095_010, w_095_015, w_095_016, w_095_017, w_095_021, w_095_025, w_095_028, w_095_029, w_095_030, w_095_031, w_095_032, w_095_034, w_095_037, w_095_040, w_095_041, w_095_042, w_095_044, w_095_045, w_095_047, w_095_048, w_095_049, w_095_051, w_095_053, w_095_055, w_095_058, w_095_059, w_095_061, w_095_063, w_095_065, w_095_067, w_095_068, w_095_069, w_095_070, w_095_072, w_095_073, w_095_075, w_095_076, w_095_079, w_095_086, w_095_089, w_095_092, w_095_093, w_095_099, w_095_102, w_095_103, w_095_104, w_095_107, w_095_108, w_095_109, w_095_111, w_095_112, w_095_113, w_095_116, w_095_118, w_095_120, w_095_121, w_095_128, w_095_129, w_095_130, w_095_132, w_095_133, w_095_134, w_095_137, w_095_139, w_095_140, w_095_145, w_095_146, w_095_147, w_095_148, w_095_152, w_095_153, w_095_154, w_095_155, w_095_162, w_095_164, w_095_167, w_095_171, w_095_172, w_095_173, w_095_176, w_095_177, w_095_178, w_095_179, w_095_180, w_095_182, w_095_184, w_095_187, w_095_189, w_095_190, w_095_193, w_095_195, w_095_198, w_095_203, w_095_204, w_095_205, w_095_206, w_095_209, w_095_211, w_095_212, w_095_213, w_095_214, w_095_215, w_095_216, w_095_219, w_095_224, w_095_225, w_095_227, w_095_229, w_095_231, w_095_232, w_095_233, w_095_235, w_095_237, w_095_238, w_095_239, w_095_240, w_095_241, w_095_244, w_095_246, w_095_249, w_095_250, w_095_252, w_095_255, w_095_257, w_095_259, w_095_261, w_095_264, w_095_265, w_095_272, w_095_273, w_095_274, w_095_275, w_095_276, w_095_277, w_095_278, w_095_279, w_095_280, w_095_284, w_095_290, w_095_292, w_095_293, w_095_294, w_095_295, w_095_297, w_095_298, w_095_299, w_095_300, w_095_301, w_095_302, w_095_304, w_095_308, w_095_309, w_095_310, w_095_312, w_095_315, w_095_317, w_095_319, w_095_321, w_095_323, w_095_328, w_095_330, w_095_331, w_095_333, w_095_334, w_095_336, w_095_337, w_095_338, w_095_342, w_095_343, w_095_344, w_095_345, w_095_346, w_095_349, w_095_351, w_095_354, w_095_355, w_095_359, w_095_360, w_095_361, w_095_362, w_095_363, w_095_365, w_095_367, w_095_368, w_095_369, w_095_370, w_095_372, w_095_373, w_095_375, w_095_376, w_095_378, w_095_379, w_095_380, w_095_381, w_095_383, w_095_388, w_095_389, w_095_390, w_095_391, w_095_394, w_095_395, w_095_398, w_095_399, w_095_400, w_095_401, w_095_402, w_095_404, w_095_406, w_095_414, w_095_415, w_095_417, w_095_420, w_095_423, w_095_425, w_095_430, w_095_431, w_095_433, w_095_434, w_095_439, w_095_440, w_095_443, w_095_445, w_095_447, w_095_448, w_095_449, w_095_450, w_095_452, w_095_455, w_095_457, w_095_458, w_095_459, w_095_460, w_095_462, w_095_465, w_095_466, w_095_467, w_095_468, w_095_469, w_095_470, w_095_471, w_095_473, w_095_474, w_095_475, w_095_477, w_095_478, w_095_480, w_095_481, w_095_483, w_095_485, w_095_486, w_095_488, w_095_491, w_095_492, w_095_493, w_095_494, w_095_496, w_095_498, w_095_502, w_095_504, w_095_506, w_095_507, w_095_509, w_095_511, w_095_512, w_095_514, w_095_515, w_095_517, w_095_520, w_095_521, w_095_523, w_095_524, w_095_525, w_095_526, w_095_531, w_095_534, w_095_535, w_095_537, w_095_538, w_095_539, w_095_540, w_095_541, w_095_545, w_095_547, w_095_549, w_095_550, w_095_552, w_095_559, w_095_560, w_095_563, w_095_567, w_095_568, w_095_571, w_095_574, w_095_578, w_095_580, w_095_582, w_095_583, w_095_584, w_095_588, w_095_589, w_095_590, w_095_591, w_095_592, w_095_593, w_095_595, w_095_597, w_095_598, w_095_599, w_095_600, w_095_602, w_095_603, w_095_605, w_095_606, w_095_611, w_095_612, w_095_613, w_095_614, w_095_616, w_095_618, w_095_620, w_095_624, w_095_627, w_095_629, w_095_630, w_095_632, w_095_635, w_095_639, w_095_644, w_095_645, w_095_650, w_095_653, w_095_654, w_095_655, w_095_656, w_095_658, w_095_659, w_095_660, w_095_661, w_095_663, w_095_664, w_095_666, w_095_667, w_095_668, w_095_671, w_095_677, w_095_680, w_095_685, w_095_686, w_095_689, w_095_690, w_095_692, w_095_693, w_095_698, w_095_699, w_095_701, w_095_705, w_095_706, w_095_707, w_095_708, w_095_711, w_095_712, w_095_713, w_095_714, w_095_717, w_095_718, w_095_719, w_095_722, w_095_723, w_095_726, w_095_729, w_095_730, w_095_732, w_095_733, w_095_735, w_095_737, w_095_738, w_095_740, w_095_747, w_095_749, w_095_750, w_095_752, w_095_753, w_095_754, w_095_755, w_095_757, w_095_758, w_095_759, w_095_760, w_095_761, w_095_762, w_095_763, w_095_764, w_095_765, w_095_768, w_095_769, w_095_772, w_095_774, w_095_775, w_095_776, w_095_777, w_095_779, w_095_780, w_095_781, w_095_782, w_095_785, w_095_786, w_095_788, w_095_793, w_095_794, w_095_795, w_095_796, w_095_798, w_095_799, w_095_801, w_095_804, w_095_805, w_095_807, w_095_809, w_095_810, w_095_813, w_095_816, w_095_817, w_095_818, w_095_819, w_095_821, w_095_823, w_095_824, w_095_826, w_095_831, w_095_833, w_095_835, w_095_836, w_095_837, w_095_838, w_095_839, w_095_843, w_095_845, w_095_847, w_095_848, w_095_850, w_095_851, w_095_853, w_095_854, w_095_856, w_095_858, w_095_859, w_095_864, w_095_865, w_095_866, w_095_869, w_095_871, w_095_875, w_095_876, w_095_877, w_095_878, w_095_881, w_095_884, w_095_889, w_095_893, w_095_894, w_095_896, w_095_898, w_095_900, w_095_901, w_095_904, w_095_905, w_095_906, w_095_909, w_095_911, w_095_912, w_095_913, w_095_914, w_095_915, w_095_916, w_095_917, w_095_918, w_095_919, w_095_920, w_095_921, w_095_923, w_095_924, w_095_928, w_095_929, w_095_930, w_095_932, w_095_936, w_095_937, w_095_938, w_095_942, w_095_943, w_095_944, w_095_945, w_095_946, w_095_947, w_095_948, w_095_949, w_095_951, w_095_952, w_095_955, w_095_958, w_095_961, w_095_963, w_095_964, w_095_965, w_095_966, w_095_968, w_095_969, w_095_970, w_095_972, w_095_973, w_095_974, w_095_975, w_095_977, w_095_980, w_095_981, w_095_983, w_095_986, w_095_988, w_095_989, w_095_990, w_095_995, w_095_998, w_095_999, w_095_1001, w_095_1002, w_095_1003, w_095_1004, w_095_1005, w_095_1007, w_095_1009, w_095_1010, w_095_1013, w_095_1016, w_095_1022, w_095_1023, w_095_1025, w_095_1026, w_095_1027, w_095_1028, w_095_1029, w_095_1030, w_095_1033, w_095_1034, w_095_1035, w_095_1039, w_095_1042, w_095_1044, w_095_1045, w_095_1047, w_095_1048, w_095_1049, w_095_1050, w_095_1051, w_095_1052, w_095_1054, w_095_1057, w_095_1058, w_095_1059, w_095_1061, w_095_1062, w_095_1064, w_095_1066, w_095_1068, w_095_1069, w_095_1070, w_095_1071, w_095_1073, w_095_1074, w_095_1075, w_095_1076, w_095_1079, w_095_1080, w_095_1084, w_095_1085, w_095_1086, w_095_1089, w_095_1091, w_095_1092, w_095_1095, w_095_1096, w_095_1097, w_095_1099, w_095_1100, w_095_1101, w_095_1102, w_095_1105, w_095_1106, w_095_1107, w_095_1109, w_095_1112, w_095_1113, w_095_1115, w_095_1116, w_095_1117, w_095_1118, w_095_1121, w_095_1122, w_095_1123, w_095_1127, w_095_1128, w_095_1132, w_095_1133, w_095_1139, w_095_1140, w_095_1142, w_095_1144, w_095_1146, w_095_1149, w_095_1151, w_095_1153, w_095_1154, w_095_1160, w_095_1161, w_095_1164, w_095_1171, w_095_1172, w_095_1173, w_095_1174, w_095_1175, w_095_1178, w_095_1179, w_095_1181, w_095_1182, w_095_1184, w_095_1186, w_095_1187, w_095_1189, w_095_1194, w_095_1196, w_095_1200, w_095_1201, w_095_1203, w_095_1207, w_095_1209, w_095_1210, w_095_1211, w_095_1212, w_095_1213, w_095_1214, w_095_1215, w_095_1216, w_095_1217, w_095_1222, w_095_1223, w_095_1224, w_095_1225, w_095_1227, w_095_1230, w_095_1231, w_095_1235, w_095_1236, w_095_1237, w_095_1238, w_095_1239, w_095_1249, w_095_1250, w_095_1251, w_095_1252, w_095_1253, w_095_1255, w_095_1256, w_095_1257, w_095_1259, w_095_1261, w_095_1262, w_095_1266, w_095_1267, w_095_1269, w_095_1270, w_095_1274, w_095_1275, w_095_1276, w_095_1277, w_095_1279, w_095_1280, w_095_1283, w_095_1285, w_095_1286, w_095_1287, w_095_1288, w_095_1290, w_095_1292, w_095_1294, w_095_1296, w_095_1299, w_095_1300, w_095_1302, w_095_1303, w_095_1304, w_095_1305, w_095_1307, w_095_1308, w_095_1309, w_095_1311, w_095_1312, w_095_1313, w_095_1316, w_095_1317, w_095_1318, w_095_1320, w_095_1322, w_095_1323, w_095_1325, w_095_1326, w_095_1327, w_095_1328, w_095_1330, w_095_1331, w_095_1332, w_095_1334, w_095_1337, w_095_1338, w_095_1339, w_095_1343, w_095_1345, w_095_1346, w_095_1354, w_095_1356, w_095_1357, w_095_1358, w_095_1359, w_095_1362, w_095_1363, w_095_1364, w_095_1365, w_095_1371, w_095_1372, w_095_1373, w_095_1374, w_095_1377, w_095_1378, w_095_1380, w_095_1383, w_095_1386, w_095_1387, w_095_1389, w_095_1393, w_095_1394, w_095_1396, w_095_1397, w_095_1398, w_095_1399, w_095_1401, w_095_1402, w_095_1403, w_095_1406, w_095_1408, w_095_1411, w_095_1414, w_095_1416, w_095_1417, w_095_1419, w_095_1421, w_095_1423, w_095_1425, w_095_1426, w_095_1427, w_095_1430, w_095_1432, w_095_1435, w_095_1436, w_095_1437, w_095_1440, w_095_1442, w_095_1444, w_095_1445, w_095_1448, w_095_1451, w_095_1452, w_095_1454, w_095_1456, w_095_1457, w_095_1461, w_095_1462, w_095_1463, w_095_1464, w_095_1466, w_095_1467, w_095_1468, w_095_1469, w_095_1472, w_095_1486, w_095_1487, w_095_1489, w_095_1490, w_095_1493, w_095_1494, w_095_1495, w_095_1496, w_095_1498, w_095_1500, w_095_1501, w_095_1504, w_095_1505, w_095_1509, w_095_1510, w_095_1512, w_095_1513, w_095_1515, w_095_1517, w_095_1520, w_095_1522, w_095_1525, w_095_1526, w_095_1527, w_095_1528, w_095_1529, w_095_1530, w_095_1532, w_095_1533, w_095_1536, w_095_1538, w_095_1540, w_095_1542, w_095_1544, w_095_1548, w_095_1550, w_095_1551, w_095_1552, w_095_1553, w_095_1554, w_095_1556, w_095_1559, w_095_1560, w_095_1561, w_095_1562, w_095_1563, w_095_1565, w_095_1566, w_095_1567, w_095_1568, w_095_1570, w_095_1571, w_095_1572, w_095_1575, w_095_1577, w_095_1581, w_095_1582, w_095_1583, w_095_1584, w_095_1585, w_095_1587, w_095_1590, w_095_1593, w_095_1596, w_095_1598, w_095_1599, w_095_1600, w_095_1601, w_095_1602, w_095_1603, w_095_1607, w_095_1608, w_095_1612, w_095_1613, w_095_1615, w_095_1616, w_095_1617, w_095_1618, w_095_1619, w_095_1626, w_095_1629, w_095_1632, w_095_1635, w_095_1638, w_095_1639, w_095_1643, w_095_1644, w_095_1645, w_095_1646, w_095_1647, w_095_1648, w_095_1649, w_095_1652, w_095_1654, w_095_1656, w_095_1657, w_095_1658, w_095_1659, w_095_1660, w_095_1661, w_095_1665, w_095_1666, w_095_1667, w_095_1668, w_095_1670, w_095_1671, w_095_1672, w_095_1673, w_095_1675, w_095_1676, w_095_1677, w_095_1679, w_095_1680, w_095_1681, w_095_1684, w_095_1685, w_095_1686, w_095_1688, w_095_1689, w_095_1690, w_095_1691, w_095_1692, w_095_1694, w_095_1695, w_095_1697, w_095_1698, w_095_1699, w_095_1700, w_095_1701, w_095_1703, w_095_1705, w_095_1707, w_095_1709, w_095_1712, w_095_1713, w_095_1714, w_095_1716, w_095_1720, w_095_1723, w_095_1724, w_095_1729, w_095_1731, w_095_1733, w_095_1735, w_095_1736, w_095_1737, w_095_1738, w_095_1739, w_095_1740, w_095_1741, w_095_1742, w_095_1744, w_095_1745, w_095_1747, w_095_1748, w_095_1749, w_095_1752, w_095_1753, w_095_1755, w_095_1756, w_095_1757, w_095_1760, w_095_1762, w_095_1764, w_095_1767, w_095_1769, w_095_1771, w_095_1774, w_095_1777, w_095_1779, w_095_1780, w_095_1783, w_095_1784, w_095_1785, w_095_1786, w_095_1787, w_095_1789, w_095_1791, w_095_1792, w_095_1793, w_095_1796, w_095_1798, w_095_1802, w_095_1806, w_095_1807, w_095_1814, w_095_1815, w_095_1817, w_095_1818, w_095_1820, w_095_1822, w_095_1823, w_095_1825, w_095_1826, w_095_1828, w_095_1830, w_095_1834, w_095_1835, w_095_1836, w_095_1837, w_095_1838, w_095_1840, w_095_1842, w_095_1843, w_095_1844, w_095_1847, w_095_1848, w_095_1852, w_095_1854, w_095_1857, w_095_1858, w_095_1863, w_095_1864, w_095_1867, w_095_1870, w_095_1872, w_095_1875, w_095_1876, w_095_1880, w_095_1881, w_095_1882, w_095_1884, w_095_1885, w_095_1887, w_095_1888, w_095_1889, w_095_1890, w_095_1893, w_095_1894, w_095_1895, w_095_1897, w_095_1903, w_095_1904, w_095_1908, w_095_1909, w_095_1913, w_095_1914, w_095_1915, w_095_1916, w_095_1917, w_095_1918, w_095_1923, w_095_1925, w_095_1929, w_095_1931, w_095_1933, w_095_1934, w_095_1935, w_095_1938, w_095_1939, w_095_1940, w_095_1941, w_095_1942, w_095_1943, w_095_1948, w_095_1949, w_095_1952, w_095_1955, w_095_1958, w_095_1959, w_095_1963, w_095_1964, w_095_1967, w_095_1969, w_095_1970, w_095_1971, w_095_1972, w_095_1973, w_095_1974, w_095_1975, w_095_1976, w_095_1978, w_095_1979, w_095_1981, w_095_1985, w_095_1986, w_095_1987, w_095_1989, w_095_1991, w_095_1993, w_095_1994, w_095_1996, w_095_1997, w_095_1998, w_095_1999, w_095_2000, w_095_2001, w_095_2003, w_095_2004, w_095_2007, w_095_2008, w_095_2009, w_095_2011, w_095_2012, w_095_2013, w_095_2015, w_095_2018, w_095_2019, w_095_2021, w_095_2022, w_095_2023, w_095_2026, w_095_2027, w_095_2029, w_095_2031, w_095_2032, w_095_2033, w_095_2034, w_095_2035, w_095_2036, w_095_2038, w_095_2039, w_095_2040, w_095_2042, w_095_2047, w_095_2048, w_095_2051, w_095_2053, w_095_2055, w_095_2056, w_095_2057, w_095_2059, w_095_2060, w_095_2061, w_095_2062, w_095_2068, w_095_2069, w_095_2070, w_095_2072, w_095_2074, w_095_2077, w_095_2078, w_095_2080, w_095_2082, w_095_2084, w_095_2085, w_095_2089, w_095_2090, w_095_2092, w_095_2093, w_095_2094, w_095_2095, w_095_2096, w_095_2097, w_095_2099, w_095_2100, w_095_2101, w_095_2103, w_095_2108, w_095_2109, w_095_2113, w_095_2114, w_095_2116, w_095_2120, w_095_2121, w_095_2123, w_095_2124, w_095_2125, w_095_2131, w_095_2132, w_095_2139, w_095_2140, w_095_2141, w_095_2145, w_095_2146, w_095_2147, w_095_2148, w_095_2153, w_095_2154, w_095_2155, w_095_2156, w_095_2158, w_095_2161, w_095_2162, w_095_2163, w_095_2164, w_095_2168, w_095_2173, w_095_2174, w_095_2175, w_095_2177, w_095_2178, w_095_2181, w_095_2182, w_095_2184, w_095_2186, w_095_2187, w_095_2188, w_095_2191, w_095_2192, w_095_2193, w_095_2195, w_095_2196, w_095_2197, w_095_2198, w_095_2199, w_095_2203, w_095_2204, w_095_2206, w_095_2208, w_095_2209, w_095_2211, w_095_2215, w_095_2217, w_095_2218, w_095_2220, w_095_2222, w_095_2223, w_095_2225, w_095_2228, w_095_2229, w_095_2231, w_095_2232, w_095_2237, w_095_2238, w_095_2240, w_095_2243, w_095_2244, w_095_2250, w_095_2252, w_095_2256, w_095_2257, w_095_2259, w_095_2261, w_095_2263, w_095_2264, w_095_2268, w_095_2269, w_095_2270, w_095_2271, w_095_2272, w_095_2273, w_095_2274, w_095_2275, w_095_2276, w_095_2277, w_095_2280, w_095_2281, w_095_2282, w_095_2284, w_095_2287, w_095_2288, w_095_2289, w_095_2291, w_095_2293, w_095_2294, w_095_2299, w_095_2304, w_095_2305, w_095_2306, w_095_2307, w_095_2310, w_095_2311, w_095_2315, w_095_2316, w_095_2317, w_095_2318, w_095_2321, w_095_2323, w_095_2325, w_095_2327, w_095_2330, w_095_2332, w_095_2336, w_095_2339, w_095_2342, w_095_2343, w_095_2344, w_095_2345, w_095_2346, w_095_2355, w_095_2356, w_095_2358, w_095_2359, w_095_2362, w_095_2365, w_095_2366, w_095_2367, w_095_2368, w_095_2369, w_095_2370, w_095_2371, w_095_2372, w_095_2373, w_095_2374, w_095_2375, w_095_2376, w_095_2379, w_095_2383, w_095_2384, w_095_2385, w_095_2386, w_095_2388, w_095_2389, w_095_2393, w_095_2394, w_095_2398, w_095_2399, w_095_2400, w_095_2404, w_095_2406, w_095_2407, w_095_2411, w_095_2412, w_095_2415, w_095_2416, w_095_2417, w_095_2418, w_095_2420, w_095_2422, w_095_2423, w_095_2424, w_095_2425, w_095_2427, w_095_2428, w_095_2430, w_095_2433, w_095_2436, w_095_2437, w_095_2438, w_095_2440, w_095_2441, w_095_2444, w_095_2446, w_095_2448, w_095_2449, w_095_2451, w_095_2452, w_095_2455, w_095_2456, w_095_2458, w_095_2459, w_095_2461, w_095_2462, w_095_2463, w_095_2464, w_095_2465, w_095_2467, w_095_2468, w_095_2469, w_095_2471, w_095_2472, w_095_2474, w_095_2475, w_095_2477, w_095_2478, w_095_2479, w_095_2483, w_095_2487, w_095_2489, w_095_2490, w_095_2491, w_095_2492, w_095_2493, w_095_2495, w_095_2496, w_095_2499, w_095_2500, w_095_2501, w_095_2502, w_095_2506, w_095_2508, w_095_2509, w_095_2511, w_095_2512, w_095_2513, w_095_2516, w_095_2517, w_095_2518, w_095_2519, w_095_2520, w_095_2521, w_095_2522, w_095_2523, w_095_2524, w_095_2525, w_095_2526, w_095_2527, w_095_2528, w_095_2529, w_095_2532, w_095_2534, w_095_2537, w_095_2538, w_095_2539, w_095_2540, w_095_2542, w_095_2543, w_095_2546, w_095_2548, w_095_2549, w_095_2550, w_095_2551, w_095_2553, w_095_2556, w_095_2558, w_095_2559, w_095_2561, w_095_2563, w_095_2565, w_095_2566, w_095_2567, w_095_2568, w_095_2569, w_095_2571, w_095_2573, w_095_2574, w_095_2575, w_095_2576, w_095_2577, w_095_2580, w_095_2581, w_095_2583, w_095_2585, w_095_2586, w_095_2588, w_095_2589, w_095_2590, w_095_2591, w_095_2592, w_095_2593, w_095_2595, w_095_2599, w_095_2600, w_095_2601, w_095_2603, w_095_2606, w_095_2607, w_095_2611, w_095_2612, w_095_2617, w_095_2618, w_095_2619, w_095_2620, w_095_2622, w_095_2623, w_095_2626, w_095_2628, w_095_2629, w_095_2630, w_095_2633, w_095_2635, w_095_2636, w_095_2639, w_095_2640, w_095_2641, w_095_2643, w_095_2644, w_095_2645, w_095_2646, w_095_2648, w_095_2650, w_095_2652, w_095_2653, w_095_2656, w_095_2657, w_095_2658, w_095_2663, w_095_2664, w_095_2666, w_095_2669, w_095_2670, w_095_2671, w_095_2672, w_095_2673, w_095_2677, w_095_2684, w_095_2685, w_095_2687, w_095_2688, w_095_2689, w_095_2691, w_095_2692, w_095_2694, w_095_2696, w_095_2697, w_095_2698, w_095_2699, w_095_2704, w_095_2710, w_095_2711, w_095_2713, w_095_2714, w_095_2719, w_095_2720, w_095_2726, w_095_2727, w_095_2730, w_095_2731, w_095_2732, w_095_2733, w_095_2736, w_095_2738, w_095_2739, w_095_2740, w_095_2741, w_095_2742, w_095_2744, w_095_2745, w_095_2748, w_095_2749, w_095_2751, w_095_2752, w_095_2755, w_095_2756, w_095_2757, w_095_2759, w_095_2761, w_095_2766, w_095_2767, w_095_2772, w_095_2774, w_095_2776, w_095_2778, w_095_2780, w_095_2781, w_095_2792, w_095_2793, w_095_2800, w_095_2803, w_095_2806, w_095_2807, w_095_2811, w_095_2816, w_095_2818, w_095_2823, w_095_2825, w_095_2826, w_095_2828, w_095_2832, w_095_2833, w_095_2834, w_095_2836, w_095_2837, w_095_2838, w_095_2839, w_095_2841, w_095_2844, w_095_2845, w_095_2848, w_095_2851, w_095_2857, w_095_2859, w_095_2860, w_095_2863, w_095_2865, w_095_2871, w_095_2875, w_095_2876, w_095_2878, w_095_2883, w_095_2885, w_095_2886, w_095_2888, w_095_2891, w_095_2893, w_095_2897, w_095_2898, w_095_2901, w_095_2905, w_095_2907, w_095_2911, w_095_2918, w_095_2919, w_095_2920, w_095_2921, w_095_2926, w_095_2929, w_095_2930, w_095_2933, w_095_2936, w_095_2943, w_095_2945, w_095_2948, w_095_2952, w_095_2953, w_095_2955, w_095_2957, w_095_2958, w_095_2964, w_095_2965, w_095_2969, w_095_2971, w_095_2972, w_095_2974, w_095_2976, w_095_2978, w_095_2979, w_095_2983, w_095_2984, w_095_2985, w_095_2993, w_095_2996, w_095_3000, w_095_3001, w_095_3005, w_095_3006, w_095_3007, w_095_3008, w_095_3010, w_095_3013, w_095_3015, w_095_3016, w_095_3020, w_095_3022, w_095_3023, w_095_3026, w_095_3033, w_095_3036, w_095_3038, w_095_3041, w_095_3044, w_095_3046, w_095_3048, w_095_3049, w_095_3051, w_095_3054, w_095_3055, w_095_3058, w_095_3061, w_095_3062, w_095_3063, w_095_3067, w_095_3068, w_095_3069, w_095_3070, w_095_3072, w_095_3074, w_095_3075, w_095_3078, w_095_3083, w_095_3084, w_095_3087, w_095_3088, w_095_3089, w_095_3090, w_095_3092, w_095_3097, w_095_3099, w_095_3105, w_095_3107, w_095_3108, w_095_3110, w_095_3112, w_095_3114, w_095_3120, w_095_3125, w_095_3127, w_095_3129, w_095_3130, w_095_3131, w_095_3135, w_095_3144, w_095_3145, w_095_3146, w_095_3147, w_095_3149, w_095_3152, w_095_3153, w_095_3155, w_095_3157, w_095_3163, w_095_3174, w_095_3177, w_095_3189, w_095_3191, w_095_3193, w_095_3194, w_095_3195, w_095_3200, w_095_3202, w_095_3204, w_095_3205, w_095_3207, w_095_3210, w_095_3211, w_095_3212, w_095_3215, w_095_3218, w_095_3220, w_095_3221, w_095_3225, w_095_3227, w_095_3229, w_095_3234, w_095_3237, w_095_3240, w_095_3241, w_095_3244, w_095_3248, w_095_3252, w_095_3259, w_095_3260, w_095_3262, w_095_3264, w_095_3266, w_095_3270, w_095_3271, w_095_3272, w_095_3273, w_095_3274, w_095_3275, w_095_3276, w_095_3277, w_095_3278, w_095_3281, w_095_3282, w_095_3283, w_095_3287, w_095_3288, w_095_3291, w_095_3292, w_095_3294, w_095_3296, w_095_3299, w_095_3300, w_095_3301, w_095_3304, w_095_3305, w_095_3306, w_095_3310, w_095_3312, w_095_3313, w_095_3314, w_095_3318, w_095_3322, w_095_3323, w_095_3325, w_095_3328, w_095_3329, w_095_3331, w_095_3336, w_095_3337, w_095_3339, w_095_3340, w_095_3343, w_095_3353, w_095_3354, w_095_3355, w_095_3356, w_095_3358, w_095_3359, w_095_3361, w_095_3362, w_095_3363, w_095_3365, w_095_3367, w_095_3371, w_095_3373, w_095_3376, w_095_3377, w_095_3379, w_095_3382, w_095_3384, w_095_3386, w_095_3387, w_095_3389, w_095_3391, w_095_3396, w_095_3398, w_095_3401, w_095_3404, w_095_3405, w_095_3406, w_095_3410, w_095_3411, w_095_3413, w_095_3414, w_095_3415, w_095_3416, w_095_3421, w_095_3423, w_095_3425, w_095_3427, w_095_3428, w_095_3429, w_095_3430, w_095_3434, w_095_3436, w_095_3438, w_095_3439, w_095_3440, w_095_3441, w_095_3442, w_095_3444, w_095_3446, w_095_3452, w_095_3455, w_095_3456, w_095_3457, w_095_3459, w_095_3464, w_095_3466, w_095_3471, w_095_3474, w_095_3475, w_095_3476, w_095_3478, w_095_3481, w_095_3482, w_095_3483, w_095_3484, w_095_3487, w_095_3488, w_095_3489, w_095_3490, w_095_3491, w_095_3492, w_095_3495, w_095_3498, w_095_3502, w_095_3503, w_095_3506, w_095_3509, w_095_3510, w_095_3512, w_095_3515, w_095_3516, w_095_3523, w_095_3524, w_095_3526, w_095_3528, w_095_3533, w_095_3537, w_095_3538, w_095_3539, w_095_3541, w_095_3543, w_095_3546, w_095_3553, w_095_3555, w_095_3556, w_095_3559, w_095_3563, w_095_3565, w_095_3569, w_095_3573, w_095_3574, w_095_3575, w_095_3577, w_095_3581, w_095_3582, w_095_3586, w_095_3588, w_095_3589, w_095_3590, w_095_3593, w_095_3599, w_095_3602, w_095_3603, w_095_3604, w_095_3605, w_095_3608, w_095_3610, w_095_3612, w_095_3616, w_095_3617;
  wire w_096_000, w_096_005, w_096_007, w_096_009, w_096_014, w_096_018, w_096_021, w_096_027, w_096_037, w_096_039, w_096_043, w_096_045, w_096_046, w_096_047, w_096_050, w_096_051, w_096_053, w_096_055, w_096_056, w_096_064, w_096_067, w_096_074, w_096_077, w_096_078, w_096_079, w_096_084, w_096_086, w_096_089, w_096_090, w_096_092, w_096_093, w_096_094, w_096_095, w_096_097, w_096_103, w_096_104, w_096_106, w_096_108, w_096_109, w_096_114, w_096_115, w_096_118, w_096_120, w_096_122, w_096_123, w_096_124, w_096_130, w_096_133, w_096_136, w_096_144, w_096_152, w_096_154, w_096_155, w_096_157, w_096_160, w_096_162, w_096_165, w_096_169, w_096_171, w_096_175, w_096_185, w_096_187, w_096_188, w_096_190, w_096_191, w_096_193, w_096_195, w_096_198, w_096_199, w_096_202, w_096_205, w_096_206, w_096_207, w_096_212, w_096_215, w_096_219, w_096_221, w_096_225, w_096_227, w_096_229, w_096_236, w_096_237, w_096_241, w_096_242, w_096_246, w_096_247, w_096_248, w_096_251, w_096_255, w_096_257, w_096_258, w_096_259, w_096_261, w_096_262, w_096_264, w_096_267, w_096_270, w_096_271, w_096_272, w_096_274, w_096_275, w_096_276, w_096_277, w_096_279, w_096_283, w_096_284, w_096_286, w_096_293, w_096_296, w_096_302, w_096_303, w_096_305, w_096_307, w_096_309, w_096_312, w_096_316, w_096_318, w_096_325, w_096_326, w_096_329, w_096_331, w_096_332, w_096_333, w_096_335, w_096_336, w_096_338, w_096_342, w_096_343, w_096_344, w_096_355, w_096_360, w_096_364, w_096_365, w_096_368, w_096_372, w_096_374, w_096_378, w_096_379, w_096_382, w_096_383, w_096_386, w_096_388, w_096_389, w_096_396, w_096_397, w_096_398, w_096_401, w_096_405, w_096_408, w_096_411, w_096_412, w_096_413, w_096_415, w_096_417, w_096_418, w_096_419, w_096_421, w_096_422, w_096_423, w_096_425, w_096_428, w_096_429, w_096_430, w_096_433, w_096_442, w_096_448, w_096_451, w_096_452, w_096_457, w_096_458, w_096_460, w_096_462, w_096_463, w_096_467, w_096_468, w_096_470, w_096_471, w_096_474, w_096_475, w_096_478, w_096_479, w_096_484, w_096_485, w_096_489, w_096_491, w_096_496, w_096_501, w_096_504, w_096_505, w_096_511, w_096_512, w_096_514, w_096_517, w_096_519, w_096_520, w_096_521, w_096_531, w_096_532, w_096_535, w_096_539, w_096_540, w_096_541, w_096_543, w_096_544, w_096_545, w_096_548, w_096_549, w_096_550, w_096_552, w_096_556, w_096_562, w_096_573, w_096_574, w_096_576, w_096_577, w_096_578, w_096_580, w_096_581, w_096_583, w_096_584, w_096_585, w_096_590, w_096_591, w_096_592, w_096_595, w_096_596, w_096_597, w_096_598, w_096_599, w_096_604, w_096_605, w_096_612, w_096_619, w_096_623, w_096_624, w_096_625, w_096_628, w_096_629, w_096_633, w_096_634, w_096_635, w_096_637, w_096_638, w_096_639, w_096_640, w_096_642, w_096_643, w_096_644, w_096_648, w_096_650, w_096_651, w_096_655, w_096_659, w_096_664, w_096_667, w_096_669, w_096_672, w_096_673, w_096_675, w_096_677, w_096_680, w_096_684, w_096_685, w_096_686, w_096_687, w_096_689, w_096_690, w_096_693, w_096_694, w_096_702, w_096_703, w_096_704, w_096_708, w_096_710, w_096_712, w_096_714, w_096_715, w_096_720, w_096_722, w_096_724, w_096_725, w_096_726, w_096_728, w_096_730, w_096_731, w_096_733, w_096_734, w_096_735, w_096_739, w_096_744, w_096_745, w_096_747, w_096_748, w_096_749, w_096_750, w_096_753, w_096_758, w_096_760, w_096_762, w_096_763, w_096_766, w_096_768, w_096_769, w_096_771, w_096_772, w_096_773, w_096_774, w_096_775, w_096_777, w_096_779, w_096_785, w_096_786, w_096_787, w_096_788, w_096_790, w_096_795, w_096_797, w_096_798, w_096_799, w_096_805, w_096_806, w_096_808, w_096_814, w_096_815, w_096_819, w_096_820, w_096_825, w_096_828, w_096_829, w_096_832, w_096_834, w_096_836, w_096_838, w_096_839, w_096_840, w_096_843, w_096_844, w_096_845, w_096_848, w_096_851, w_096_853, w_096_855, w_096_858, w_096_859, w_096_865, w_096_866, w_096_870, w_096_872, w_096_873, w_096_874, w_096_875, w_096_877, w_096_880, w_096_881, w_096_882, w_096_884, w_096_885, w_096_886, w_096_890, w_096_892, w_096_893, w_096_897, w_096_905, w_096_906, w_096_907, w_096_911, w_096_914, w_096_915, w_096_921, w_096_925, w_096_933, w_096_934, w_096_938, w_096_939, w_096_940, w_096_941, w_096_942, w_096_944, w_096_947, w_096_948, w_096_949, w_096_954, w_096_956, w_096_957, w_096_961, w_096_965, w_096_970, w_096_972, w_096_975, w_096_981, w_096_982, w_096_983, w_096_986, w_096_992, w_096_997, w_096_998, w_096_999, w_096_1001, w_096_1002, w_096_1010, w_096_1014, w_096_1015, w_096_1020, w_096_1022, w_096_1023, w_096_1025, w_096_1027, w_096_1028, w_096_1029, w_096_1030, w_096_1035, w_096_1038, w_096_1040, w_096_1041, w_096_1044, w_096_1045, w_096_1046, w_096_1048, w_096_1051, w_096_1053, w_096_1054, w_096_1058, w_096_1062, w_096_1071, w_096_1074, w_096_1077, w_096_1078, w_096_1080, w_096_1083, w_096_1086, w_096_1089, w_096_1096, w_096_1098, w_096_1099, w_096_1100, w_096_1102, w_096_1103, w_096_1104, w_096_1106, w_096_1111, w_096_1112, w_096_1113, w_096_1115, w_096_1116, w_096_1118, w_096_1119, w_096_1121, w_096_1123, w_096_1125, w_096_1126, w_096_1133, w_096_1140, w_096_1142, w_096_1146, w_096_1148, w_096_1150, w_096_1155, w_096_1157, w_096_1159, w_096_1160, w_096_1162, w_096_1165, w_096_1167, w_096_1168, w_096_1169, w_096_1170, w_096_1171, w_096_1175, w_096_1180, w_096_1181, w_096_1183, w_096_1187, w_096_1188, w_096_1190, w_096_1192, w_096_1194, w_096_1195, w_096_1196, w_096_1197, w_096_1201, w_096_1203, w_096_1206, w_096_1208, w_096_1210, w_096_1211, w_096_1213, w_096_1217, w_096_1219, w_096_1222, w_096_1224, w_096_1225, w_096_1226, w_096_1237, w_096_1238, w_096_1239, w_096_1240, w_096_1244, w_096_1245, w_096_1246, w_096_1247, w_096_1252, w_096_1254, w_096_1259, w_096_1261, w_096_1265, w_096_1266, w_096_1267, w_096_1269, w_096_1271, w_096_1273, w_096_1275, w_096_1279, w_096_1281, w_096_1283, w_096_1284, w_096_1285, w_096_1286, w_096_1289, w_096_1293, w_096_1295, w_096_1296, w_096_1297, w_096_1299, w_096_1303, w_096_1304, w_096_1305, w_096_1306, w_096_1309, w_096_1315, w_096_1318, w_096_1330, w_096_1331, w_096_1333, w_096_1334, w_096_1335, w_096_1336, w_096_1339, w_096_1340, w_096_1347, w_096_1348, w_096_1353, w_096_1354, w_096_1356, w_096_1358, w_096_1359, w_096_1361, w_096_1366, w_096_1373, w_096_1375, w_096_1376, w_096_1379, w_096_1380, w_096_1382, w_096_1383, w_096_1384, w_096_1388, w_096_1389, w_096_1390, w_096_1393, w_096_1394, w_096_1395, w_096_1397, w_096_1399, w_096_1401, w_096_1402, w_096_1403, w_096_1405, w_096_1408, w_096_1410, w_096_1411, w_096_1412, w_096_1413, w_096_1416, w_096_1417, w_096_1418, w_096_1420, w_096_1421, w_096_1422, w_096_1423, w_096_1434, w_096_1441, w_096_1442, w_096_1449, w_096_1451, w_096_1452, w_096_1453, w_096_1455, w_096_1458, w_096_1459, w_096_1460, w_096_1462, w_096_1465, w_096_1469, w_096_1470, w_096_1472, w_096_1477, w_096_1479, w_096_1481, w_096_1484, w_096_1485, w_096_1489, w_096_1492, w_096_1495, w_096_1498, w_096_1500, w_096_1502, w_096_1504, w_096_1506, w_096_1510, w_096_1511, w_096_1515, w_096_1517, w_096_1519, w_096_1520, w_096_1523, w_096_1524, w_096_1526, w_096_1527, w_096_1528, w_096_1529, w_096_1531, w_096_1532, w_096_1533, w_096_1534, w_096_1535, w_096_1537, w_096_1538, w_096_1543, w_096_1546, w_096_1551, w_096_1557, w_096_1561, w_096_1563, w_096_1565, w_096_1566, w_096_1567, w_096_1569, w_096_1570, w_096_1571, w_096_1572, w_096_1573, w_096_1575, w_096_1578, w_096_1580, w_096_1584, w_096_1585, w_096_1586, w_096_1588, w_096_1590, w_096_1591, w_096_1592, w_096_1593, w_096_1595, w_096_1598, w_096_1604, w_096_1608, w_096_1612, w_096_1614, w_096_1618, w_096_1621, w_096_1623, w_096_1624, w_096_1625, w_096_1627, w_096_1631, w_096_1633, w_096_1635, w_096_1636, w_096_1637, w_096_1638, w_096_1641, w_096_1642, w_096_1644, w_096_1646, w_096_1648, w_096_1649, w_096_1651, w_096_1653, w_096_1656, w_096_1657, w_096_1658, w_096_1660, w_096_1661, w_096_1664, w_096_1666, w_096_1668, w_096_1671, w_096_1673, w_096_1674, w_096_1678, w_096_1682, w_096_1685, w_096_1686, w_096_1691, w_096_1692, w_096_1693, w_096_1695, w_096_1697, w_096_1698, w_096_1699, w_096_1701, w_096_1702, w_096_1703, w_096_1704, w_096_1707, w_096_1708, w_096_1710, w_096_1712, w_096_1714, w_096_1715, w_096_1716, w_096_1717, w_096_1719, w_096_1721, w_096_1725, w_096_1726, w_096_1728, w_096_1730, w_096_1731, w_096_1733, w_096_1735, w_096_1736, w_096_1737, w_096_1739, w_096_1741, w_096_1743, w_096_1744, w_096_1746, w_096_1747, w_096_1754, w_096_1757, w_096_1762, w_096_1764, w_096_1766, w_096_1767, w_096_1768, w_096_1771, w_096_1773, w_096_1774, w_096_1775, w_096_1779, w_096_1781, w_096_1783, w_096_1787, w_096_1789, w_096_1791, w_096_1793, w_096_1798, w_096_1801, w_096_1802, w_096_1804, w_096_1805, w_096_1807, w_096_1809, w_096_1811, w_096_1812, w_096_1813, w_096_1814, w_096_1815, w_096_1816, w_096_1818, w_096_1819, w_096_1822, w_096_1824, w_096_1827, w_096_1830, w_096_1831, w_096_1832, w_096_1836, w_096_1838, w_096_1839, w_096_1842, w_096_1843, w_096_1844, w_096_1845, w_096_1848, w_096_1849, w_096_1850, w_096_1853, w_096_1854, w_096_1858, w_096_1860, w_096_1866, w_096_1867, w_096_1868, w_096_1869, w_096_1870, w_096_1872, w_096_1877, w_096_1881, w_096_1882, w_096_1887, w_096_1889, w_096_1893, w_096_1895, w_096_1896, w_096_1897, w_096_1898, w_096_1899, w_096_1904, w_096_1905, w_096_1912, w_096_1914, w_096_1917, w_096_1918, w_096_1920, w_096_1928, w_096_1929, w_096_1931, w_096_1933, w_096_1934, w_096_1938, w_096_1940, w_096_1943, w_096_1946, w_096_1949, w_096_1951, w_096_1952, w_096_1954, w_096_1955, w_096_1959, w_096_1964, w_096_1965, w_096_1967, w_096_1968, w_096_1969, w_096_1973, w_096_1974, w_096_1979, w_096_1980, w_096_1981, w_096_1985, w_096_1987, w_096_1989, w_096_1993, w_096_1995, w_096_1998, w_096_2006, w_096_2008, w_096_2009, w_096_2014, w_096_2016, w_096_2017, w_096_2018, w_096_2020, w_096_2021, w_096_2023, w_096_2026, w_096_2030, w_096_2033, w_096_2035, w_096_2037, w_096_2044, w_096_2045, w_096_2047, w_096_2049, w_096_2050, w_096_2051, w_096_2054, w_096_2057, w_096_2059, w_096_2060, w_096_2065, w_096_2071, w_096_2072, w_096_2074, w_096_2075, w_096_2076, w_096_2078, w_096_2080, w_096_2081, w_096_2085, w_096_2086, w_096_2087, w_096_2088, w_096_2090, w_096_2092, w_096_2097, w_096_2102, w_096_2106, w_096_2109, w_096_2111, w_096_2114, w_096_2118, w_096_2119, w_096_2121, w_096_2123, w_096_2124, w_096_2128, w_096_2130, w_096_2134, w_096_2136, w_096_2140, w_096_2141, w_096_2146, w_096_2151, w_096_2153, w_096_2154, w_096_2158, w_096_2159, w_096_2160, w_096_2162, w_096_2166, w_096_2167, w_096_2170, w_096_2171, w_096_2173, w_096_2174, w_096_2177, w_096_2182, w_096_2183, w_096_2186, w_096_2189, w_096_2194, w_096_2197, w_096_2200, w_096_2202, w_096_2205, w_096_2211, w_096_2213, w_096_2215, w_096_2221, w_096_2222, w_096_2223, w_096_2227, w_096_2229, w_096_2230, w_096_2231, w_096_2233, w_096_2239, w_096_2244, w_096_2247, w_096_2248, w_096_2253, w_096_2257, w_096_2258, w_096_2259, w_096_2264, w_096_2266, w_096_2269, w_096_2270, w_096_2278, w_096_2284, w_096_2285, w_096_2287, w_096_2288, w_096_2291, w_096_2299, w_096_2302, w_096_2305, w_096_2306, w_096_2307, w_096_2312, w_096_2313, w_096_2316, w_096_2317, w_096_2318, w_096_2326, w_096_2333, w_096_2334, w_096_2338, w_096_2339, w_096_2341, w_096_2342, w_096_2343, w_096_2345, w_096_2351, w_096_2352, w_096_2355, w_096_2356, w_096_2359, w_096_2360, w_096_2361, w_096_2364, w_096_2365, w_096_2367, w_096_2368, w_096_2370, w_096_2371, w_096_2372, w_096_2373, w_096_2374, w_096_2378, w_096_2382, w_096_2385, w_096_2386, w_096_2394, w_096_2395, w_096_2397, w_096_2402, w_096_2403, w_096_2405, w_096_2412, w_096_2414, w_096_2428, w_096_2429, w_096_2431, w_096_2434, w_096_2435, w_096_2436, w_096_2438, w_096_2439, w_096_2448, w_096_2449, w_096_2450, w_096_2452, w_096_2456, w_096_2458, w_096_2459, w_096_2460, w_096_2464, w_096_2468, w_096_2469, w_096_2471, w_096_2472, w_096_2473, w_096_2477, w_096_2479, w_096_2482, w_096_2484, w_096_2486, w_096_2487, w_096_2488, w_096_2490, w_096_2494, w_096_2497, w_096_2498, w_096_2500, w_096_2501, w_096_2503, w_096_2505, w_096_2507, w_096_2510, w_096_2511, w_096_2512, w_096_2513, w_096_2516, w_096_2518, w_096_2519, w_096_2520, w_096_2522, w_096_2524, w_096_2525, w_096_2533, w_096_2537, w_096_2540, w_096_2542, w_096_2544, w_096_2546, w_096_2548, w_096_2549, w_096_2551, w_096_2552, w_096_2564, w_096_2565, w_096_2566, w_096_2569, w_096_2571, w_096_2574, w_096_2580, w_096_2582, w_096_2586, w_096_2588, w_096_2593, w_096_2594, w_096_2596, w_096_2597, w_096_2599, w_096_2601, w_096_2602, w_096_2607, w_096_2609, w_096_2610, w_096_2611, w_096_2612, w_096_2613, w_096_2615, w_096_2616, w_096_2617, w_096_2620, w_096_2623, w_096_2626, w_096_2630, w_096_2632, w_096_2634, w_096_2638, w_096_2640, w_096_2643, w_096_2644, w_096_2645, w_096_2647, w_096_2649, w_096_2657, w_096_2659, w_096_2660, w_096_2663, w_096_2664, w_096_2665, w_096_2667, w_096_2668, w_096_2670, w_096_2671, w_096_2678, w_096_2679, w_096_2686, w_096_2698, w_096_2701, w_096_2704, w_096_2707, w_096_2708, w_096_2710, w_096_2716, w_096_2720, w_096_2727, w_096_2734, w_096_2737, w_096_2746, w_096_2747, w_096_2753, w_096_2754, w_096_2755, w_096_2756, w_096_2757, w_096_2759, w_096_2765, w_096_2766, w_096_2767, w_096_2771, w_096_2772, w_096_2777, w_096_2779, w_096_2781, w_096_2784, w_096_2786, w_096_2794, w_096_2797, w_096_2800, w_096_2805, w_096_2806, w_096_2809, w_096_2811, w_096_2815, w_096_2825, w_096_2831, w_096_2832, w_096_2834, w_096_2837, w_096_2838, w_096_2840, w_096_2841, w_096_2842, w_096_2847, w_096_2851, w_096_2855, w_096_2856, w_096_2857, w_096_2860, w_096_2861, w_096_2864, w_096_2866, w_096_2868, w_096_2869, w_096_2876, w_096_2882, w_096_2886, w_096_2887, w_096_2888, w_096_2890, w_096_2898, w_096_2899, w_096_2900, w_096_2901, w_096_2907, w_096_2909, w_096_2912, w_096_2913, w_096_2915, w_096_2917, w_096_2918, w_096_2919, w_096_2920, w_096_2926, w_096_2928, w_096_2929, w_096_2930, w_096_2934, w_096_2935, w_096_2937, w_096_2941, w_096_2942, w_096_2946, w_096_2948, w_096_2949, w_096_2952, w_096_2957, w_096_2963, w_096_2964, w_096_2970, w_096_2974, w_096_2981, w_096_2985, w_096_2986, w_096_2991, w_096_2994, w_096_3002, w_096_3003, w_096_3004, w_096_3009, w_096_3013, w_096_3015, w_096_3018, w_096_3024, w_096_3029, w_096_3032, w_096_3039, w_096_3042, w_096_3043, w_096_3044, w_096_3045, w_096_3055, w_096_3062, w_096_3063, w_096_3069, w_096_3073, w_096_3077, w_096_3080, w_096_3083, w_096_3090, w_096_3094, w_096_3095, w_096_3096, w_096_3097, w_096_3098, w_096_3100, w_096_3104, w_096_3107, w_096_3109, w_096_3110, w_096_3111, w_096_3113, w_096_3114, w_096_3115, w_096_3116, w_096_3117, w_096_3119, w_096_3120, w_096_3121, w_096_3127, w_096_3132, w_096_3133, w_096_3137, w_096_3141, w_096_3143, w_096_3150, w_096_3154, w_096_3156, w_096_3157, w_096_3161, w_096_3162, w_096_3163, w_096_3168, w_096_3174, w_096_3175, w_096_3176, w_096_3178, w_096_3184, w_096_3185, w_096_3187, w_096_3188, w_096_3190, w_096_3193, w_096_3194, w_096_3195, w_096_3196, w_096_3197, w_096_3199, w_096_3203, w_096_3205, w_096_3206, w_096_3208, w_096_3209, w_096_3211, w_096_3213, w_096_3214, w_096_3222, w_096_3226, w_096_3228, w_096_3229, w_096_3230, w_096_3231, w_096_3232, w_096_3233, w_096_3236, w_096_3238, w_096_3247, w_096_3248, w_096_3250, w_096_3251, w_096_3255, w_096_3259, w_096_3261, w_096_3262, w_096_3263, w_096_3265, w_096_3269, w_096_3270, w_096_3271, w_096_3272, w_096_3274, w_096_3275, w_096_3277, w_096_3278, w_096_3281, w_096_3282, w_096_3285, w_096_3286, w_096_3287, w_096_3289, w_096_3294, w_096_3300, w_096_3301, w_096_3304, w_096_3313, w_096_3315, w_096_3316, w_096_3320, w_096_3322, w_096_3328, w_096_3330, w_096_3334, w_096_3338, w_096_3339, w_096_3340, w_096_3341, w_096_3342, w_096_3343, w_096_3345, w_096_3346, w_096_3354, w_096_3359, w_096_3360, w_096_3361, w_096_3362, w_096_3365, w_096_3366, w_096_3374, w_096_3375, w_096_3376, w_096_3378, w_096_3379, w_096_3382, w_096_3383, w_096_3384, w_096_3386, w_096_3390, w_096_3393, w_096_3406, w_096_3412, w_096_3414, w_096_3418, w_096_3420, w_096_3421, w_096_3424, w_096_3425, w_096_3426, w_096_3428, w_096_3430, w_096_3432, w_096_3436, w_096_3437, w_096_3438, w_096_3440, w_096_3441, w_096_3445, w_096_3452, w_096_3455, w_096_3456, w_096_3461, w_096_3462, w_096_3463, w_096_3464, w_096_3465, w_096_3467, w_096_3468, w_096_3470, w_096_3477, w_096_3478, w_096_3480, w_096_3484, w_096_3485, w_096_3486, w_096_3487, w_096_3489, w_096_3493, w_096_3494, w_096_3495, w_096_3496, w_096_3498, w_096_3500, w_096_3502, w_096_3503, w_096_3508, w_096_3510, w_096_3511, w_096_3513, w_096_3514, w_096_3516, w_096_3519, w_096_3521, w_096_3522, w_096_3523, w_096_3529, w_096_3530, w_096_3531, w_096_3532, w_096_3534, w_096_3536, w_096_3537, w_096_3538, w_096_3540, w_096_3541, w_096_3542, w_096_3543, w_096_3545, w_096_3546, w_096_3547, w_096_3555, w_096_3556, w_096_3559, w_096_3561, w_096_3565, w_096_3566, w_096_3568, w_096_3573, w_096_3577, w_096_3586, w_096_3594, w_096_3598, w_096_3601, w_096_3609, w_096_3611, w_096_3612, w_096_3613, w_096_3617, w_096_3622, w_096_3624, w_096_3625, w_096_3630, w_096_3635, w_096_3638, w_096_3642, w_096_3649, w_096_3650, w_096_3651, w_096_3653, w_096_3657, w_096_3659, w_096_3660, w_096_3665, w_096_3667, w_096_3670, w_096_3671, w_096_3672, w_096_3691, w_096_3698, w_096_3703, w_096_3706, w_096_3707, w_096_3711, w_096_3719, w_096_3728, w_096_3730, w_096_3743, w_096_3749, w_096_3753, w_096_3759, w_096_3769, w_096_3777, w_096_3780, w_096_3783, w_096_3787, w_096_3790, w_096_3792, w_096_3794, w_096_3799, w_096_3809, w_096_3812, w_096_3815, w_096_3816, w_096_3817, w_096_3819, w_096_3820, w_096_3821, w_096_3825, w_096_3833, w_096_3835, w_096_3837, w_096_3839, w_096_3843, w_096_3848, w_096_3850, w_096_3852, w_096_3857, w_096_3858, w_096_3860, w_096_3863, w_096_3880, w_096_3883, w_096_3892, w_096_3896, w_096_3901, w_096_3906, w_096_3911, w_096_3914, w_096_3916, w_096_3918, w_096_3922, w_096_3923, w_096_3932, w_096_3935, w_096_3940, w_096_3942, w_096_3951, w_096_3959, w_096_3961, w_096_3968, w_096_3972, w_096_3974, w_096_3975, w_096_3978, w_096_3982, w_096_3985, w_096_3986, w_096_3987, w_096_3998, w_096_3999, w_096_4004, w_096_4006, w_096_4010, w_096_4015, w_096_4016, w_096_4017, w_096_4028, w_096_4031, w_096_4036, w_096_4038, w_096_4047, w_096_4050, w_096_4051, w_096_4054, w_096_4056, w_096_4067, w_096_4070, w_096_4071, w_096_4072, w_096_4073, w_096_4081, w_096_4085, w_096_4088, w_096_4093, w_096_4101, w_096_4102, w_096_4110, w_096_4111, w_096_4114, w_096_4119, w_096_4123, w_096_4124, w_096_4125, w_096_4126, w_096_4130, w_096_4142, w_096_4143, w_096_4147, w_096_4148, w_096_4159, w_096_4161, w_096_4171, w_096_4176, w_096_4178, w_096_4179, w_096_4181, w_096_4194, w_096_4199, w_096_4210, w_096_4215, w_096_4220, w_096_4224, w_096_4234, w_096_4239, w_096_4241, w_096_4243, w_096_4245, w_096_4249, w_096_4250, w_096_4251, w_096_4256, w_096_4258, w_096_4264, w_096_4266, w_096_4281, w_096_4282, w_096_4289, w_096_4293, w_096_4296, w_096_4299, w_096_4303, w_096_4309, w_096_4320, w_096_4321, w_096_4325, w_096_4328, w_096_4332, w_096_4335, w_096_4337, w_096_4342, w_096_4344, w_096_4346, w_096_4364, w_096_4365, w_096_4366, w_096_4367, w_096_4369, w_096_4371, w_096_4376, w_096_4377, w_096_4379, w_096_4382, w_096_4384, w_096_4392, w_096_4394, w_096_4400, w_096_4405, w_096_4408, w_096_4413, w_096_4416, w_096_4417, w_096_4426, w_096_4427, w_096_4438, w_096_4442, w_096_4449, w_096_4458, w_096_4464, w_096_4475, w_096_4481, w_096_4483, w_096_4484, w_096_4490, w_096_4491, w_096_4492, w_096_4494, w_096_4499, w_096_4503, w_096_4506, w_096_4509, w_096_4510, w_096_4514, w_096_4524, w_096_4527, w_096_4529, w_096_4530, w_096_4532, w_096_4533, w_096_4543, w_096_4545, w_096_4546, w_096_4553, w_096_4557, w_096_4559, w_096_4560, w_096_4562, w_096_4570, w_096_4576, w_096_4600, w_096_4604, w_096_4616, w_096_4618, w_096_4621, w_096_4623, w_096_4624, w_096_4626, w_096_4637, w_096_4638, w_096_4642, w_096_4654, w_096_4658, w_096_4659, w_096_4660, w_096_4663, w_096_4665, w_096_4667, w_096_4673, w_096_4678, w_096_4681, w_096_4685, w_096_4686, w_096_4688, w_096_4696, w_096_4702, w_096_4704, w_096_4705, w_096_4707, w_096_4713, w_096_4720, w_096_4722, w_096_4726, w_096_4727, w_096_4732, w_096_4744, w_096_4749, w_096_4750, w_096_4753, w_096_4758, w_096_4759, w_096_4762, w_096_4764, w_096_4765, w_096_4772, w_096_4778, w_096_4782, w_096_4783, w_096_4786, w_096_4807, w_096_4812, w_096_4815, w_096_4817, w_096_4819, w_096_4822, w_096_4823, w_096_4828, w_096_4830, w_096_4843, w_096_4845, w_096_4848, w_096_4852, w_096_4854, w_096_4858, w_096_4866, w_096_4867, w_096_4869, w_096_4872, w_096_4875, w_096_4883, w_096_4886, w_096_4892, w_096_4901, w_096_4902, w_096_4909, w_096_4911, w_096_4914, w_096_4917, w_096_4918, w_096_4926, w_096_4946, w_096_4960, w_096_4962, w_096_4968, w_096_4969, w_096_4974, w_096_4979, w_096_4981, w_096_4984, w_096_4988, w_096_4991, w_096_4996, w_096_4998, w_096_4999, w_096_5007, w_096_5013, w_096_5023, w_096_5024, w_096_5030, w_096_5059, w_096_5060, w_096_5072, w_096_5074, w_096_5082, w_096_5083, w_096_5088, w_096_5091, w_096_5094, w_096_5104, w_096_5128, w_096_5131, w_096_5134, w_096_5136, w_096_5141, w_096_5146, w_096_5147, w_096_5151, w_096_5155, w_096_5164, w_096_5166, w_096_5167, w_096_5168, w_096_5170, w_096_5174, w_096_5176, w_096_5183, w_096_5193, w_096_5196, w_096_5203, w_096_5206, w_096_5208, w_096_5212, w_096_5216, w_096_5219, w_096_5230, w_096_5241, w_096_5245, w_096_5247, w_096_5253, w_096_5259, w_096_5261, w_096_5269, w_096_5272, w_096_5289, w_096_5291, w_096_5300, w_096_5302, w_096_5307, w_096_5308, w_096_5312, w_096_5313, w_096_5319, w_096_5322, w_096_5323, w_096_5324, w_096_5327, w_096_5329, w_096_5331, w_096_5335, w_096_5338, w_096_5339, w_096_5341, w_096_5345, w_096_5348, w_096_5355, w_096_5361, w_096_5366, w_096_5377, w_096_5379, w_096_5382, w_096_5383, w_096_5384, w_096_5386, w_096_5393, w_096_5396, w_096_5397, w_096_5399, w_096_5400, w_096_5410, w_096_5415, w_096_5417, w_096_5419, w_096_5420, w_096_5429, w_096_5430, w_096_5433, w_096_5434, w_096_5438, w_096_5440, w_096_5450, w_096_5452, w_096_5461, w_096_5469, w_096_5470, w_096_5474, w_096_5476, w_096_5485, w_096_5487, w_096_5492, w_096_5498, w_096_5499, w_096_5503, w_096_5506, w_096_5509, w_096_5519, w_096_5520, w_096_5530, w_096_5537, w_096_5538, w_096_5540, w_096_5542, w_096_5550, w_096_5558, w_096_5562, w_096_5565, w_096_5570, w_096_5571, w_096_5573, w_096_5574, w_096_5575, w_096_5584, w_096_5592, w_096_5596, w_096_5599, w_096_5601, w_096_5602, w_096_5603, w_096_5605, w_096_5607, w_096_5608, w_096_5618, w_096_5623, w_096_5624, w_096_5638, w_096_5639, w_096_5641, w_096_5644, w_096_5648, w_096_5651, w_096_5658, w_096_5660, w_096_5663, w_096_5665, w_096_5666, w_096_5669, w_096_5674, w_096_5676, w_096_5678, w_096_5680, w_096_5683, w_096_5685, w_096_5686, w_096_5687, w_096_5702, w_096_5718, w_096_5722, w_096_5728, w_096_5731, w_096_5734, w_096_5737, w_096_5740, w_096_5752, w_096_5754, w_096_5762, w_096_5764, w_096_5770, w_096_5771, w_096_5780, w_096_5787, w_096_5792, w_096_5795, w_096_5796, w_096_5798, w_096_5812, w_096_5820, w_096_5821, w_096_5824, w_096_5832, w_096_5833, w_096_5842, w_096_5849, w_096_5864, w_096_5867, w_096_5868, w_096_5871, w_096_5873, w_096_5882, w_096_5884, w_096_5887, w_096_5892, w_096_5902, w_096_5905, w_096_5907, w_096_5909, w_096_5924, w_096_5925, w_096_5946, w_096_5948, w_096_5950, w_096_5954, w_096_5961, w_096_5964, w_096_5969, w_096_5972, w_096_5973, w_096_5977, w_096_5991, w_096_5993, w_096_5997, w_096_5999, w_096_6005, w_096_6006, w_096_6008, w_096_6012, w_096_6015, w_096_6026, w_096_6028, w_096_6032, w_096_6037, w_096_6038, w_096_6040, w_096_6044, w_096_6046, w_096_6055, w_096_6056, w_096_6057, w_096_6063, w_096_6072, w_096_6075, w_096_6082, w_096_6083, w_096_6084, w_096_6093, w_096_6095, w_096_6096, w_096_6099, w_096_6100, w_096_6101, w_096_6105, w_096_6109, w_096_6117, w_096_6119, w_096_6124, w_096_6126, w_096_6127, w_096_6135, w_096_6140, w_096_6141, w_096_6146, w_096_6151, w_096_6155, w_096_6164, w_096_6166, w_096_6171, w_096_6177, w_096_6191, w_096_6192, w_096_6197, w_096_6199, w_096_6200, w_096_6207, w_096_6209, w_096_6211, w_096_6216, w_096_6217, w_096_6218, w_096_6222, w_096_6223, w_096_6238, w_096_6240, w_096_6242, w_096_6244, w_096_6252, w_096_6253, w_096_6254, w_096_6258, w_096_6260, w_096_6265, w_096_6270, w_096_6275, w_096_6276, w_096_6282, w_096_6287, w_096_6290, w_096_6291, w_096_6292, w_096_6297, w_096_6298, w_096_6302, w_096_6303, w_096_6306, w_096_6312, w_096_6318, w_096_6320, w_096_6321, w_096_6324, w_096_6328, w_096_6341, w_096_6342, w_096_6344, w_096_6349, w_096_6351, w_096_6357, w_096_6362, w_096_6374, w_096_6375, w_096_6377, w_096_6379, w_096_6393, w_096_6405, w_096_6406, w_096_6411, w_096_6415, w_096_6418, w_096_6419, w_096_6422, w_096_6427, w_096_6429, w_096_6431, w_096_6433, w_096_6437, w_096_6440, w_096_6447, w_096_6457;
  wire w_097_000, w_097_003, w_097_004, w_097_007, w_097_008, w_097_015, w_097_019, w_097_021, w_097_029, w_097_034, w_097_045, w_097_048, w_097_051, w_097_053, w_097_060, w_097_061, w_097_062, w_097_064, w_097_066, w_097_067, w_097_070, w_097_071, w_097_074, w_097_078, w_097_080, w_097_084, w_097_085, w_097_088, w_097_090, w_097_094, w_097_095, w_097_098, w_097_101, w_097_104, w_097_106, w_097_109, w_097_113, w_097_116, w_097_117, w_097_120, w_097_127, w_097_128, w_097_131, w_097_132, w_097_133, w_097_142, w_097_143, w_097_144, w_097_146, w_097_152, w_097_159, w_097_165, w_097_166, w_097_167, w_097_171, w_097_172, w_097_174, w_097_178, w_097_183, w_097_186, w_097_189, w_097_192, w_097_194, w_097_195, w_097_196, w_097_203, w_097_208, w_097_209, w_097_211, w_097_214, w_097_216, w_097_218, w_097_221, w_097_222, w_097_224, w_097_231, w_097_233, w_097_237, w_097_240, w_097_243, w_097_246, w_097_251, w_097_255, w_097_260, w_097_261, w_097_264, w_097_266, w_097_267, w_097_269, w_097_270, w_097_272, w_097_274, w_097_275, w_097_277, w_097_279, w_097_281, w_097_282, w_097_285, w_097_286, w_097_287, w_097_288, w_097_291, w_097_292, w_097_299, w_097_300, w_097_302, w_097_304, w_097_306, w_097_307, w_097_308, w_097_313, w_097_321, w_097_323, w_097_325, w_097_331, w_097_335, w_097_337, w_097_338, w_097_345, w_097_346, w_097_348, w_097_349, w_097_354, w_097_356, w_097_357, w_097_359, w_097_361, w_097_367, w_097_375, w_097_377, w_097_380, w_097_383, w_097_387, w_097_391, w_097_395, w_097_397, w_097_398, w_097_405, w_097_423, w_097_424, w_097_427, w_097_428, w_097_431, w_097_433, w_097_441, w_097_442, w_097_443, w_097_446, w_097_452, w_097_453, w_097_456, w_097_459, w_097_461, w_097_462, w_097_463, w_097_466, w_097_468, w_097_469, w_097_475, w_097_477, w_097_478, w_097_479, w_097_481, w_097_484, w_097_485, w_097_489, w_097_491, w_097_496, w_097_497, w_097_498, w_097_501, w_097_504, w_097_506, w_097_507, w_097_513, w_097_515, w_097_524, w_097_525, w_097_526, w_097_527, w_097_529, w_097_533, w_097_535, w_097_541, w_097_548, w_097_549, w_097_556, w_097_562, w_097_564, w_097_566, w_097_567, w_097_569, w_097_576, w_097_580, w_097_584, w_097_585, w_097_586, w_097_587, w_097_588, w_097_591, w_097_592, w_097_593, w_097_594, w_097_595, w_097_596, w_097_597, w_097_601, w_097_604, w_097_609, w_097_615, w_097_619, w_097_620, w_097_621, w_097_622, w_097_626, w_097_628, w_097_633, w_097_634, w_097_635, w_097_636, w_097_638, w_097_643, w_097_645, w_097_649, w_097_650, w_097_652, w_097_656, w_097_660, w_097_663, w_097_665, w_097_666, w_097_667, w_097_668, w_097_676, w_097_680, w_097_683, w_097_684, w_097_688, w_097_690, w_097_699, w_097_705, w_097_707, w_097_709, w_097_713, w_097_716, w_097_722, w_097_724, w_097_725, w_097_727, w_097_731, w_097_745, w_097_750, w_097_754, w_097_758, w_097_761, w_097_763, w_097_764, w_097_769, w_097_772, w_097_775, w_097_785, w_097_793, w_097_794, w_097_800, w_097_803, w_097_805, w_097_809, w_097_815, w_097_818, w_097_820, w_097_824, w_097_825, w_097_830, w_097_835, w_097_841, w_097_842, w_097_843, w_097_857, w_097_860, w_097_863, w_097_865, w_097_867, w_097_876, w_097_879, w_097_882, w_097_891, w_097_892, w_097_895, w_097_896, w_097_897, w_097_906, w_097_908, w_097_909, w_097_913, w_097_920, w_097_925, w_097_937, w_097_938, w_097_947, w_097_948, w_097_953, w_097_954, w_097_956, w_097_957, w_097_961, w_097_968, w_097_975, w_097_977, w_097_978, w_097_980, w_097_983, w_097_985, w_097_990, w_097_992, w_097_994, w_097_1003, w_097_1004, w_097_1006, w_097_1007, w_097_1008, w_097_1023, w_097_1024, w_097_1025, w_097_1028, w_097_1029, w_097_1033, w_097_1038, w_097_1042, w_097_1051, w_097_1063, w_097_1066, w_097_1070, w_097_1071, w_097_1073, w_097_1078, w_097_1079, w_097_1082, w_097_1090, w_097_1099, w_097_1106, w_097_1111, w_097_1115, w_097_1116, w_097_1124, w_097_1131, w_097_1139, w_097_1142, w_097_1145, w_097_1150, w_097_1152, w_097_1154, w_097_1161, w_097_1163, w_097_1168, w_097_1169, w_097_1176, w_097_1179, w_097_1188, w_097_1200, w_097_1201, w_097_1203, w_097_1211, w_097_1220, w_097_1222, w_097_1224, w_097_1228, w_097_1232, w_097_1234, w_097_1241, w_097_1243, w_097_1245, w_097_1256, w_097_1257, w_097_1258, w_097_1262, w_097_1264, w_097_1265, w_097_1269, w_097_1282, w_097_1288, w_097_1292, w_097_1299, w_097_1301, w_097_1302, w_097_1306, w_097_1315, w_097_1324, w_097_1328, w_097_1333, w_097_1341, w_097_1354, w_097_1355, w_097_1359, w_097_1360, w_097_1364, w_097_1366, w_097_1371, w_097_1374, w_097_1376, w_097_1379, w_097_1380, w_097_1381, w_097_1385, w_097_1389, w_097_1391, w_097_1400, w_097_1401, w_097_1405, w_097_1410, w_097_1412, w_097_1414, w_097_1418, w_097_1419, w_097_1420, w_097_1421, w_097_1427, w_097_1433, w_097_1443, w_097_1445, w_097_1454, w_097_1455, w_097_1466, w_097_1483, w_097_1484, w_097_1488, w_097_1492, w_097_1494, w_097_1498, w_097_1502, w_097_1506, w_097_1509, w_097_1510, w_097_1511, w_097_1517, w_097_1519, w_097_1525, w_097_1530, w_097_1531, w_097_1542, w_097_1544, w_097_1546, w_097_1556, w_097_1558, w_097_1560, w_097_1563, w_097_1567, w_097_1569, w_097_1573, w_097_1580, w_097_1581, w_097_1585, w_097_1597, w_097_1607, w_097_1608, w_097_1614, w_097_1629, w_097_1634, w_097_1637, w_097_1642, w_097_1645, w_097_1646, w_097_1652, w_097_1656, w_097_1661, w_097_1662, w_097_1671, w_097_1677, w_097_1679, w_097_1680, w_097_1686, w_097_1691, w_097_1692, w_097_1694, w_097_1701, w_097_1703, w_097_1713, w_097_1714, w_097_1719, w_097_1720, w_097_1721, w_097_1722, w_097_1741, w_097_1742, w_097_1749, w_097_1753, w_097_1756, w_097_1761, w_097_1765, w_097_1769, w_097_1770, w_097_1774, w_097_1777, w_097_1778, w_097_1782, w_097_1792, w_097_1803, w_097_1810, w_097_1812, w_097_1813, w_097_1814, w_097_1818, w_097_1836, w_097_1843, w_097_1845, w_097_1853, w_097_1855, w_097_1858, w_097_1859, w_097_1861, w_097_1875, w_097_1879, w_097_1881, w_097_1882, w_097_1889, w_097_1894, w_097_1897, w_097_1902, w_097_1904, w_097_1908, w_097_1914, w_097_1917, w_097_1926, w_097_1940, w_097_1942, w_097_1952, w_097_1963, w_097_1964, w_097_1965, w_097_1966, w_097_1969, w_097_1974, w_097_1978, w_097_1987, w_097_1988, w_097_2009, w_097_2013, w_097_2014, w_097_2025, w_097_2027, w_097_2029, w_097_2046, w_097_2049, w_097_2054, w_097_2061, w_097_2064, w_097_2070, w_097_2071, w_097_2073, w_097_2078, w_097_2080, w_097_2081, w_097_2083, w_097_2097, w_097_2098, w_097_2109, w_097_2110, w_097_2114, w_097_2118, w_097_2129, w_097_2133, w_097_2135, w_097_2140, w_097_2147, w_097_2149, w_097_2150, w_097_2153, w_097_2155, w_097_2157, w_097_2164, w_097_2165, w_097_2166, w_097_2179, w_097_2183, w_097_2188, w_097_2189, w_097_2199, w_097_2204, w_097_2205, w_097_2209, w_097_2214, w_097_2215, w_097_2224, w_097_2227, w_097_2234, w_097_2236, w_097_2241, w_097_2244, w_097_2246, w_097_2248, w_097_2249, w_097_2251, w_097_2266, w_097_2267, w_097_2268, w_097_2271, w_097_2273, w_097_2275, w_097_2276, w_097_2278, w_097_2280, w_097_2282, w_097_2284, w_097_2287, w_097_2293, w_097_2296, w_097_2306, w_097_2309, w_097_2312, w_097_2318, w_097_2320, w_097_2328, w_097_2334, w_097_2337, w_097_2339, w_097_2344, w_097_2349, w_097_2350, w_097_2362, w_097_2373, w_097_2374, w_097_2379, w_097_2393, w_097_2405, w_097_2406, w_097_2432, w_097_2448, w_097_2449, w_097_2452, w_097_2454, w_097_2474, w_097_2475, w_097_2478, w_097_2484, w_097_2485, w_097_2505, w_097_2516, w_097_2517, w_097_2522, w_097_2528, w_097_2529, w_097_2538, w_097_2541, w_097_2542, w_097_2546, w_097_2547, w_097_2549, w_097_2554, w_097_2556, w_097_2562, w_097_2564, w_097_2568, w_097_2569, w_097_2577, w_097_2579, w_097_2585, w_097_2587, w_097_2588, w_097_2589, w_097_2592, w_097_2594, w_097_2596, w_097_2597, w_097_2598, w_097_2603, w_097_2616, w_097_2627, w_097_2631, w_097_2643, w_097_2645, w_097_2647, w_097_2648, w_097_2649, w_097_2652, w_097_2653, w_097_2654, w_097_2659, w_097_2670, w_097_2676, w_097_2677, w_097_2679, w_097_2687, w_097_2688, w_097_2695, w_097_2696, w_097_2699, w_097_2702, w_097_2705, w_097_2707, w_097_2713, w_097_2715, w_097_2719, w_097_2722, w_097_2725, w_097_2727, w_097_2732, w_097_2735, w_097_2740, w_097_2741, w_097_2744, w_097_2745, w_097_2746, w_097_2750, w_097_2753, w_097_2755, w_097_2766, w_097_2774, w_097_2775, w_097_2776, w_097_2779, w_097_2786, w_097_2787, w_097_2789, w_097_2792, w_097_2800, w_097_2801, w_097_2808, w_097_2810, w_097_2817, w_097_2820, w_097_2822, w_097_2823, w_097_2824, w_097_2841, w_097_2855, w_097_2856, w_097_2859, w_097_2861, w_097_2878, w_097_2880, w_097_2884, w_097_2888, w_097_2889, w_097_2890, w_097_2891, w_097_2892, w_097_2907, w_097_2916, w_097_2918, w_097_2921, w_097_2928, w_097_2930, w_097_2931, w_097_2932, w_097_2938, w_097_2939, w_097_2945, w_097_2947, w_097_2948, w_097_2955, w_097_2964, w_097_2965, w_097_2976, w_097_2978, w_097_2981, w_097_2982, w_097_2986, w_097_2994, w_097_2995, w_097_3003, w_097_3009, w_097_3014, w_097_3025, w_097_3029, w_097_3032, w_097_3033, w_097_3045, w_097_3046, w_097_3047, w_097_3049, w_097_3053, w_097_3061, w_097_3064, w_097_3067, w_097_3069, w_097_3072, w_097_3073, w_097_3079, w_097_3087, w_097_3090, w_097_3095, w_097_3096, w_097_3097, w_097_3100, w_097_3107, w_097_3109, w_097_3116, w_097_3117, w_097_3118, w_097_3119, w_097_3121, w_097_3125, w_097_3126, w_097_3128, w_097_3130, w_097_3132, w_097_3143, w_097_3146, w_097_3151, w_097_3154, w_097_3157, w_097_3164, w_097_3169, w_097_3171, w_097_3176, w_097_3180, w_097_3182, w_097_3187, w_097_3193, w_097_3194, w_097_3196, w_097_3202, w_097_3204, w_097_3207, w_097_3208, w_097_3210, w_097_3211, w_097_3218, w_097_3220, w_097_3227, w_097_3233, w_097_3235, w_097_3238, w_097_3248, w_097_3249, w_097_3260, w_097_3265, w_097_3269, w_097_3271, w_097_3274, w_097_3275, w_097_3276, w_097_3277, w_097_3283, w_097_3285, w_097_3286, w_097_3288, w_097_3289, w_097_3290, w_097_3302, w_097_3305, w_097_3310, w_097_3316, w_097_3318, w_097_3322, w_097_3330, w_097_3332, w_097_3343, w_097_3346, w_097_3348, w_097_3351, w_097_3355, w_097_3359, w_097_3369, w_097_3376, w_097_3385, w_097_3387, w_097_3396, w_097_3399, w_097_3402, w_097_3415, w_097_3416, w_097_3420, w_097_3436, w_097_3438, w_097_3446, w_097_3453, w_097_3460, w_097_3465, w_097_3472, w_097_3489, w_097_3496, w_097_3498, w_097_3502, w_097_3508, w_097_3514, w_097_3518, w_097_3527, w_097_3529, w_097_3536, w_097_3537, w_097_3538, w_097_3541, w_097_3548, w_097_3562, w_097_3572, w_097_3574, w_097_3588, w_097_3590, w_097_3596, w_097_3597, w_097_3605, w_097_3616, w_097_3620, w_097_3621, w_097_3624, w_097_3628, w_097_3629, w_097_3635, w_097_3642, w_097_3643, w_097_3647, w_097_3653, w_097_3656, w_097_3672, w_097_3674, w_097_3677, w_097_3680, w_097_3682, w_097_3690, w_097_3695, w_097_3696, w_097_3704, w_097_3712, w_097_3715, w_097_3718, w_097_3720, w_097_3729, w_097_3730, w_097_3734, w_097_3736, w_097_3737, w_097_3743, w_097_3744, w_097_3745, w_097_3747, w_097_3748, w_097_3750, w_097_3753, w_097_3758, w_097_3760, w_097_3764, w_097_3765, w_097_3772, w_097_3782, w_097_3787, w_097_3802, w_097_3804, w_097_3806, w_097_3808, w_097_3809, w_097_3812, w_097_3814, w_097_3816, w_097_3823, w_097_3824, w_097_3829, w_097_3834, w_097_3844, w_097_3845, w_097_3849, w_097_3851, w_097_3859, w_097_3869, w_097_3875, w_097_3878, w_097_3879, w_097_3880, w_097_3885, w_097_3888, w_097_3889, w_097_3890, w_097_3896, w_097_3897, w_097_3900, w_097_3902, w_097_3918, w_097_3921, w_097_3928, w_097_3930, w_097_3931, w_097_3933, w_097_3934, w_097_3940, w_097_3951, w_097_3952, w_097_3953, w_097_3966, w_097_3967, w_097_3969, w_097_3973, w_097_3977, w_097_3979, w_097_3980, w_097_3981, w_097_3998, w_097_4001, w_097_4002, w_097_4006, w_097_4007, w_097_4008, w_097_4010, w_097_4013, w_097_4023, w_097_4025, w_097_4030, w_097_4035, w_097_4036, w_097_4037, w_097_4038, w_097_4044, w_097_4052, w_097_4054, w_097_4056, w_097_4057, w_097_4060, w_097_4067, w_097_4081, w_097_4087, w_097_4090, w_097_4094, w_097_4095, w_097_4106, w_097_4112, w_097_4115, w_097_4126, w_097_4127, w_097_4131, w_097_4133, w_097_4138, w_097_4149, w_097_4157, w_097_4161, w_097_4162, w_097_4166, w_097_4187, w_097_4192, w_097_4193, w_097_4204, w_097_4222, w_097_4226, w_097_4228, w_097_4235, w_097_4240, w_097_4245, w_097_4246, w_097_4247, w_097_4250, w_097_4253, w_097_4254, w_097_4258, w_097_4266, w_097_4269, w_097_4276, w_097_4281, w_097_4282, w_097_4284, w_097_4292, w_097_4308, w_097_4311, w_097_4314, w_097_4319, w_097_4320, w_097_4321, w_097_4330, w_097_4337, w_097_4339, w_097_4340, w_097_4341, w_097_4348, w_097_4349, w_097_4354, w_097_4355, w_097_4358, w_097_4366, w_097_4389, w_097_4390, w_097_4395, w_097_4396, w_097_4397, w_097_4399, w_097_4402, w_097_4411, w_097_4416, w_097_4423, w_097_4424, w_097_4431, w_097_4432, w_097_4435, w_097_4437, w_097_4445, w_097_4454, w_097_4455, w_097_4456, w_097_4472, w_097_4476, w_097_4478, w_097_4484, w_097_4485, w_097_4489, w_097_4493, w_097_4495, w_097_4500, w_097_4502, w_097_4508, w_097_4518, w_097_4519, w_097_4522, w_097_4527, w_097_4530, w_097_4533, w_097_4544, w_097_4548, w_097_4554, w_097_4556, w_097_4562, w_097_4564, w_097_4565, w_097_4567, w_097_4569, w_097_4579, w_097_4580, w_097_4583, w_097_4586, w_097_4588, w_097_4594, w_097_4602, w_097_4603, w_097_4604, w_097_4610, w_097_4614, w_097_4615, w_097_4616, w_097_4621, w_097_4624, w_097_4635, w_097_4641, w_097_4647, w_097_4655, w_097_4662, w_097_4670, w_097_4671, w_097_4673, w_097_4675, w_097_4676, w_097_4684, w_097_4688, w_097_4690, w_097_4694, w_097_4702, w_097_4703, w_097_4706, w_097_4708, w_097_4709, w_097_4719, w_097_4721, w_097_4727, w_097_4730, w_097_4734, w_097_4738, w_097_4747, w_097_4750, w_097_4751, w_097_4757, w_097_4759, w_097_4761, w_097_4763, w_097_4766, w_097_4768, w_097_4770, w_097_4776, w_097_4782, w_097_4784, w_097_4788, w_097_4792, w_097_4797, w_097_4802, w_097_4804, w_097_4808, w_097_4811, w_097_4812, w_097_4813, w_097_4820, w_097_4828, w_097_4829, w_097_4848, w_097_4862, w_097_4865, w_097_4878, w_097_4887, w_097_4895, w_097_4901, w_097_4909, w_097_4910, w_097_4911, w_097_4933, w_097_4934, w_097_4938, w_097_4942, w_097_4945, w_097_4948, w_097_4955, w_097_4971, w_097_4976, w_097_4987, w_097_4988, w_097_4990, w_097_4992, w_097_4993, w_097_4995, w_097_4998, w_097_5008, w_097_5010, w_097_5022, w_097_5023, w_097_5026, w_097_5028, w_097_5030, w_097_5032, w_097_5033, w_097_5037, w_097_5038, w_097_5044, w_097_5052, w_097_5056, w_097_5059, w_097_5060, w_097_5073, w_097_5077, w_097_5080, w_097_5084, w_097_5087, w_097_5088, w_097_5089, w_097_5090, w_097_5093, w_097_5099, w_097_5100, w_097_5111, w_097_5112, w_097_5115, w_097_5118, w_097_5125, w_097_5127, w_097_5130, w_097_5134, w_097_5137, w_097_5144, w_097_5148, w_097_5151, w_097_5153, w_097_5161, w_097_5162, w_097_5168, w_097_5171, w_097_5173, w_097_5174, w_097_5181, w_097_5200, w_097_5201, w_097_5203, w_097_5204, w_097_5205, w_097_5209, w_097_5210, w_097_5213, w_097_5218, w_097_5220, w_097_5221, w_097_5222, w_097_5223, w_097_5228, w_097_5241, w_097_5245, w_097_5256, w_097_5259, w_097_5270, w_097_5275, w_097_5285, w_097_5290, w_097_5291, w_097_5292, w_097_5293, w_097_5296, w_097_5307, w_097_5309, w_097_5316, w_097_5321, w_097_5323, w_097_5325, w_097_5326, w_097_5329, w_097_5330, w_097_5332, w_097_5341, w_097_5344, w_097_5347, w_097_5354, w_097_5355, w_097_5356, w_097_5361, w_097_5370, w_097_5374, w_097_5375, w_097_5380, w_097_5382, w_097_5384, w_097_5387, w_097_5391, w_097_5392, w_097_5395, w_097_5397, w_097_5406, w_097_5407, w_097_5411, w_097_5412, w_097_5413, w_097_5414, w_097_5422, w_097_5425, w_097_5428, w_097_5432, w_097_5433, w_097_5442, w_097_5446, w_097_5452, w_097_5454, w_097_5459, w_097_5463, w_097_5464, w_097_5471, w_097_5477, w_097_5480, w_097_5481, w_097_5482, w_097_5483, w_097_5487, w_097_5491, w_097_5504, w_097_5508, w_097_5509, w_097_5523, w_097_5528, w_097_5531, w_097_5539, w_097_5540, w_097_5541, w_097_5543, w_097_5544, w_097_5552, w_097_5556, w_097_5562, w_097_5577, w_097_5581, w_097_5583, w_097_5584, w_097_5585, w_097_5588, w_097_5589, w_097_5593, w_097_5611, w_097_5616, w_097_5617, w_097_5618, w_097_5619, w_097_5625, w_097_5627, w_097_5634, w_097_5635, w_097_5636, w_097_5645, w_097_5649, w_097_5653, w_097_5659, w_097_5661, w_097_5667, w_097_5668, w_097_5669, w_097_5674, w_097_5677, w_097_5679, w_097_5681, w_097_5683, w_097_5684, w_097_5685, w_097_5686, w_097_5688, w_097_5690, w_097_5693, w_097_5694, w_097_5695, w_097_5705, w_097_5713, w_097_5719, w_097_5727, w_097_5734, w_097_5741, w_097_5745, w_097_5757, w_097_5758, w_097_5760, w_097_5762, w_097_5764, w_097_5767, w_097_5769, w_097_5780, w_097_5781, w_097_5782, w_097_5783, w_097_5794, w_097_5796, w_097_5797, w_097_5801, w_097_5802, w_097_5803, w_097_5811, w_097_5816, w_097_5819, w_097_5834, w_097_5845, w_097_5856, w_097_5868, w_097_5869, w_097_5870, w_097_5872, w_097_5873, w_097_5879, w_097_5881, w_097_5884, w_097_5894, w_097_5904, w_097_5905, w_097_5909, w_097_5913, w_097_5914, w_097_5916, w_097_5918, w_097_5919, w_097_5920, w_097_5922, w_097_5927, w_097_5932, w_097_5934, w_097_5935, w_097_5938, w_097_5955, w_097_5960, w_097_5961, w_097_5964, w_097_5966, w_097_5970, w_097_5975, w_097_5977, w_097_5981, w_097_5989, w_097_6005, w_097_6009, w_097_6012, w_097_6015, w_097_6017, w_097_6019, w_097_6020, w_097_6025, w_097_6033, w_097_6046, w_097_6049, w_097_6050, w_097_6064, w_097_6069, w_097_6070, w_097_6075, w_097_6084, w_097_6087, w_097_6090, w_097_6093, w_097_6097, w_097_6111, w_097_6115, w_097_6116, w_097_6117, w_097_6118, w_097_6124, w_097_6127, w_097_6129, w_097_6130, w_097_6133, w_097_6136, w_097_6145, w_097_6146, w_097_6148, w_097_6155, w_097_6160, w_097_6161, w_097_6163, w_097_6172, w_097_6173, w_097_6174, w_097_6176, w_097_6181, w_097_6182, w_097_6184, w_097_6185, w_097_6187, w_097_6189, w_097_6191, w_097_6193, w_097_6194, w_097_6198, w_097_6201, w_097_6202, w_097_6204, w_097_6205, w_097_6206, w_097_6209, w_097_6212, w_097_6217, w_097_6222, w_097_6234, w_097_6236, w_097_6237, w_097_6243, w_097_6245, w_097_6248, w_097_6250, w_097_6252, w_097_6257, w_097_6276, w_097_6277, w_097_6290, w_097_6293, w_097_6299, w_097_6302, w_097_6303, w_097_6306, w_097_6314, w_097_6315, w_097_6322, w_097_6323, w_097_6329, w_097_6333, w_097_6337, w_097_6339, w_097_6340, w_097_6342, w_097_6351, w_097_6359, w_097_6361, w_097_6370, w_097_6372, w_097_6386, w_097_6391, w_097_6406, w_097_6416, w_097_6425, w_097_6428, w_097_6429, w_097_6435, w_097_6438, w_097_6442, w_097_6446, w_097_6449, w_097_6451, w_097_6455, w_097_6457, w_097_6461, w_097_6468, w_097_6472, w_097_6474, w_097_6475, w_097_6477, w_097_6483, w_097_6485, w_097_6497, w_097_6509, w_097_6512, w_097_6513, w_097_6518, w_097_6522, w_097_6524, w_097_6526, w_097_6530, w_097_6532, w_097_6533, w_097_6534, w_097_6537, w_097_6538, w_097_6546, w_097_6551, w_097_6554, w_097_6558, w_097_6562, w_097_6563, w_097_6567, w_097_6571, w_097_6572, w_097_6573, w_097_6578, w_097_6583, w_097_6598, w_097_6599, w_097_6600, w_097_6610, w_097_6612, w_097_6620, w_097_6621, w_097_6626, w_097_6627, w_097_6629, w_097_6632, w_097_6633, w_097_6634, w_097_6641, w_097_6647, w_097_6651, w_097_6657, w_097_6674, w_097_6679, w_097_6684, w_097_6689, w_097_6694, w_097_6708, w_097_6711, w_097_6713, w_097_6715, w_097_6720, w_097_6724, w_097_6733, w_097_6735, w_097_6738, w_097_6740, w_097_6745, w_097_6747, w_097_6751, w_097_6753, w_097_6754, w_097_6760, w_097_6764, w_097_6765, w_097_6771, w_097_6772, w_097_6775, w_097_6779, w_097_6784, w_097_6794, w_097_6807, w_097_6808, w_097_6810, w_097_6811, w_097_6819, w_097_6822, w_097_6824, w_097_6825, w_097_6826, w_097_6827, w_097_6829, w_097_6830, w_097_6836, w_097_6837, w_097_6840, w_097_6842, w_097_6843, w_097_6845, w_097_6849, w_097_6851, w_097_6858, w_097_6859, w_097_6862, w_097_6867, w_097_6869, w_097_6873, w_097_6877, w_097_6878, w_097_6882, w_097_6884, w_097_6889, w_097_6891, w_097_6896, w_097_6899, w_097_6904, w_097_6908, w_097_6910, w_097_6915, w_097_6917, w_097_6920, w_097_6928, w_097_6929, w_097_6930, w_097_6933, w_097_6940, w_097_6942, w_097_6945, w_097_6946, w_097_6949, w_097_6951, w_097_6953, w_097_6954, w_097_6955, w_097_6956, w_097_6965, w_097_6967, w_097_6968, w_097_6971, w_097_6990, w_097_6999, w_097_7012, w_097_7016, w_097_7024, w_097_7028, w_097_7035, w_097_7040, w_097_7048, w_097_7049, w_097_7052, w_097_7053, w_097_7055, w_097_7061, w_097_7063, w_097_7072, w_097_7073, w_097_7078, w_097_7081, w_097_7092, w_097_7097, w_097_7102, w_097_7113, w_097_7116, w_097_7121, w_097_7122, w_097_7126, w_097_7127, w_097_7146, w_097_7154, w_097_7156, w_097_7158, w_097_7161, w_097_7163, w_097_7164, w_097_7169, w_097_7170, w_097_7171, w_097_7172, w_097_7173, w_097_7190, w_097_7200, w_097_7211, w_097_7221, w_097_7232, w_097_7233, w_097_7237, w_097_7243, w_097_7244, w_097_7250, w_097_7255, w_097_7260, w_097_7262, w_097_7265, w_097_7266, w_097_7274, w_097_7275, w_097_7291, w_097_7292, w_097_7302, w_097_7319, w_097_7322, w_097_7325, w_097_7327, w_097_7337, w_097_7338, w_097_7341, w_097_7344, w_097_7351, w_097_7357, w_097_7358, w_097_7361, w_097_7364, w_097_7372, w_097_7381, w_097_7382, w_097_7383, w_097_7387, w_097_7392, w_097_7399, w_097_7402, w_097_7404, w_097_7408, w_097_7410, w_097_7417, w_097_7419, w_097_7427, w_097_7433, w_097_7436, w_097_7440, w_097_7443, w_097_7446, w_097_7450, w_097_7451, w_097_7454, w_097_7456, w_097_7459, w_097_7460, w_097_7463, w_097_7469, w_097_7475, w_097_7479, w_097_7481, w_097_7485, w_097_7486, w_097_7495, w_097_7497, w_097_7499, w_097_7503, w_097_7504, w_097_7505, w_097_7508, w_097_7512, w_097_7519, w_097_7530, w_097_7534, w_097_7536, w_097_7537, w_097_7538, w_097_7539, w_097_7542, w_097_7554, w_097_7555, w_097_7560, w_097_7562, w_097_7567, w_097_7570, w_097_7572, w_097_7580, w_097_7587, w_097_7588, w_097_7602, w_097_7605, w_097_7610, w_097_7612, w_097_7616, w_097_7617, w_097_7618, w_097_7620, w_097_7628, w_097_7629, w_097_7635, w_097_7640, w_097_7641, w_097_7642, w_097_7644, w_097_7648, w_097_7649, w_097_7650, w_097_7652, w_097_7653, w_097_7666, w_097_7668, w_097_7669, w_097_7672, w_097_7683, w_097_7685, w_097_7687, w_097_7688, w_097_7691, w_097_7702, w_097_7705, w_097_7718, w_097_7728, w_097_7731, w_097_7742, w_097_7746, w_097_7747, w_097_7754, w_097_7757, w_097_7767, w_097_7775, w_097_7784, w_097_7787, w_097_7792, w_097_7794, w_097_7795, w_097_7797, w_097_7810, w_097_7811, w_097_7816, w_097_7817, w_097_7826, w_097_7827, w_097_7828, w_097_7832, w_097_7835, w_097_7838, w_097_7845, w_097_7852, w_097_7856, w_097_7863, w_097_7870, w_097_7871, w_097_7884, w_097_7889, w_097_7897, w_097_7904, w_097_7908, w_097_7911, w_097_7913, w_097_7916, w_097_7917, w_097_7925, w_097_7926, w_097_7927, w_097_7928, w_097_7936, w_097_7938, w_097_7939, w_097_7952, w_097_7953, w_097_7958, w_097_7959, w_097_7961, w_097_7962, w_097_7974, w_097_7979, w_097_7982, w_097_7983, w_097_7985, w_097_7988, w_097_7993, w_097_7996, w_097_7997, w_097_8005, w_097_8010, w_097_8015, w_097_8018, w_097_8019, w_097_8037, w_097_8044, w_097_8045, w_097_8054, w_097_8059, w_097_8060, w_097_8065, w_097_8067, w_097_8069, w_097_8084, w_097_8090, w_097_8092, w_097_8093, w_097_8099, w_097_8103, w_097_8110, w_097_8114, w_097_8117, w_097_8123, w_097_8128, w_097_8136, w_097_8142, w_097_8144, w_097_8145, w_097_8148, w_097_8151, w_097_8162, w_097_8165, w_097_8171, w_097_8175, w_097_8186, w_097_8189, w_097_8191, w_097_8194, w_097_8196, w_097_8197, w_097_8198, w_097_8201, w_097_8202, w_097_8203, w_097_8206, w_097_8216, w_097_8217, w_097_8224, w_097_8226, w_097_8229, w_097_8231, w_097_8237, w_097_8240, w_097_8243, w_097_8245, w_097_8248, w_097_8253, w_097_8255, w_097_8257, w_097_8262, w_097_8277, w_097_8279, w_097_8280, w_097_8282, w_097_8293, w_097_8300, w_097_8301, w_097_8304, w_097_8306, w_097_8307, w_097_8308, w_097_8312, w_097_8313, w_097_8314, w_097_8321, w_097_8331, w_097_8332, w_097_8335, w_097_8348, w_097_8354, w_097_8357, w_097_8359, w_097_8364, w_097_8378, w_097_8379, w_097_8390, w_097_8392, w_097_8406, w_097_8416, w_097_8427, w_097_8434, w_097_8435, w_097_8441, w_097_8447, w_097_8452, w_097_8454, w_097_8458, w_097_8465, w_097_8473, w_097_8474, w_097_8476, w_097_8482, w_097_8491, w_097_8493, w_097_8494, w_097_8498, w_097_8504, w_097_8509, w_097_8512, w_097_8517, w_097_8519, w_097_8529, w_097_8533, w_097_8537, w_097_8546, w_097_8548, w_097_8551, w_097_8556, w_097_8558, w_097_8560, w_097_8561, w_097_8562, w_097_8570, w_097_8574, w_097_8576, w_097_8577, w_097_8579, w_097_8585, w_097_8586, w_097_8590, w_097_8595, w_097_8605, w_097_8610, w_097_8614, w_097_8616, w_097_8620, w_097_8621, w_097_8623, w_097_8624, w_097_8629, w_097_8630, w_097_8638, w_097_8644, w_097_8647, w_097_8649, w_097_8655, w_097_8667, w_097_8668, w_097_8671, w_097_8674, w_097_8678, w_097_8686, w_097_8688, w_097_8690, w_097_8698, w_097_8702, w_097_8707, w_097_8712, w_097_8716, w_097_8717, w_097_8721, w_097_8725, w_097_8727, w_097_8728, w_097_8738, w_097_8740, w_097_8745, w_097_8752, w_097_8753, w_097_8759, w_097_8765, w_097_8772, w_097_8773, w_097_8779, w_097_8784, w_097_8793, w_097_8797, w_097_8809, w_097_8811, w_097_8819, w_097_8822, w_097_8836, w_097_8838, w_097_8839, w_097_8840, w_097_8843, w_097_8854, w_097_8858, w_097_8860, w_097_8866, w_097_8867, w_097_8870, w_097_8874, w_097_8877, w_097_8891, w_097_8893, w_097_8903, w_097_8906, w_097_8909, w_097_8914, w_097_8925, w_097_8932, w_097_8939, w_097_8945, w_097_8958, w_097_8963, w_097_8975, w_097_8977, w_097_8978, w_097_8984, w_097_8985, w_097_8986, w_097_8987, w_097_8988, w_097_8990, w_097_8991, w_097_9001, w_097_9002, w_097_9003, w_097_9005, w_097_9006, w_097_9015, w_097_9027, w_097_9030, w_097_9032, w_097_9034, w_097_9035, w_097_9045, w_097_9053, w_097_9066, w_097_9070, w_097_9079, w_097_9081, w_097_9084, w_097_9088, w_097_9093, w_097_9104, w_097_9107, w_097_9109, w_097_9115, w_097_9121, w_097_9131, w_097_9133, w_097_9138, w_097_9139, w_097_9141, w_097_9150, w_097_9152, w_097_9156, w_097_9160, w_097_9161, w_097_9165, w_097_9166, w_097_9175, w_097_9176, w_097_9178, w_097_9180, w_097_9182, w_097_9185, w_097_9203, w_097_9205, w_097_9209, w_097_9211, w_097_9214, w_097_9217, w_097_9220, w_097_9225, w_097_9229, w_097_9230, w_097_9231, w_097_9233, w_097_9234, w_097_9235, w_097_9239, w_097_9242, w_097_9247, w_097_9249, w_097_9257, w_097_9261, w_097_9263, w_097_9264, w_097_9267, w_097_9272, w_097_9277, w_097_9282, w_097_9289, w_097_9299, w_097_9304, w_097_9308, w_097_9311, w_097_9323, w_097_9328, w_097_9330;
  wire w_098_003, w_098_005, w_098_007, w_098_008, w_098_009, w_098_010, w_098_012, w_098_017, w_098_022, w_098_024, w_098_025, w_098_035, w_098_037, w_098_040, w_098_045, w_098_050, w_098_053, w_098_055, w_098_056, w_098_058, w_098_060, w_098_061, w_098_062, w_098_064, w_098_067, w_098_069, w_098_071, w_098_075, w_098_076, w_098_078, w_098_081, w_098_082, w_098_086, w_098_087, w_098_089, w_098_091, w_098_097, w_098_101, w_098_102, w_098_103, w_098_106, w_098_107, w_098_109, w_098_111, w_098_113, w_098_116, w_098_119, w_098_120, w_098_121, w_098_122, w_098_124, w_098_134, w_098_135, w_098_136, w_098_138, w_098_139, w_098_142, w_098_143, w_098_148, w_098_149, w_098_150, w_098_153, w_098_154, w_098_155, w_098_157, w_098_159, w_098_160, w_098_161, w_098_170, w_098_172, w_098_178, w_098_181, w_098_182, w_098_189, w_098_191, w_098_192, w_098_194, w_098_197, w_098_199, w_098_200, w_098_201, w_098_203, w_098_205, w_098_207, w_098_209, w_098_213, w_098_214, w_098_222, w_098_225, w_098_230, w_098_232, w_098_238, w_098_239, w_098_241, w_098_246, w_098_249, w_098_250, w_098_252, w_098_255, w_098_261, w_098_262, w_098_269, w_098_270, w_098_271, w_098_272, w_098_279, w_098_282, w_098_284, w_098_287, w_098_288, w_098_289, w_098_292, w_098_293, w_098_294, w_098_298, w_098_299, w_098_300, w_098_301, w_098_304, w_098_307, w_098_309, w_098_311, w_098_314, w_098_315, w_098_316, w_098_318, w_098_319, w_098_323, w_098_324, w_098_328, w_098_329, w_098_330, w_098_333, w_098_341, w_098_343, w_098_344, w_098_350, w_098_352, w_098_353, w_098_358, w_098_359, w_098_364, w_098_367, w_098_371, w_098_375, w_098_376, w_098_378, w_098_379, w_098_380, w_098_382, w_098_384, w_098_385, w_098_386, w_098_387, w_098_389, w_098_394, w_098_395, w_098_397, w_098_398, w_098_400, w_098_401, w_098_402, w_098_403, w_098_404, w_098_407, w_098_408, w_098_411, w_098_413, w_098_415, w_098_417, w_098_419, w_098_420, w_098_421, w_098_422, w_098_424, w_098_425, w_098_429, w_098_430, w_098_431, w_098_432, w_098_434, w_098_436, w_098_437, w_098_439, w_098_445, w_098_447, w_098_449, w_098_450, w_098_457, w_098_466, w_098_487, w_098_494, w_098_499, w_098_502, w_098_504, w_098_507, w_098_511, w_098_513, w_098_516, w_098_518, w_098_520, w_098_522, w_098_525, w_098_531, w_098_532, w_098_534, w_098_538, w_098_543, w_098_544, w_098_548, w_098_550, w_098_551, w_098_558, w_098_560, w_098_563, w_098_569, w_098_573, w_098_578, w_098_583, w_098_586, w_098_601, w_098_607, w_098_609, w_098_611, w_098_616, w_098_617, w_098_626, w_098_628, w_098_629, w_098_632, w_098_636, w_098_639, w_098_658, w_098_660, w_098_665, w_098_667, w_098_668, w_098_678, w_098_682, w_098_683, w_098_684, w_098_689, w_098_690, w_098_696, w_098_703, w_098_706, w_098_710, w_098_712, w_098_717, w_098_728, w_098_731, w_098_735, w_098_738, w_098_739, w_098_743, w_098_745, w_098_752, w_098_756, w_098_757, w_098_758, w_098_763, w_098_766, w_098_774, w_098_775, w_098_781, w_098_804, w_098_806, w_098_807, w_098_808, w_098_810, w_098_812, w_098_816, w_098_818, w_098_821, w_098_822, w_098_834, w_098_845, w_098_850, w_098_858, w_098_860, w_098_862, w_098_871, w_098_875, w_098_876, w_098_878, w_098_879, w_098_880, w_098_884, w_098_885, w_098_888, w_098_889, w_098_895, w_098_899, w_098_900, w_098_903, w_098_912, w_098_937, w_098_940, w_098_941, w_098_947, w_098_953, w_098_963, w_098_964, w_098_966, w_098_967, w_098_968, w_098_971, w_098_980, w_098_989, w_098_996, w_098_999, w_098_1000, w_098_1005, w_098_1007, w_098_1010, w_098_1012, w_098_1015, w_098_1023, w_098_1029, w_098_1036, w_098_1039, w_098_1040, w_098_1041, w_098_1044, w_098_1051, w_098_1057, w_098_1061, w_098_1066, w_098_1067, w_098_1068, w_098_1070, w_098_1073, w_098_1074, w_098_1076, w_098_1081, w_098_1085, w_098_1088, w_098_1093, w_098_1099, w_098_1101, w_098_1103, w_098_1104, w_098_1110, w_098_1120, w_098_1125, w_098_1128, w_098_1130, w_098_1131, w_098_1145, w_098_1147, w_098_1148, w_098_1155, w_098_1156, w_098_1161, w_098_1165, w_098_1167, w_098_1177, w_098_1179, w_098_1199, w_098_1209, w_098_1214, w_098_1215, w_098_1216, w_098_1217, w_098_1237, w_098_1238, w_098_1244, w_098_1251, w_098_1252, w_098_1253, w_098_1259, w_098_1262, w_098_1264, w_098_1268, w_098_1271, w_098_1275, w_098_1283, w_098_1288, w_098_1298, w_098_1301, w_098_1315, w_098_1318, w_098_1320, w_098_1322, w_098_1323, w_098_1328, w_098_1329, w_098_1333, w_098_1334, w_098_1337, w_098_1340, w_098_1350, w_098_1354, w_098_1362, w_098_1363, w_098_1364, w_098_1366, w_098_1371, w_098_1372, w_098_1375, w_098_1376, w_098_1377, w_098_1378, w_098_1379, w_098_1385, w_098_1387, w_098_1396, w_098_1400, w_098_1408, w_098_1410, w_098_1413, w_098_1423, w_098_1425, w_098_1427, w_098_1434, w_098_1436, w_098_1441, w_098_1444, w_098_1446, w_098_1449, w_098_1460, w_098_1465, w_098_1474, w_098_1476, w_098_1480, w_098_1484, w_098_1492, w_098_1494, w_098_1502, w_098_1504, w_098_1508, w_098_1513, w_098_1522, w_098_1524, w_098_1532, w_098_1547, w_098_1549, w_098_1558, w_098_1560, w_098_1567, w_098_1568, w_098_1573, w_098_1575, w_098_1576, w_098_1579, w_098_1584, w_098_1588, w_098_1592, w_098_1609, w_098_1614, w_098_1619, w_098_1620, w_098_1621, w_098_1628, w_098_1630, w_098_1640, w_098_1643, w_098_1650, w_098_1652, w_098_1654, w_098_1656, w_098_1663, w_098_1665, w_098_1685, w_098_1687, w_098_1693, w_098_1694, w_098_1698, w_098_1703, w_098_1712, w_098_1713, w_098_1715, w_098_1717, w_098_1724, w_098_1726, w_098_1728, w_098_1742, w_098_1750, w_098_1756, w_098_1758, w_098_1765, w_098_1775, w_098_1787, w_098_1790, w_098_1795, w_098_1797, w_098_1802, w_098_1806, w_098_1816, w_098_1818, w_098_1820, w_098_1829, w_098_1830, w_098_1831, w_098_1837, w_098_1838, w_098_1848, w_098_1850, w_098_1858, w_098_1860, w_098_1861, w_098_1866, w_098_1871, w_098_1874, w_098_1883, w_098_1886, w_098_1888, w_098_1892, w_098_1893, w_098_1896, w_098_1897, w_098_1899, w_098_1900, w_098_1906, w_098_1908, w_098_1912, w_098_1923, w_098_1928, w_098_1931, w_098_1942, w_098_1948, w_098_1950, w_098_1954, w_098_1956, w_098_1957, w_098_1968, w_098_1969, w_098_1970, w_098_1971, w_098_1974, w_098_1978, w_098_1984, w_098_1989, w_098_1992, w_098_1994, w_098_1996, w_098_2001, w_098_2004, w_098_2005, w_098_2013, w_098_2016, w_098_2032, w_098_2033, w_098_2034, w_098_2035, w_098_2049, w_098_2053, w_098_2054, w_098_2059, w_098_2063, w_098_2066, w_098_2071, w_098_2074, w_098_2085, w_098_2089, w_098_2091, w_098_2094, w_098_2096, w_098_2099, w_098_2101, w_098_2104, w_098_2106, w_098_2108, w_098_2109, w_098_2112, w_098_2115, w_098_2133, w_098_2144, w_098_2153, w_098_2158, w_098_2165, w_098_2175, w_098_2176, w_098_2177, w_098_2181, w_098_2188, w_098_2196, w_098_2198, w_098_2204, w_098_2210, w_098_2216, w_098_2223, w_098_2227, w_098_2236, w_098_2238, w_098_2239, w_098_2241, w_098_2242, w_098_2245, w_098_2251, w_098_2252, w_098_2255, w_098_2262, w_098_2274, w_098_2275, w_098_2277, w_098_2283, w_098_2284, w_098_2285, w_098_2288, w_098_2290, w_098_2297, w_098_2301, w_098_2302, w_098_2305, w_098_2306, w_098_2308, w_098_2310, w_098_2312, w_098_2316, w_098_2330, w_098_2331, w_098_2333, w_098_2338, w_098_2341, w_098_2342, w_098_2348, w_098_2353, w_098_2356, w_098_2363, w_098_2372, w_098_2384, w_098_2388, w_098_2390, w_098_2392, w_098_2402, w_098_2403, w_098_2408, w_098_2410, w_098_2416, w_098_2422, w_098_2429, w_098_2437, w_098_2441, w_098_2445, w_098_2449, w_098_2451, w_098_2455, w_098_2457, w_098_2458, w_098_2467, w_098_2469, w_098_2470, w_098_2482, w_098_2484, w_098_2486, w_098_2487, w_098_2492, w_098_2497, w_098_2507, w_098_2518, w_098_2530, w_098_2532, w_098_2560, w_098_2561, w_098_2563, w_098_2571, w_098_2574, w_098_2584, w_098_2589, w_098_2590, w_098_2603, w_098_2612, w_098_2614, w_098_2616, w_098_2625, w_098_2629, w_098_2630, w_098_2639, w_098_2643, w_098_2644, w_098_2645, w_098_2647, w_098_2649, w_098_2653, w_098_2659, w_098_2666, w_098_2667, w_098_2669, w_098_2670, w_098_2681, w_098_2691, w_098_2692, w_098_2701, w_098_2702, w_098_2706, w_098_2708, w_098_2721, w_098_2722, w_098_2731, w_098_2734, w_098_2742, w_098_2750, w_098_2753, w_098_2759, w_098_2762, w_098_2764, w_098_2768, w_098_2769, w_098_2773, w_098_2780, w_098_2781, w_098_2786, w_098_2787, w_098_2788, w_098_2789, w_098_2790, w_098_2792, w_098_2812, w_098_2813, w_098_2818, w_098_2820, w_098_2821, w_098_2822, w_098_2827, w_098_2830, w_098_2831, w_098_2833, w_098_2834, w_098_2836, w_098_2846, w_098_2850, w_098_2860, w_098_2861, w_098_2862, w_098_2863, w_098_2864, w_098_2869, w_098_2878, w_098_2881, w_098_2889, w_098_2890, w_098_2894, w_098_2896, w_098_2901, w_098_2908, w_098_2918, w_098_2926, w_098_2928, w_098_2938, w_098_2939, w_098_2941, w_098_2942, w_098_2945, w_098_2947, w_098_2949, w_098_2952, w_098_2955, w_098_2958, w_098_2964, w_098_2967, w_098_2968, w_098_2970, w_098_2972, w_098_2974, w_098_2978, w_098_2979, w_098_2981, w_098_2987, w_098_2997, w_098_3000, w_098_3001, w_098_3003, w_098_3015, w_098_3016, w_098_3022, w_098_3023, w_098_3029, w_098_3036, w_098_3043, w_098_3045, w_098_3047, w_098_3054, w_098_3055, w_098_3059, w_098_3060, w_098_3067, w_098_3068, w_098_3079, w_098_3080, w_098_3084, w_098_3094, w_098_3098, w_098_3104, w_098_3106, w_098_3109, w_098_3112, w_098_3118, w_098_3119, w_098_3120, w_098_3125, w_098_3131, w_098_3132, w_098_3144, w_098_3150, w_098_3151, w_098_3160, w_098_3161, w_098_3164, w_098_3165, w_098_3171, w_098_3173, w_098_3179, w_098_3180, w_098_3190, w_098_3192, w_098_3198, w_098_3209, w_098_3210, w_098_3215, w_098_3229, w_098_3230, w_098_3231, w_098_3239, w_098_3246, w_098_3248, w_098_3249, w_098_3251, w_098_3255, w_098_3262, w_098_3263, w_098_3265, w_098_3267, w_098_3284, w_098_3293, w_098_3294, w_098_3301, w_098_3308, w_098_3309, w_098_3314, w_098_3315, w_098_3316, w_098_3320, w_098_3321, w_098_3328, w_098_3329, w_098_3332, w_098_3335, w_098_3343, w_098_3344, w_098_3347, w_098_3349, w_098_3350, w_098_3360, w_098_3374, w_098_3378, w_098_3379, w_098_3381, w_098_3394, w_098_3403, w_098_3412, w_098_3414, w_098_3415, w_098_3416, w_098_3424, w_098_3432, w_098_3433, w_098_3439, w_098_3440, w_098_3447, w_098_3459, w_098_3465, w_098_3467, w_098_3468, w_098_3472, w_098_3474, w_098_3479, w_098_3481, w_098_3484, w_098_3490, w_098_3491, w_098_3496, w_098_3505, w_098_3517, w_098_3523, w_098_3531, w_098_3537, w_098_3538, w_098_3541, w_098_3544, w_098_3545, w_098_3548, w_098_3551, w_098_3552, w_098_3557, w_098_3559, w_098_3562, w_098_3568, w_098_3570, w_098_3575, w_098_3578, w_098_3580, w_098_3585, w_098_3586, w_098_3592, w_098_3595, w_098_3596, w_098_3597, w_098_3600, w_098_3602, w_098_3608, w_098_3610, w_098_3611, w_098_3612, w_098_3618, w_098_3621, w_098_3622, w_098_3625, w_098_3626, w_098_3628, w_098_3634, w_098_3641, w_098_3642, w_098_3644, w_098_3654, w_098_3657, w_098_3658, w_098_3662, w_098_3663, w_098_3665, w_098_3670, w_098_3690, w_098_3701, w_098_3710, w_098_3716, w_098_3719, w_098_3723, w_098_3726, w_098_3727, w_098_3731, w_098_3732, w_098_3735, w_098_3737, w_098_3746, w_098_3757, w_098_3761, w_098_3766, w_098_3768, w_098_3772, w_098_3787, w_098_3792, w_098_3793, w_098_3794, w_098_3802, w_098_3803, w_098_3810, w_098_3813, w_098_3816, w_098_3822, w_098_3827, w_098_3835, w_098_3836, w_098_3844, w_098_3845, w_098_3847, w_098_3850, w_098_3853, w_098_3868, w_098_3869, w_098_3871, w_098_3880, w_098_3881, w_098_3883, w_098_3884, w_098_3886, w_098_3892, w_098_3895, w_098_3905, w_098_3914, w_098_3927, w_098_3938, w_098_3952, w_098_3954, w_098_3955, w_098_3972, w_098_3974, w_098_3977, w_098_3980, w_098_3982, w_098_3986, w_098_3988, w_098_3993, w_098_4000, w_098_4001, w_098_4002, w_098_4007, w_098_4011, w_098_4014, w_098_4020, w_098_4022, w_098_4026, w_098_4028, w_098_4030, w_098_4035, w_098_4037, w_098_4038, w_098_4041, w_098_4046, w_098_4054, w_098_4056, w_098_4059, w_098_4081, w_098_4085, w_098_4087, w_098_4091, w_098_4098, w_098_4099, w_098_4108, w_098_4119, w_098_4127, w_098_4132, w_098_4133, w_098_4137, w_098_4142, w_098_4143, w_098_4149, w_098_4162, w_098_4165, w_098_4169, w_098_4182, w_098_4183, w_098_4189, w_098_4191, w_098_4193, w_098_4196, w_098_4197, w_098_4199, w_098_4206, w_098_4208, w_098_4217, w_098_4229, w_098_4233, w_098_4238, w_098_4240, w_098_4242, w_098_4244, w_098_4246, w_098_4247, w_098_4251, w_098_4255, w_098_4256, w_098_4258, w_098_4261, w_098_4274, w_098_4275, w_098_4277, w_098_4280, w_098_4282, w_098_4287, w_098_4291, w_098_4292, w_098_4297, w_098_4306, w_098_4307, w_098_4310, w_098_4311, w_098_4319, w_098_4327, w_098_4328, w_098_4333, w_098_4335, w_098_4339, w_098_4348, w_098_4352, w_098_4353, w_098_4355, w_098_4357, w_098_4358, w_098_4366, w_098_4367, w_098_4368, w_098_4370, w_098_4372, w_098_4373, w_098_4374, w_098_4379, w_098_4382, w_098_4383, w_098_4388, w_098_4403, w_098_4404, w_098_4416, w_098_4420, w_098_4423, w_098_4428, w_098_4442, w_098_4443, w_098_4447, w_098_4451, w_098_4452, w_098_4458, w_098_4462, w_098_4466, w_098_4473, w_098_4475, w_098_4476, w_098_4478, w_098_4480, w_098_4486, w_098_4500, w_098_4502, w_098_4517, w_098_4519, w_098_4520, w_098_4525, w_098_4535, w_098_4537, w_098_4538, w_098_4545, w_098_4547, w_098_4550, w_098_4552, w_098_4560, w_098_4561, w_098_4563, w_098_4566, w_098_4570, w_098_4572, w_098_4576, w_098_4577, w_098_4579, w_098_4582, w_098_4583, w_098_4587, w_098_4590, w_098_4598, w_098_4599, w_098_4601, w_098_4604, w_098_4609, w_098_4618, w_098_4625, w_098_4626, w_098_4633, w_098_4634, w_098_4636, w_098_4640, w_098_4641, w_098_4642, w_098_4645, w_098_4653, w_098_4667, w_098_4672, w_098_4681, w_098_4698, w_098_4706, w_098_4717, w_098_4718, w_098_4720, w_098_4725, w_098_4729, w_098_4731, w_098_4732, w_098_4735, w_098_4736, w_098_4740, w_098_4741, w_098_4749, w_098_4754, w_098_4758, w_098_4762, w_098_4763, w_098_4766, w_098_4769, w_098_4774, w_098_4778, w_098_4782, w_098_4788, w_098_4796, w_098_4802, w_098_4809, w_098_4810, w_098_4815, w_098_4816, w_098_4818, w_098_4822, w_098_4828, w_098_4831, w_098_4832, w_098_4833, w_098_4835, w_098_4844, w_098_4845, w_098_4846, w_098_4860, w_098_4861, w_098_4863, w_098_4868, w_098_4870, w_098_4880, w_098_4882, w_098_4884, w_098_4888, w_098_4889, w_098_4903, w_098_4911, w_098_4912, w_098_4914, w_098_4918, w_098_4919, w_098_4922, w_098_4925, w_098_4926, w_098_4927, w_098_4928, w_098_4932, w_098_4933, w_098_4940, w_098_4953, w_098_4954, w_098_4955, w_098_4956, w_098_4961, w_098_4962, w_098_4964, w_098_4968, w_098_4969, w_098_4978, w_098_4985, w_098_4995, w_098_4998, w_098_5008, w_098_5009, w_098_5012, w_098_5024, w_098_5025, w_098_5026, w_098_5027, w_098_5030, w_098_5037, w_098_5040, w_098_5045, w_098_5047, w_098_5051, w_098_5052, w_098_5053, w_098_5054, w_098_5056, w_098_5071, w_098_5079, w_098_5080, w_098_5084, w_098_5089, w_098_5090, w_098_5091, w_098_5092, w_098_5094, w_098_5126, w_098_5132, w_098_5133, w_098_5137, w_098_5142, w_098_5149, w_098_5154, w_098_5157, w_098_5158, w_098_5159, w_098_5160, w_098_5166, w_098_5172, w_098_5174, w_098_5183, w_098_5193, w_098_5209, w_098_5212, w_098_5213, w_098_5217, w_098_5220, w_098_5229, w_098_5230, w_098_5240, w_098_5243, w_098_5247, w_098_5252, w_098_5253, w_098_5255, w_098_5257, w_098_5265, w_098_5267, w_098_5269, w_098_5275, w_098_5279, w_098_5288, w_098_5290, w_098_5294, w_098_5306, w_098_5314, w_098_5316, w_098_5319, w_098_5323, w_098_5325, w_098_5334, w_098_5341, w_098_5343, w_098_5346, w_098_5352, w_098_5358, w_098_5361, w_098_5365, w_098_5371, w_098_5375, w_098_5376, w_098_5379, w_098_5380, w_098_5381, w_098_5384, w_098_5387, w_098_5393, w_098_5396, w_098_5403, w_098_5405, w_098_5406, w_098_5409, w_098_5413, w_098_5414, w_098_5417, w_098_5421, w_098_5426, w_098_5429, w_098_5438, w_098_5439, w_098_5441, w_098_5447, w_098_5450, w_098_5467, w_098_5469, w_098_5476, w_098_5478, w_098_5482, w_098_5508, w_098_5509, w_098_5510, w_098_5512, w_098_5513, w_098_5515, w_098_5516, w_098_5517, w_098_5527, w_098_5531, w_098_5533, w_098_5537, w_098_5538, w_098_5540, w_098_5543, w_098_5551, w_098_5552, w_098_5557, w_098_5569, w_098_5572, w_098_5579, w_098_5581, w_098_5590, w_098_5594, w_098_5595, w_098_5599, w_098_5605, w_098_5608, w_098_5614, w_098_5615, w_098_5618, w_098_5619, w_098_5624, w_098_5628, w_098_5632, w_098_5635, w_098_5638, w_098_5643, w_098_5645, w_098_5648, w_098_5657, w_098_5659, w_098_5663, w_098_5671, w_098_5675, w_098_5679, w_098_5685, w_098_5688, w_098_5692, w_098_5696, w_098_5698, w_098_5699, w_098_5707, w_098_5708, w_098_5714, w_098_5717, w_098_5720, w_098_5721, w_098_5725, w_098_5727, w_098_5728, w_098_5742, w_098_5745, w_098_5750, w_098_5752, w_098_5754, w_098_5756, w_098_5760, w_098_5766, w_098_5772, w_098_5779, w_098_5783, w_098_5786, w_098_5789, w_098_5797, w_098_5811, w_098_5821, w_098_5823, w_098_5828, w_098_5833, w_098_5837, w_098_5838, w_098_5841, w_098_5842, w_098_5849, w_098_5855, w_098_5857, w_098_5866, w_098_5868, w_098_5869, w_098_5872, w_098_5879, w_098_5882, w_098_5883, w_098_5890, w_098_5891, w_098_5892, w_098_5894, w_098_5906, w_098_5920, w_098_5922, w_098_5924, w_098_5927, w_098_5934, w_098_5941, w_098_5948, w_098_5949, w_098_5950, w_098_5957, w_098_5964, w_098_5965, w_098_5970, w_098_5973, w_098_5977, w_098_5980, w_098_5985, w_098_6004, w_098_6011, w_098_6013, w_098_6014, w_098_6025, w_098_6037, w_098_6038, w_098_6042, w_098_6043, w_098_6046, w_098_6053, w_098_6056, w_098_6066, w_098_6067, w_098_6068, w_098_6069, w_098_6070, w_098_6079, w_098_6082, w_098_6084, w_098_6087, w_098_6090, w_098_6109, w_098_6110, w_098_6112, w_098_6114, w_098_6117, w_098_6118, w_098_6125, w_098_6131, w_098_6132, w_098_6133, w_098_6134, w_098_6135, w_098_6155, w_098_6156, w_098_6163, w_098_6165, w_098_6170, w_098_6171, w_098_6181, w_098_6191, w_098_6194, w_098_6196, w_098_6200, w_098_6203, w_098_6207, w_098_6209, w_098_6211, w_098_6212, w_098_6216, w_098_6219, w_098_6220, w_098_6221, w_098_6223, w_098_6226, w_098_6236, w_098_6244, w_098_6250, w_098_6253, w_098_6271, w_098_6275, w_098_6277, w_098_6280, w_098_6284, w_098_6290, w_098_6291, w_098_6292, w_098_6305, w_098_6319, w_098_6324, w_098_6325, w_098_6326, w_098_6327, w_098_6328, w_098_6333, w_098_6334, w_098_6356, w_098_6357, w_098_6361, w_098_6368, w_098_6378, w_098_6380, w_098_6382, w_098_6384, w_098_6385, w_098_6390, w_098_6391, w_098_6394, w_098_6406, w_098_6410, w_098_6417, w_098_6418, w_098_6425, w_098_6430, w_098_6433, w_098_6435, w_098_6438, w_098_6445, w_098_6455, w_098_6461, w_098_6462, w_098_6482, w_098_6486, w_098_6492, w_098_6494, w_098_6496, w_098_6498, w_098_6503, w_098_6506, w_098_6507, w_098_6508, w_098_6509, w_098_6516, w_098_6519, w_098_6523, w_098_6524, w_098_6526, w_098_6536, w_098_6539, w_098_6541, w_098_6549, w_098_6551, w_098_6555, w_098_6556, w_098_6558, w_098_6562, w_098_6578, w_098_6581, w_098_6582, w_098_6585, w_098_6590, w_098_6596, w_098_6604, w_098_6611, w_098_6612, w_098_6614, w_098_6615, w_098_6618, w_098_6619, w_098_6622, w_098_6623, w_098_6627, w_098_6628, w_098_6629, w_098_6647, w_098_6655, w_098_6657, w_098_6659, w_098_6663, w_098_6671, w_098_6672, w_098_6677, w_098_6678, w_098_6682, w_098_6695, w_098_6709, w_098_6711, w_098_6722, w_098_6723, w_098_6725, w_098_6730, w_098_6732, w_098_6738, w_098_6743, w_098_6744, w_098_6745, w_098_6746, w_098_6747, w_098_6752, w_098_6755, w_098_6757, w_098_6770, w_098_6800, w_098_6817, w_098_6818, w_098_6820, w_098_6823, w_098_6826, w_098_6837, w_098_6838, w_098_6839, w_098_6841, w_098_6848, w_098_6855, w_098_6858, w_098_6859, w_098_6860, w_098_6861, w_098_6862, w_098_6865, w_098_6867, w_098_6869, w_098_6872, w_098_6896, w_098_6899, w_098_6910, w_098_6912, w_098_6921, w_098_6924, w_098_6925, w_098_6931, w_098_6936, w_098_6938, w_098_6941, w_098_6942, w_098_6946, w_098_6959, w_098_6960, w_098_6961, w_098_6962, w_098_6976, w_098_6977, w_098_6993, w_098_6998, w_098_7006, w_098_7022, w_098_7023, w_098_7026, w_098_7034, w_098_7041, w_098_7043, w_098_7049, w_098_7052, w_098_7058, w_098_7069, w_098_7070, w_098_7075, w_098_7079, w_098_7089, w_098_7091, w_098_7097, w_098_7103, w_098_7110, w_098_7114, w_098_7116, w_098_7129, w_098_7131, w_098_7132, w_098_7136, w_098_7137, w_098_7145, w_098_7146, w_098_7150, w_098_7155, w_098_7156, w_098_7157, w_098_7163, w_098_7179, w_098_7190, w_098_7193, w_098_7199, w_098_7209, w_098_7212, w_098_7217, w_098_7222, w_098_7223, w_098_7227, w_098_7230, w_098_7247, w_098_7248, w_098_7252, w_098_7259, w_098_7265, w_098_7266, w_098_7268, w_098_7271, w_098_7273, w_098_7274, w_098_7275, w_098_7294, w_098_7301, w_098_7303, w_098_7304, w_098_7309, w_098_7312, w_098_7314, w_098_7321, w_098_7323, w_098_7327, w_098_7329, w_098_7331, w_098_7338, w_098_7345, w_098_7350, w_098_7353, w_098_7357, w_098_7362, w_098_7377, w_098_7385, w_098_7386, w_098_7387, w_098_7388, w_098_7394, w_098_7396, w_098_7397, w_098_7400, w_098_7413, w_098_7424, w_098_7427, w_098_7437, w_098_7447, w_098_7457, w_098_7462, w_098_7465, w_098_7466, w_098_7467, w_098_7474, w_098_7475, w_098_7477, w_098_7480, w_098_7482, w_098_7486, w_098_7489, w_098_7495, w_098_7496, w_098_7498, w_098_7499, w_098_7506, w_098_7517, w_098_7519, w_098_7524, w_098_7527, w_098_7530, w_098_7537, w_098_7555, w_098_7563, w_098_7566, w_098_7574, w_098_7579, w_098_7581, w_098_7582, w_098_7588, w_098_7591, w_098_7594, w_098_7595, w_098_7596, w_098_7600, w_098_7612, w_098_7614, w_098_7616, w_098_7620, w_098_7621, w_098_7622, w_098_7627, w_098_7633, w_098_7635, w_098_7640, w_098_7643, w_098_7644, w_098_7649, w_098_7654, w_098_7655, w_098_7659, w_098_7663, w_098_7668, w_098_7674, w_098_7680, w_098_7686, w_098_7692, w_098_7700, w_098_7704, w_098_7707, w_098_7713, w_098_7718, w_098_7730, w_098_7734, w_098_7735, w_098_7742, w_098_7751, w_098_7756, w_098_7761, w_098_7764, w_098_7770, w_098_7771, w_098_7773, w_098_7779, w_098_7781, w_098_7782, w_098_7787, w_098_7793, w_098_7795, w_098_7799, w_098_7805, w_098_7812, w_098_7813, w_098_7815, w_098_7830, w_098_7835, w_098_7839, w_098_7846, w_098_7852, w_098_7856, w_098_7857, w_098_7858, w_098_7860, w_098_7862, w_098_7866, w_098_7873, w_098_7876, w_098_7877, w_098_7881, w_098_7888, w_098_7894, w_098_7897, w_098_7907, w_098_7909, w_098_7910, w_098_7914, w_098_7918, w_098_7920, w_098_7922, w_098_7923, w_098_7924, w_098_7930, w_098_7933, w_098_7937, w_098_7940, w_098_7943, w_098_7945, w_098_7946, w_098_7955, w_098_7960, w_098_7961, w_098_7975, w_098_7976, w_098_7979, w_098_7982, w_098_7986, w_098_7989, w_098_7991, w_098_7996, w_098_8004, w_098_8011, w_098_8016, w_098_8018, w_098_8028, w_098_8029, w_098_8031, w_098_8035, w_098_8037, w_098_8044, w_098_8047, w_098_8049, w_098_8055, w_098_8056, w_098_8057, w_098_8059, w_098_8066, w_098_8094, w_098_8099, w_098_8100, w_098_8104, w_098_8106, w_098_8108, w_098_8111, w_098_8116, w_098_8117, w_098_8122, w_098_8124, w_098_8125, w_098_8127, w_098_8131, w_098_8132, w_098_8133, w_098_8137, w_098_8152, w_098_8161, w_098_8165, w_098_8166, w_098_8170, w_098_8172, w_098_8176, w_098_8178, w_098_8180, w_098_8182, w_098_8183, w_098_8186, w_098_8188, w_098_8203, w_098_8215, w_098_8219, w_098_8223, w_098_8224, w_098_8225, w_098_8227, w_098_8237, w_098_8242, w_098_8244, w_098_8245, w_098_8246, w_098_8247, w_098_8250, w_098_8257, w_098_8270, w_098_8283, w_098_8284, w_098_8287, w_098_8288, w_098_8306, w_098_8314, w_098_8324, w_098_8327, w_098_8332, w_098_8335, w_098_8344, w_098_8346, w_098_8355, w_098_8356, w_098_8378, w_098_8380, w_098_8391, w_098_8401, w_098_8406, w_098_8407, w_098_8413, w_098_8416, w_098_8418, w_098_8422, w_098_8425, w_098_8427, w_098_8435, w_098_8436, w_098_8439, w_098_8440, w_098_8444, w_098_8451, w_098_8453, w_098_8458, w_098_8460, w_098_8462, w_098_8463, w_098_8476, w_098_8478, w_098_8479, w_098_8481, w_098_8482, w_098_8484, w_098_8488, w_098_8490, w_098_8492, w_098_8502, w_098_8503, w_098_8506, w_098_8507, w_098_8508, w_098_8510, w_098_8519, w_098_8521, w_098_8528, w_098_8531, w_098_8535, w_098_8538, w_098_8543, w_098_8544, w_098_8545, w_098_8551, w_098_8552, w_098_8555, w_098_8559, w_098_8561, w_098_8566, w_098_8582, w_098_8583, w_098_8592, w_098_8596, w_098_8602, w_098_8603, w_098_8606, w_098_8610, w_098_8620, w_098_8625, w_098_8633, w_098_8635, w_098_8638, w_098_8640, w_098_8642, w_098_8656, w_098_8668, w_098_8669, w_098_8671, w_098_8672, w_098_8676, w_098_8681, w_098_8686, w_098_8692, w_098_8694, w_098_8700, w_098_8703, w_098_8705, w_098_8715, w_098_8716, w_098_8717, w_098_8719, w_098_8731, w_098_8734, w_098_8745, w_098_8751, w_098_8753, w_098_8754, w_098_8764, w_098_8772, w_098_8773, w_098_8786, w_098_8787, w_098_8789, w_098_8794, w_098_8797, w_098_8801, w_098_8807, w_098_8821, w_098_8830, w_098_8835, w_098_8837, w_098_8842, w_098_8848, w_098_8849, w_098_8851, w_098_8853, w_098_8863, w_098_8865, w_098_8868, w_098_8877, w_098_8879, w_098_8880, w_098_8882, w_098_8890, w_098_8891, w_098_8895, w_098_8897, w_098_8899, w_098_8902, w_098_8908, w_098_8909, w_098_8911, w_098_8914, w_098_8920, w_098_8933, w_098_8936, w_098_8937, w_098_8939, w_098_8941, w_098_8945, w_098_8951, w_098_8955, w_098_8961, w_098_8967, w_098_8970, w_098_8972, w_098_8993, w_098_8998, w_098_9002, w_098_9007, w_098_9012, w_098_9013, w_098_9014, w_098_9015, w_098_9017, w_098_9018, w_098_9028, w_098_9032, w_098_9039, w_098_9048, w_098_9051, w_098_9052, w_098_9067, w_098_9068, w_098_9071, w_098_9075, w_098_9078, w_098_9081, w_098_9086, w_098_9088, w_098_9095, w_098_9100, w_098_9109, w_098_9112, w_098_9115, w_098_9123, w_098_9131, w_098_9132, w_098_9134, w_098_9145, w_098_9164, w_098_9168, w_098_9172, w_098_9174, w_098_9176, w_098_9178, w_098_9184, w_098_9199, w_098_9206, w_098_9207, w_098_9217, w_098_9219, w_098_9222, w_098_9231, w_098_9234, w_098_9239, w_098_9242, w_098_9245, w_098_9247, w_098_9253, w_098_9261, w_098_9262, w_098_9269, w_098_9272, w_098_9273, w_098_9279, w_098_9280, w_098_9286, w_098_9291, w_098_9294, w_098_9295, w_098_9303, w_098_9306, w_098_9308, w_098_9310, w_098_9318, w_098_9330, w_098_9331, w_098_9332, w_098_9336, w_098_9337, w_098_9342, w_098_9343, w_098_9350, w_098_9359, w_098_9360, w_098_9362, w_098_9371, w_098_9374, w_098_9377, w_098_9381, w_098_9384, w_098_9386, w_098_9399, w_098_9401, w_098_9402, w_098_9404, w_098_9407, w_098_9420, w_098_9421, w_098_9422, w_098_9438, w_098_9442, w_098_9449, w_098_9454, w_098_9455, w_098_9458, w_098_9468, w_098_9474, w_098_9476, w_098_9480, w_098_9483, w_098_9484, w_098_9492, w_098_9498, w_098_9502, w_098_9504, w_098_9506, w_098_9507, w_098_9513, w_098_9521, w_098_9536, w_098_9548;
  wire w_099_000, w_099_007, w_099_009, w_099_013, w_099_014, w_099_017, w_099_018, w_099_020, w_099_023, w_099_031, w_099_033, w_099_039, w_099_043, w_099_044, w_099_045, w_099_047, w_099_048, w_099_049, w_099_052, w_099_060, w_099_061, w_099_063, w_099_065, w_099_066, w_099_067, w_099_068, w_099_074, w_099_076, w_099_077, w_099_081, w_099_084, w_099_085, w_099_090, w_099_093, w_099_094, w_099_095, w_099_096, w_099_099, w_099_105, w_099_106, w_099_110, w_099_111, w_099_113, w_099_117, w_099_121, w_099_122, w_099_123, w_099_124, w_099_128, w_099_132, w_099_133, w_099_134, w_099_135, w_099_137, w_099_138, w_099_139, w_099_142, w_099_146, w_099_148, w_099_150, w_099_152, w_099_153, w_099_154, w_099_155, w_099_156, w_099_158, w_099_163, w_099_166, w_099_168, w_099_170, w_099_173, w_099_175, w_099_176, w_099_180, w_099_183, w_099_184, w_099_185, w_099_186, w_099_190, w_099_191, w_099_195, w_099_198, w_099_202, w_099_205, w_099_208, w_099_217, w_099_218, w_099_221, w_099_223, w_099_224, w_099_227, w_099_231, w_099_234, w_099_236, w_099_248, w_099_249, w_099_250, w_099_251, w_099_258, w_099_260, w_099_263, w_099_271, w_099_273, w_099_274, w_099_275, w_099_278, w_099_281, w_099_283, w_099_285, w_099_288, w_099_289, w_099_292, w_099_293, w_099_294, w_099_295, w_099_298, w_099_299, w_099_304, w_099_313, w_099_315, w_099_316, w_099_317, w_099_321, w_099_325, w_099_329, w_099_331, w_099_332, w_099_333, w_099_337, w_099_339, w_099_342, w_099_345, w_099_348, w_099_350, w_099_354, w_099_356, w_099_357, w_099_361, w_099_365, w_099_372, w_099_375, w_099_377, w_099_379, w_099_382, w_099_383, w_099_385, w_099_388, w_099_391, w_099_397, w_099_403, w_099_404, w_099_405, w_099_406, w_099_408, w_099_409, w_099_412, w_099_415, w_099_416, w_099_419, w_099_421, w_099_430, w_099_433, w_099_437, w_099_443, w_099_448, w_099_451, w_099_452, w_099_456, w_099_457, w_099_458, w_099_462, w_099_464, w_099_465, w_099_474, w_099_475, w_099_478, w_099_481, w_099_482, w_099_487, w_099_488, w_099_489, w_099_495, w_099_496, w_099_497, w_099_498, w_099_499, w_099_501, w_099_505, w_099_506, w_099_507, w_099_511, w_099_515, w_099_516, w_099_517, w_099_519, w_099_529, w_099_531, w_099_532, w_099_534, w_099_540, w_099_544, w_099_551, w_099_552, w_099_553, w_099_554, w_099_556, w_099_560, w_099_561, w_099_562, w_099_563, w_099_564, w_099_569, w_099_573, w_099_576, w_099_578, w_099_581, w_099_583, w_099_584, w_099_585, w_099_588, w_099_593, w_099_595, w_099_596, w_099_597, w_099_599, w_099_606, w_099_607, w_099_611, w_099_612, w_099_613, w_099_617, w_099_618, w_099_619, w_099_621, w_099_626, w_099_627, w_099_629, w_099_630, w_099_634, w_099_635, w_099_638, w_099_640, w_099_643, w_099_645, w_099_646, w_099_647, w_099_649, w_099_654, w_099_656, w_099_662, w_099_664, w_099_666, w_099_667, w_099_669, w_099_672, w_099_673, w_099_675, w_099_676, w_099_678, w_099_679, w_099_685, w_099_692, w_099_694, w_099_699, w_099_703, w_099_708, w_099_715, w_099_717, w_099_719, w_099_720, w_099_721, w_099_726, w_099_727, w_099_728, w_099_734, w_099_735, w_099_736, w_099_740, w_099_742, w_099_743, w_099_745, w_099_746, w_099_749, w_099_750, w_099_751, w_099_752, w_099_755, w_099_760, w_099_761, w_099_763, w_099_765, w_099_766, w_099_767, w_099_769, w_099_770, w_099_773, w_099_777, w_099_784, w_099_785, w_099_788, w_099_790, w_099_791, w_099_792, w_099_793, w_099_794, w_099_795, w_099_798, w_099_799, w_099_804, w_099_808, w_099_809, w_099_811, w_099_814, w_099_819, w_099_820, w_099_821, w_099_826, w_099_827, w_099_828, w_099_829, w_099_836, w_099_839, w_099_840, w_099_843, w_099_857, w_099_862, w_099_864, w_099_865, w_099_866, w_099_867, w_099_869, w_099_870, w_099_871, w_099_875, w_099_878, w_099_885, w_099_888, w_099_894, w_099_896, w_099_898, w_099_905, w_099_906, w_099_907, w_099_910, w_099_911, w_099_912, w_099_913, w_099_915, w_099_916, w_099_918, w_099_920, w_099_923, w_099_927, w_099_929, w_099_931, w_099_933, w_099_935, w_099_939, w_099_941, w_099_944, w_099_945, w_099_947, w_099_948, w_099_951, w_099_952, w_099_954, w_099_957, w_099_959, w_099_960, w_099_962, w_099_963, w_099_964, w_099_965, w_099_969, w_099_970, w_099_971, w_099_979, w_099_981, w_099_983, w_099_984, w_099_986, w_099_989, w_099_990, w_099_991, w_099_992, w_099_1002, w_099_1005, w_099_1008, w_099_1010, w_099_1012, w_099_1013, w_099_1015, w_099_1016, w_099_1017, w_099_1019, w_099_1021, w_099_1025, w_099_1026, w_099_1027, w_099_1029, w_099_1030, w_099_1037, w_099_1040, w_099_1042, w_099_1045, w_099_1047, w_099_1048, w_099_1051, w_099_1055, w_099_1056, w_099_1057, w_099_1061, w_099_1063, w_099_1066, w_099_1071, w_099_1074, w_099_1076, w_099_1077, w_099_1079, w_099_1080, w_099_1087, w_099_1088, w_099_1091, w_099_1093, w_099_1096, w_099_1099, w_099_1107, w_099_1109, w_099_1110, w_099_1125, w_099_1128, w_099_1130, w_099_1131, w_099_1133, w_099_1136, w_099_1137, w_099_1139, w_099_1141, w_099_1145, w_099_1148, w_099_1151, w_099_1156, w_099_1157, w_099_1159, w_099_1161, w_099_1162, w_099_1168, w_099_1171, w_099_1176, w_099_1180, w_099_1184, w_099_1188, w_099_1189, w_099_1200, w_099_1207, w_099_1209, w_099_1210, w_099_1213, w_099_1215, w_099_1216, w_099_1217, w_099_1218, w_099_1221, w_099_1223, w_099_1225, w_099_1229, w_099_1231, w_099_1234, w_099_1241, w_099_1243, w_099_1247, w_099_1254, w_099_1255, w_099_1256, w_099_1260, w_099_1262, w_099_1263, w_099_1264, w_099_1267, w_099_1269, w_099_1271, w_099_1272, w_099_1273, w_099_1275, w_099_1279, w_099_1283, w_099_1285, w_099_1291, w_099_1293, w_099_1295, w_099_1298, w_099_1299, w_099_1304, w_099_1305, w_099_1312, w_099_1313, w_099_1314, w_099_1318, w_099_1319, w_099_1320, w_099_1321, w_099_1322, w_099_1323, w_099_1326, w_099_1330, w_099_1331, w_099_1332, w_099_1335, w_099_1338, w_099_1342, w_099_1344, w_099_1348, w_099_1349, w_099_1350, w_099_1353, w_099_1355, w_099_1359, w_099_1360, w_099_1365, w_099_1367, w_099_1369, w_099_1370, w_099_1372, w_099_1380, w_099_1382, w_099_1383, w_099_1384, w_099_1392, w_099_1401, w_099_1402, w_099_1404, w_099_1408, w_099_1409, w_099_1416, w_099_1417, w_099_1418, w_099_1422, w_099_1423, w_099_1424, w_099_1427, w_099_1428, w_099_1433, w_099_1435, w_099_1438, w_099_1441, w_099_1442, w_099_1444, w_099_1445, w_099_1449, w_099_1451, w_099_1452, w_099_1453, w_099_1455, w_099_1463, w_099_1464, w_099_1465, w_099_1466, w_099_1468, w_099_1473, w_099_1474, w_099_1475, w_099_1476, w_099_1481, w_099_1483, w_099_1484, w_099_1488, w_099_1489, w_099_1492, w_099_1499, w_099_1501, w_099_1503, w_099_1504, w_099_1506, w_099_1508, w_099_1511, w_099_1514, w_099_1515, w_099_1516, w_099_1522, w_099_1523, w_099_1529, w_099_1531, w_099_1538, w_099_1539, w_099_1540, w_099_1544, w_099_1547, w_099_1548, w_099_1549, w_099_1550, w_099_1551, w_099_1558, w_099_1559, w_099_1560, w_099_1561, w_099_1564, w_099_1565, w_099_1568, w_099_1570, w_099_1585, w_099_1587, w_099_1588, w_099_1589, w_099_1591, w_099_1596, w_099_1598, w_099_1599, w_099_1600, w_099_1601, w_099_1602, w_099_1607, w_099_1611, w_099_1614, w_099_1617, w_099_1625, w_099_1628, w_099_1631, w_099_1634, w_099_1635, w_099_1636, w_099_1637, w_099_1638, w_099_1642, w_099_1649, w_099_1650, w_099_1651, w_099_1654, w_099_1655, w_099_1658, w_099_1659, w_099_1663, w_099_1665, w_099_1666, w_099_1669, w_099_1670, w_099_1671, w_099_1672, w_099_1674, w_099_1679, w_099_1681, w_099_1684, w_099_1685, w_099_1686, w_099_1688, w_099_1689, w_099_1690, w_099_1691, w_099_1693, w_099_1694, w_099_1698, w_099_1699, w_099_1703, w_099_1705, w_099_1713, w_099_1717, w_099_1724, w_099_1726, w_099_1730, w_099_1733, w_099_1734, w_099_1736, w_099_1737, w_099_1738, w_099_1740, w_099_1749, w_099_1751, w_099_1753, w_099_1754, w_099_1755, w_099_1759, w_099_1760, w_099_1761, w_099_1767, w_099_1774, w_099_1776, w_099_1777, w_099_1779, w_099_1780, w_099_1781, w_099_1782, w_099_1783, w_099_1784, w_099_1789, w_099_1790, w_099_1799, w_099_1801, w_099_1802, w_099_1808, w_099_1813, w_099_1816, w_099_1820, w_099_1822, w_099_1823, w_099_1827, w_099_1828, w_099_1829, w_099_1831, w_099_1833, w_099_1834, w_099_1836, w_099_1839, w_099_1840, w_099_1841, w_099_1847, w_099_1862, w_099_1864, w_099_1868, w_099_1871, w_099_1875, w_099_1878, w_099_1881, w_099_1885, w_099_1890, w_099_1894, w_099_1902, w_099_1905, w_099_1908, w_099_1909, w_099_1913, w_099_1917, w_099_1920, w_099_1922, w_099_1929, w_099_1931, w_099_1932, w_099_1941, w_099_1943, w_099_1945, w_099_1946, w_099_1949, w_099_1951, w_099_1952, w_099_1961, w_099_1962, w_099_1963, w_099_1967, w_099_1982, w_099_1984, w_099_1997, w_099_2004, w_099_2006, w_099_2007, w_099_2008, w_099_2010, w_099_2012, w_099_2013, w_099_2020, w_099_2022, w_099_2024, w_099_2033, w_099_2043, w_099_2044, w_099_2045, w_099_2051, w_099_2052, w_099_2055, w_099_2057, w_099_2060, w_099_2064, w_099_2065, w_099_2069, w_099_2070, w_099_2083, w_099_2084, w_099_2088, w_099_2089, w_099_2090, w_099_2091, w_099_2095, w_099_2097, w_099_2099, w_099_2102, w_099_2108, w_099_2109, w_099_2110, w_099_2112, w_099_2120, w_099_2128, w_099_2132, w_099_2133, w_099_2136, w_099_2138, w_099_2145, w_099_2146, w_099_2147, w_099_2148, w_099_2155, w_099_2157, w_099_2167, w_099_2169, w_099_2170, w_099_2178, w_099_2179, w_099_2181, w_099_2183, w_099_2185, w_099_2197, w_099_2205, w_099_2220, w_099_2222, w_099_2232, w_099_2235, w_099_2237, w_099_2240, w_099_2246, w_099_2252, w_099_2263, w_099_2266, w_099_2273, w_099_2282, w_099_2284, w_099_2285, w_099_2288, w_099_2294, w_099_2295, w_099_2297, w_099_2299, w_099_2300, w_099_2302, w_099_2306, w_099_2308, w_099_2311, w_099_2322, w_099_2326, w_099_2327, w_099_2328, w_099_2341, w_099_2345, w_099_2346, w_099_2347, w_099_2349, w_099_2350, w_099_2351, w_099_2353, w_099_2357, w_099_2364, w_099_2365, w_099_2386, w_099_2391, w_099_2398, w_099_2415, w_099_2416, w_099_2420, w_099_2422, w_099_2427, w_099_2428, w_099_2429, w_099_2430, w_099_2441, w_099_2442, w_099_2444, w_099_2448, w_099_2454, w_099_2456, w_099_2458, w_099_2463, w_099_2464, w_099_2467, w_099_2468, w_099_2473, w_099_2474, w_099_2477, w_099_2486, w_099_2490, w_099_2500, w_099_2501, w_099_2510, w_099_2512, w_099_2528, w_099_2529, w_099_2536, w_099_2539, w_099_2541, w_099_2552, w_099_2553, w_099_2559, w_099_2567, w_099_2569, w_099_2576, w_099_2577, w_099_2583, w_099_2586, w_099_2589, w_099_2590, w_099_2591, w_099_2610, w_099_2615, w_099_2629, w_099_2632, w_099_2635, w_099_2637, w_099_2642, w_099_2648, w_099_2651, w_099_2656, w_099_2658, w_099_2662, w_099_2665, w_099_2674, w_099_2676, w_099_2682, w_099_2686, w_099_2687, w_099_2688, w_099_2694, w_099_2699, w_099_2707, w_099_2715, w_099_2730, w_099_2733, w_099_2735, w_099_2736, w_099_2737, w_099_2738, w_099_2747, w_099_2749, w_099_2761, w_099_2768, w_099_2771, w_099_2780, w_099_2785, w_099_2789, w_099_2792, w_099_2794, w_099_2795, w_099_2823, w_099_2825, w_099_2827, w_099_2828, w_099_2840, w_099_2854, w_099_2855, w_099_2863, w_099_2872, w_099_2874, w_099_2878, w_099_2880, w_099_2883, w_099_2888, w_099_2895, w_099_2907, w_099_2913, w_099_2914, w_099_2915, w_099_2917, w_099_2918, w_099_2922, w_099_2923, w_099_2924, w_099_2928, w_099_2931, w_099_2932, w_099_2933, w_099_2936, w_099_2939, w_099_2940, w_099_2959, w_099_2966, w_099_2969, w_099_2971, w_099_2974, w_099_2985, w_099_2986, w_099_2989, w_099_2991, w_099_2993, w_099_3002, w_099_3007, w_099_3012, w_099_3015, w_099_3029, w_099_3032, w_099_3033, w_099_3043, w_099_3045, w_099_3047, w_099_3048, w_099_3050, w_099_3053, w_099_3063, w_099_3064, w_099_3068, w_099_3074, w_099_3075, w_099_3079, w_099_3080, w_099_3081, w_099_3092, w_099_3097, w_099_3100, w_099_3111, w_099_3112, w_099_3114, w_099_3118, w_099_3119, w_099_3123, w_099_3129, w_099_3131, w_099_3137, w_099_3145, w_099_3147, w_099_3150, w_099_3152, w_099_3160, w_099_3168, w_099_3182, w_099_3188, w_099_3199, w_099_3210, w_099_3211, w_099_3224, w_099_3229, w_099_3243, w_099_3247, w_099_3262, w_099_3264, w_099_3270, w_099_3279, w_099_3286, w_099_3294, w_099_3296, w_099_3299, w_099_3301, w_099_3302, w_099_3306, w_099_3307, w_099_3308, w_099_3310, w_099_3318, w_099_3326, w_099_3339, w_099_3343, w_099_3349, w_099_3351, w_099_3354, w_099_3358, w_099_3359, w_099_3361, w_099_3364, w_099_3365, w_099_3383, w_099_3384, w_099_3386, w_099_3388, w_099_3398, w_099_3401, w_099_3408, w_099_3409, w_099_3411, w_099_3419, w_099_3428, w_099_3431, w_099_3435, w_099_3439, w_099_3448, w_099_3450, w_099_3458, w_099_3462, w_099_3466, w_099_3469, w_099_3472, w_099_3473, w_099_3474, w_099_3482, w_099_3483, w_099_3484, w_099_3487, w_099_3488, w_099_3494, w_099_3496, w_099_3498, w_099_3502, w_099_3506, w_099_3507, w_099_3510, w_099_3513, w_099_3516, w_099_3526, w_099_3534, w_099_3536, w_099_3539, w_099_3541, w_099_3543, w_099_3545, w_099_3548, w_099_3549, w_099_3550, w_099_3552, w_099_3572, w_099_3578, w_099_3582, w_099_3584, w_099_3587, w_099_3599, w_099_3606, w_099_3623, w_099_3635, w_099_3639, w_099_3648, w_099_3649, w_099_3651, w_099_3652, w_099_3657, w_099_3661, w_099_3666, w_099_3667, w_099_3668, w_099_3674, w_099_3679, w_099_3689, w_099_3690, w_099_3703, w_099_3704, w_099_3705, w_099_3708, w_099_3709, w_099_3710, w_099_3712, w_099_3713, w_099_3714, w_099_3716, w_099_3722, w_099_3723, w_099_3730, w_099_3763, w_099_3775, w_099_3778, w_099_3785, w_099_3791, w_099_3795, w_099_3796, w_099_3807, w_099_3814, w_099_3819, w_099_3824, w_099_3826, w_099_3834, w_099_3851, w_099_3854, w_099_3855, w_099_3862, w_099_3863, w_099_3864, w_099_3865, w_099_3876, w_099_3878, w_099_3880, w_099_3882, w_099_3891, w_099_3894, w_099_3897, w_099_3901, w_099_3904, w_099_3909, w_099_3910, w_099_3919, w_099_3922, w_099_3923, w_099_3926, w_099_3937, w_099_3939, w_099_3942, w_099_3948, w_099_3960, w_099_3963, w_099_3970, w_099_3985, w_099_3987, w_099_3990, w_099_3991, w_099_3995, w_099_3999, w_099_4002, w_099_4019, w_099_4024, w_099_4027, w_099_4028, w_099_4032, w_099_4035, w_099_4043, w_099_4045, w_099_4051, w_099_4053, w_099_4058, w_099_4059, w_099_4064, w_099_4072, w_099_4075, w_099_4076, w_099_4077, w_099_4079, w_099_4080, w_099_4086, w_099_4087, w_099_4088, w_099_4089, w_099_4092, w_099_4096, w_099_4100, w_099_4102, w_099_4103, w_099_4107, w_099_4114, w_099_4118, w_099_4124, w_099_4127, w_099_4133, w_099_4137, w_099_4139, w_099_4147, w_099_4150, w_099_4156, w_099_4157, w_099_4160, w_099_4171, w_099_4173, w_099_4175, w_099_4184, w_099_4186, w_099_4192, w_099_4194, w_099_4195, w_099_4196, w_099_4205, w_099_4206, w_099_4207, w_099_4211, w_099_4212, w_099_4224, w_099_4226, w_099_4227, w_099_4234, w_099_4238, w_099_4243, w_099_4250, w_099_4253, w_099_4255, w_099_4256, w_099_4257, w_099_4260, w_099_4272, w_099_4277, w_099_4278, w_099_4280, w_099_4285, w_099_4286, w_099_4287, w_099_4294, w_099_4296, w_099_4297, w_099_4299, w_099_4304, w_099_4305, w_099_4315, w_099_4322, w_099_4332, w_099_4333, w_099_4344, w_099_4345, w_099_4353, w_099_4355, w_099_4356, w_099_4364, w_099_4365, w_099_4370, w_099_4374, w_099_4375, w_099_4379, w_099_4382, w_099_4384, w_099_4386, w_099_4387, w_099_4389, w_099_4391, w_099_4394, w_099_4395, w_099_4403, w_099_4406, w_099_4408, w_099_4413, w_099_4417, w_099_4419, w_099_4420, w_099_4424, w_099_4428, w_099_4430, w_099_4431, w_099_4432, w_099_4440, w_099_4442, w_099_4444, w_099_4452, w_099_4454, w_099_4456, w_099_4457, w_099_4459, w_099_4460, w_099_4468, w_099_4470, w_099_4474, w_099_4475, w_099_4480, w_099_4484, w_099_4485, w_099_4491, w_099_4495, w_099_4496, w_099_4498, w_099_4505, w_099_4511, w_099_4514, w_099_4522, w_099_4526, w_099_4545, w_099_4547, w_099_4549, w_099_4550, w_099_4557, w_099_4566, w_099_4573, w_099_4576, w_099_4578, w_099_4583, w_099_4586, w_099_4588, w_099_4592, w_099_4594, w_099_4603, w_099_4607, w_099_4626, w_099_4640, w_099_4643, w_099_4648, w_099_4659, w_099_4661, w_099_4664, w_099_4666, w_099_4668, w_099_4679, w_099_4681, w_099_4683, w_099_4688, w_099_4692, w_099_4696, w_099_4697, w_099_4702, w_099_4704, w_099_4710, w_099_4713, w_099_4727, w_099_4732, w_099_4733, w_099_4735, w_099_4740, w_099_4748, w_099_4755, w_099_4756, w_099_4762, w_099_4763, w_099_4766, w_099_4771, w_099_4772, w_099_4776, w_099_4777, w_099_4780, w_099_4783, w_099_4785, w_099_4788, w_099_4789, w_099_4792, w_099_4795, w_099_4805, w_099_4809, w_099_4810, w_099_4813, w_099_4814, w_099_4817, w_099_4824, w_099_4829, w_099_4834, w_099_4836, w_099_4837, w_099_4840, w_099_4843, w_099_4845, w_099_4847, w_099_4849, w_099_4851, w_099_4857, w_099_4863, w_099_4864, w_099_4867, w_099_4877, w_099_4884, w_099_4886, w_099_4888, w_099_4889, w_099_4895, w_099_4903, w_099_4906, w_099_4908, w_099_4909, w_099_4910, w_099_4916, w_099_4919, w_099_4921, w_099_4923, w_099_4934, w_099_4937, w_099_4939, w_099_4945, w_099_4951, w_099_4954, w_099_4956, w_099_4964, w_099_4966, w_099_4970, w_099_4972, w_099_4974, w_099_4984, w_099_4987, w_099_4988, w_099_4999, w_099_5000, w_099_5003, w_099_5006, w_099_5009, w_099_5012, w_099_5021, w_099_5023, w_099_5030, w_099_5042, w_099_5046, w_099_5051, w_099_5052, w_099_5056, w_099_5057, w_099_5069, w_099_5071, w_099_5072, w_099_5078, w_099_5087, w_099_5091, w_099_5093, w_099_5095, w_099_5102, w_099_5104, w_099_5105, w_099_5107, w_099_5116, w_099_5124, w_099_5131, w_099_5135, w_099_5141, w_099_5143, w_099_5146, w_099_5147, w_099_5148, w_099_5149, w_099_5151, w_099_5156, w_099_5158, w_099_5165, w_099_5167, w_099_5184, w_099_5194, w_099_5196, w_099_5197, w_099_5214, w_099_5219, w_099_5221, w_099_5226, w_099_5233, w_099_5235, w_099_5236, w_099_5251, w_099_5252, w_099_5254, w_099_5256, w_099_5265, w_099_5270, w_099_5277, w_099_5280, w_099_5282, w_099_5283, w_099_5289, w_099_5294, w_099_5295, w_099_5299, w_099_5303, w_099_5304, w_099_5308, w_099_5309, w_099_5312, w_099_5319, w_099_5325, w_099_5332, w_099_5338, w_099_5340, w_099_5349, w_099_5353, w_099_5355, w_099_5356, w_099_5360, w_099_5362, w_099_5365, w_099_5369, w_099_5370, w_099_5372, w_099_5375, w_099_5376, w_099_5382, w_099_5385, w_099_5388, w_099_5397, w_099_5400, w_099_5407, w_099_5409, w_099_5414, w_099_5420, w_099_5424, w_099_5425, w_099_5428, w_099_5440, w_099_5444, w_099_5446, w_099_5456, w_099_5463, w_099_5466, w_099_5468, w_099_5476, w_099_5485, w_099_5486, w_099_5490, w_099_5495, w_099_5503, w_099_5522, w_099_5532, w_099_5546, w_099_5555, w_099_5557, w_099_5559, w_099_5564, w_099_5566, w_099_5570, w_099_5572, w_099_5581, w_099_5583, w_099_5588, w_099_5590, w_099_5603, w_099_5606, w_099_5608, w_099_5611, w_099_5617, w_099_5621, w_099_5640, w_099_5649, w_099_5669, w_099_5679, w_099_5684, w_099_5689, w_099_5694, w_099_5695, w_099_5697, w_099_5705, w_099_5708, w_099_5711, w_099_5720, w_099_5728, w_099_5731, w_099_5733, w_099_5737, w_099_5747, w_099_5748, w_099_5749, w_099_5750, w_099_5754, w_099_5755, w_099_5757, w_099_5758, w_099_5760, w_099_5766, w_099_5767, w_099_5768, w_099_5770, w_099_5776, w_099_5779, w_099_5792, w_099_5797, w_099_5798, w_099_5801, w_099_5813, w_099_5814, w_099_5824, w_099_5825, w_099_5826, w_099_5834, w_099_5841, w_099_5850, w_099_5854, w_099_5855, w_099_5856, w_099_5866, w_099_5871, w_099_5873, w_099_5875, w_099_5883, w_099_5884, w_099_5895, w_099_5898, w_099_5907, w_099_5915, w_099_5922, w_099_5929, w_099_5932, w_099_5939, w_099_5944, w_099_5954, w_099_5956, w_099_5959, w_099_5968, w_099_5970, w_099_5973, w_099_5974, w_099_5978, w_099_5982, w_099_5989, w_099_5992, w_099_5997, w_099_5999, w_099_6004, w_099_6007, w_099_6016, w_099_6024, w_099_6028, w_099_6030, w_099_6035, w_099_6037, w_099_6043, w_099_6045, w_099_6051, w_099_6052, w_099_6066, w_099_6067, w_099_6070, w_099_6081, w_099_6093, w_099_6094, w_099_6095, w_099_6099, w_099_6102, w_099_6105, w_099_6112, w_099_6113, w_099_6116, w_099_6117, w_099_6120, w_099_6130, w_099_6135, w_099_6136, w_099_6145, w_099_6147, w_099_6157, w_099_6159, w_099_6163, w_099_6164, w_099_6172, w_099_6173, w_099_6175, w_099_6181, w_099_6184, w_099_6189, w_099_6190, w_099_6194, w_099_6203, w_099_6209, w_099_6210, w_099_6217, w_099_6219, w_099_6220, w_099_6223, w_099_6224, w_099_6227, w_099_6229, w_099_6235, w_099_6246, w_099_6247, w_099_6256, w_099_6258, w_099_6259, w_099_6272, w_099_6273, w_099_6275, w_099_6276, w_099_6278, w_099_6286, w_099_6293, w_099_6298, w_099_6299, w_099_6300, w_099_6309, w_099_6312, w_099_6319, w_099_6333, w_099_6339, w_099_6343, w_099_6347, w_099_6354, w_099_6356, w_099_6365, w_099_6369, w_099_6370, w_099_6372, w_099_6377, w_099_6380, w_099_6383, w_099_6386, w_099_6408, w_099_6414, w_099_6419, w_099_6426, w_099_6430, w_099_6432, w_099_6440, w_099_6445, w_099_6446, w_099_6449, w_099_6469, w_099_6472, w_099_6473, w_099_6474, w_099_6481, w_099_6485, w_099_6486, w_099_6492, w_099_6495, w_099_6504, w_099_6512, w_099_6516, w_099_6520, w_099_6528, w_099_6531, w_099_6533, w_099_6540, w_099_6543, w_099_6547, w_099_6549, w_099_6551, w_099_6552, w_099_6558, w_099_6562, w_099_6567, w_099_6569, w_099_6574, w_099_6577, w_099_6578, w_099_6581, w_099_6584, w_099_6592, w_099_6593, w_099_6595, w_099_6596, w_099_6597, w_099_6600, w_099_6607, w_099_6611, w_099_6620, w_099_6626, w_099_6628, w_099_6629, w_099_6630, w_099_6636, w_099_6645, w_099_6651, w_099_6658, w_099_6662, w_099_6668, w_099_6672, w_099_6675, w_099_6679, w_099_6682, w_099_6686, w_099_6689, w_099_6690, w_099_6692, w_099_6694, w_099_6710, w_099_6712, w_099_6714, w_099_6719, w_099_6722, w_099_6724, w_099_6726, w_099_6733, w_099_6735, w_099_6738, w_099_6741, w_099_6745, w_099_6755, w_099_6757, w_099_6762, w_099_6773, w_099_6781, w_099_6784, w_099_6790, w_099_6801, w_099_6806, w_099_6811, w_099_6813, w_099_6814, w_099_6816, w_099_6817, w_099_6821, w_099_6831, w_099_6836, w_099_6837, w_099_6839, w_099_6844, w_099_6846, w_099_6848, w_099_6850, w_099_6859, w_099_6863, w_099_6867, w_099_6868, w_099_6876, w_099_6879, w_099_6881, w_099_6890, w_099_6896, w_099_6901, w_099_6905, w_099_6908, w_099_6909, w_099_6911, w_099_6914, w_099_6916, w_099_6920, w_099_6923, w_099_6926, w_099_6927, w_099_6931, w_099_6937, w_099_6938, w_099_6942, w_099_6944, w_099_6957, w_099_6961, w_099_6966, w_099_6969, w_099_6971, w_099_6972, w_099_6974, w_099_6976, w_099_6977, w_099_6978, w_099_6981, w_099_6984, w_099_6985, w_099_6998, w_099_7003, w_099_7008, w_099_7009, w_099_7013, w_099_7014, w_099_7018, w_099_7026, w_099_7037, w_099_7050, w_099_7056, w_099_7058, w_099_7064, w_099_7071, w_099_7074, w_099_7075, w_099_7076, w_099_7084, w_099_7091, w_099_7092, w_099_7107, w_099_7111, w_099_7115, w_099_7118, w_099_7120, w_099_7123, w_099_7129, w_099_7130, w_099_7142, w_099_7156, w_099_7164, w_099_7166, w_099_7175, w_099_7179, w_099_7189, w_099_7190, w_099_7201, w_099_7203, w_099_7204, w_099_7207, w_099_7209, w_099_7210, w_099_7211, w_099_7216, w_099_7231, w_099_7233, w_099_7237, w_099_7238, w_099_7242, w_099_7243, w_099_7247, w_099_7254, w_099_7256, w_099_7284, w_099_7294, w_099_7296, w_099_7298, w_099_7316, w_099_7322, w_099_7328, w_099_7330, w_099_7331, w_099_7333, w_099_7339, w_099_7340, w_099_7347, w_099_7348, w_099_7349, w_099_7350, w_099_7362, w_099_7369, w_099_7370, w_099_7374, w_099_7378, w_099_7382, w_099_7383, w_099_7386, w_099_7387, w_099_7388, w_099_7390, w_099_7395, w_099_7401, w_099_7421, w_099_7426, w_099_7429, w_099_7434, w_099_7435, w_099_7449, w_099_7450, w_099_7464, w_099_7467, w_099_7480, w_099_7482, w_099_7485, w_099_7486, w_099_7488, w_099_7492, w_099_7496, w_099_7506, w_099_7507, w_099_7514, w_099_7516, w_099_7523, w_099_7525, w_099_7527, w_099_7530, w_099_7535, w_099_7542, w_099_7551, w_099_7553, w_099_7560, w_099_7564, w_099_7565, w_099_7566, w_099_7572, w_099_7581, w_099_7582, w_099_7586, w_099_7588, w_099_7594, w_099_7595, w_099_7605, w_099_7607, w_099_7612, w_099_7617, w_099_7619, w_099_7628, w_099_7634, w_099_7638, w_099_7646, w_099_7647, w_099_7650, w_099_7662, w_099_7670, w_099_7671, w_099_7673, w_099_7684, w_099_7689, w_099_7699, w_099_7711, w_099_7712, w_099_7715, w_099_7720, w_099_7734, w_099_7737, w_099_7742, w_099_7751, w_099_7754, w_099_7764, w_099_7766, w_099_7768, w_099_7769, w_099_7777, w_099_7781, w_099_7786, w_099_7792, w_099_7798, w_099_7802, w_099_7805, w_099_7809, w_099_7815, w_099_7822, w_099_7833, w_099_7836, w_099_7837, w_099_7844, w_099_7847, w_099_7861, w_099_7868, w_099_7874, w_099_7878, w_099_7880, w_099_7900, w_099_7902, w_099_7904, w_099_7905, w_099_7906, w_099_7909, w_099_7928, w_099_7934, w_099_7937, w_099_7943, w_099_7950, w_099_7954, w_099_7960, w_099_7961, w_099_7966, w_099_7970, w_099_7984, w_099_7989, w_099_8005, w_099_8012, w_099_8013, w_099_8014, w_099_8020, w_099_8021, w_099_8040, w_099_8042, w_099_8043, w_099_8048, w_099_8051, w_099_8054, w_099_8056, w_099_8066, w_099_8068, w_099_8079, w_099_8085, w_099_8092, w_099_8097, w_099_8103, w_099_8105, w_099_8108, w_099_8109, w_099_8110, w_099_8111, w_099_8114, w_099_8119, w_099_8120, w_099_8122, w_099_8123, w_099_8125, w_099_8127, w_099_8142, w_099_8143, w_099_8155;
  wire w_100_005, w_100_007, w_100_009, w_100_012, w_100_015, w_100_021, w_100_022, w_100_025, w_100_039, w_100_040, w_100_047, w_100_048, w_100_054, w_100_055, w_100_056, w_100_057, w_100_060, w_100_064, w_100_070, w_100_072, w_100_076, w_100_077, w_100_080, w_100_081, w_100_086, w_100_087, w_100_090, w_100_093, w_100_094, w_100_096, w_100_098, w_100_099, w_100_100, w_100_103, w_100_109, w_100_112, w_100_113, w_100_114, w_100_117, w_100_120, w_100_123, w_100_124, w_100_128, w_100_130, w_100_132, w_100_134, w_100_136, w_100_137, w_100_139, w_100_140, w_100_141, w_100_146, w_100_149, w_100_151, w_100_152, w_100_155, w_100_159, w_100_160, w_100_163, w_100_169, w_100_174, w_100_176, w_100_178, w_100_180, w_100_182, w_100_186, w_100_187, w_100_193, w_100_203, w_100_208, w_100_212, w_100_218, w_100_220, w_100_222, w_100_223, w_100_226, w_100_232, w_100_234, w_100_236, w_100_237, w_100_247, w_100_250, w_100_251, w_100_254, w_100_255, w_100_256, w_100_257, w_100_260, w_100_262, w_100_263, w_100_265, w_100_267, w_100_273, w_100_274, w_100_278, w_100_280, w_100_282, w_100_291, w_100_292, w_100_296, w_100_297, w_100_299, w_100_300, w_100_305, w_100_307, w_100_317, w_100_318, w_100_319, w_100_323, w_100_327, w_100_328, w_100_331, w_100_332, w_100_335, w_100_337, w_100_338, w_100_342, w_100_346, w_100_350, w_100_351, w_100_353, w_100_354, w_100_355, w_100_357, w_100_358, w_100_359, w_100_360, w_100_361, w_100_369, w_100_371, w_100_374, w_100_375, w_100_380, w_100_385, w_100_395, w_100_397, w_100_401, w_100_405, w_100_407, w_100_411, w_100_412, w_100_414, w_100_416, w_100_417, w_100_418, w_100_419, w_100_420, w_100_427, w_100_431, w_100_433, w_100_437, w_100_438, w_100_443, w_100_447, w_100_449, w_100_452, w_100_455, w_100_456, w_100_458, w_100_460, w_100_462, w_100_466, w_100_469, w_100_470, w_100_473, w_100_477, w_100_479, w_100_480, w_100_482, w_100_489, w_100_491, w_100_494, w_100_495, w_100_496, w_100_497, w_100_498, w_100_500, w_100_503, w_100_504, w_100_506, w_100_508, w_100_513, w_100_517, w_100_518, w_100_519, w_100_520, w_100_522, w_100_525, w_100_529, w_100_530, w_100_532, w_100_546, w_100_551, w_100_554, w_100_557, w_100_561, w_100_563, w_100_565, w_100_567, w_100_568, w_100_571, w_100_572, w_100_574, w_100_580, w_100_583, w_100_584, w_100_585, w_100_586, w_100_593, w_100_602, w_100_604, w_100_610, w_100_611, w_100_613, w_100_615, w_100_616, w_100_618, w_100_621, w_100_623, w_100_624, w_100_625, w_100_631, w_100_634, w_100_635, w_100_639, w_100_642, w_100_644, w_100_647, w_100_650, w_100_651, w_100_652, w_100_653, w_100_654, w_100_656, w_100_657, w_100_659, w_100_662, w_100_664, w_100_665, w_100_666, w_100_667, w_100_668, w_100_670, w_100_673, w_100_676, w_100_677, w_100_678, w_100_681, w_100_684, w_100_686, w_100_689, w_100_690, w_100_691, w_100_695, w_100_697, w_100_700, w_100_705, w_100_708, w_100_715, w_100_719, w_100_721, w_100_726, w_100_727, w_100_728, w_100_730, w_100_731, w_100_732, w_100_734, w_100_736, w_100_737, w_100_741, w_100_743, w_100_745, w_100_748, w_100_749, w_100_752, w_100_753, w_100_755, w_100_758, w_100_761, w_100_767, w_100_769, w_100_770, w_100_771, w_100_773, w_100_775, w_100_776, w_100_781, w_100_782, w_100_784, w_100_787, w_100_788, w_100_789, w_100_790, w_100_791, w_100_793, w_100_795, w_100_798, w_100_804, w_100_808, w_100_816, w_100_817, w_100_820, w_100_821, w_100_823, w_100_828, w_100_834, w_100_835, w_100_838, w_100_840, w_100_841, w_100_842, w_100_843, w_100_844, w_100_845, w_100_846, w_100_847, w_100_848, w_100_851, w_100_853, w_100_855, w_100_856, w_100_857, w_100_858, w_100_860, w_100_862, w_100_868, w_100_869, w_100_871, w_100_875, w_100_876, w_100_877, w_100_882, w_100_883, w_100_886, w_100_887, w_100_888, w_100_890, w_100_892, w_100_893, w_100_894, w_100_899, w_100_902, w_100_903, w_100_906, w_100_909, w_100_910, w_100_911, w_100_916, w_100_917, w_100_921, w_100_925, w_100_930, w_100_934, w_100_935, w_100_937, w_100_938, w_100_941, w_100_942, w_100_943, w_100_945, w_100_946, w_100_950, w_100_954, w_100_955, w_100_957, w_100_961, w_100_964, w_100_965, w_100_966, w_100_968, w_100_969, w_100_976, w_100_977, w_100_978, w_100_979, w_100_980, w_100_983, w_100_985, w_100_986, w_100_988, w_100_989, w_100_991, w_100_996, w_100_1001, w_100_1005, w_100_1008, w_100_1009, w_100_1010, w_100_1011, w_100_1012, w_100_1013, w_100_1015, w_100_1016, w_100_1017, w_100_1018, w_100_1020, w_100_1024, w_100_1025, w_100_1026, w_100_1032, w_100_1036, w_100_1039, w_100_1041, w_100_1042, w_100_1044, w_100_1049, w_100_1053, w_100_1054, w_100_1056, w_100_1057, w_100_1058, w_100_1060, w_100_1061, w_100_1069, w_100_1070, w_100_1075, w_100_1077, w_100_1078, w_100_1080, w_100_1081, w_100_1082, w_100_1085, w_100_1088, w_100_1089, w_100_1091, w_100_1092, w_100_1093, w_100_1095, w_100_1096, w_100_1101, w_100_1102, w_100_1110, w_100_1120, w_100_1129, w_100_1131, w_100_1134, w_100_1140, w_100_1145, w_100_1146, w_100_1156, w_100_1159, w_100_1161, w_100_1165, w_100_1174, w_100_1175, w_100_1183, w_100_1191, w_100_1196, w_100_1201, w_100_1221, w_100_1223, w_100_1225, w_100_1232, w_100_1233, w_100_1234, w_100_1240, w_100_1244, w_100_1247, w_100_1253, w_100_1262, w_100_1265, w_100_1266, w_100_1268, w_100_1274, w_100_1278, w_100_1286, w_100_1293, w_100_1306, w_100_1310, w_100_1313, w_100_1315, w_100_1316, w_100_1319, w_100_1322, w_100_1338, w_100_1343, w_100_1349, w_100_1354, w_100_1358, w_100_1360, w_100_1364, w_100_1365, w_100_1366, w_100_1370, w_100_1371, w_100_1375, w_100_1376, w_100_1377, w_100_1380, w_100_1382, w_100_1384, w_100_1389, w_100_1391, w_100_1394, w_100_1403, w_100_1404, w_100_1406, w_100_1411, w_100_1414, w_100_1419, w_100_1421, w_100_1422, w_100_1424, w_100_1427, w_100_1428, w_100_1433, w_100_1435, w_100_1438, w_100_1441, w_100_1448, w_100_1452, w_100_1457, w_100_1458, w_100_1464, w_100_1465, w_100_1467, w_100_1473, w_100_1477, w_100_1480, w_100_1482, w_100_1485, w_100_1486, w_100_1490, w_100_1496, w_100_1498, w_100_1507, w_100_1510, w_100_1518, w_100_1519, w_100_1532, w_100_1536, w_100_1537, w_100_1541, w_100_1542, w_100_1551, w_100_1566, w_100_1567, w_100_1572, w_100_1577, w_100_1581, w_100_1586, w_100_1587, w_100_1590, w_100_1591, w_100_1593, w_100_1599, w_100_1606, w_100_1607, w_100_1611, w_100_1612, w_100_1613, w_100_1620, w_100_1622, w_100_1628, w_100_1631, w_100_1634, w_100_1642, w_100_1643, w_100_1644, w_100_1647, w_100_1652, w_100_1656, w_100_1673, w_100_1677, w_100_1690, w_100_1692, w_100_1697, w_100_1703, w_100_1709, w_100_1711, w_100_1719, w_100_1720, w_100_1725, w_100_1732, w_100_1737, w_100_1740, w_100_1741, w_100_1742, w_100_1744, w_100_1748, w_100_1749, w_100_1751, w_100_1755, w_100_1756, w_100_1758, w_100_1766, w_100_1768, w_100_1777, w_100_1778, w_100_1781, w_100_1792, w_100_1793, w_100_1795, w_100_1801, w_100_1808, w_100_1816, w_100_1818, w_100_1820, w_100_1821, w_100_1829, w_100_1831, w_100_1832, w_100_1837, w_100_1838, w_100_1841, w_100_1845, w_100_1848, w_100_1853, w_100_1855, w_100_1858, w_100_1865, w_100_1867, w_100_1888, w_100_1889, w_100_1892, w_100_1896, w_100_1897, w_100_1900, w_100_1901, w_100_1913, w_100_1925, w_100_1926, w_100_1931, w_100_1935, w_100_1936, w_100_1939, w_100_1943, w_100_1945, w_100_1947, w_100_1950, w_100_1955, w_100_1967, w_100_1976, w_100_1979, w_100_1980, w_100_1986, w_100_1987, w_100_1996, w_100_1997, w_100_1999, w_100_2008, w_100_2009, w_100_2012, w_100_2016, w_100_2026, w_100_2028, w_100_2029, w_100_2036, w_100_2041, w_100_2051, w_100_2060, w_100_2066, w_100_2076, w_100_2078, w_100_2085, w_100_2090, w_100_2101, w_100_2113, w_100_2117, w_100_2119, w_100_2126, w_100_2130, w_100_2133, w_100_2138, w_100_2140, w_100_2146, w_100_2147, w_100_2148, w_100_2153, w_100_2164, w_100_2167, w_100_2169, w_100_2171, w_100_2172, w_100_2173, w_100_2176, w_100_2178, w_100_2181, w_100_2191, w_100_2192, w_100_2193, w_100_2203, w_100_2206, w_100_2207, w_100_2210, w_100_2214, w_100_2215, w_100_2217, w_100_2220, w_100_2226, w_100_2235, w_100_2238, w_100_2243, w_100_2249, w_100_2252, w_100_2253, w_100_2260, w_100_2263, w_100_2265, w_100_2267, w_100_2273, w_100_2277, w_100_2278, w_100_2289, w_100_2290, w_100_2293, w_100_2295, w_100_2296, w_100_2300, w_100_2303, w_100_2304, w_100_2310, w_100_2314, w_100_2320, w_100_2326, w_100_2338, w_100_2342, w_100_2343, w_100_2347, w_100_2349, w_100_2350, w_100_2363, w_100_2365, w_100_2366, w_100_2372, w_100_2375, w_100_2380, w_100_2381, w_100_2390, w_100_2400, w_100_2402, w_100_2403, w_100_2417, w_100_2424, w_100_2428, w_100_2429, w_100_2431, w_100_2432, w_100_2435, w_100_2437, w_100_2445, w_100_2451, w_100_2453, w_100_2454, w_100_2455, w_100_2456, w_100_2469, w_100_2472, w_100_2475, w_100_2478, w_100_2479, w_100_2486, w_100_2487, w_100_2491, w_100_2493, w_100_2500, w_100_2502, w_100_2505, w_100_2509, w_100_2513, w_100_2522, w_100_2529, w_100_2538, w_100_2540, w_100_2542, w_100_2544, w_100_2550, w_100_2566, w_100_2571, w_100_2574, w_100_2575, w_100_2577, w_100_2595, w_100_2598, w_100_2599, w_100_2601, w_100_2603, w_100_2607, w_100_2612, w_100_2615, w_100_2619, w_100_2622, w_100_2623, w_100_2627, w_100_2629, w_100_2631, w_100_2635, w_100_2636, w_100_2643, w_100_2644, w_100_2648, w_100_2654, w_100_2655, w_100_2659, w_100_2662, w_100_2665, w_100_2670, w_100_2671, w_100_2672, w_100_2692, w_100_2704, w_100_2710, w_100_2730, w_100_2732, w_100_2740, w_100_2755, w_100_2756, w_100_2762, w_100_2763, w_100_2764, w_100_2765, w_100_2767, w_100_2770, w_100_2773, w_100_2774, w_100_2775, w_100_2778, w_100_2785, w_100_2808, w_100_2823, w_100_2825, w_100_2831, w_100_2833, w_100_2843, w_100_2845, w_100_2847, w_100_2848, w_100_2849, w_100_2857, w_100_2859, w_100_2861, w_100_2868, w_100_2870, w_100_2872, w_100_2876, w_100_2877, w_100_2878, w_100_2888, w_100_2900, w_100_2905, w_100_2908, w_100_2913, w_100_2915, w_100_2923, w_100_2932, w_100_2935, w_100_2941, w_100_2950, w_100_2953, w_100_2956, w_100_2962, w_100_2967, w_100_2970, w_100_2975, w_100_2980, w_100_2986, w_100_2988, w_100_2997, w_100_3002, w_100_3005, w_100_3011, w_100_3018, w_100_3023, w_100_3026, w_100_3027, w_100_3028, w_100_3033, w_100_3034, w_100_3037, w_100_3038, w_100_3047, w_100_3050, w_100_3051, w_100_3082, w_100_3092, w_100_3094, w_100_3099, w_100_3107, w_100_3112, w_100_3113, w_100_3116, w_100_3123, w_100_3131, w_100_3137, w_100_3144, w_100_3147, w_100_3150, w_100_3158, w_100_3165, w_100_3166, w_100_3174, w_100_3179, w_100_3185, w_100_3186, w_100_3187, w_100_3188, w_100_3196, w_100_3204, w_100_3206, w_100_3212, w_100_3218, w_100_3219, w_100_3227, w_100_3228, w_100_3233, w_100_3237, w_100_3241, w_100_3242, w_100_3253, w_100_3255, w_100_3258, w_100_3259, w_100_3260, w_100_3264, w_100_3270, w_100_3271, w_100_3273, w_100_3277, w_100_3282, w_100_3286, w_100_3287, w_100_3295, w_100_3301, w_100_3302, w_100_3303, w_100_3319, w_100_3320, w_100_3323, w_100_3327, w_100_3332, w_100_3335, w_100_3337, w_100_3342, w_100_3349, w_100_3350, w_100_3352, w_100_3353, w_100_3354, w_100_3360, w_100_3370, w_100_3379, w_100_3391, w_100_3398, w_100_3400, w_100_3401, w_100_3406, w_100_3413, w_100_3414, w_100_3415, w_100_3418, w_100_3422, w_100_3434, w_100_3455, w_100_3457, w_100_3464, w_100_3466, w_100_3473, w_100_3474, w_100_3479, w_100_3484, w_100_3490, w_100_3492, w_100_3507, w_100_3523, w_100_3531, w_100_3534, w_100_3535, w_100_3542, w_100_3545, w_100_3549, w_100_3559, w_100_3562, w_100_3563, w_100_3566, w_100_3569, w_100_3571, w_100_3578, w_100_3581, w_100_3599, w_100_3601, w_100_3602, w_100_3604, w_100_3611, w_100_3616, w_100_3627, w_100_3631, w_100_3633, w_100_3639, w_100_3641, w_100_3645, w_100_3648, w_100_3650, w_100_3653, w_100_3655, w_100_3657, w_100_3658, w_100_3670, w_100_3673, w_100_3675, w_100_3676, w_100_3677, w_100_3679, w_100_3686, w_100_3694, w_100_3699, w_100_3712, w_100_3717, w_100_3721, w_100_3724, w_100_3730, w_100_3733, w_100_3741, w_100_3744, w_100_3757, w_100_3760, w_100_3770, w_100_3772, w_100_3781, w_100_3795, w_100_3797, w_100_3804, w_100_3807, w_100_3810, w_100_3813, w_100_3816, w_100_3819, w_100_3821, w_100_3823, w_100_3824, w_100_3826, w_100_3832, w_100_3834, w_100_3839, w_100_3844, w_100_3847, w_100_3854, w_100_3862, w_100_3863, w_100_3872, w_100_3876, w_100_3885, w_100_3889, w_100_3895, w_100_3901, w_100_3903, w_100_3906, w_100_3926, w_100_3928, w_100_3939, w_100_3948, w_100_3954, w_100_3958, w_100_3961, w_100_3963, w_100_3966, w_100_3971, w_100_3974, w_100_3977, w_100_3978, w_100_3994, w_100_3997, w_100_3999, w_100_4000, w_100_4016, w_100_4018, w_100_4021, w_100_4030, w_100_4031, w_100_4032, w_100_4036, w_100_4041, w_100_4044, w_100_4045, w_100_4048, w_100_4050, w_100_4051, w_100_4053, w_100_4054, w_100_4056, w_100_4057, w_100_4067, w_100_4073, w_100_4074, w_100_4086, w_100_4089, w_100_4091, w_100_4093, w_100_4094, w_100_4096, w_100_4099, w_100_4120, w_100_4121, w_100_4126, w_100_4127, w_100_4128, w_100_4132, w_100_4133, w_100_4134, w_100_4144, w_100_4146, w_100_4159, w_100_4160, w_100_4161, w_100_4162, w_100_4163, w_100_4169, w_100_4170, w_100_4175, w_100_4180, w_100_4181, w_100_4183, w_100_4186, w_100_4192, w_100_4196, w_100_4199, w_100_4204, w_100_4215, w_100_4216, w_100_4220, w_100_4221, w_100_4223, w_100_4226, w_100_4231, w_100_4234, w_100_4243, w_100_4247, w_100_4248, w_100_4262, w_100_4263, w_100_4270, w_100_4278, w_100_4288, w_100_4319, w_100_4320, w_100_4326, w_100_4328, w_100_4340, w_100_4343, w_100_4347, w_100_4356, w_100_4369, w_100_4371, w_100_4374, w_100_4376, w_100_4377, w_100_4391, w_100_4397, w_100_4400, w_100_4403, w_100_4425, w_100_4428, w_100_4440, w_100_4441, w_100_4450, w_100_4451, w_100_4452, w_100_4464, w_100_4466, w_100_4467, w_100_4472, w_100_4479, w_100_4486, w_100_4491, w_100_4494, w_100_4501, w_100_4508, w_100_4512, w_100_4513, w_100_4521, w_100_4537, w_100_4545, w_100_4550, w_100_4556, w_100_4557, w_100_4560, w_100_4562, w_100_4573, w_100_4574, w_100_4575, w_100_4576, w_100_4581, w_100_4584, w_100_4586, w_100_4587, w_100_4590, w_100_4612, w_100_4620, w_100_4621, w_100_4622, w_100_4623, w_100_4625, w_100_4634, w_100_4636, w_100_4640, w_100_4641, w_100_4646, w_100_4650, w_100_4658, w_100_4661, w_100_4666, w_100_4667, w_100_4668, w_100_4673, w_100_4675, w_100_4678, w_100_4688, w_100_4690, w_100_4695, w_100_4703, w_100_4704, w_100_4709, w_100_4711, w_100_4718, w_100_4719, w_100_4720, w_100_4725, w_100_4726, w_100_4732, w_100_4751, w_100_4753, w_100_4757, w_100_4759, w_100_4760, w_100_4772, w_100_4773, w_100_4775, w_100_4777, w_100_4780, w_100_4792, w_100_4793, w_100_4800, w_100_4803, w_100_4804, w_100_4806, w_100_4807, w_100_4815, w_100_4817, w_100_4823, w_100_4830, w_100_4832, w_100_4838, w_100_4839, w_100_4846, w_100_4850, w_100_4853, w_100_4862, w_100_4865, w_100_4871, w_100_4874, w_100_4881, w_100_4885, w_100_4890, w_100_4894, w_100_4899, w_100_4905, w_100_4911, w_100_4913, w_100_4915, w_100_4924, w_100_4927, w_100_4938, w_100_4940, w_100_4942, w_100_4949, w_100_4958, w_100_4959, w_100_4961, w_100_4963, w_100_4964, w_100_4968, w_100_4969, w_100_4972, w_100_4973, w_100_4974, w_100_4990, w_100_4993, w_100_4996, w_100_4997, w_100_4998, w_100_5000, w_100_5008, w_100_5012, w_100_5017, w_100_5024, w_100_5028, w_100_5037, w_100_5043, w_100_5048, w_100_5051, w_100_5054, w_100_5064, w_100_5067, w_100_5086, w_100_5088, w_100_5090, w_100_5096, w_100_5106, w_100_5110, w_100_5112, w_100_5117, w_100_5118, w_100_5123, w_100_5127, w_100_5129, w_100_5146, w_100_5150, w_100_5152, w_100_5155, w_100_5157, w_100_5160, w_100_5162, w_100_5165, w_100_5166, w_100_5168, w_100_5169, w_100_5170, w_100_5173, w_100_5183, w_100_5184, w_100_5192, w_100_5193, w_100_5200, w_100_5207, w_100_5210, w_100_5220, w_100_5222, w_100_5227, w_100_5229, w_100_5239, w_100_5242, w_100_5247, w_100_5248, w_100_5253, w_100_5257, w_100_5258, w_100_5259, w_100_5266, w_100_5271, w_100_5272, w_100_5276, w_100_5285, w_100_5304, w_100_5305, w_100_5306, w_100_5308, w_100_5313, w_100_5316, w_100_5317, w_100_5322, w_100_5323, w_100_5327, w_100_5333, w_100_5339, w_100_5341, w_100_5352, w_100_5359, w_100_5360, w_100_5361, w_100_5367, w_100_5368, w_100_5372, w_100_5373, w_100_5377, w_100_5381, w_100_5394, w_100_5401, w_100_5403, w_100_5404, w_100_5406, w_100_5407, w_100_5412, w_100_5418, w_100_5419, w_100_5422, w_100_5423, w_100_5424, w_100_5428, w_100_5430, w_100_5437, w_100_5440, w_100_5441, w_100_5442, w_100_5450, w_100_5456, w_100_5464, w_100_5475, w_100_5477, w_100_5478, w_100_5481, w_100_5482, w_100_5484, w_100_5485, w_100_5486, w_100_5487, w_100_5488, w_100_5492, w_100_5493, w_100_5508, w_100_5510, w_100_5513, w_100_5515, w_100_5524, w_100_5536, w_100_5542, w_100_5548, w_100_5553, w_100_5559, w_100_5572, w_100_5573, w_100_5585, w_100_5594, w_100_5602, w_100_5608, w_100_5609, w_100_5618, w_100_5619, w_100_5622, w_100_5626, w_100_5631, w_100_5632, w_100_5633, w_100_5640, w_100_5652, w_100_5653, w_100_5654, w_100_5658, w_100_5660, w_100_5662, w_100_5666, w_100_5667, w_100_5673, w_100_5674, w_100_5688, w_100_5689, w_100_5692, w_100_5693, w_100_5695, w_100_5699, w_100_5701, w_100_5708, w_100_5721, w_100_5732, w_100_5743, w_100_5755, w_100_5758, w_100_5763, w_100_5764, w_100_5766, w_100_5767, w_100_5775, w_100_5777, w_100_5779, w_100_5793, w_100_5796, w_100_5800, w_100_5801, w_100_5804, w_100_5811, w_100_5815, w_100_5820, w_100_5824, w_100_5825, w_100_5827, w_100_5830, w_100_5846, w_100_5850, w_100_5853, w_100_5857, w_100_5859, w_100_5861, w_100_5862, w_100_5869, w_100_5871, w_100_5873, w_100_5876, w_100_5886, w_100_5891, w_100_5895, w_100_5902, w_100_5911, w_100_5912, w_100_5915, w_100_5916, w_100_5930, w_100_5931, w_100_5942, w_100_5944, w_100_5946, w_100_5950, w_100_5955, w_100_5961, w_100_5975, w_100_5976, w_100_5979, w_100_5981, w_100_5982, w_100_5985, w_100_5987, w_100_5993, w_100_5994, w_100_5996, w_100_5997, w_100_6005, w_100_6007, w_100_6009, w_100_6012, w_100_6017, w_100_6019, w_100_6021, w_100_6024, w_100_6026, w_100_6027, w_100_6038, w_100_6039, w_100_6045, w_100_6055, w_100_6059, w_100_6060, w_100_6061, w_100_6064, w_100_6065, w_100_6068, w_100_6070, w_100_6078, w_100_6084, w_100_6086, w_100_6087, w_100_6089, w_100_6091, w_100_6096, w_100_6100, w_100_6102, w_100_6111, w_100_6114, w_100_6122, w_100_6125, w_100_6129, w_100_6138, w_100_6140, w_100_6144, w_100_6154, w_100_6158, w_100_6166, w_100_6168, w_100_6176, w_100_6177, w_100_6179, w_100_6182, w_100_6184, w_100_6189, w_100_6191, w_100_6192, w_100_6204, w_100_6211, w_100_6212, w_100_6213, w_100_6219, w_100_6221, w_100_6222, w_100_6226, w_100_6229, w_100_6245, w_100_6251, w_100_6253, w_100_6256, w_100_6261, w_100_6265, w_100_6267, w_100_6270, w_100_6271, w_100_6272, w_100_6283, w_100_6284, w_100_6285, w_100_6287, w_100_6296, w_100_6299, w_100_6305, w_100_6306, w_100_6309, w_100_6317, w_100_6319, w_100_6324, w_100_6328, w_100_6329, w_100_6331, w_100_6335, w_100_6342, w_100_6350, w_100_6359, w_100_6360, w_100_6368, w_100_6382, w_100_6395, w_100_6398, w_100_6400, w_100_6402, w_100_6414, w_100_6415, w_100_6416, w_100_6431, w_100_6434, w_100_6439, w_100_6449, w_100_6450, w_100_6451, w_100_6453, w_100_6454, w_100_6462, w_100_6467, w_100_6469, w_100_6470, w_100_6472, w_100_6481, w_100_6486, w_100_6490, w_100_6505, w_100_6507, w_100_6509, w_100_6510, w_100_6515, w_100_6519, w_100_6529, w_100_6535, w_100_6547, w_100_6551, w_100_6553, w_100_6554, w_100_6557, w_100_6559, w_100_6563, w_100_6570, w_100_6572, w_100_6587, w_100_6595, w_100_6598, w_100_6600, w_100_6604, w_100_6606, w_100_6609, w_100_6610, w_100_6613, w_100_6614, w_100_6617, w_100_6618, w_100_6622, w_100_6626, w_100_6628, w_100_6636, w_100_6640, w_100_6644, w_100_6651, w_100_6655, w_100_6662, w_100_6668, w_100_6669, w_100_6670, w_100_6672, w_100_6679, w_100_6681, w_100_6690, w_100_6693, w_100_6698, w_100_6703, w_100_6718, w_100_6719, w_100_6726, w_100_6730, w_100_6732, w_100_6737, w_100_6739, w_100_6754, w_100_6755, w_100_6763, w_100_6767, w_100_6770, w_100_6773, w_100_6775, w_100_6780, w_100_6783, w_100_6785, w_100_6787, w_100_6790, w_100_6791, w_100_6794, w_100_6795, w_100_6806, w_100_6808, w_100_6813, w_100_6821, w_100_6823, w_100_6828, w_100_6833, w_100_6838, w_100_6853, w_100_6869, w_100_6880, w_100_6882, w_100_6893, w_100_6897, w_100_6900, w_100_6920, w_100_6929, w_100_6931, w_100_6936, w_100_6940, w_100_6946, w_100_6952, w_100_6958, w_100_6971, w_100_6974, w_100_6978, w_100_6979, w_100_6984, w_100_6991, w_100_6993, w_100_6995, w_100_6999, w_100_7011, w_100_7013, w_100_7025, w_100_7028, w_100_7029, w_100_7031, w_100_7033, w_100_7034, w_100_7041, w_100_7046, w_100_7047, w_100_7050, w_100_7061, w_100_7064, w_100_7066, w_100_7073, w_100_7082, w_100_7104, w_100_7105, w_100_7106, w_100_7108, w_100_7109, w_100_7123, w_100_7125, w_100_7129, w_100_7135, w_100_7140, w_100_7149, w_100_7152, w_100_7155, w_100_7156, w_100_7157, w_100_7160, w_100_7166, w_100_7169, w_100_7174, w_100_7181, w_100_7184, w_100_7186, w_100_7187, w_100_7191, w_100_7196, w_100_7207, w_100_7208, w_100_7214, w_100_7218, w_100_7233, w_100_7240, w_100_7253, w_100_7255, w_100_7258, w_100_7259, w_100_7261, w_100_7265, w_100_7267, w_100_7272, w_100_7278, w_100_7280, w_100_7283, w_100_7296, w_100_7299, w_100_7301, w_100_7304, w_100_7305, w_100_7321, w_100_7326, w_100_7328, w_100_7336, w_100_7348, w_100_7361, w_100_7366, w_100_7373, w_100_7375, w_100_7383, w_100_7391, w_100_7393, w_100_7395, w_100_7402, w_100_7407, w_100_7413, w_100_7415, w_100_7416, w_100_7418, w_100_7420, w_100_7421, w_100_7423, w_100_7425, w_100_7449, w_100_7472, w_100_7484, w_100_7485, w_100_7486, w_100_7496, w_100_7501, w_100_7511, w_100_7533, w_100_7535, w_100_7536, w_100_7546, w_100_7547, w_100_7548, w_100_7552, w_100_7555, w_100_7559, w_100_7564, w_100_7566, w_100_7573, w_100_7574, w_100_7576, w_100_7582, w_100_7583, w_100_7586, w_100_7589, w_100_7593, w_100_7605, w_100_7606, w_100_7608, w_100_7609, w_100_7613, w_100_7623, w_100_7629, w_100_7632, w_100_7633, w_100_7638, w_100_7643, w_100_7648, w_100_7650, w_100_7658, w_100_7667, w_100_7680, w_100_7682, w_100_7684, w_100_7687, w_100_7688, w_100_7689, w_100_7696, w_100_7701, w_100_7704, w_100_7705, w_100_7709, w_100_7712, w_100_7716, w_100_7718, w_100_7720, w_100_7726, w_100_7727, w_100_7730, w_100_7733, w_100_7734, w_100_7748, w_100_7749, w_100_7752, w_100_7762, w_100_7767, w_100_7772, w_100_7773, w_100_7775, w_100_7788, w_100_7792, w_100_7797, w_100_7802, w_100_7803, w_100_7804, w_100_7812, w_100_7815, w_100_7817, w_100_7821, w_100_7831, w_100_7841, w_100_7848, w_100_7854, w_100_7865, w_100_7867, w_100_7868, w_100_7870, w_100_7887, w_100_7897, w_100_7902, w_100_7904, w_100_7907, w_100_7910, w_100_7911, w_100_7916, w_100_7922, w_100_7928, w_100_7929, w_100_7935, w_100_7936, w_100_7937, w_100_7942, w_100_7945, w_100_7947, w_100_7949, w_100_7954, w_100_7957, w_100_7959, w_100_7961, w_100_7965, w_100_7968, w_100_7973, w_100_7977, w_100_7980, w_100_7982, w_100_7983, w_100_7985, w_100_7986, w_100_7992, w_100_8007, w_100_8043, w_100_8046, w_100_8047, w_100_8053, w_100_8058, w_100_8059, w_100_8060, w_100_8061, w_100_8068, w_100_8082, w_100_8089, w_100_8097, w_100_8106, w_100_8112, w_100_8117, w_100_8126, w_100_8134, w_100_8136, w_100_8137, w_100_8138, w_100_8163, w_100_8176, w_100_8178, w_100_8179, w_100_8189, w_100_8190, w_100_8195, w_100_8198, w_100_8201, w_100_8216, w_100_8235, w_100_8238, w_100_8244, w_100_8257, w_100_8262, w_100_8263, w_100_8266, w_100_8274, w_100_8275, w_100_8278, w_100_8283, w_100_8284, w_100_8298, w_100_8302, w_100_8309, w_100_8314, w_100_8321, w_100_8322, w_100_8323, w_100_8325, w_100_8331, w_100_8352, w_100_8356, w_100_8363, w_100_8365, w_100_8371, w_100_8373, w_100_8377, w_100_8378, w_100_8380, w_100_8386, w_100_8393, w_100_8397, w_100_8404, w_100_8407, w_100_8413, w_100_8419, w_100_8426, w_100_8430, w_100_8435, w_100_8447, w_100_8455, w_100_8459, w_100_8474, w_100_8483, w_100_8496, w_100_8500, w_100_8502, w_100_8516, w_100_8529, w_100_8534, w_100_8536, w_100_8549, w_100_8552, w_100_8558, w_100_8560, w_100_8562, w_100_8566, w_100_8569, w_100_8570, w_100_8572, w_100_8585, w_100_8586, w_100_8590, w_100_8592, w_100_8596, w_100_8599, w_100_8603, w_100_8606, w_100_8609, w_100_8612, w_100_8613, w_100_8620, w_100_8626, w_100_8627, w_100_8637, w_100_8642, w_100_8643, w_100_8644, w_100_8645, w_100_8646, w_100_8652, w_100_8654, w_100_8676, w_100_8681, w_100_8689, w_100_8705, w_100_8706, w_100_8716, w_100_8720, w_100_8729, w_100_8733, w_100_8746, w_100_8752, w_100_8754, w_100_8768, w_100_8769, w_100_8770, w_100_8773, w_100_8774, w_100_8776, w_100_8777, w_100_8780, w_100_8794, w_100_8795, w_100_8796, w_100_8800, w_100_8808, w_100_8816, w_100_8819, w_100_8822, w_100_8825, w_100_8832, w_100_8838, w_100_8840, w_100_8844, w_100_8853, w_100_8863, w_100_8866, w_100_8869, w_100_8870, w_100_8872, w_100_8873, w_100_8881;
  wire w_101_000, w_101_002, w_101_004, w_101_005, w_101_006, w_101_007, w_101_010, w_101_012, w_101_014, w_101_016, w_101_017, w_101_018, w_101_021, w_101_022, w_101_023, w_101_024, w_101_027, w_101_029, w_101_030, w_101_031, w_101_035, w_101_036, w_101_038, w_101_039, w_101_040, w_101_041, w_101_042, w_101_044, w_101_046, w_101_050, w_101_051, w_101_052, w_101_053, w_101_054, w_101_057, w_101_058, w_101_060, w_101_061, w_101_062, w_101_063, w_101_065, w_101_066, w_101_068, w_101_073, w_101_074, w_101_076, w_101_078, w_101_079, w_101_082, w_101_084, w_101_086, w_101_089, w_101_091, w_101_092, w_101_093, w_101_094, w_101_095, w_101_102, w_101_103, w_101_105, w_101_107, w_101_109, w_101_111, w_101_117, w_101_119, w_101_123, w_101_125, w_101_127, w_101_128, w_101_129, w_101_133, w_101_135, w_101_136, w_101_137, w_101_139, w_101_140, w_101_142, w_101_144, w_101_146, w_101_147, w_101_148, w_101_150, w_101_152, w_101_159, w_101_163, w_101_164, w_101_165, w_101_167, w_101_168, w_101_169, w_101_171, w_101_172, w_101_173, w_101_175, w_101_176, w_101_178, w_101_180, w_101_182, w_101_183, w_101_184, w_101_186, w_101_187, w_101_188, w_101_191, w_101_192, w_101_196, w_101_197, w_101_198, w_101_199, w_101_203, w_101_205, w_101_206, w_101_207, w_101_208, w_101_209, w_101_210, w_101_211, w_101_213, w_101_214, w_101_215, w_101_219, w_101_220, w_101_221, w_101_222, w_101_227, w_101_231, w_101_233, w_101_234, w_101_235, w_101_236, w_101_238, w_101_240, w_101_246, w_101_251, w_101_252, w_101_253, w_101_254, w_101_264, w_101_268, w_101_269, w_101_270, w_101_271, w_101_272, w_101_273, w_101_276, w_101_277, w_101_286, w_101_287, w_101_289, w_101_292, w_101_296, w_101_298, w_101_299, w_101_301, w_101_302, w_101_304, w_101_306, w_101_307, w_101_308, w_101_309, w_101_310, w_101_312, w_101_315, w_101_317, w_101_319, w_101_320, w_101_321, w_101_322, w_101_323, w_101_328, w_101_329, w_101_330, w_101_333, w_101_334, w_101_335, w_101_338, w_101_340, w_101_346, w_101_348, w_101_351, w_101_352, w_101_353, w_101_354, w_101_355, w_101_356, w_101_358, w_101_360, w_101_361, w_101_362, w_101_364, w_101_366, w_101_368, w_101_369, w_101_371, w_101_375, w_101_376, w_101_378, w_101_382, w_101_383, w_101_386, w_101_392, w_101_396, w_101_398, w_101_399, w_101_400, w_101_401, w_101_402, w_101_403, w_101_404, w_101_408, w_101_409, w_101_412, w_101_415, w_101_416, w_101_418, w_101_420, w_101_421, w_101_422, w_101_424, w_101_429, w_101_431, w_101_432, w_101_435, w_101_436, w_101_437, w_101_439, w_101_441, w_101_448, w_101_449, w_101_450, w_101_451, w_101_453, w_101_454, w_101_456, w_101_457, w_101_459, w_101_463, w_101_465, w_101_466, w_101_467, w_101_470, w_101_476, w_101_478, w_101_479, w_101_481, w_101_483, w_101_486, w_101_487, w_101_490, w_101_494, w_101_495, w_101_496, w_101_497, w_101_501, w_101_503, w_101_505, w_101_508, w_101_509, w_101_511, w_101_512, w_101_513, w_101_514, w_101_515, w_101_516, w_101_517, w_101_518, w_101_522, w_101_524, w_101_525, w_101_526, w_101_530, w_101_537, w_101_538, w_101_540, w_101_541, w_101_544, w_101_545, w_101_546, w_101_547, w_101_551, w_101_552, w_101_554, w_101_557, w_101_558, w_101_559, w_101_560, w_101_562, w_101_566, w_101_567, w_101_569, w_101_570, w_101_571, w_101_576, w_101_578, w_101_579, w_101_580, w_101_583, w_101_586, w_101_589, w_101_591, w_101_595, w_101_597, w_101_598, w_101_601, w_101_602, w_101_605, w_101_606, w_101_609, w_101_610, w_101_614, w_101_615, w_101_617, w_101_620, w_101_621, w_101_622, w_101_623, w_101_624, w_101_625, w_101_630, w_101_631, w_101_632, w_101_634, w_101_635, w_101_636, w_101_640, w_101_641, w_101_643, w_101_644, w_101_647, w_101_649, w_101_650, w_101_651, w_101_652, w_101_653, w_101_654, w_101_655, w_101_656, w_101_658, w_101_661, w_101_666, w_101_667, w_101_668, w_101_672, w_101_673, w_101_676, w_101_679, w_101_683, w_101_685, w_101_686, w_101_687, w_101_689, w_101_690, w_101_691, w_101_693, w_101_697, w_101_702, w_101_705, w_101_709, w_101_710, w_101_711, w_101_715, w_101_716, w_101_717, w_101_719, w_101_720, w_101_722, w_101_725, w_101_726, w_101_727, w_101_730, w_101_733, w_101_735, w_101_738, w_101_741, w_101_743, w_101_749, w_101_750, w_101_752, w_101_754, w_101_756, w_101_761, w_101_768, w_101_770, w_101_771, w_101_777, w_101_778, w_101_779, w_101_780, w_101_782, w_101_784, w_101_785, w_101_788, w_101_791, w_101_792, w_101_796, w_101_797, w_101_798, w_101_800, w_101_801, w_101_802, w_101_805, w_101_806, w_101_807, w_101_809, w_101_812, w_101_814, w_101_823, w_101_825, w_101_827, w_101_828, w_101_831, w_101_832, w_101_835, w_101_837, w_101_838, w_101_839, w_101_842, w_101_843, w_101_844, w_101_845, w_101_847, w_101_849, w_101_850, w_101_851, w_101_852, w_101_855, w_101_856, w_101_858, w_101_859, w_101_863, w_101_871, w_101_874, w_101_875, w_101_876, w_101_877, w_101_879, w_101_880, w_101_881, w_101_884, w_101_887, w_101_896, w_101_903, w_101_905, w_101_909, w_101_910, w_101_911, w_101_913, w_101_915, w_101_916, w_101_917, w_101_918, w_101_920, w_101_922, w_101_923, w_101_924, w_101_926, w_101_927, w_101_930, w_101_931, w_101_933, w_101_935, w_101_936, w_101_938, w_101_939, w_101_940, w_101_942, w_101_946, w_101_947, w_101_949, w_101_950, w_101_952, w_101_953, w_101_954, w_101_955, w_101_957, w_101_959, w_101_960, w_101_961, w_101_964, w_101_966, w_101_967, w_101_968, w_101_970, w_101_972, w_101_973, w_101_975, w_101_984, w_101_985, w_101_986, w_101_987, w_101_989, w_101_990, w_101_993, w_101_996, w_101_999, w_101_1002, w_101_1004, w_101_1005, w_101_1006, w_101_1007, w_101_1012, w_101_1013, w_101_1015, w_101_1017, w_101_1019, w_101_1020, w_101_1021, w_101_1022, w_101_1023, w_101_1026, w_101_1027, w_101_1030, w_101_1031, w_101_1032, w_101_1033, w_101_1035, w_101_1039, w_101_1040, w_101_1041, w_101_1047, w_101_1049, w_101_1050, w_101_1052, w_101_1054, w_101_1064, w_101_1067, w_101_1069, w_101_1071, w_101_1074, w_101_1075, w_101_1078, w_101_1083, w_101_1084, w_101_1086, w_101_1089, w_101_1091, w_101_1092, w_101_1093, w_101_1094, w_101_1095, w_101_1099, w_101_1101, w_101_1102, w_101_1108, w_101_1112, w_101_1114, w_101_1115, w_101_1118, w_101_1119, w_101_1125, w_101_1129, w_101_1131, w_101_1132, w_101_1139, w_101_1144, w_101_1147, w_101_1149, w_101_1151, w_101_1160, w_101_1168, w_101_1169, w_101_1171, w_101_1173, w_101_1174, w_101_1177, w_101_1178, w_101_1179, w_101_1180, w_101_1182, w_101_1184, w_101_1186, w_101_1187, w_101_1189, w_101_1193, w_101_1196, w_101_1199, w_101_1200, w_101_1202, w_101_1209, w_101_1219, w_101_1220, w_101_1221, w_101_1224, w_101_1225, w_101_1227, w_101_1228, w_101_1230, w_101_1232, w_101_1235, w_101_1238, w_101_1240, w_101_1241, w_101_1246, w_101_1247, w_101_1250, w_101_1252, w_101_1260, w_101_1264, w_101_1273, w_101_1275, w_101_1279, w_101_1280, w_101_1283, w_101_1284, w_101_1287, w_101_1289, w_101_1294, w_101_1304, w_101_1306, w_101_1309, w_101_1311, w_101_1315, w_101_1317, w_101_1320, w_101_1321, w_101_1323, w_101_1328, w_101_1330, w_101_1333, w_101_1335, w_101_1341, w_101_1342, w_101_1345, w_101_1349, w_101_1355, w_101_1356, w_101_1359, w_101_1362, w_101_1363, w_101_1366, w_101_1369, w_101_1370, w_101_1371, w_101_1374, w_101_1375, w_101_1376, w_101_1377, w_101_1382, w_101_1385, w_101_1386, w_101_1390, w_101_1391, w_101_1395, w_101_1396, w_101_1398, w_101_1400, w_101_1401, w_101_1408, w_101_1410, w_101_1411, w_101_1413, w_101_1415, w_101_1419, w_101_1420, w_101_1423, w_101_1426, w_101_1427, w_101_1433, w_101_1434, w_101_1437, w_101_1439, w_101_1441, w_101_1443, w_101_1448, w_101_1449, w_101_1452, w_101_1457, w_101_1458, w_101_1461, w_101_1463, w_101_1468, w_101_1469, w_101_1470, w_101_1471, w_101_1474, w_101_1475, w_101_1479, w_101_1485, w_101_1488, w_101_1489, w_101_1495, w_101_1499, w_101_1503, w_101_1504, w_101_1505, w_101_1508, w_101_1511, w_101_1512, w_101_1517, w_101_1520, w_101_1521, w_101_1524, w_101_1525, w_101_1527, w_101_1529, w_101_1530, w_101_1537, w_101_1539, w_101_1541, w_101_1542, w_101_1545, w_101_1546, w_101_1548, w_101_1549, w_101_1550, w_101_1551, w_101_1552, w_101_1553, w_101_1554, w_101_1555, w_101_1556, w_101_1559, w_101_1560, w_101_1561, w_101_1568, w_101_1569, w_101_1571, w_101_1574, w_101_1576, w_101_1577, w_101_1578, w_101_1583, w_101_1586, w_101_1588, w_101_1592, w_101_1593, w_101_1594, w_101_1595, w_101_1598, w_101_1599, w_101_1600, w_101_1605, w_101_1606, w_101_1609, w_101_1611, w_101_1613, w_101_1615, w_101_1617, w_101_1620, w_101_1621, w_101_1622, w_101_1625, w_101_1630, w_101_1632, w_101_1638, w_101_1640, w_101_1641, w_101_1642, w_101_1643, w_101_1644, w_101_1646, w_101_1649, w_101_1650, w_101_1651, w_101_1652, w_101_1655, w_101_1657, w_101_1658, w_101_1660, w_101_1661, w_101_1662, w_101_1665, w_101_1667, w_101_1669, w_101_1671, w_101_1676, w_101_1677, w_101_1681, w_101_1685, w_101_1686, w_101_1691, w_101_1692, w_101_1695, w_101_1696, w_101_1701, w_101_1702, w_101_1704, w_101_1707, w_101_1708, w_101_1710, w_101_1714, w_101_1715, w_101_1717, w_101_1719, w_101_1722, w_101_1723, w_101_1728, w_101_1734, w_101_1735, w_101_1737, w_101_1743, w_101_1746, w_101_1747, w_101_1748, w_101_1753, w_101_1756, w_101_1759, w_101_1760, w_101_1762, w_101_1763, w_101_1764, w_101_1765, w_101_1766, w_101_1771, w_101_1776, w_101_1777, w_101_1779, w_101_1781, w_101_1783, w_101_1786, w_101_1788, w_101_1792, w_101_1793, w_101_1794, w_101_1795, w_101_1796, w_101_1797, w_101_1798, w_101_1800, w_101_1801, w_101_1804, w_101_1805, w_101_1806, w_101_1808, w_101_1810, w_101_1814, w_101_1815, w_101_1819, w_101_1823, w_101_1825, w_101_1828, w_101_1835, w_101_1836, w_101_1842, w_101_1844, w_101_1846, w_101_1849, w_101_1850, w_101_1854, w_101_1856, w_101_1857, w_101_1859, w_101_1863, w_101_1864, w_101_1869, w_101_1870, w_101_1872, w_101_1873, w_101_1879, w_101_1886, w_101_1889, w_101_1892, w_101_1900, w_101_1914, w_101_1916, w_101_1919, w_101_1922, w_101_1925, w_101_1930, w_101_1931, w_101_1933, w_101_1935, w_101_1936, w_101_1937, w_101_1939, w_101_1941, w_101_1944, w_101_1946, w_101_1947, w_101_1953, w_101_1956, w_101_1958, w_101_1959, w_101_1960, w_101_1961, w_101_1965, w_101_1967, w_101_1969, w_101_1972, w_101_1973, w_101_1974, w_101_1975, w_101_1976, w_101_1980, w_101_1981, w_101_1987, w_101_1988, w_101_1989, w_101_1999, w_101_2000, w_101_2003, w_101_2006, w_101_2008, w_101_2011, w_101_2015, w_101_2016, w_101_2021, w_101_2024, w_101_2037, w_101_2038, w_101_2039, w_101_2041, w_101_2042, w_101_2043, w_101_2045, w_101_2046, w_101_2047, w_101_2049, w_101_2052, w_101_2053, w_101_2057, w_101_2061, w_101_2063, w_101_2066, w_101_2068, w_101_2069, w_101_2079, w_101_2080, w_101_2084, w_101_2086, w_101_2087, w_101_2090, w_101_2091, w_101_2094, w_101_2095, w_101_2096, w_101_2097, w_101_2098, w_101_2099, w_101_2104, w_101_2108, w_101_2109, w_101_2110, w_101_2115, w_101_2116, w_101_2119, w_101_2120, w_101_2122, w_101_2123, w_101_2124, w_101_2130, w_101_2134, w_101_2140, w_101_2143, w_101_2145, w_101_2148, w_101_2155, w_101_2158, w_101_2162, w_101_2164, w_101_2165, w_101_2167, w_101_2168, w_101_2170, w_101_2172, w_101_2173, w_101_2175, w_101_2183, w_101_2187, w_101_2188, w_101_2191, w_101_2194, w_101_2195, w_101_2201, w_101_2204, w_101_2205, w_101_2213, w_101_2216, w_101_2218, w_101_2219, w_101_2220, w_101_2227, w_101_2228, w_101_2238, w_101_2241, w_101_2248, w_101_2249, w_101_2250, w_101_2251, w_101_2253, w_101_2254, w_101_2255, w_101_2258, w_101_2260, w_101_2265, w_101_2267, w_101_2268, w_101_2269, w_101_2271, w_101_2275, w_101_2277, w_101_2280, w_101_2281, w_101_2283, w_101_2287, w_101_2289, w_101_2290, w_101_2291, w_101_2295, w_101_2296, w_101_2299, w_101_2300, w_101_2301, w_101_2303, w_101_2304, w_101_2307, w_101_2314, w_101_2316, w_101_2323, w_101_2324, w_101_2329, w_101_2332, w_101_2333, w_101_2334, w_101_2335, w_101_2337, w_101_2338, w_101_2339, w_101_2340, w_101_2341, w_101_2346, w_101_2347, w_101_2348, w_101_2350, w_101_2353, w_101_2354, w_101_2363, w_101_2364, w_101_2365, w_101_2368, w_101_2372, w_101_2374, w_101_2375, w_101_2380, w_101_2382, w_101_2384, w_101_2390, w_101_2391, w_101_2392, w_101_2394, w_101_2399, w_101_2402, w_101_2403, w_101_2404, w_101_2412, w_101_2414, w_101_2418, w_101_2419, w_101_2425, w_101_2429, w_101_2432, w_101_2436, w_101_2440, w_101_2443, w_101_2444, w_101_2446, w_101_2448, w_101_2454, w_101_2459, w_101_2461, w_101_2462, w_101_2463, w_101_2464, w_101_2465, w_101_2474, w_101_2477, w_101_2478, w_101_2481, w_101_2484, w_101_2493, w_101_2495, w_101_2496, w_101_2497, w_101_2498, w_101_2500, w_101_2501, w_101_2503, w_101_2506, w_101_2514, w_101_2517, w_101_2518, w_101_2519, w_101_2520, w_101_2521, w_101_2523, w_101_2531, w_101_2536, w_101_2537, w_101_2540, w_101_2543, w_101_2547, w_101_2548, w_101_2549, w_101_2550, w_101_2551, w_101_2555, w_101_2556, w_101_2561, w_101_2564, w_101_2570, w_101_2571, w_101_2573, w_101_2574, w_101_2581, w_101_2583, w_101_2587, w_101_2588, w_101_2592, w_101_2593, w_101_2598, w_101_2600, w_101_2606, w_101_2609, w_101_2610, w_101_2612, w_101_2614, w_101_2615, w_101_2618, w_101_2619, w_101_2620, w_101_2623, w_101_2626, w_101_2627, w_101_2631, w_101_2633, w_101_2634, w_101_2635, w_101_2638, w_101_2640, w_101_2643, w_101_2645, w_101_2648, w_101_2649, w_101_2656, w_101_2658, w_101_2662, w_101_2663, w_101_2665, w_101_2668, w_101_2670, w_101_2672, w_101_2674, w_101_2675, w_101_2676, w_101_2680, w_101_2682, w_101_2683, w_101_2685, w_101_2686, w_101_2692, w_101_2695, w_101_2696, w_101_2698, w_101_2711, w_101_2717, w_101_2719, w_101_2722, w_101_2724, w_101_2725, w_101_2729, w_101_2730, w_101_2736, w_101_2738, w_101_2739, w_101_2740, w_101_2741, w_101_2745, w_101_2747, w_101_2749, w_101_2750, w_101_2751, w_101_2753, w_101_2754, w_101_2757, w_101_2758, w_101_2759, w_101_2760, w_101_2763, w_101_2764, w_101_2765, w_101_2767, w_101_2769, w_101_2771, w_101_2772, w_101_2773, w_101_2774, w_101_2776, w_101_2779, w_101_2783, w_101_2785, w_101_2786, w_101_2792, w_101_2793, w_101_2796, w_101_2797, w_101_2798, w_101_2801, w_101_2803, w_101_2812, w_101_2814, w_101_2815, w_101_2816, w_101_2817, w_101_2818, w_101_2822, w_101_2824, w_101_2827, w_101_2829, w_101_2831, w_101_2832, w_101_2837, w_101_2840, w_101_2842, w_101_2845, w_101_2847, w_101_2849, w_101_2850, w_101_2853, w_101_2856, w_101_2857, w_101_2860, w_101_2866, w_101_2869, w_101_2870, w_101_2871, w_101_2872, w_101_2873, w_101_2875, w_101_2878, w_101_2881, w_101_2884, w_101_2887, w_101_2892, w_101_2893, w_101_2896, w_101_2897, w_101_2902, w_101_2904, w_101_2909, w_101_2910, w_101_2912, w_101_2913, w_101_2914, w_101_2916, w_101_2918, w_101_2920, w_101_2922, w_101_2923, w_101_2935, w_101_2943, w_101_2949, w_101_2955, w_101_2956, w_101_2958, w_101_2961, w_101_2963, w_101_2965, w_101_2966, w_101_2968, w_101_2970, w_101_2971, w_101_2972, w_101_2977, w_101_2984, w_101_2985, w_101_2986, w_101_2990, w_101_2991, w_101_2995, w_101_3000, w_101_3003, w_101_3004, w_101_3005, w_101_3010, w_101_3011, w_101_3018, w_101_3020, w_101_3025, w_101_3029, w_101_3031, w_101_3034, w_101_3040, w_101_3042, w_101_3043, w_101_3044, w_101_3050, w_101_3053, w_101_3055, w_101_3056, w_101_3060, w_101_3062, w_101_3063, w_101_3064, w_101_3068, w_101_3070, w_101_3072, w_101_3073, w_101_3075, w_101_3076, w_101_3084, w_101_3085, w_101_3088, w_101_3090, w_101_3093, w_101_3095, w_101_3100, w_101_3101, w_101_3106, w_101_3108, w_101_3111, w_101_3113, w_101_3116, w_101_3120, w_101_3123, w_101_3127, w_101_3129, w_101_3130, w_101_3134, w_101_3137, w_101_3138, w_101_3140, w_101_3141, w_101_3143, w_101_3145, w_101_3151, w_101_3155, w_101_3156, w_101_3157, w_101_3164, w_101_3168, w_101_3171, w_101_3172, w_101_3173, w_101_3175, w_101_3177, w_101_3178, w_101_3180, w_101_3182, w_101_3183, w_101_3184, w_101_3185, w_101_3187, w_101_3196, w_101_3198, w_101_3201, w_101_3202, w_101_3205, w_101_3206, w_101_3207, w_101_3209, w_101_3212, w_101_3216, w_101_3220, w_101_3221, w_101_3224, w_101_3226, w_101_3229, w_101_3230, w_101_3233, w_101_3238, w_101_3240, w_101_3241, w_101_3244, w_101_3248, w_101_3249, w_101_3250, w_101_3251, w_101_3252, w_101_3254, w_101_3256, w_101_3257, w_101_3261, w_101_3263, w_101_3265, w_101_3266, w_101_3267, w_101_3276, w_101_3277, w_101_3279, w_101_3282, w_101_3285, w_101_3286, w_101_3290, w_101_3291, w_101_3292, w_101_3293, w_101_3294, w_101_3299, w_101_3301, w_101_3304, w_101_3305, w_101_3307, w_101_3316, w_101_3318, w_101_3320, w_101_3322, w_101_3326, w_101_3330, w_101_3331, w_101_3336, w_101_3340, w_101_3348, w_101_3351, w_101_3357, w_101_3361, w_101_3363, w_101_3365, w_101_3368, w_101_3369, w_101_3376, w_101_3378, w_101_3384, w_101_3389, w_101_3391, w_101_3393, w_101_3394, w_101_3395, w_101_3396, w_101_3402, w_101_3414, w_101_3418, w_101_3419, w_101_3423, w_101_3424, w_101_3426, w_101_3429, w_101_3430, w_101_3432, w_101_3435, w_101_3436, w_101_3437, w_101_3438, w_101_3439, w_101_3441, w_101_3444, w_101_3449, w_101_3456, w_101_3459, w_101_3463, w_101_3465, w_101_3468, w_101_3470, w_101_3480, w_101_3481, w_101_3483, w_101_3484, w_101_3485, w_101_3486, w_101_3494, w_101_3496, w_101_3499, w_101_3502, w_101_3504, w_101_3509, w_101_3513, w_101_3514, w_101_3517, w_101_3522, w_101_3526, w_101_3532, w_101_3535, w_101_3544, w_101_3547, w_101_3550, w_101_3551, w_101_3560, w_101_3563, w_101_3567, w_101_3568, w_101_3569, w_101_3570, w_101_3573, w_101_3579, w_101_3580, w_101_3582, w_101_3584, w_101_3588, w_101_3599, w_101_3601, w_101_3602, w_101_3604, w_101_3606, w_101_3607, w_101_3610, w_101_3611, w_101_3613, w_101_3615, w_101_3617, w_101_3624, w_101_3628, w_101_3629, w_101_3635, w_101_3639, w_101_3640, w_101_3641, w_101_3643, w_101_3644, w_101_3645, w_101_3650, w_101_3651, w_101_3653, w_101_3657, w_101_3660, w_101_3661, w_101_3665, w_101_3670, w_101_3671, w_101_3676, w_101_3680, w_101_3681, w_101_3683, w_101_3688, w_101_3690, w_101_3693, w_101_3694, w_101_3699, w_101_3701, w_101_3704, w_101_3707, w_101_3708, w_101_3709, w_101_3710, w_101_3711, w_101_3716, w_101_3719, w_101_3720, w_101_3721, w_101_3724, w_101_3730, w_101_3731, w_101_3734, w_101_3736, w_101_3739, w_101_3740, w_101_3747, w_101_3749, w_101_3758, w_101_3760, w_101_3764, w_101_3765, w_101_3771, w_101_3772, w_101_3778, w_101_3780, w_101_3781, w_101_3782, w_101_3784, w_101_3785, w_101_3786, w_101_3788, w_101_3789, w_101_3790, w_101_3792, w_101_3797, w_101_3799, w_101_3800, w_101_3808, w_101_3812, w_101_3813, w_101_3819, w_101_3820, w_101_3822, w_101_3825, w_101_3830, w_101_3831, w_101_3832, w_101_3833, w_101_3834, w_101_3837, w_101_3840, w_101_3841, w_101_3842, w_101_3845, w_101_3846, w_101_3848, w_101_3851, w_101_3857, w_101_3859, w_101_3860, w_101_3861, w_101_3865, w_101_3868, w_101_3872, w_101_3874, w_101_3875, w_101_3877, w_101_3886, w_101_3890, w_101_3892, w_101_3893, w_101_3897, w_101_3907, w_101_3909, w_101_3913, w_101_3919, w_101_3921, w_101_3922, w_101_3924, w_101_3929, w_101_3937, w_101_3939, w_101_3943, w_101_3948, w_101_3949, w_101_3951, w_101_3952, w_101_3953, w_101_3958, w_101_3960, w_101_3962, w_101_3964, w_101_3965, w_101_3966, w_101_3967, w_101_3968, w_101_3969, w_101_3971, w_101_3972, w_101_3975, w_101_3977, w_101_3978, w_101_3980, w_101_3983, w_101_3986, w_101_3987, w_101_3989, w_101_3993, w_101_3994, w_101_3998, w_101_4000, w_101_4001, w_101_4002, w_101_4003, w_101_4009, w_101_4012, w_101_4014, w_101_4016, w_101_4018, w_101_4025, w_101_4028, w_101_4031, w_101_4032, w_101_4038, w_101_4040, w_101_4041, w_101_4043, w_101_4047, w_101_4048, w_101_4049, w_101_4050, w_101_4051, w_101_4052, w_101_4057, w_101_4058, w_101_4060, w_101_4065, w_101_4068, w_101_4069, w_101_4070, w_101_4071, w_101_4079, w_101_4082, w_101_4083, w_101_4084, w_101_4087, w_101_4090, w_101_4092, w_101_4093, w_101_4100, w_101_4102, w_101_4105, w_101_4106, w_101_4109, w_101_4111, w_101_4114, w_101_4116, w_101_4119, w_101_4120, w_101_4121, w_101_4125, w_101_4127, w_101_4128, w_101_4131, w_101_4136, w_101_4139, w_101_4140, w_101_4144, w_101_4150, w_101_4158, w_101_4159, w_101_4167, w_101_4170, w_101_4172, w_101_4173, w_101_4176, w_101_4186, w_101_4188, w_101_4194, w_101_4197, w_101_4199, w_101_4201, w_101_4203, w_101_4205, w_101_4206, w_101_4207, w_101_4211, w_101_4213, w_101_4214, w_101_4221, w_101_4224, w_101_4225, w_101_4227, w_101_4228, w_101_4231, w_101_4232, w_101_4234, w_101_4235, w_101_4239, w_101_4243, w_101_4244, w_101_4248, w_101_4249, w_101_4250, w_101_4251, w_101_4254, w_101_4255, w_101_4256, w_101_4257, w_101_4258, w_101_4262, w_101_4263, w_101_4267, w_101_4269, w_101_4273, w_101_4275, w_101_4277, w_101_4279, w_101_4285, w_101_4286, w_101_4287, w_101_4292, w_101_4293, w_101_4294, w_101_4301, w_101_4307, w_101_4308, w_101_4310, w_101_4313, w_101_4314, w_101_4317, w_101_4318, w_101_4321, w_101_4322, w_101_4325, w_101_4328, w_101_4329, w_101_4334, w_101_4335, w_101_4337, w_101_4338, w_101_4339, w_101_4341, w_101_4343, w_101_4344, w_101_4345, w_101_4348, w_101_4352, w_101_4354, w_101_4358, w_101_4359, w_101_4363, w_101_4367, w_101_4370, w_101_4372, w_101_4377, w_101_4392, w_101_4393, w_101_4397, w_101_4398, w_101_4403, w_101_4406, w_101_4407, w_101_4412, w_101_4414, w_101_4419, w_101_4422, w_101_4424, w_101_4431, w_101_4438, w_101_4441, w_101_4446, w_101_4447, w_101_4448, w_101_4453, w_101_4454, w_101_4455, w_101_4456, w_101_4457, w_101_4460, w_101_4462, w_101_4468, w_101_4470, w_101_4471, w_101_4473, w_101_4474, w_101_4475;
  wire w_102_000, w_102_001, w_102_002, w_102_003, w_102_004, w_102_005, w_102_006, w_102_008, w_102_010, w_102_011, w_102_012, w_102_013, w_102_014, w_102_016, w_102_017, w_102_018, w_102_019, w_102_020, w_102_021, w_102_022, w_102_023, w_102_024, w_102_025, w_102_027, w_102_028, w_102_029, w_102_030, w_102_031, w_102_032, w_102_033, w_102_034, w_102_035, w_102_036, w_102_037, w_102_038, w_102_039, w_102_040, w_102_041, w_102_045, w_102_046, w_102_047, w_102_048, w_102_049, w_102_050, w_102_051, w_102_052, w_102_053, w_102_054, w_102_058, w_102_060, w_102_061, w_102_063, w_102_065, w_102_066, w_102_067, w_102_068, w_102_069, w_102_070, w_102_072, w_102_075, w_102_076, w_102_079, w_102_080, w_102_081, w_102_083, w_102_084, w_102_085, w_102_086, w_102_087, w_102_088, w_102_089, w_102_090, w_102_091, w_102_092, w_102_094, w_102_095, w_102_096, w_102_097, w_102_102, w_102_103, w_102_105, w_102_108, w_102_111, w_102_112, w_102_113, w_102_114, w_102_115, w_102_116, w_102_117, w_102_118, w_102_119, w_102_121, w_102_122, w_102_123, w_102_124, w_102_125, w_102_126, w_102_127, w_102_129, w_102_130, w_102_131, w_102_132, w_102_133, w_102_135, w_102_136, w_102_137, w_102_138, w_102_139, w_102_140, w_102_141, w_102_142, w_102_143, w_102_144, w_102_146, w_102_147, w_102_148, w_102_149, w_102_150, w_102_151, w_102_154, w_102_156, w_102_159, w_102_160, w_102_163, w_102_165, w_102_166, w_102_168, w_102_169, w_102_171, w_102_173, w_102_174, w_102_176, w_102_177, w_102_179, w_102_180, w_102_181, w_102_182, w_102_183, w_102_185, w_102_187, w_102_188, w_102_189, w_102_191, w_102_192, w_102_193, w_102_194, w_102_195, w_102_196, w_102_197, w_102_198, w_102_199, w_102_200, w_102_201, w_102_202, w_102_203, w_102_205, w_102_206, w_102_207, w_102_209, w_102_210, w_102_211, w_102_212, w_102_213, w_102_216, w_102_217, w_102_218, w_102_219, w_102_220, w_102_223, w_102_225, w_102_226, w_102_227, w_102_228, w_102_229, w_102_230, w_102_232, w_102_233, w_102_234, w_102_235, w_102_237, w_102_238, w_102_239, w_102_240, w_102_242, w_102_243, w_102_244, w_102_247, w_102_249, w_102_250, w_102_252, w_102_253, w_102_256, w_102_257, w_102_258, w_102_261, w_102_264, w_102_265, w_102_266, w_102_268, w_102_269, w_102_271, w_102_272, w_102_273, w_102_274, w_102_276, w_102_277, w_102_279, w_102_281, w_102_283, w_102_284, w_102_285, w_102_286, w_102_287, w_102_288, w_102_289, w_102_290, w_102_291, w_102_292, w_102_297, w_102_299, w_102_300, w_102_301, w_102_303, w_102_305, w_102_307, w_102_309, w_102_310, w_102_311, w_102_312, w_102_313, w_102_314, w_102_317, w_102_318, w_102_320, w_102_321, w_102_322, w_102_323, w_102_324, w_102_325, w_102_326, w_102_327, w_102_328, w_102_331, w_102_332, w_102_333, w_102_334, w_102_335, w_102_336, w_102_339, w_102_340, w_102_345, w_102_346, w_102_347, w_102_349, w_102_350, w_102_353, w_102_354, w_102_356, w_102_358, w_102_360, w_102_361, w_102_362, w_102_363, w_102_364, w_102_367, w_102_368, w_102_369, w_102_371, w_102_372, w_102_373, w_102_375, w_102_376, w_102_377, w_102_379, w_102_380, w_102_382, w_102_386, w_102_387, w_102_389, w_102_391, w_102_392, w_102_393, w_102_394, w_102_396, w_102_397, w_102_399, w_102_400, w_102_401, w_102_402, w_102_404, w_102_405, w_102_407, w_102_408, w_102_410, w_102_412, w_102_414, w_102_416, w_102_417, w_102_418, w_102_421, w_102_422, w_102_423, w_102_424, w_102_425, w_102_426, w_102_429, w_102_432, w_102_434, w_102_435, w_102_436, w_102_437, w_102_438, w_102_441, w_102_445, w_102_446, w_102_447, w_102_448, w_102_449, w_102_450, w_102_452, w_102_453, w_102_454, w_102_456, w_102_457, w_102_458, w_102_459, w_102_460, w_102_461, w_102_463, w_102_465, w_102_466, w_102_468, w_102_470, w_102_472, w_102_474, w_102_475, w_102_476, w_102_477, w_102_478, w_102_479, w_102_480, w_102_481, w_102_485, w_102_490, w_102_492, w_102_495, w_102_499, w_102_504, w_102_505, w_102_506, w_102_507, w_102_508, w_102_509, w_102_510, w_102_511, w_102_512, w_102_514, w_102_515, w_102_518, w_102_519, w_102_520, w_102_524, w_102_525, w_102_526, w_102_531, w_102_532, w_102_535, w_102_537, w_102_538, w_102_539, w_102_540, w_102_541, w_102_542, w_102_543, w_102_544, w_102_545, w_102_546, w_102_547, w_102_549, w_102_551, w_102_552, w_102_554, w_102_555, w_102_556, w_102_558, w_102_559, w_102_563, w_102_565, w_102_566, w_102_567, w_102_568, w_102_570, w_102_571, w_102_572, w_102_573, w_102_574, w_102_575, w_102_576, w_102_577, w_102_578, w_102_581, w_102_582, w_102_583, w_102_585, w_102_592, w_102_593, w_102_595, w_102_597, w_102_599, w_102_600, w_102_601, w_102_602, w_102_604, w_102_605, w_102_606, w_102_608, w_102_610, w_102_611, w_102_612, w_102_613, w_102_615, w_102_616, w_102_620, w_102_622, w_102_623, w_102_624, w_102_625, w_102_627, w_102_629, w_102_631, w_102_633, w_102_640, w_102_642, w_102_643, w_102_645, w_102_646, w_102_648, w_102_649, w_102_650, w_102_651, w_102_652, w_102_653, w_102_654, w_102_655, w_102_659, w_102_660, w_102_662, w_102_663, w_102_668, w_102_669, w_102_670, w_102_672, w_102_675, w_102_676, w_102_679, w_102_682, w_102_684, w_102_687, w_102_689, w_102_691, w_102_692, w_102_694, w_102_695, w_102_696, w_102_697, w_102_699, w_102_701, w_102_703, w_102_704, w_102_706, w_102_707, w_102_710, w_102_712, w_102_714, w_102_715, w_102_716, w_102_719, w_102_721, w_102_724, w_102_725, w_102_726, w_102_729, w_102_730, w_102_731, w_102_732, w_102_733, w_102_735, w_102_737, w_102_739, w_102_740, w_102_744, w_102_745, w_102_748, w_102_751, w_102_752, w_102_753, w_102_755, w_102_761, w_102_763, w_102_764, w_102_766, w_102_767, w_102_769, w_102_770, w_102_774, w_102_775, w_102_778, w_102_779, w_102_781, w_102_783, w_102_785, w_102_787, w_102_789, w_102_791, w_102_792, w_102_793, w_102_794, w_102_796, w_102_797, w_102_798, w_102_799, w_102_800, w_102_801, w_102_802, w_102_803, w_102_804, w_102_806, w_102_807, w_102_809, w_102_811, w_102_813, w_102_814, w_102_815, w_102_817, w_102_818, w_102_819, w_102_820, w_102_821, w_102_822, w_102_824, w_102_827, w_102_828, w_102_829, w_102_830, w_102_833, w_102_834, w_102_835, w_102_836, w_102_839, w_102_841, w_102_842, w_102_844, w_102_845, w_102_850, w_102_851, w_102_852, w_102_853, w_102_854, w_102_857, w_102_858, w_102_859, w_102_864, w_102_865, w_102_866, w_102_867, w_102_868, w_102_870, w_102_871, w_102_875, w_102_878, w_102_880, w_102_881, w_102_882, w_102_883, w_102_885, w_102_886, w_102_888, w_102_890, w_102_891, w_102_892, w_102_893, w_102_895, w_102_896, w_102_897, w_102_900, w_102_901, w_102_902, w_102_903, w_102_904, w_102_906, w_102_908, w_102_909, w_102_912, w_102_913, w_102_914, w_102_915, w_102_918, w_102_919, w_102_920, w_102_921, w_102_922, w_102_923, w_102_924, w_102_925, w_102_927, w_102_929, w_102_930, w_102_931, w_102_933, w_102_934, w_102_935, w_102_936, w_102_937, w_102_938, w_102_939, w_102_940, w_102_941, w_102_942, w_102_943, w_102_946, w_102_947, w_102_949, w_102_950, w_102_952, w_102_954, w_102_956, w_102_957, w_102_959, w_102_960, w_102_963, w_102_964, w_102_966, w_102_967, w_102_968, w_102_970, w_102_971, w_102_972, w_102_973, w_102_976, w_102_977, w_102_979, w_102_980, w_102_983, w_102_985, w_102_986, w_102_987, w_102_988, w_102_992, w_102_993, w_102_994, w_102_995, w_102_996, w_102_999, w_102_1001, w_102_1002, w_102_1004, w_102_1006, w_102_1007, w_102_1008, w_102_1009, w_102_1010, w_102_1012, w_102_1013, w_102_1014, w_102_1015, w_102_1017, w_102_1018, w_102_1019, w_102_1022, w_102_1025, w_102_1026, w_102_1029, w_102_1030, w_102_1031, w_102_1033, w_102_1034, w_102_1036, w_102_1037, w_102_1038, w_102_1039, w_102_1040, w_102_1043, w_102_1044, w_102_1045, w_102_1046, w_102_1049, w_102_1050, w_102_1051, w_102_1052, w_102_1053, w_102_1055, w_102_1057, w_102_1060, w_102_1062, w_102_1066, w_102_1068, w_102_1069, w_102_1070, w_102_1071, w_102_1072, w_102_1073, w_102_1074, w_102_1075, w_102_1077, w_102_1080, w_102_1083, w_102_1084, w_102_1085, w_102_1087, w_102_1089, w_102_1090, w_102_1092, w_102_1095, w_102_1096, w_102_1099, w_102_1100, w_102_1105, w_102_1106, w_102_1107, w_102_1108, w_102_1111, w_102_1112, w_102_1115, w_102_1116, w_102_1117, w_102_1118, w_102_1119, w_102_1120, w_102_1121, w_102_1122, w_102_1123, w_102_1124, w_102_1125, w_102_1126, w_102_1127, w_102_1129, w_102_1130, w_102_1132, w_102_1133, w_102_1135, w_102_1137, w_102_1139, w_102_1140, w_102_1141, w_102_1146, w_102_1147, w_102_1148, w_102_1149, w_102_1152, w_102_1155, w_102_1156, w_102_1158, w_102_1160, w_102_1161, w_102_1164, w_102_1165, w_102_1166, w_102_1167, w_102_1168, w_102_1169, w_102_1170, w_102_1173, w_102_1174, w_102_1176, w_102_1177, w_102_1179, w_102_1183, w_102_1184, w_102_1187, w_102_1188, w_102_1189, w_102_1191, w_102_1192, w_102_1193, w_102_1195, w_102_1196, w_102_1197, w_102_1198, w_102_1199, w_102_1200, w_102_1201, w_102_1202, w_102_1204, w_102_1205, w_102_1208, w_102_1209, w_102_1211, w_102_1214, w_102_1216, w_102_1217, w_102_1218, w_102_1220, w_102_1223, w_102_1224, w_102_1225, w_102_1227, w_102_1230, w_102_1234, w_102_1235, w_102_1237, w_102_1238, w_102_1240, w_102_1243, w_102_1244, w_102_1245, w_102_1246, w_102_1247, w_102_1248, w_102_1249, w_102_1250, w_102_1251, w_102_1252, w_102_1253, w_102_1255, w_102_1257, w_102_1258, w_102_1259, w_102_1260, w_102_1261, w_102_1262, w_102_1264, w_102_1265, w_102_1267, w_102_1268, w_102_1271, w_102_1274, w_102_1275, w_102_1277, w_102_1279, w_102_1280, w_102_1281, w_102_1282, w_102_1283, w_102_1290, w_102_1292, w_102_1293, w_102_1294, w_102_1295, w_102_1296, w_102_1297, w_102_1299, w_102_1301, w_102_1302, w_102_1303, w_102_1306, w_102_1309, w_102_1311, w_102_1312, w_102_1315, w_102_1318, w_102_1319, w_102_1320, w_102_1322, w_102_1323, w_102_1324, w_102_1325, w_102_1326, w_102_1327, w_102_1328, w_102_1329, w_102_1330, w_102_1334, w_102_1336, w_102_1338, w_102_1339, w_102_1341, w_102_1342, w_102_1347, w_102_1349, w_102_1350, w_102_1351, w_102_1354, w_102_1355, w_102_1358, w_102_1362, w_102_1363, w_102_1364, w_102_1365, w_102_1368, w_102_1370, w_102_1371, w_102_1373, w_102_1374, w_102_1375, w_102_1376, w_102_1377, w_102_1379, w_102_1380, w_102_1381, w_102_1382, w_102_1384, w_102_1387, w_102_1388, w_102_1389, w_102_1391, w_102_1392, w_102_1394, w_102_1395, w_102_1397, w_102_1398, w_102_1400, w_102_1401, w_102_1406, w_102_1407, w_102_1410, w_102_1411, w_102_1415, w_102_1416, w_102_1418, w_102_1420, w_102_1422, w_102_1423, w_102_1424, w_102_1425, w_102_1426, w_102_1427, w_102_1428, w_102_1431, w_102_1433, w_102_1435, w_102_1436, w_102_1437, w_102_1438, w_102_1439, w_102_1440, w_102_1442, w_102_1443, w_102_1444, w_102_1445, w_102_1448, w_102_1449, w_102_1450, w_102_1452, w_102_1455, w_102_1457, w_102_1458, w_102_1459, w_102_1461, w_102_1462, w_102_1463, w_102_1464, w_102_1466, w_102_1469, w_102_1471, w_102_1472, w_102_1473, w_102_1474, w_102_1475, w_102_1477, w_102_1479, w_102_1481, w_102_1482, w_102_1483, w_102_1485, w_102_1486, w_102_1489, w_102_1492, w_102_1494, w_102_1495, w_102_1497, w_102_1498, w_102_1500, w_102_1501, w_102_1503, w_102_1504, w_102_1505, w_102_1506, w_102_1509, w_102_1513, w_102_1514, w_102_1515, w_102_1519, w_102_1521, w_102_1522, w_102_1524, w_102_1526, w_102_1527, w_102_1528, w_102_1529, w_102_1530, w_102_1533, w_102_1535, w_102_1539, w_102_1540, w_102_1542, w_102_1543, w_102_1544, w_102_1547, w_102_1549, w_102_1553, w_102_1556, w_102_1557, w_102_1558, w_102_1559, w_102_1561, w_102_1562, w_102_1563, w_102_1564, w_102_1565, w_102_1567, w_102_1571, w_102_1572, w_102_1573, w_102_1574, w_102_1575, w_102_1576, w_102_1577, w_102_1578, w_102_1579, w_102_1582, w_102_1583, w_102_1585, w_102_1586, w_102_1589, w_102_1590, w_102_1593, w_102_1594, w_102_1595, w_102_1598, w_102_1599, w_102_1600, w_102_1601, w_102_1602, w_102_1603, w_102_1604, w_102_1605, w_102_1607, w_102_1608, w_102_1609, w_102_1610, w_102_1613, w_102_1614, w_102_1615, w_102_1616, w_102_1617, w_102_1621, w_102_1622, w_102_1624, w_102_1625, w_102_1627, w_102_1629, w_102_1630, w_102_1633, w_102_1634, w_102_1635, w_102_1637, w_102_1638, w_102_1640, w_102_1641, w_102_1642, w_102_1645, w_102_1646, w_102_1647, w_102_1648, w_102_1649, w_102_1650, w_102_1652, w_102_1653, w_102_1654, w_102_1656, w_102_1657, w_102_1658, w_102_1659, w_102_1660, w_102_1662, w_102_1663, w_102_1665, w_102_1666, w_102_1668, w_102_1670, w_102_1671, w_102_1672, w_102_1673, w_102_1674, w_102_1678, w_102_1679, w_102_1680, w_102_1681, w_102_1682, w_102_1683, w_102_1684, w_102_1685, w_102_1687, w_102_1689, w_102_1690, w_102_1693, w_102_1695, w_102_1700, w_102_1702, w_102_1703, w_102_1704, w_102_1705, w_102_1706, w_102_1707, w_102_1708, w_102_1709, w_102_1712, w_102_1713, w_102_1715, w_102_1716, w_102_1717, w_102_1719, w_102_1721, w_102_1722, w_102_1725, w_102_1727, w_102_1728, w_102_1729, w_102_1730, w_102_1731, w_102_1732, w_102_1734, w_102_1735, w_102_1737, w_102_1738, w_102_1739, w_102_1740, w_102_1741, w_102_1742, w_102_1743, w_102_1744, w_102_1745, w_102_1747, w_102_1748, w_102_1749, w_102_1750, w_102_1754, w_102_1756, w_102_1757, w_102_1759, w_102_1761, w_102_1762, w_102_1763, w_102_1764, w_102_1766, w_102_1767, w_102_1768, w_102_1769, w_102_1772, w_102_1773, w_102_1775, w_102_1776, w_102_1777, w_102_1779, w_102_1781, w_102_1783, w_102_1785, w_102_1787, w_102_1788, w_102_1790, w_102_1791, w_102_1792, w_102_1793, w_102_1794, w_102_1797, w_102_1798, w_102_1800, w_102_1801, w_102_1803, w_102_1805, w_102_1806, w_102_1807, w_102_1808, w_102_1809, w_102_1810, w_102_1811, w_102_1812, w_102_1813, w_102_1816, w_102_1817, w_102_1818, w_102_1822, w_102_1823, w_102_1824, w_102_1825, w_102_1828, w_102_1829, w_102_1831, w_102_1832, w_102_1833, w_102_1834, w_102_1839, w_102_1843, w_102_1846, w_102_1848, w_102_1849, w_102_1850, w_102_1852, w_102_1853, w_102_1855, w_102_1856, w_102_1857, w_102_1860, w_102_1861, w_102_1862, w_102_1863, w_102_1864, w_102_1865, w_102_1867, w_102_1868, w_102_1869, w_102_1870, w_102_1872, w_102_1873, w_102_1874, w_102_1875, w_102_1876, w_102_1877, w_102_1878, w_102_1879, w_102_1880, w_102_1881, w_102_1883, w_102_1885, w_102_1886, w_102_1888, w_102_1889, w_102_1890, w_102_1892, w_102_1894, w_102_1897, w_102_1898, w_102_1899, w_102_1902, w_102_1903, w_102_1904, w_102_1905, w_102_1906, w_102_1908, w_102_1909, w_102_1910, w_102_1911, w_102_1912, w_102_1913, w_102_1914, w_102_1916, w_102_1919, w_102_1920, w_102_1921, w_102_1922, w_102_1923, w_102_1924, w_102_1926, w_102_1930, w_102_1931, w_102_1932, w_102_1933, w_102_1934, w_102_1935, w_102_1936, w_102_1937, w_102_1938, w_102_1942, w_102_1943, w_102_1946, w_102_1947, w_102_1948, w_102_1950, w_102_1952, w_102_1954, w_102_1955, w_102_1956, w_102_1957, w_102_1960, w_102_1961, w_102_1962, w_102_1963, w_102_1964, w_102_1965, w_102_1967, w_102_1968, w_102_1969, w_102_1972, w_102_1973, w_102_1975, w_102_1979, w_102_1980, w_102_1983, w_102_1984, w_102_1985, w_102_1986, w_102_1988, w_102_1990, w_102_1992, w_102_1993, w_102_1996, w_102_1999, w_102_2000, w_102_2001, w_102_2003, w_102_2005, w_102_2006, w_102_2007, w_102_2008, w_102_2012, w_102_2013, w_102_2014, w_102_2015, w_102_2016, w_102_2017, w_102_2018, w_102_2019, w_102_2020, w_102_2023, w_102_2024, w_102_2026, w_102_2027, w_102_2029, w_102_2030, w_102_2031, w_102_2033, w_102_2034, w_102_2035, w_102_2036, w_102_2038, w_102_2040, w_102_2043, w_102_2044, w_102_2045, w_102_2046, w_102_2048, w_102_2049, w_102_2050, w_102_2052, w_102_2053, w_102_2058, w_102_2059, w_102_2061, w_102_2066, w_102_2067, w_102_2068, w_102_2069, w_102_2070, w_102_2071, w_102_2073, w_102_2074, w_102_2075, w_102_2076, w_102_2078, w_102_2081, w_102_2084, w_102_2085, w_102_2086, w_102_2088, w_102_2089, w_102_2090, w_102_2092, w_102_2093, w_102_2094, w_102_2095, w_102_2096, w_102_2099, w_102_2100, w_102_2105, w_102_2106, w_102_2107, w_102_2109, w_102_2111, w_102_2113, w_102_2114, w_102_2115, w_102_2116, w_102_2118, w_102_2119, w_102_2120, w_102_2121, w_102_2122, w_102_2123, w_102_2124, w_102_2125, w_102_2126, w_102_2128, w_102_2129, w_102_2130, w_102_2132, w_102_2133, w_102_2136, w_102_2137, w_102_2138, w_102_2140, w_102_2141, w_102_2144, w_102_2147, w_102_2148, w_102_2149, w_102_2151, w_102_2152, w_102_2153, w_102_2154, w_102_2155, w_102_2158, w_102_2159, w_102_2161, w_102_2163, w_102_2164, w_102_2166, w_102_2167, w_102_2168, w_102_2170, w_102_2171, w_102_2175, w_102_2176, w_102_2177, w_102_2178, w_102_2179, w_102_2180, w_102_2181, w_102_2183, w_102_2185, w_102_2187, w_102_2188, w_102_2189, w_102_2190, w_102_2195, w_102_2196, w_102_2197, w_102_2199, w_102_2203, w_102_2204, w_102_2206, w_102_2209, w_102_2210, w_102_2212, w_102_2213, w_102_2214, w_102_2215, w_102_2217, w_102_2218, w_102_2220, w_102_2221, w_102_2222, w_102_2225, w_102_2226, w_102_2230, w_102_2231, w_102_2232, w_102_2233, w_102_2234, w_102_2235, w_102_2236, w_102_2237, w_102_2238, w_102_2239, w_102_2240, w_102_2241, w_102_2242, w_102_2243, w_102_2244, w_102_2246, w_102_2247, w_102_2251, w_102_2252, w_102_2253, w_102_2255, w_102_2256, w_102_2258, w_102_2259, w_102_2260, w_102_2261, w_102_2264, w_102_2266, w_102_2267, w_102_2269, w_102_2271, w_102_2272, w_102_2273, w_102_2274, w_102_2276, w_102_2278, w_102_2279, w_102_2280, w_102_2282, w_102_2283, w_102_2284, w_102_2285, w_102_2286, w_102_2288, w_102_2289, w_102_2290, w_102_2292, w_102_2295, w_102_2296, w_102_2297, w_102_2298, w_102_2300, w_102_2305, w_102_2308, w_102_2313, w_102_2314, w_102_2315, w_102_2317, w_102_2319, w_102_2320, w_102_2322, w_102_2323, w_102_2326, w_102_2327, w_102_2328, w_102_2329, w_102_2333, w_102_2334, w_102_2338, w_102_2341, w_102_2342, w_102_2344, w_102_2345, w_102_2347, w_102_2348, w_102_2349, w_102_2352, w_102_2354, w_102_2356, w_102_2357, w_102_2359, w_102_2360, w_102_2361, w_102_2362, w_102_2363, w_102_2366, w_102_2367, w_102_2368, w_102_2369, w_102_2370, w_102_2373, w_102_2374, w_102_2375, w_102_2377, w_102_2378, w_102_2379, w_102_2380, w_102_2382, w_102_2383, w_102_2384, w_102_2385, w_102_2386, w_102_2387, w_102_2388, w_102_2391, w_102_2392, w_102_2394, w_102_2395, w_102_2396, w_102_2398, w_102_2399, w_102_2400, w_102_2402, w_102_2403, w_102_2404;
  wire w_103_000, w_103_001, w_103_002, w_103_003, w_103_004, w_103_005, w_103_006, w_103_007, w_103_008, w_103_009, w_103_011, w_103_012, w_103_013, w_103_014, w_103_015, w_103_016, w_103_017, w_103_018, w_103_019, w_103_020, w_103_021, w_103_022, w_103_023, w_103_024, w_103_025, w_103_026, w_103_027, w_103_028, w_103_029, w_103_030, w_103_031, w_103_032, w_103_033, w_103_034, w_103_035, w_103_036, w_103_037, w_103_038, w_103_039, w_103_040, w_103_041, w_103_042, w_103_043, w_103_044, w_103_045, w_103_046, w_103_047, w_103_048, w_103_049, w_103_050, w_103_051, w_103_052, w_103_053, w_103_054, w_103_055, w_103_056, w_103_057, w_103_058, w_103_059, w_103_060, w_103_061, w_103_062, w_103_063, w_103_064, w_103_065, w_103_066, w_103_067, w_103_068, w_103_069, w_103_070, w_103_071, w_103_072, w_103_073, w_103_074, w_103_075, w_103_076, w_103_077, w_103_078, w_103_079, w_103_080, w_103_081, w_103_082, w_103_083, w_103_084, w_103_085, w_103_086, w_103_087, w_103_089, w_103_090, w_103_091, w_103_092, w_103_093, w_103_094, w_103_095, w_103_096, w_103_097, w_103_098, w_103_099, w_103_100, w_103_101, w_103_102, w_103_103, w_103_104, w_103_105, w_103_106, w_103_107, w_103_108, w_103_109, w_103_110, w_103_111, w_103_112, w_103_114, w_103_115, w_103_116, w_103_117, w_103_118, w_103_119, w_103_120, w_103_121, w_103_122, w_103_123, w_103_124, w_103_125, w_103_126, w_103_127, w_103_128, w_103_129, w_103_130, w_103_131, w_103_132, w_103_133, w_103_134, w_103_135, w_103_137, w_103_138, w_103_139, w_103_140, w_103_141, w_103_142, w_103_143, w_103_144, w_103_145, w_103_146, w_103_147, w_103_148, w_103_149, w_103_150, w_103_151, w_103_152, w_103_153, w_103_154, w_103_155, w_103_156, w_103_157, w_103_158, w_103_159, w_103_160, w_103_161, w_103_163, w_103_164, w_103_165, w_103_166, w_103_167, w_103_168, w_103_169, w_103_170, w_103_172, w_103_174, w_103_175, w_103_176, w_103_177, w_103_179, w_103_180, w_103_181, w_103_182, w_103_183, w_103_184, w_103_185, w_103_186, w_103_187, w_103_189, w_103_190, w_103_191, w_103_193, w_103_194, w_103_195, w_103_196, w_103_197, w_103_198, w_103_199, w_103_200, w_103_201, w_103_202, w_103_203, w_103_205, w_103_206, w_103_207, w_103_208, w_103_209, w_103_210, w_103_211, w_103_212, w_103_213, w_103_214, w_103_215, w_103_216, w_103_217, w_103_218, w_103_219, w_103_220, w_103_221, w_103_222, w_103_223, w_103_224, w_103_225, w_103_226, w_103_227, w_103_228, w_103_229, w_103_230, w_103_231, w_103_232, w_103_233, w_103_234, w_103_235, w_103_236, w_103_237, w_103_238, w_103_239, w_103_240, w_103_241, w_103_242, w_103_243, w_103_244, w_103_245, w_103_246, w_103_247, w_103_248, w_103_249, w_103_250, w_103_251, w_103_252, w_103_253, w_103_254, w_103_255, w_103_257, w_103_258, w_103_259, w_103_260, w_103_261, w_103_262, w_103_263, w_103_264, w_103_265, w_103_266, w_103_268, w_103_269, w_103_270, w_103_271, w_103_272, w_103_273, w_103_274, w_103_275, w_103_276, w_103_277, w_103_278, w_103_279, w_103_280, w_103_281, w_103_283, w_103_284, w_103_285, w_103_286, w_103_287, w_103_288, w_103_289, w_103_290, w_103_292, w_103_294, w_103_295, w_103_297, w_103_298, w_103_299, w_103_300, w_103_301, w_103_302, w_103_303, w_103_304, w_103_305, w_103_306, w_103_307, w_103_308, w_103_309, w_103_310, w_103_311, w_103_312, w_103_313, w_103_314, w_103_315, w_103_316, w_103_317, w_103_318, w_103_319, w_103_321, w_103_322, w_103_323, w_103_324, w_103_325, w_103_326, w_103_327, w_103_328, w_103_329, w_103_330, w_103_331, w_103_332, w_103_333, w_103_334, w_103_335, w_103_337, w_103_338, w_103_339, w_103_340, w_103_341, w_103_342, w_103_343, w_103_344, w_103_345, w_103_346, w_103_347, w_103_348, w_103_349, w_103_350, w_103_351, w_103_352, w_103_353, w_103_354, w_103_356, w_103_357, w_103_358, w_103_359, w_103_360, w_103_361, w_103_362, w_103_363, w_103_364, w_103_365, w_103_366, w_103_367, w_103_368, w_103_369, w_103_370, w_103_371, w_103_372, w_103_373, w_103_374, w_103_375, w_103_376, w_103_377, w_103_378, w_103_379, w_103_380, w_103_381, w_103_383, w_103_384, w_103_385, w_103_386, w_103_387, w_103_388, w_103_389, w_103_390, w_103_391, w_103_392, w_103_394, w_103_395, w_103_396, w_103_397, w_103_398, w_103_399, w_103_400, w_103_401, w_103_402, w_103_403, w_103_404, w_103_405, w_103_406, w_103_407, w_103_408, w_103_409, w_103_410, w_103_411, w_103_412, w_103_413, w_103_414, w_103_415, w_103_416, w_103_417, w_103_418, w_103_419, w_103_420, w_103_421, w_103_422, w_103_423, w_103_424, w_103_425, w_103_427, w_103_428, w_103_429, w_103_430, w_103_431, w_103_432, w_103_433, w_103_434, w_103_435, w_103_436, w_103_437, w_103_438, w_103_439, w_103_440, w_103_441, w_103_442, w_103_443, w_103_444, w_103_445, w_103_446, w_103_447, w_103_449, w_103_450, w_103_451, w_103_453, w_103_454, w_103_455, w_103_456, w_103_457, w_103_458, w_103_459, w_103_460, w_103_461, w_103_462, w_103_463, w_103_464, w_103_465, w_103_466, w_103_467, w_103_469, w_103_470, w_103_471, w_103_472, w_103_473, w_103_474, w_103_475, w_103_476, w_103_477, w_103_478, w_103_479, w_103_481, w_103_482, w_103_483, w_103_485, w_103_486, w_103_487, w_103_488, w_103_489, w_103_490, w_103_491, w_103_492, w_103_493, w_103_494, w_103_496, w_103_497, w_103_499, w_103_500, w_103_501, w_103_502, w_103_503, w_103_504, w_103_505, w_103_506, w_103_507, w_103_508, w_103_509, w_103_510, w_103_511, w_103_512, w_103_513, w_103_514, w_103_515, w_103_516, w_103_517, w_103_518, w_103_519, w_103_520, w_103_521, w_103_522, w_103_523, w_103_524, w_103_525, w_103_526, w_103_527, w_103_528, w_103_529, w_103_530, w_103_531, w_103_532, w_103_533, w_103_534, w_103_535, w_103_536, w_103_537, w_103_538, w_103_539, w_103_540, w_103_541, w_103_542, w_103_543, w_103_544, w_103_545, w_103_546, w_103_547, w_103_548, w_103_549, w_103_550, w_103_551, w_103_552, w_103_553, w_103_554, w_103_555, w_103_556, w_103_557, w_103_558, w_103_559, w_103_560, w_103_561, w_103_562, w_103_563, w_103_564, w_103_565, w_103_566, w_103_568, w_103_569, w_103_570, w_103_571, w_103_572, w_103_573, w_103_574, w_103_575, w_103_576, w_103_577, w_103_579, w_103_580, w_103_581, w_103_582, w_103_583, w_103_585, w_103_587, w_103_588, w_103_589, w_103_590, w_103_591, w_103_592, w_103_593, w_103_594, w_103_595, w_103_596, w_103_597, w_103_598, w_103_599, w_103_600, w_103_601, w_103_603, w_103_604, w_103_605, w_103_606, w_103_607, w_103_608, w_103_609, w_103_610, w_103_611, w_103_612, w_103_613, w_103_614, w_103_615, w_103_616, w_103_617, w_103_618, w_103_619, w_103_620, w_103_621, w_103_622, w_103_623, w_103_624, w_103_625, w_103_626, w_103_628, w_103_629, w_103_630, w_103_631, w_103_632, w_103_635, w_103_636, w_103_637, w_103_638, w_103_639, w_103_640, w_103_641, w_103_642, w_103_643, w_103_644, w_103_645, w_103_646, w_103_647, w_103_648, w_103_649, w_103_650, w_103_651, w_103_652, w_103_653, w_103_654, w_103_655, w_103_657, w_103_658, w_103_660, w_103_661, w_103_662, w_103_663, w_103_664, w_103_665, w_103_666, w_103_667, w_103_668, w_103_669, w_103_670, w_103_671, w_103_672, w_103_674, w_103_675, w_103_676, w_103_678, w_103_679, w_103_680, w_103_681, w_103_682, w_103_683, w_103_684, w_103_685, w_103_686, w_103_687, w_103_688, w_103_689, w_103_690, w_103_691, w_103_692, w_103_693, w_103_694, w_103_695, w_103_696, w_103_697, w_103_698, w_103_699, w_103_700, w_103_701, w_103_702, w_103_703, w_103_704, w_103_705, w_103_706, w_103_707, w_103_708, w_103_709, w_103_710, w_103_711, w_103_712, w_103_713, w_103_714, w_103_715, w_103_716, w_103_717, w_103_718, w_103_719, w_103_720, w_103_721, w_103_722, w_103_723, w_103_724, w_103_725, w_103_726, w_103_727, w_103_728, w_103_729, w_103_730, w_103_731, w_103_733, w_103_734, w_103_735, w_103_736, w_103_737, w_103_738, w_103_739, w_103_740, w_103_741, w_103_742, w_103_743, w_103_744, w_103_745, w_103_746, w_103_747, w_103_748, w_103_749, w_103_750, w_103_751, w_103_752, w_103_753, w_103_754, w_103_756, w_103_757, w_103_758, w_103_759, w_103_760, w_103_761, w_103_762, w_103_763, w_103_764, w_103_765, w_103_766, w_103_767, w_103_768, w_103_769, w_103_770, w_103_771, w_103_772, w_103_773, w_103_774, w_103_775, w_103_776, w_103_777, w_103_778, w_103_779, w_103_780, w_103_781, w_103_782, w_103_783, w_103_784, w_103_785, w_103_786, w_103_787, w_103_788, w_103_789, w_103_790, w_103_792, w_103_793, w_103_794, w_103_795, w_103_796, w_103_797, w_103_798, w_103_799, w_103_800, w_103_801, w_103_802, w_103_803, w_103_804, w_103_805, w_103_806, w_103_807, w_103_808, w_103_809, w_103_810, w_103_811, w_103_812, w_103_813, w_103_814, w_103_815, w_103_816, w_103_817, w_103_818, w_103_819, w_103_820, w_103_822, w_103_823, w_103_824, w_103_825, w_103_826, w_103_827;
  wire w_104_001, w_104_003, w_104_004, w_104_005, w_104_007, w_104_008, w_104_011, w_104_013, w_104_015, w_104_016, w_104_018, w_104_019, w_104_020, w_104_021, w_104_022, w_104_023, w_104_024, w_104_026, w_104_028, w_104_029, w_104_030, w_104_031, w_104_033, w_104_034, w_104_036, w_104_038, w_104_039, w_104_040, w_104_041, w_104_042, w_104_046, w_104_048, w_104_049, w_104_050, w_104_051, w_104_052, w_104_053, w_104_054, w_104_056, w_104_059, w_104_061, w_104_063, w_104_064, w_104_065, w_104_066, w_104_070, w_104_071, w_104_073, w_104_075, w_104_076, w_104_078, w_104_080, w_104_082, w_104_083, w_104_085, w_104_087, w_104_088, w_104_090, w_104_091, w_104_092, w_104_093, w_104_094, w_104_095, w_104_096, w_104_097, w_104_098, w_104_100, w_104_102, w_104_103, w_104_105, w_104_106, w_104_108, w_104_111, w_104_112, w_104_114, w_104_116, w_104_118, w_104_119, w_104_122, w_104_124, w_104_125, w_104_126, w_104_127, w_104_128, w_104_129, w_104_130, w_104_131, w_104_132, w_104_134, w_104_135, w_104_137, w_104_139, w_104_141, w_104_142, w_104_143, w_104_144, w_104_145, w_104_147, w_104_148, w_104_149, w_104_150, w_104_151, w_104_156, w_104_157, w_104_158, w_104_159, w_104_160, w_104_162, w_104_163, w_104_164, w_104_165, w_104_166, w_104_168, w_104_169, w_104_171, w_104_173, w_104_174, w_104_175, w_104_176, w_104_181, w_104_183, w_104_185, w_104_186, w_104_187, w_104_188, w_104_189, w_104_190, w_104_191, w_104_192, w_104_193, w_104_194, w_104_195, w_104_197, w_104_198, w_104_200, w_104_201, w_104_202, w_104_203, w_104_204, w_104_205, w_104_208, w_104_209, w_104_210, w_104_212, w_104_213, w_104_214, w_104_216, w_104_217, w_104_219, w_104_221, w_104_222, w_104_223, w_104_225, w_104_226, w_104_227, w_104_229, w_104_231, w_104_232, w_104_234, w_104_235, w_104_238, w_104_239, w_104_240, w_104_241, w_104_242, w_104_244, w_104_248, w_104_251, w_104_252, w_104_255, w_104_256, w_104_258, w_104_260, w_104_262, w_104_263, w_104_264, w_104_265, w_104_266, w_104_268, w_104_270, w_104_272, w_104_273, w_104_274, w_104_276, w_104_278, w_104_279, w_104_281, w_104_284, w_104_285, w_104_286, w_104_287, w_104_289, w_104_290, w_104_291, w_104_294, w_104_296, w_104_299, w_104_300, w_104_301, w_104_302, w_104_303, w_104_306, w_104_307, w_104_308, w_104_310, w_104_312, w_104_313, w_104_314, w_104_317, w_104_318, w_104_321, w_104_322, w_104_323, w_104_326, w_104_328, w_104_330, w_104_332, w_104_333, w_104_335, w_104_336, w_104_338, w_104_340, w_104_342, w_104_343, w_104_344, w_104_345, w_104_346, w_104_348, w_104_350, w_104_353, w_104_354, w_104_356, w_104_357, w_104_358, w_104_360, w_104_361, w_104_362, w_104_363, w_104_364, w_104_365, w_104_366, w_104_368, w_104_370, w_104_371, w_104_373, w_104_376, w_104_378, w_104_381, w_104_382, w_104_383, w_104_385, w_104_386, w_104_387, w_104_388, w_104_389, w_104_390, w_104_391, w_104_392, w_104_393, w_104_395, w_104_396, w_104_397, w_104_398, w_104_400, w_104_401, w_104_402, w_104_403, w_104_404, w_104_406, w_104_407, w_104_408, w_104_409, w_104_410, w_104_411, w_104_412, w_104_414, w_104_415, w_104_419, w_104_423, w_104_425, w_104_426, w_104_428, w_104_429, w_104_431, w_104_433, w_104_434, w_104_435, w_104_439, w_104_442, w_104_443, w_104_446, w_104_447, w_104_448, w_104_450, w_104_452, w_104_453, w_104_454, w_104_455, w_104_459, w_104_460, w_104_462, w_104_463, w_104_465, w_104_466, w_104_467, w_104_470, w_104_471, w_104_473, w_104_475, w_104_476, w_104_477, w_104_480, w_104_482, w_104_485, w_104_486, w_104_487, w_104_488, w_104_489, w_104_491, w_104_493, w_104_496, w_104_498, w_104_499, w_104_500, w_104_501, w_104_502, w_104_505, w_104_506, w_104_507, w_104_509, w_104_510, w_104_512, w_104_513, w_104_517, w_104_520, w_104_521, w_104_523, w_104_533, w_104_536, w_104_539, w_104_540, w_104_541, w_104_545, w_104_546, w_104_548, w_104_550, w_104_552, w_104_553, w_104_558, w_104_559, w_104_561, w_104_562, w_104_563, w_104_564, w_104_565, w_104_566, w_104_567, w_104_570, w_104_571, w_104_572, w_104_574, w_104_575, w_104_577, w_104_579, w_104_581, w_104_582, w_104_583, w_104_585, w_104_586, w_104_587, w_104_589, w_104_590, w_104_592, w_104_594, w_104_595, w_104_598, w_104_600, w_104_602, w_104_603, w_104_604, w_104_607, w_104_610, w_104_612, w_104_613, w_104_618, w_104_619, w_104_620, w_104_622, w_104_624, w_104_625, w_104_626, w_104_627, w_104_628, w_104_630, w_104_632, w_104_633, w_104_635, w_104_637, w_104_638, w_104_639, w_104_640, w_104_641, w_104_642, w_104_645, w_104_648, w_104_649, w_104_652, w_104_655, w_104_657, w_104_658, w_104_659, w_104_660, w_104_661, w_104_662, w_104_665, w_104_666, w_104_667, w_104_668, w_104_669, w_104_673, w_104_674, w_104_679, w_104_684, w_104_685, w_104_687, w_104_689, w_104_690, w_104_692, w_104_693, w_104_695, w_104_696, w_104_697, w_104_699, w_104_700, w_104_704, w_104_705, w_104_706, w_104_707, w_104_708, w_104_709, w_104_711, w_104_712, w_104_713, w_104_714, w_104_715, w_104_716, w_104_717, w_104_718, w_104_719, w_104_720, w_104_723, w_104_725, w_104_726, w_104_727, w_104_728, w_104_730, w_104_732, w_104_733, w_104_734, w_104_735, w_104_736, w_104_737, w_104_738, w_104_739, w_104_740, w_104_741, w_104_742, w_104_744, w_104_745, w_104_753, w_104_755, w_104_756, w_104_757, w_104_759, w_104_762, w_104_764, w_104_771, w_104_772, w_104_773, w_104_774, w_104_776, w_104_778, w_104_779, w_104_780, w_104_781, w_104_783, w_104_784, w_104_785, w_104_788, w_104_790, w_104_792, w_104_794, w_104_795, w_104_796, w_104_800, w_104_802, w_104_803, w_104_804, w_104_807, w_104_809, w_104_811, w_104_812, w_104_813, w_104_814, w_104_816, w_104_819, w_104_821, w_104_824, w_104_825, w_104_827, w_104_829, w_104_831, w_104_832, w_104_833, w_104_835, w_104_836, w_104_837, w_104_838, w_104_840, w_104_842, w_104_845, w_104_846, w_104_848, w_104_853, w_104_854, w_104_855, w_104_858, w_104_859, w_104_860, w_104_861, w_104_862, w_104_863, w_104_864, w_104_868, w_104_869, w_104_870, w_104_871, w_104_873, w_104_874, w_104_875, w_104_877, w_104_880, w_104_881, w_104_885, w_104_886, w_104_888, w_104_889, w_104_890, w_104_891, w_104_892, w_104_893, w_104_895, w_104_897, w_104_898, w_104_899, w_104_902, w_104_903, w_104_904, w_104_906, w_104_907, w_104_908, w_104_910, w_104_911, w_104_914, w_104_915, w_104_918, w_104_919, w_104_921, w_104_923, w_104_925, w_104_926, w_104_927, w_104_928, w_104_930, w_104_932, w_104_934, w_104_935, w_104_936, w_104_940, w_104_942, w_104_943, w_104_944, w_104_945, w_104_946, w_104_947, w_104_948, w_104_950, w_104_951, w_104_952, w_104_955, w_104_957, w_104_959, w_104_962, w_104_964, w_104_966, w_104_967, w_104_968, w_104_969, w_104_972, w_104_979, w_104_980, w_104_981, w_104_983, w_104_984, w_104_985, w_104_986, w_104_987, w_104_988, w_104_989, w_104_991, w_104_992, w_104_993, w_104_995, w_104_998, w_104_999, w_104_1003, w_104_1004, w_104_1007, w_104_1010, w_104_1011, w_104_1012, w_104_1015, w_104_1017, w_104_1020, w_104_1021, w_104_1023, w_104_1024, w_104_1029, w_104_1031, w_104_1032, w_104_1035, w_104_1036, w_104_1037, w_104_1038, w_104_1039, w_104_1042, w_104_1043, w_104_1045, w_104_1046, w_104_1050, w_104_1051, w_104_1052, w_104_1053, w_104_1057, w_104_1059, w_104_1060, w_104_1062, w_104_1064, w_104_1065, w_104_1066, w_104_1068, w_104_1069, w_104_1071, w_104_1072, w_104_1073, w_104_1074, w_104_1075, w_104_1077, w_104_1078, w_104_1079, w_104_1080, w_104_1081, w_104_1082, w_104_1083, w_104_1084, w_104_1088, w_104_1089, w_104_1090, w_104_1094, w_104_1096, w_104_1097, w_104_1098, w_104_1099, w_104_1102, w_104_1103, w_104_1107, w_104_1108, w_104_1109, w_104_1110, w_104_1112, w_104_1113, w_104_1115, w_104_1117, w_104_1118, w_104_1119, w_104_1120, w_104_1121, w_104_1126, w_104_1127, w_104_1128, w_104_1130, w_104_1131, w_104_1132, w_104_1133, w_104_1135, w_104_1138, w_104_1139, w_104_1140, w_104_1141, w_104_1143, w_104_1144, w_104_1147, w_104_1150, w_104_1152, w_104_1153, w_104_1154, w_104_1155, w_104_1157, w_104_1163, w_104_1166, w_104_1170, w_104_1171, w_104_1172, w_104_1173, w_104_1176, w_104_1177, w_104_1178, w_104_1181, w_104_1182, w_104_1183, w_104_1184, w_104_1185, w_104_1187, w_104_1188, w_104_1191, w_104_1192, w_104_1193, w_104_1194, w_104_1197, w_104_1198, w_104_1199, w_104_1203, w_104_1204, w_104_1206, w_104_1207, w_104_1208, w_104_1211, w_104_1214, w_104_1215, w_104_1216, w_104_1218, w_104_1219, w_104_1220, w_104_1221, w_104_1222, w_104_1223, w_104_1225, w_104_1226, w_104_1227, w_104_1228, w_104_1230, w_104_1232, w_104_1233, w_104_1235, w_104_1237, w_104_1238, w_104_1239, w_104_1241, w_104_1242, w_104_1243, w_104_1244, w_104_1245, w_104_1246, w_104_1247, w_104_1248, w_104_1249, w_104_1251, w_104_1252, w_104_1253, w_104_1256, w_104_1257, w_104_1258, w_104_1259, w_104_1260, w_104_1261, w_104_1262, w_104_1263, w_104_1265, w_104_1267, w_104_1268, w_104_1269, w_104_1271, w_104_1272, w_104_1273, w_104_1275, w_104_1276, w_104_1277, w_104_1278, w_104_1279, w_104_1282, w_104_1283, w_104_1285, w_104_1292, w_104_1293, w_104_1294, w_104_1298, w_104_1299, w_104_1300, w_104_1302, w_104_1303, w_104_1304, w_104_1306, w_104_1307, w_104_1308, w_104_1309, w_104_1314, w_104_1315, w_104_1316, w_104_1317, w_104_1320, w_104_1321, w_104_1326, w_104_1329, w_104_1330, w_104_1331, w_104_1332, w_104_1334, w_104_1337, w_104_1338, w_104_1340, w_104_1341, w_104_1342, w_104_1343, w_104_1344, w_104_1350, w_104_1351, w_104_1352, w_104_1354, w_104_1358, w_104_1359, w_104_1362, w_104_1364, w_104_1365, w_104_1366, w_104_1369, w_104_1370, w_104_1373, w_104_1374, w_104_1376, w_104_1377, w_104_1378, w_104_1380, w_104_1382, w_104_1384, w_104_1386, w_104_1387, w_104_1389, w_104_1390, w_104_1391, w_104_1392, w_104_1394, w_104_1396, w_104_1397, w_104_1399, w_104_1403, w_104_1406, w_104_1407, w_104_1411, w_104_1415, w_104_1416, w_104_1418, w_104_1419, w_104_1421, w_104_1423, w_104_1424, w_104_1428, w_104_1434, w_104_1435, w_104_1439, w_104_1440, w_104_1441, w_104_1442, w_104_1443, w_104_1445, w_104_1447, w_104_1448, w_104_1449, w_104_1450, w_104_1451, w_104_1453, w_104_1454, w_104_1455, w_104_1456, w_104_1457, w_104_1459, w_104_1460, w_104_1461, w_104_1463, w_104_1466, w_104_1469, w_104_1470, w_104_1471, w_104_1472, w_104_1474, w_104_1475, w_104_1476, w_104_1479, w_104_1480, w_104_1481, w_104_1483, w_104_1484, w_104_1485, w_104_1487, w_104_1488, w_104_1489, w_104_1490, w_104_1491, w_104_1493, w_104_1494, w_104_1495, w_104_1499, w_104_1500, w_104_1504, w_104_1505, w_104_1506, w_104_1508, w_104_1509, w_104_1511, w_104_1514, w_104_1516, w_104_1518, w_104_1522, w_104_1523, w_104_1524, w_104_1525, w_104_1526, w_104_1527, w_104_1528, w_104_1530, w_104_1531, w_104_1533, w_104_1534, w_104_1537, w_104_1539, w_104_1540, w_104_1541, w_104_1542, w_104_1544, w_104_1547, w_104_1548, w_104_1550, w_104_1551, w_104_1552, w_104_1553, w_104_1554, w_104_1557, w_104_1558, w_104_1559, w_104_1560, w_104_1561, w_104_1562, w_104_1563, w_104_1564, w_104_1565, w_104_1567, w_104_1569, w_104_1572, w_104_1573, w_104_1574, w_104_1575, w_104_1576, w_104_1578, w_104_1579, w_104_1581, w_104_1582, w_104_1584, w_104_1585, w_104_1587, w_104_1588, w_104_1590, w_104_1591, w_104_1592, w_104_1593, w_104_1595, w_104_1596, w_104_1600, w_104_1601, w_104_1603, w_104_1604, w_104_1607, w_104_1608, w_104_1610, w_104_1611, w_104_1612, w_104_1615, w_104_1616, w_104_1617, w_104_1618, w_104_1619, w_104_1623, w_104_1624, w_104_1629, w_104_1633, w_104_1634, w_104_1635, w_104_1636, w_104_1638, w_104_1640, w_104_1641, w_104_1642, w_104_1643, w_104_1644, w_104_1646, w_104_1648, w_104_1649, w_104_1650, w_104_1651, w_104_1654, w_104_1656, w_104_1657, w_104_1658, w_104_1660, w_104_1661, w_104_1662, w_104_1663, w_104_1664, w_104_1665, w_104_1668, w_104_1670, w_104_1674, w_104_1675, w_104_1676, w_104_1678, w_104_1679, w_104_1680, w_104_1682, w_104_1684, w_104_1685, w_104_1686, w_104_1688, w_104_1690, w_104_1691, w_104_1692, w_104_1696, w_104_1699, w_104_1706, w_104_1710, w_104_1713, w_104_1715, w_104_1716, w_104_1717, w_104_1718, w_104_1719, w_104_1720, w_104_1724, w_104_1725, w_104_1726, w_104_1728, w_104_1729, w_104_1731, w_104_1732, w_104_1733, w_104_1736, w_104_1737, w_104_1739, w_104_1740, w_104_1741, w_104_1745, w_104_1748, w_104_1750, w_104_1751, w_104_1754, w_104_1759, w_104_1761, w_104_1765, w_104_1767, w_104_1775, w_104_1778, w_104_1780, w_104_1782, w_104_1783, w_104_1784, w_104_1786, w_104_1787, w_104_1790, w_104_1792, w_104_1793, w_104_1794, w_104_1795, w_104_1796, w_104_1797, w_104_1798, w_104_1799, w_104_1800, w_104_1801, w_104_1804, w_104_1806, w_104_1807, w_104_1808, w_104_1811, w_104_1812, w_104_1813, w_104_1814, w_104_1815, w_104_1816, w_104_1818, w_104_1819, w_104_1820, w_104_1821, w_104_1823, w_104_1824, w_104_1826, w_104_1828, w_104_1830, w_104_1832, w_104_1833, w_104_1835, w_104_1836, w_104_1837, w_104_1839, w_104_1840, w_104_1841, w_104_1842, w_104_1844, w_104_1845, w_104_1846, w_104_1847, w_104_1848, w_104_1849, w_104_1852, w_104_1853, w_104_1854, w_104_1855, w_104_1857, w_104_1858, w_104_1860, w_104_1861, w_104_1864, w_104_1865, w_104_1866, w_104_1867, w_104_1868, w_104_1870, w_104_1871, w_104_1873, w_104_1874, w_104_1875, w_104_1876, w_104_1878, w_104_1879, w_104_1880, w_104_1881, w_104_1883, w_104_1884, w_104_1885, w_104_1886, w_104_1887, w_104_1888, w_104_1891, w_104_1893, w_104_1894, w_104_1895, w_104_1896, w_104_1897, w_104_1898, w_104_1901, w_104_1904, w_104_1905, w_104_1906, w_104_1908, w_104_1910, w_104_1911, w_104_1912, w_104_1914, w_104_1916, w_104_1918, w_104_1919, w_104_1920, w_104_1921, w_104_1922, w_104_1923, w_104_1925, w_104_1927, w_104_1928, w_104_1929, w_104_1930, w_104_1934, w_104_1935, w_104_1936, w_104_1939, w_104_1940, w_104_1943, w_104_1944, w_104_1945, w_104_1946, w_104_1948, w_104_1949, w_104_1950, w_104_1951, w_104_1952, w_104_1953, w_104_1954, w_104_1955, w_104_1957, w_104_1960, w_104_1962, w_104_1964, w_104_1966, w_104_1970, w_104_1971, w_104_1973, w_104_1974, w_104_1978, w_104_1980, w_104_1981, w_104_1983, w_104_1984, w_104_1985, w_104_1986, w_104_1988, w_104_1989, w_104_1990, w_104_1993, w_104_1996, w_104_1997, w_104_1998, w_104_2001, w_104_2004, w_104_2005, w_104_2006, w_104_2011, w_104_2012, w_104_2013, w_104_2014, w_104_2015, w_104_2016, w_104_2018, w_104_2020, w_104_2023, w_104_2024, w_104_2025, w_104_2026, w_104_2027, w_104_2029, w_104_2030, w_104_2031, w_104_2032, w_104_2033, w_104_2034, w_104_2036, w_104_2039, w_104_2040, w_104_2041, w_104_2043, w_104_2044, w_104_2045, w_104_2046, w_104_2048, w_104_2049, w_104_2050, w_104_2051, w_104_2052, w_104_2053, w_104_2056, w_104_2060, w_104_2061, w_104_2062, w_104_2063, w_104_2064, w_104_2065, w_104_2066, w_104_2068, w_104_2069, w_104_2074, w_104_2075, w_104_2076, w_104_2079, w_104_2080, w_104_2082, w_104_2084, w_104_2085, w_104_2087, w_104_2088, w_104_2090, w_104_2091, w_104_2093, w_104_2094, w_104_2095, w_104_2096, w_104_2097, w_104_2098, w_104_2099, w_104_2101, w_104_2105, w_104_2106, w_104_2107, w_104_2108, w_104_2110, w_104_2112, w_104_2118, w_104_2120, w_104_2122, w_104_2125, w_104_2126, w_104_2129, w_104_2130, w_104_2133, w_104_2135, w_104_2136, w_104_2137, w_104_2140, w_104_2141, w_104_2142, w_104_2145, w_104_2147, w_104_2150, w_104_2151, w_104_2152, w_104_2154, w_104_2156, w_104_2157, w_104_2158, w_104_2160, w_104_2161, w_104_2162, w_104_2165, w_104_2166, w_104_2167, w_104_2168, w_104_2169, w_104_2170, w_104_2171, w_104_2172, w_104_2173, w_104_2176, w_104_2178, w_104_2181, w_104_2183, w_104_2185, w_104_2186, w_104_2187, w_104_2189, w_104_2191, w_104_2192, w_104_2193, w_104_2194, w_104_2195, w_104_2198, w_104_2199, w_104_2200, w_104_2201, w_104_2202, w_104_2203, w_104_2204, w_104_2206, w_104_2212, w_104_2214, w_104_2215, w_104_2216, w_104_2217, w_104_2218, w_104_2222, w_104_2223, w_104_2224, w_104_2226, w_104_2227, w_104_2228, w_104_2229, w_104_2230, w_104_2231, w_104_2232, w_104_2233, w_104_2236, w_104_2237, w_104_2238, w_104_2240, w_104_2241, w_104_2242, w_104_2244, w_104_2245, w_104_2246, w_104_2247, w_104_2248, w_104_2249, w_104_2250, w_104_2251, w_104_2253, w_104_2254, w_104_2256, w_104_2257, w_104_2258, w_104_2259, w_104_2260, w_104_2261, w_104_2263, w_104_2264, w_104_2265, w_104_2268, w_104_2269, w_104_2273, w_104_2275, w_104_2276, w_104_2280, w_104_2281, w_104_2282, w_104_2283, w_104_2284, w_104_2285, w_104_2286, w_104_2287, w_104_2288, w_104_2291, w_104_2292, w_104_2293, w_104_2295, w_104_2296, w_104_2298, w_104_2299, w_104_2300, w_104_2301, w_104_2302, w_104_2303, w_104_2305, w_104_2307, w_104_2308, w_104_2309, w_104_2310, w_104_2312, w_104_2313, w_104_2315, w_104_2317, w_104_2319, w_104_2324, w_104_2325, w_104_2326, w_104_2327, w_104_2328, w_104_2330, w_104_2332, w_104_2334, w_104_2335, w_104_2340, w_104_2343, w_104_2346, w_104_2349, w_104_2351, w_104_2352, w_104_2353, w_104_2355, w_104_2356, w_104_2357, w_104_2358, w_104_2359, w_104_2360, w_104_2361, w_104_2362, w_104_2364, w_104_2366, w_104_2367, w_104_2368, w_104_2369, w_104_2370, w_104_2375, w_104_2376, w_104_2378, w_104_2379, w_104_2381, w_104_2384, w_104_2387, w_104_2389, w_104_2390, w_104_2391, w_104_2392, w_104_2393, w_104_2397, w_104_2398, w_104_2400, w_104_2401, w_104_2403, w_104_2404, w_104_2405, w_104_2408, w_104_2409, w_104_2411, w_104_2412, w_104_2413, w_104_2414, w_104_2419, w_104_2420, w_104_2424, w_104_2427, w_104_2429, w_104_2431, w_104_2432, w_104_2433, w_104_2435, w_104_2436, w_104_2437, w_104_2438, w_104_2441, w_104_2444, w_104_2446, w_104_2447, w_104_2448, w_104_2449, w_104_2450, w_104_2451, w_104_2458, w_104_2461;
  wire w_105_001, w_105_003, w_105_014, w_105_016, w_105_019, w_105_020, w_105_021, w_105_023, w_105_026, w_105_030, w_105_034, w_105_035, w_105_038, w_105_040, w_105_042, w_105_043, w_105_049, w_105_053, w_105_055, w_105_056, w_105_057, w_105_058, w_105_060, w_105_064, w_105_065, w_105_067, w_105_068, w_105_070, w_105_071, w_105_072, w_105_073, w_105_074, w_105_077, w_105_078, w_105_079, w_105_080, w_105_082, w_105_090, w_105_092, w_105_097, w_105_100, w_105_103, w_105_106, w_105_110, w_105_113, w_105_117, w_105_119, w_105_123, w_105_124, w_105_125, w_105_126, w_105_127, w_105_128, w_105_131, w_105_134, w_105_135, w_105_137, w_105_138, w_105_144, w_105_150, w_105_151, w_105_157, w_105_159, w_105_162, w_105_164, w_105_165, w_105_168, w_105_171, w_105_175, w_105_180, w_105_181, w_105_182, w_105_183, w_105_191, w_105_193, w_105_197, w_105_200, w_105_208, w_105_212, w_105_213, w_105_215, w_105_217, w_105_219, w_105_221, w_105_227, w_105_229, w_105_233, w_105_235, w_105_241, w_105_242, w_105_246, w_105_252, w_105_253, w_105_258, w_105_261, w_105_266, w_105_267, w_105_268, w_105_270, w_105_275, w_105_277, w_105_278, w_105_283, w_105_284, w_105_286, w_105_288, w_105_289, w_105_291, w_105_292, w_105_295, w_105_302, w_105_307, w_105_311, w_105_312, w_105_316, w_105_317, w_105_319, w_105_320, w_105_325, w_105_328, w_105_329, w_105_330, w_105_334, w_105_337, w_105_341, w_105_343, w_105_347, w_105_348, w_105_350, w_105_351, w_105_354, w_105_363, w_105_364, w_105_366, w_105_370, w_105_371, w_105_374, w_105_376, w_105_377, w_105_383, w_105_386, w_105_387, w_105_391, w_105_396, w_105_399, w_105_402, w_105_404, w_105_406, w_105_407, w_105_412, w_105_413, w_105_415, w_105_417, w_105_418, w_105_422, w_105_423, w_105_424, w_105_426, w_105_427, w_105_428, w_105_429, w_105_431, w_105_434, w_105_435, w_105_436, w_105_441, w_105_444, w_105_445, w_105_447, w_105_451, w_105_452, w_105_455, w_105_462, w_105_465, w_105_466, w_105_470, w_105_473, w_105_479, w_105_480, w_105_481, w_105_483, w_105_484, w_105_485, w_105_488, w_105_491, w_105_493, w_105_494, w_105_495, w_105_500, w_105_504, w_105_510, w_105_511, w_105_513, w_105_514, w_105_524, w_105_525, w_105_526, w_105_527, w_105_535, w_105_536, w_105_537, w_105_539, w_105_541, w_105_542, w_105_545, w_105_547, w_105_550, w_105_551, w_105_553, w_105_554, w_105_557, w_105_559, w_105_563, w_105_568, w_105_569, w_105_570, w_105_571, w_105_572, w_105_577, w_105_578, w_105_579, w_105_580, w_105_581, w_105_583, w_105_584, w_105_585, w_105_588, w_105_589, w_105_590, w_105_592, w_105_596, w_105_598, w_105_603, w_105_606, w_105_619, w_105_622, w_105_623, w_105_627, w_105_629, w_105_630, w_105_632, w_105_635, w_105_636, w_105_640, w_105_646, w_105_654, w_105_655, w_105_658, w_105_662, w_105_668, w_105_671, w_105_673, w_105_676, w_105_677, w_105_679, w_105_680, w_105_681, w_105_683, w_105_688, w_105_692, w_105_694, w_105_695, w_105_700, w_105_701, w_105_702, w_105_703, w_105_704, w_105_705, w_105_708, w_105_709, w_105_712, w_105_713, w_105_716, w_105_719, w_105_720, w_105_721, w_105_730, w_105_731, w_105_732, w_105_734, w_105_739, w_105_744, w_105_746, w_105_749, w_105_757, w_105_759, w_105_761, w_105_764, w_105_767, w_105_768, w_105_769, w_105_771, w_105_772, w_105_776, w_105_781, w_105_791, w_105_796, w_105_798, w_105_800, w_105_801, w_105_804, w_105_805, w_105_811, w_105_814, w_105_818, w_105_823, w_105_827, w_105_829, w_105_831, w_105_834, w_105_837, w_105_843, w_105_845, w_105_846, w_105_848, w_105_852, w_105_853, w_105_855, w_105_858, w_105_861, w_105_866, w_105_867, w_105_868, w_105_869, w_105_871, w_105_872, w_105_873, w_105_875, w_105_877, w_105_878, w_105_879, w_105_882, w_105_884, w_105_890, w_105_892, w_105_893, w_105_895, w_105_900, w_105_903, w_105_904, w_105_906, w_105_907, w_105_909, w_105_910, w_105_923, w_105_927, w_105_931, w_105_934, w_105_935, w_105_936, w_105_939, w_105_940, w_105_941, w_105_942, w_105_946, w_105_950, w_105_951, w_105_953, w_105_954, w_105_955, w_105_958, w_105_960, w_105_965, w_105_967, w_105_969, w_105_972, w_105_975, w_105_976, w_105_980, w_105_984, w_105_985, w_105_987, w_105_991, w_105_993, w_105_996, w_105_1000, w_105_1007, w_105_1009, w_105_1013, w_105_1014, w_105_1015, w_105_1019, w_105_1024, w_105_1025, w_105_1027, w_105_1029, w_105_1031, w_105_1034, w_105_1037, w_105_1046, w_105_1050, w_105_1051, w_105_1052, w_105_1055, w_105_1058, w_105_1059, w_105_1060, w_105_1062, w_105_1063, w_105_1064, w_105_1065, w_105_1069, w_105_1073, w_105_1074, w_105_1077, w_105_1081, w_105_1086, w_105_1093, w_105_1094, w_105_1096, w_105_1097, w_105_1099, w_105_1101, w_105_1102, w_105_1103, w_105_1105, w_105_1111, w_105_1114, w_105_1115, w_105_1122, w_105_1123, w_105_1124, w_105_1127, w_105_1129, w_105_1131, w_105_1134, w_105_1135, w_105_1137, w_105_1142, w_105_1147, w_105_1149, w_105_1151, w_105_1153, w_105_1154, w_105_1156, w_105_1159, w_105_1161, w_105_1166, w_105_1170, w_105_1171, w_105_1172, w_105_1174, w_105_1176, w_105_1178, w_105_1184, w_105_1188, w_105_1190, w_105_1196, w_105_1197, w_105_1199, w_105_1200, w_105_1203, w_105_1206, w_105_1211, w_105_1213, w_105_1215, w_105_1219, w_105_1221, w_105_1226, w_105_1228, w_105_1229, w_105_1230, w_105_1239, w_105_1240, w_105_1241, w_105_1246, w_105_1251, w_105_1253, w_105_1254, w_105_1257, w_105_1262, w_105_1264, w_105_1267, w_105_1277, w_105_1278, w_105_1280, w_105_1281, w_105_1282, w_105_1283, w_105_1292, w_105_1295, w_105_1297, w_105_1299, w_105_1301, w_105_1304, w_105_1305, w_105_1306, w_105_1307, w_105_1308, w_105_1311, w_105_1312, w_105_1313, w_105_1315, w_105_1316, w_105_1326, w_105_1327, w_105_1328, w_105_1330, w_105_1331, w_105_1332, w_105_1333, w_105_1335, w_105_1337, w_105_1339, w_105_1340, w_105_1342, w_105_1346, w_105_1350, w_105_1351, w_105_1352, w_105_1353, w_105_1357, w_105_1359, w_105_1361, w_105_1363, w_105_1364, w_105_1365, w_105_1371, w_105_1372, w_105_1376, w_105_1380, w_105_1382, w_105_1383, w_105_1385, w_105_1387, w_105_1388, w_105_1389, w_105_1392, w_105_1394, w_105_1396, w_105_1403, w_105_1405, w_105_1408, w_105_1410, w_105_1411, w_105_1412, w_105_1414, w_105_1415, w_105_1418, w_105_1421, w_105_1425, w_105_1433, w_105_1438, w_105_1440, w_105_1443, w_105_1444, w_105_1448, w_105_1451, w_105_1457, w_105_1458, w_105_1462, w_105_1468, w_105_1470, w_105_1474, w_105_1477, w_105_1482, w_105_1484, w_105_1486, w_105_1488, w_105_1490, w_105_1491, w_105_1493, w_105_1494, w_105_1495, w_105_1501, w_105_1509, w_105_1519, w_105_1522, w_105_1523, w_105_1526, w_105_1529, w_105_1541, w_105_1549, w_105_1551, w_105_1556, w_105_1559, w_105_1560, w_105_1561, w_105_1563, w_105_1571, w_105_1573, w_105_1574, w_105_1578, w_105_1580, w_105_1581, w_105_1582, w_105_1583, w_105_1586, w_105_1587, w_105_1589, w_105_1592, w_105_1600, w_105_1601, w_105_1603, w_105_1604, w_105_1605, w_105_1612, w_105_1614, w_105_1616, w_105_1624, w_105_1627, w_105_1628, w_105_1630, w_105_1631, w_105_1634, w_105_1637, w_105_1639, w_105_1641, w_105_1647, w_105_1648, w_105_1650, w_105_1651, w_105_1655, w_105_1657, w_105_1662, w_105_1663, w_105_1665, w_105_1674, w_105_1679, w_105_1684, w_105_1685, w_105_1691, w_105_1694, w_105_1695, w_105_1696, w_105_1698, w_105_1701, w_105_1703, w_105_1704, w_105_1708, w_105_1711, w_105_1712, w_105_1713, w_105_1717, w_105_1720, w_105_1723, w_105_1726, w_105_1727, w_105_1728, w_105_1729, w_105_1736, w_105_1738, w_105_1744, w_105_1745, w_105_1753, w_105_1760, w_105_1765, w_105_1769, w_105_1770, w_105_1772, w_105_1773, w_105_1775, w_105_1779, w_105_1783, w_105_1784, w_105_1786, w_105_1790, w_105_1791, w_105_1797, w_105_1806, w_105_1810, w_105_1814, w_105_1816, w_105_1818, w_105_1819, w_105_1820, w_105_1830, w_105_1832, w_105_1833, w_105_1836, w_105_1837, w_105_1839, w_105_1841, w_105_1843, w_105_1845, w_105_1846, w_105_1853, w_105_1854, w_105_1855, w_105_1857, w_105_1862, w_105_1864, w_105_1865, w_105_1867, w_105_1872, w_105_1877, w_105_1879, w_105_1882, w_105_1885, w_105_1888, w_105_1890, w_105_1896, w_105_1898, w_105_1899, w_105_1904, w_105_1912, w_105_1913, w_105_1918, w_105_1921, w_105_1923, w_105_1936, w_105_1937, w_105_1939, w_105_1941, w_105_1944, w_105_1945, w_105_1946, w_105_1951, w_105_1955, w_105_1959, w_105_1966, w_105_1967, w_105_1969, w_105_1970, w_105_1974, w_105_1977, w_105_1978, w_105_1979, w_105_1993, w_105_1996, w_105_2007, w_105_2008, w_105_2010, w_105_2011, w_105_2013, w_105_2014, w_105_2017, w_105_2019, w_105_2021, w_105_2027, w_105_2028, w_105_2037, w_105_2038, w_105_2039, w_105_2040, w_105_2041, w_105_2046, w_105_2048, w_105_2050, w_105_2053, w_105_2054, w_105_2056, w_105_2064, w_105_2066, w_105_2067, w_105_2071, w_105_2074, w_105_2076, w_105_2078, w_105_2081, w_105_2085, w_105_2086, w_105_2087, w_105_2088, w_105_2092, w_105_2094, w_105_2095, w_105_2096, w_105_2101, w_105_2102, w_105_2103, w_105_2104, w_105_2115, w_105_2117, w_105_2119, w_105_2122, w_105_2126, w_105_2127, w_105_2130, w_105_2132, w_105_2135, w_105_2137, w_105_2145, w_105_2146, w_105_2147, w_105_2150, w_105_2157, w_105_2158, w_105_2162, w_105_2166, w_105_2168, w_105_2170, w_105_2173, w_105_2174, w_105_2180, w_105_2181, w_105_2182, w_105_2194, w_105_2197, w_105_2198, w_105_2201, w_105_2207, w_105_2209, w_105_2212, w_105_2214, w_105_2215, w_105_2216, w_105_2217, w_105_2218, w_105_2219, w_105_2221, w_105_2223, w_105_2225, w_105_2226, w_105_2229, w_105_2231, w_105_2236, w_105_2239, w_105_2240, w_105_2241, w_105_2245, w_105_2247, w_105_2248, w_105_2249, w_105_2250, w_105_2254, w_105_2255, w_105_2256, w_105_2257, w_105_2262, w_105_2263, w_105_2266, w_105_2267, w_105_2269, w_105_2274, w_105_2275, w_105_2278, w_105_2285, w_105_2287, w_105_2292, w_105_2295, w_105_2298, w_105_2300, w_105_2303, w_105_2304, w_105_2306, w_105_2309, w_105_2316, w_105_2319, w_105_2321, w_105_2327, w_105_2328, w_105_2329, w_105_2331, w_105_2333, w_105_2334, w_105_2337, w_105_2338, w_105_2343, w_105_2344, w_105_2348, w_105_2352, w_105_2354, w_105_2356, w_105_2357, w_105_2358, w_105_2362, w_105_2365, w_105_2366, w_105_2368, w_105_2370, w_105_2371, w_105_2374, w_105_2380, w_105_2384, w_105_2388, w_105_2389, w_105_2392, w_105_2393, w_105_2394, w_105_2398, w_105_2400, w_105_2403, w_105_2415, w_105_2423, w_105_2424, w_105_2425, w_105_2428, w_105_2429, w_105_2431, w_105_2433, w_105_2436, w_105_2439, w_105_2440, w_105_2441, w_105_2442, w_105_2445, w_105_2446, w_105_2447, w_105_2448, w_105_2450, w_105_2453, w_105_2456, w_105_2459, w_105_2460, w_105_2462, w_105_2463, w_105_2464, w_105_2468, w_105_2469, w_105_2471, w_105_2476, w_105_2477, w_105_2478, w_105_2480, w_105_2481, w_105_2483, w_105_2487, w_105_2500, w_105_2505, w_105_2507, w_105_2510, w_105_2514, w_105_2516, w_105_2517, w_105_2523, w_105_2527, w_105_2528, w_105_2531, w_105_2533, w_105_2540, w_105_2541, w_105_2543, w_105_2544, w_105_2545, w_105_2546, w_105_2548, w_105_2552, w_105_2556, w_105_2559, w_105_2561, w_105_2565, w_105_2566, w_105_2567, w_105_2571, w_105_2578, w_105_2581, w_105_2583, w_105_2592, w_105_2593, w_105_2594, w_105_2596, w_105_2599, w_105_2603, w_105_2606, w_105_2607, w_105_2609, w_105_2614, w_105_2618, w_105_2621, w_105_2623, w_105_2627, w_105_2631, w_105_2639, w_105_2643, w_105_2644, w_105_2646, w_105_2647, w_105_2656, w_105_2666, w_105_2675, w_105_2677, w_105_2679, w_105_2685, w_105_2713, w_105_2719, w_105_2720, w_105_2730, w_105_2733, w_105_2739, w_105_2741, w_105_2745, w_105_2751, w_105_2754, w_105_2779, w_105_2787, w_105_2788, w_105_2798, w_105_2799, w_105_2800, w_105_2803, w_105_2808, w_105_2810, w_105_2812, w_105_2816, w_105_2821, w_105_2831, w_105_2832, w_105_2837, w_105_2853, w_105_2867, w_105_2876, w_105_2880, w_105_2884, w_105_2886, w_105_2895, w_105_2907, w_105_2909, w_105_2916, w_105_2920, w_105_2934, w_105_2936, w_105_2937, w_105_2938, w_105_2945, w_105_2947, w_105_2953, w_105_2961, w_105_2962, w_105_2972, w_105_2973, w_105_2977, w_105_2979, w_105_2983, w_105_2985, w_105_2986, w_105_2990, w_105_3000, w_105_3003, w_105_3006, w_105_3007, w_105_3008, w_105_3015, w_105_3017, w_105_3018, w_105_3020, w_105_3023, w_105_3025, w_105_3031, w_105_3035, w_105_3036, w_105_3043, w_105_3046, w_105_3049, w_105_3053, w_105_3055, w_105_3056, w_105_3063, w_105_3067, w_105_3075, w_105_3078, w_105_3080, w_105_3081, w_105_3082, w_105_3088, w_105_3091, w_105_3092, w_105_3096, w_105_3105, w_105_3108, w_105_3112, w_105_3122, w_105_3123, w_105_3131, w_105_3132, w_105_3137, w_105_3142, w_105_3146, w_105_3147, w_105_3160, w_105_3164, w_105_3167, w_105_3170, w_105_3178, w_105_3179, w_105_3187, w_105_3189, w_105_3194, w_105_3197, w_105_3205, w_105_3207, w_105_3212, w_105_3214, w_105_3221, w_105_3229, w_105_3231, w_105_3237, w_105_3238, w_105_3240, w_105_3245, w_105_3246, w_105_3249, w_105_3251, w_105_3252, w_105_3265, w_105_3268, w_105_3274, w_105_3280, w_105_3283, w_105_3297, w_105_3300, w_105_3305, w_105_3313, w_105_3314, w_105_3320, w_105_3329, w_105_3331, w_105_3333, w_105_3338, w_105_3339, w_105_3346, w_105_3347, w_105_3349, w_105_3350, w_105_3357, w_105_3365, w_105_3366, w_105_3368, w_105_3369, w_105_3371, w_105_3377, w_105_3388, w_105_3392, w_105_3399, w_105_3401, w_105_3408, w_105_3410, w_105_3417, w_105_3421, w_105_3425, w_105_3426, w_105_3429, w_105_3434, w_105_3437, w_105_3440, w_105_3441, w_105_3443, w_105_3449, w_105_3457, w_105_3459, w_105_3460, w_105_3462, w_105_3478, w_105_3481, w_105_3488, w_105_3506, w_105_3515, w_105_3516, w_105_3535, w_105_3543, w_105_3544, w_105_3545, w_105_3548, w_105_3557, w_105_3559, w_105_3563, w_105_3567, w_105_3568, w_105_3570, w_105_3572, w_105_3577, w_105_3583, w_105_3590, w_105_3594, w_105_3595, w_105_3600, w_105_3601, w_105_3604, w_105_3608, w_105_3621, w_105_3622, w_105_3633, w_105_3635, w_105_3675, w_105_3681, w_105_3685, w_105_3688, w_105_3694, w_105_3697, w_105_3699, w_105_3705, w_105_3709, w_105_3714, w_105_3716, w_105_3719, w_105_3725, w_105_3726, w_105_3728, w_105_3734, w_105_3735, w_105_3744, w_105_3748, w_105_3750, w_105_3752, w_105_3753, w_105_3758, w_105_3767, w_105_3773, w_105_3774, w_105_3784, w_105_3789, w_105_3790, w_105_3793, w_105_3798, w_105_3800, w_105_3803, w_105_3810, w_105_3812, w_105_3813, w_105_3821, w_105_3822, w_105_3828, w_105_3837, w_105_3842, w_105_3849, w_105_3856, w_105_3859, w_105_3863, w_105_3867, w_105_3876, w_105_3885, w_105_3891, w_105_3894, w_105_3895, w_105_3897, w_105_3900, w_105_3903, w_105_3905, w_105_3906, w_105_3907, w_105_3911, w_105_3912, w_105_3914, w_105_3915, w_105_3920, w_105_3922, w_105_3924, w_105_3931, w_105_3938, w_105_3944, w_105_3948, w_105_3951, w_105_3955, w_105_3964, w_105_3974, w_105_3983, w_105_3988, w_105_3989, w_105_4001, w_105_4011, w_105_4015, w_105_4017, w_105_4020, w_105_4026, w_105_4033, w_105_4035, w_105_4036, w_105_4041, w_105_4044, w_105_4046, w_105_4053, w_105_4061, w_105_4070, w_105_4071, w_105_4074, w_105_4083, w_105_4088, w_105_4094, w_105_4095, w_105_4096, w_105_4101, w_105_4104, w_105_4106, w_105_4109, w_105_4125, w_105_4129, w_105_4161, w_105_4164, w_105_4167, w_105_4170, w_105_4173, w_105_4181, w_105_4182, w_105_4191, w_105_4193, w_105_4197, w_105_4204, w_105_4205, w_105_4214, w_105_4215, w_105_4224, w_105_4228, w_105_4246, w_105_4247, w_105_4260, w_105_4265, w_105_4269, w_105_4276, w_105_4278, w_105_4280, w_105_4282, w_105_4284, w_105_4289, w_105_4294, w_105_4298, w_105_4304, w_105_4310, w_105_4334, w_105_4338, w_105_4339, w_105_4347, w_105_4350, w_105_4361, w_105_4366, w_105_4372, w_105_4377, w_105_4378, w_105_4381, w_105_4382, w_105_4387, w_105_4391, w_105_4395, w_105_4397, w_105_4408, w_105_4409, w_105_4417, w_105_4424, w_105_4425, w_105_4435, w_105_4440, w_105_4442, w_105_4453, w_105_4454, w_105_4456, w_105_4465, w_105_4474, w_105_4475, w_105_4478, w_105_4480, w_105_4486, w_105_4495, w_105_4497, w_105_4508, w_105_4517, w_105_4528, w_105_4547, w_105_4548, w_105_4549, w_105_4550, w_105_4551, w_105_4565, w_105_4575, w_105_4576, w_105_4579, w_105_4580, w_105_4584, w_105_4590, w_105_4594, w_105_4610, w_105_4614, w_105_4618, w_105_4627, w_105_4634, w_105_4635, w_105_4636, w_105_4640, w_105_4651, w_105_4652, w_105_4654, w_105_4657, w_105_4678, w_105_4680, w_105_4681, w_105_4687, w_105_4697, w_105_4698, w_105_4711, w_105_4715, w_105_4716, w_105_4721, w_105_4726, w_105_4730, w_105_4732, w_105_4737, w_105_4740, w_105_4748, w_105_4749, w_105_4750, w_105_4762, w_105_4763, w_105_4767, w_105_4769, w_105_4773, w_105_4779, w_105_4782, w_105_4783, w_105_4784, w_105_4787, w_105_4791, w_105_4796, w_105_4817, w_105_4823, w_105_4825, w_105_4830, w_105_4832, w_105_4833, w_105_4836, w_105_4846, w_105_4848, w_105_4854, w_105_4861, w_105_4862, w_105_4866, w_105_4871, w_105_4876, w_105_4877, w_105_4878, w_105_4881, w_105_4883, w_105_4886, w_105_4888, w_105_4891, w_105_4895, w_105_4897, w_105_4909, w_105_4916, w_105_4920, w_105_4922, w_105_4924, w_105_4930, w_105_4931, w_105_4932, w_105_4935, w_105_4936, w_105_4937, w_105_4938, w_105_4942, w_105_4949, w_10