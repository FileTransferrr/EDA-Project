package dsim_vpi_pkg;
typedef chandle vpiHandle;
localparam vpiAlways = 1;
localparam vpiAssignStmt = 2;
localparam vpiAssignment = 3;
localparam vpiBegin = 4;
localparam vpiCase = 5;
localparam vpiCaseItem = 6;
localparam vpiConstant = 7;
localparam vpiContAssign = 8;
localparam vpiDeassign = 9;
localparam vpiDefParam = 10;
localparam vpiDelayControl = 11;
localparam vpiDisable = 12;
localparam vpiEventControl = 13;
localparam vpiEventStmt = 14;
localparam vpiFor = 15;
localparam vpiForce = 16;
localparam vpiForever = 17;
localparam vpiFork = 18;
localparam vpiFuncCall = 19;
localparam vpiFunction = 20;
localparam vpiGate = 21;
localparam vpiIf = 22;
localparam vpiIfElse = 23;
localparam vpiInitial = 24;
localparam vpiIntegerVar = 25;
localparam vpiInterModPath = 26;
localparam vpiIterator = 27;
localparam vpiIODecl = 28;
localparam vpiMemory = 29;
localparam vpiMemoryWord = 30;
localparam vpiModPath = 31;
localparam vpiModule = 32;
localparam vpiNamedBegin = 33;
localparam vpiNamedEvent = 34;
localparam vpiNamedFork = 35;
localparam vpiNet = 36;
localparam vpiNetBit = 37;
localparam vpiNullStmt = 38;
localparam vpiOperation = 39;
localparam vpiParamAssign = 40;
localparam vpiParameter = 41;
localparam vpiPartSelect = 42;
localparam vpiPathTerm = 43;
localparam vpiPort = 44;
localparam vpiPortBit = 45;
localparam vpiPrimTerm = 46;
localparam vpiRealVar = 47;
localparam vpiReg = 48;
localparam vpiRegBit = 49;
localparam vpiRelease = 50;
localparam vpiRepeat = 51;
localparam vpiRepeatControl = 52;
localparam vpiSchedEvent = 53;
localparam vpiSpecParam = 54;
localparam vpiSwitch = 55;
localparam vpiSysFuncCall = 56;
localparam vpiSysTaskCall = 57;
localparam vpiTableEntry = 58;
localparam vpiTask = 59;
localparam vpiTaskCall = 60;
localparam vpiTchk = 61;
localparam vpiTchkTerm = 62;
localparam vpiTimeVar = 63;
localparam vpiTimeQueue = 64;
localparam vpiUdp = 65;
localparam vpiUdpDefn = 66;
localparam vpiUserSystf = 67;
localparam vpiVarSelect = 68;
localparam vpiWait = 69;
localparam vpiWhile = 70;
localparam vpiAttribute = 105;
localparam vpiBitSelect = 106;
localparam vpiCallback = 107;
localparam vpiDelayTerm = 108;
localparam vpiDelayDevice = 109;
localparam vpiFrame = 110;
localparam vpiGateArray = 111;
localparam vpiModuleArray = 112;
localparam vpiPrimitiveArray = 113;
localparam vpiNetArray = 114;
localparam vpiRange = 115;
localparam vpiRegArray = 116;
localparam vpiSwitchArray = 117;
localparam vpiUdpArray = 118;
localparam vpiContAssignBit = 128;
localparam vpiNamedEventArray = 129;
localparam vpiIndexedPartSelect = 130;
localparam vpiGenScopeArray = 133;
localparam vpiGenScope = 134;
localparam vpiGenVar = 135;
localparam vpiCondition = 71;
localparam vpiDelay = 72;
localparam vpiElseStmt = 73;
localparam vpiForIncStmt = 74;
localparam vpiForInitStmt = 75;
localparam vpiHighConn = 76;
localparam vpiLhs = 77;
localparam vpiIndex = 78;
localparam vpiLeftRange = 79;
localparam vpiLowConn = 80;
localparam vpiParent = 81;
localparam vpiRhs = 82;
localparam vpiRightRange = 83;
localparam vpiScope = 84;
localparam vpiSysTfCall = 85;
localparam vpiTchkDataTerm = 86;
localparam vpiTchkNotifier = 87;
localparam vpiTchkRefTerm = 88;
localparam vpiArgument = 89;
localparam vpiBit = 90;
localparam vpiDriver = 91;
localparam vpiInternalScope = 92;
localparam vpiLoad = 93;
localparam vpiModDataPathIn = 94;
localparam vpiModPathIn = 95;
localparam vpiModPathOut = 96;
localparam vpiOperand = 97;
localparam vpiPortInst = 98;
localparam vpiProcess = 99;
localparam vpiVariables = 100;
localparam vpiUse = 101;
localparam vpiExpr = 102;
localparam vpiPrimitive = 103;
localparam vpiStmt = 104;
localparam vpiActiveTimeFormat = 119;
localparam vpiInTerm = 120;
localparam vpiInstanceArray = 121;
localparam vpiLocalDriver = 122;
localparam vpiLocalLoad = 123;
localparam vpiOutTerm = 124;
localparam vpiPorts = 125;
localparam vpiSimNet = 126;
localparam vpiTaskFunc = 127;
localparam vpiBaseExpr = 131;
localparam vpiWidthExpr = 132;
localparam vpiType = 1;
localparam vpiName = 2;
localparam vpiFullName = 3;
localparam vpiSize = 4;
localparam vpiFile = 5;
localparam vpiLineNo = 6;
localparam vpiTopModule = 7;
localparam vpiCellInstance = 8;
localparam vpiDefName = 9;
localparam vpiProtected = 10;
localparam vpiTimeUnit = 11;
localparam vpiTimePrecision = 12;
localparam vpiDefNetType = 13;
localparam vpiUnconnDrive = 14;
localparam vpiHighZ = 1;
localparam vpiPull1 = 2;
localparam vpiPull0 = 3;
localparam vpiDefFile = 15;
localparam vpiDefLineNo = 16;
localparam vpiDefDelayMode = 47;
localparam vpiDelayModeNone = 1;
localparam vpiDelayModePath = 2;
localparam vpiDelayModeDistrib = 3;
localparam vpiDelayModeUnit = 4;
localparam vpiDelayModeZero = 5;
localparam vpiDelayModeMTM = 6;
localparam vpiDefDecayTime = 48;
localparam vpiScalar = 17;
localparam vpiVector = 18;
localparam vpiExplicitName = 19;
localparam vpiDirection = 20;
localparam vpiInput = 1;
localparam vpiOutput = 2;
localparam vpiInout = 3;
localparam vpiMixedIO = 4;
localparam vpiNoDirection = 5;
localparam vpiConnByName = 21;
localparam vpiNetType = 22;
localparam vpiWire = 1;
localparam vpiWand = 2;
localparam vpiWor = 3;
localparam vpiTri = 4;
localparam vpiTri0 = 5;
localparam vpiTri1 = 6;
localparam vpiTriReg = 7;
localparam vpiTriAnd = 8;
localparam vpiTriOr = 9;
localparam vpiSupply1 = 10;
localparam vpiSupply0 = 11;
localparam vpiNone = 12;
localparam vpiUwire = 13;
localparam vpiExplicitScalared = 23;
localparam vpiExplicitVectored = 24;
localparam vpiExpanded = 25;
localparam vpiImplicitDecl = 26;
localparam vpiChargeStrength = 27;
localparam vpiArray = 28;
localparam vpiPortIndex = 29;
localparam vpiTermIndex = 30;
localparam vpiStrength0 = 31;
localparam vpiStrength1 = 32;
localparam vpiPrimType = 33;
localparam vpiAndPrim = 1;
localparam vpiNandPrim = 2;
localparam vpiNorPrim = 3;
localparam vpiOrPrim = 4;
localparam vpiXorPrim = 5;
localparam vpiXnorPrim = 6;
localparam vpiBufPrim = 7;
localparam vpiNotPrim = 8;
localparam vpiBufif0Prim = 9;
localparam vpiBufif1Prim = 10;
localparam vpiNotif0Prim = 11;
localparam vpiNotif1Prim = 12;
localparam vpiNmosPrim = 13;
localparam vpiPmosPrim = 14;
localparam vpiCmosPrim = 15;
localparam vpiRnmosPrim = 16;
localparam vpiRpmosPrim = 17;
localparam vpiRcmosPrim = 18;
localparam vpiRtranPrim = 19;
localparam vpiRtranif0Prim = 20;
localparam vpiRtranif1Prim = 21;
localparam vpiTranPrim = 22;
localparam vpiTranif0Prim = 23;
localparam vpiTranif1Prim = 24;
localparam vpiPullupPrim = 25;
localparam vpiPulldownPrim = 26;
localparam vpiSeqPrim = 27;
localparam vpiCombPrim = 28;
localparam vpiPolarity = 34;
localparam vpiDataPolarity = 35;
localparam vpiPositive = 1;
localparam vpiNegative = 2;
localparam vpiUnknown = 3;
localparam vpiEdge = 36;
localparam vpiNoEdge = 0;
localparam vpiEdge01 = 0;
localparam vpiEdge10 = 0;
localparam vpiEdge0x = 0;
localparam vpiEdgex1 = 0;
localparam vpiEdge1x = 0;
localparam vpiEdgex0 = 0;
localparam vpiPathType = 37;
localparam vpiPathFull = 1;
localparam vpiPathParallel = 2;
localparam vpiTchkType = 38;
localparam vpiSetup = 1;
localparam vpiHold = 2;
localparam vpiPeriod = 3;
localparam vpiWidth = 4;
localparam vpiSkew = 5;
localparam vpiRecovery = 6;
localparam vpiNoChange = 7;
localparam vpiSetupHold = 8;
localparam vpiFullskew = 9;
localparam vpiRecrem = 10;
localparam vpiRemoval = 11;
localparam vpiTimeskew = 12;
localparam vpiOpType = 39;
localparam vpiMinusOp = 1;
localparam vpiPlusOp = 2;
localparam vpiNotOp = 3;
localparam vpiBitNegOp = 4;
localparam vpiUnaryAndOp = 5;
localparam vpiUnaryNandOp = 6;
localparam vpiUnaryOrOp = 7;
localparam vpiUnaryNorOp = 8;
localparam vpiUnaryXorOp = 9;
localparam vpiUnaryXNorOp = 10;
localparam vpiSubOp = 11;
localparam vpiDivOp = 12;
localparam vpiModOp = 13;
localparam vpiEqOp = 14;
localparam vpiNeqOp = 15;
localparam vpiCaseEqOp = 16;
localparam vpiCaseNeqOp = 17;
localparam vpiGtOp = 18;
localparam vpiGeOp = 19;
localparam vpiLtOp = 20;
localparam vpiLeOp = 21;
localparam vpiLShiftOp = 22;
localparam vpiRShiftOp = 23;
localparam vpiAddOp = 24;
localparam vpiMultOp = 25;
localparam vpiLogAndOp = 26;
localparam vpiLogOrOp = 27;
localparam vpiBitAndOp = 28;
localparam vpiBitOrOp = 29;
localparam vpiBitXorOp = 30;
localparam vpiBitXNorOp = 31;
localparam vpiConditionOp = 32;
localparam vpiConcatOp = 33;
localparam vpiMultiConcatOp = 34;
localparam vpiEventOrOp = 35;
localparam vpiNullOp = 36;
localparam vpiListOp = 37;
localparam vpiMinTypMaxOp = 38;
localparam vpiPosedgeOp = 39;
localparam vpiNegedgeOp = 40;
localparam vpiArithLShiftOp = 41;
localparam vpiArithRShiftOp = 42;
localparam vpiPowerOp = 43;
localparam vpiConstType = 40;
localparam vpiDecConst = 1;
localparam vpiRealConst = 2;
localparam vpiBinaryConst = 3;
localparam vpiOctConst = 4;
localparam vpiHexConst = 5;
localparam vpiStringConst = 6;
localparam vpiIntConst = 7;
localparam vpiBlocking = 41;
localparam vpiCaseType = 42;
localparam vpiCaseExact = 1;
localparam vpiCaseX = 2;
localparam vpiCaseZ = 3;
localparam vpiNetDeclAssign = 43;
localparam vpiFuncType = 44;
localparam vpiIntFunc = 1;
localparam vpiRealFunc = 2;
localparam vpiTimeFunc = 3;
localparam vpiSizedFunc = 4;
localparam vpiSizedSignedFunc = 5;
localparam vpiUserDefn = 45;
localparam vpiScheduled = 46;
localparam vpiActive = 49;
localparam vpiAutomatic = 50;
localparam vpiCell = 51;
localparam vpiConfig = 52;
localparam vpiConstantSelect = 53;
localparam vpiDecompile = 54;
localparam vpiDefAttribute = 55;
localparam vpiDelayType = 56;
localparam vpiModPathDelay = 1;
localparam vpiInterModPathDelay = 2;
localparam vpiMIPDelay = 3;
localparam vpiIteratorType = 57;
localparam vpiLibrary = 58;
localparam vpiMultiArray = 59;
localparam vpiOffset = 60;
localparam vpiResolvedNetType = 61;
localparam vpiSaveRestartID = 62;
localparam vpiSaveRestartLocation = 63;
localparam vpiValid = 64;
localparam vpiSigned = 65;
localparam vpiLocalParam = 70;
localparam vpiModPathHasIfNone = 71;
localparam vpiIndexedPartSelectType = 72;
localparam vpiPosIndexed = 1;
localparam vpiNegIndexed = 2;
localparam vpiIsMemory = 73;
localparam vpiIsProtected = 74;
localparam vpiStop = 66;
localparam vpiFinish = 67;
localparam vpiReset = 68;
localparam vpiSetInteractiveScope = 69;
localparam vpiScaledRealTime = 1;
localparam vpiSimTime = 2;
localparam vpiSuppressTime = 3;
localparam vpiSupplyDrive = 0;
localparam vpiStrongDrive = 0;
localparam vpiPullDrive = 0;
localparam vpiWeakDrive = 0;
localparam vpiLargeCharge = 0;
localparam vpiMediumCharge = 0;
localparam vpiSmallCharge = 0;
localparam vpiHiZ = 0;
localparam vpiBinStrVal = 1;
localparam vpiOctStrVal = 2;
localparam vpiDecStrVal = 3;
localparam vpiHexStrVal = 4;
localparam vpiScalarVal = 5;
localparam vpiIntVal = 6;
localparam vpiRealVal = 7;
localparam vpiStringVal = 8;
localparam vpiVectorVal = 9;
localparam vpiStrengthVal = 10;
localparam vpiTimeVal = 11;
localparam vpiObjTypeVal = 12;
localparam vpiSuppressVal = 13;
localparam vpiNoDelay = 1;
localparam vpiInertialDelay = 2;
localparam vpiTransportDelay = 3;
localparam vpiPureTransportDelay = 4;
localparam vpiForceFlag = 5;
localparam vpiReleaseFlag = 6;
localparam vpiCancelEvent = 7;
localparam vpiReturnEvent = 0;
localparam vpi0 = 0;
localparam vpi1 = 1;
localparam vpiZ = 2;
localparam vpiX = 3;
localparam vpiH = 4;
localparam vpiL = 5;
localparam vpiDontCare = 6;
localparam vpiSysTask = 1;
localparam vpiSysFunc = 2;
localparam vpiCompile = 1;
localparam vpiPLI = 2;
localparam vpiRun = 3;
localparam vpiNotice = 1;
localparam vpiWarning = 2;
localparam vpiError = 3;
localparam vpiSystem = 4;
localparam vpiInternal = 5;
localparam cbValueChange = 1;
localparam cbStmt = 2;
localparam cbForce = 3;
localparam cbRelease = 4;
localparam cbAtStartOfSimTime = 5;
localparam cbReadWriteSynch = 6;
localparam cbReadOnlySynch = 7;
localparam cbNextSimTime = 8;
localparam cbAfterDelay = 9;
localparam cbEndOfCompile = 10;
localparam cbStartOfSimulation = 11;
localparam cbEndOfSimulation = 12;
localparam cbError = 13;
localparam cbTchkViolation = 14;
localparam cbStartOfSave = 15;
localparam cbEndOfSave = 16;
localparam cbStartOfRestart = 17;
localparam cbEndOfRestart = 18;
localparam cbStartOfReset = 19;
localparam cbEndOfReset = 20;
localparam cbEnterInteractive = 21;
localparam cbExitInteractive = 22;
localparam cbInteractiveScopeChange = 23;
localparam cbUnresolvedSystf = 24;
localparam cbAssign = 25;
localparam cbDeassign = 26;
localparam cbDisable = 27;
localparam cbPLIError = 28;
localparam cbSignal = 29;
localparam cbNBASynch = 30;
localparam cbAtEndOfSimTime = 31;
localparam vpiPackage = 600;
localparam vpiInterface = 601;
localparam vpiProgram = 602;
localparam vpiInterfaceArray = 603;
localparam vpiProgramArray = 604;
localparam vpiTypespec = 605;
localparam vpiModport = 606;
localparam vpiInterfaceTfDecl = 607;
localparam vpiRefObj = 608;
localparam vpiTypeParameter = 609;
localparam vpiLongIntVar = 610;
localparam vpiShortIntVar = 611;
localparam vpiIntVar = 612;
localparam vpiShortRealVar = 613;
localparam vpiByteVar = 614;
localparam vpiClassVar = 615;
localparam vpiStringVar = 616;
localparam vpiEnumVar = 617;
localparam vpiStructVar = 618;
localparam vpiUnionVar = 619;
localparam vpiBitVar = 620;
localparam vpiClassObj = 621;
localparam vpiChandleVar = 622;
localparam vpiPackedArrayVar = 623;
localparam vpiVirtualInterfaceVar = 728;
localparam vpiLongIntTypespec = 625;
localparam vpiShortRealTypespec = 626;
localparam vpiByteTypespec = 627;
localparam vpiShortIntTypespec = 628;
localparam vpiIntTypespec = 629;
localparam vpiClassTypespec = 630;
localparam vpiStringTypespec = 631;
localparam vpiChandleTypespec = 632;
localparam vpiEnumTypespec = 633;
localparam vpiEnumConst = 634;
localparam vpiIntegerTypespec = 635;
localparam vpiTimeTypespec = 636;
localparam vpiRealTypespec = 637;
localparam vpiStructTypespec = 638;
localparam vpiUnionTypespec = 639;
localparam vpiBitTypespec = 640;
localparam vpiLogicTypespec = 641;
localparam vpiArrayTypespec = 642;
localparam vpiVoidTypespec = 643;
localparam vpiTypespecMember = 644;
localparam vpiPackedArrayTypespec = 692;
localparam vpiSequenceTypespec = 696;
localparam vpiPropertyTypespec = 697;
localparam vpiEventTypespec = 698;
localparam vpiInterfaceTypespec = 906;
localparam vpiClockingBlock = 650;
localparam vpiClockingIODecl = 651;
localparam vpiClassDefn = 652;
localparam vpiConstraint = 653;
localparam vpiConstraintOrdering = 654;
localparam vpiDistItem = 645;
localparam vpiAliasStmt = 646;
localparam vpiThread = 647;
localparam vpiMethodFuncCall = 648;
localparam vpiMethodTaskCall = 649;
localparam vpiAssert = 686;
localparam vpiAssume = 687;
localparam vpiCover = 688;
localparam vpiRestrict = 901;
localparam vpiDisableCondition = 689;
localparam vpiClockingEvent = 690;
localparam vpiPropertyDecl = 655;
localparam vpiPropertySpec = 656;
localparam vpiPropertyExpr = 657;
localparam vpiMulticlockSequenceExpr = 658;
localparam vpiClockedSeq = 659;
localparam vpiClockedProp = 902;
localparam vpiPropertyInst = 660;
localparam vpiSequenceDecl = 661;
localparam vpiCaseProperty = 662;
localparam vpiCasePropertyItem = 905;
localparam vpiSequenceInst = 664;
localparam vpiImmediateAssert = 665;
localparam vpiImmediateAssume = 694;
localparam vpiImmediateCover = 695;
localparam vpiReturn = 666;
localparam vpiAnyPattern = 667;
localparam vpiTaggedPattern = 668;
localparam vpiStructPattern = 669;
localparam vpiDoWhile = 670;
localparam vpiOrderedWait = 671;
localparam vpiWaitFork = 672;
localparam vpiDisableFork = 673;
localparam vpiExpectStmt = 674;
localparam vpiForeachStmt = 675;
localparam vpiReturnStmt = 691;
localparam vpiFinal = 676;
localparam vpiExtends = 677;
localparam vpiDistribution = 678;
localparam vpiSeqFormalDecl = 679;
localparam vpiPropFormalDecl = 699;
localparam vpiEnumNet = 680;
localparam vpiIntegerNet = 681;
localparam vpiTimeNet = 682;
localparam vpiStructNet = 683;
localparam vpiBreak = 684;
localparam vpiContinue = 685;
localparam vpiPackedArrayNet = 693;
localparam vpiConstraintExpr = 747;
localparam vpiElseConst = 748;
localparam vpiImplication = 749;
localparam vpiConstrIf = 738;
localparam vpiConstrIfElse = 739;
localparam vpiConstrForEach = 736;
localparam vpiSoftDisable = 733;
localparam vpiLetDecl = 903;
localparam vpiLetExpr = 904;
localparam vpiActual = 700;
localparam vpiTypedefAlias = 701;
localparam vpiIndexTypespec = 702;
localparam vpiBaseTypespec = 703;
localparam vpiElemTypespec = 704;
localparam vpiInputSkew = 706;
localparam vpiOutputSkew = 707;
localparam vpiGlobalClocking = 708;
localparam vpiDefaultClocking = 709;
localparam vpiDefaultDisableIff = 710;
localparam vpiOrigin = 713;
localparam vpiPrefix = 714;
localparam vpiWith = 715;
localparam vpiProperty = 718;
localparam vpiValueRange = 720;
localparam vpiPattern = 721;
localparam vpiWeight = 722;
localparam vpiConstraintItem = 746;
localparam vpiTypedef = 725;
localparam vpiImport = 726;
localparam vpiDerivedClasses = 727;
localparam vpiMethods = 730;
localparam vpiSolveBefore = 731;
localparam vpiSolveAfter = 732;
localparam vpiWaitingProcesses = 734;
localparam vpiMessages = 735;
localparam vpiLoopVars = 737;
localparam vpiConcurrentAssertions = 740;
localparam vpiMatchItem = 741;
localparam vpiMember = 742;
localparam vpiElement = 743;
localparam vpiAssertion = 744;
localparam vpiInstance = 745;
localparam vpiTop = 600;
localparam vpiUnit = 602;
localparam vpiJoinType = 603;
localparam vpiJoin = 0;
localparam vpiJoinNone = 1;
localparam vpiJoinAny = 2;
localparam vpiAccessType = 604;
localparam vpiForkJoinAcc = 1;
localparam vpiExternAcc = 2;
localparam vpiDPIExportAcc = 3;
localparam vpiDPIImportAcc = 4;
localparam vpiArrayType = 606;
localparam vpiStaticArray = 1;
localparam vpiDynamicArray = 2;
localparam vpiAssocArray = 3;
localparam vpiQueueArray = 4;
localparam vpiArrayMember = 607;
localparam vpiIsRandomized = 608;
localparam vpiLocalVarDecls = 609;
localparam vpiOpStrong = 656;
localparam vpiRandType = 610;
localparam vpiNotRand = 1;
localparam vpiRand = 2;
localparam vpiRandC = 3;
localparam vpiPortType = 611;
localparam vpiInterfacePort = 1;
localparam vpiModportPort = 2;
localparam vpiConstantVariable = 612;
localparam vpiStructUnionMember = 615;
localparam vpiVisibility = 620;
localparam vpiPublicVis = 1;
localparam vpiProtectedVis = 2;
localparam vpiLocalVis = 3;
localparam vpiOneStepConst = 9;
localparam vpiUnboundedConst = 10;
localparam vpiNullConst = 11;
localparam vpiAlwaysType = 624;
localparam vpiAlwaysComb = 2;
localparam vpiAlwaysFF = 3;
localparam vpiAlwaysLatch = 4;
localparam vpiDistType = 625;
localparam vpiEqualDist = 1;
localparam vpiDivDist = 2;
localparam vpiPacked = 630;
localparam vpiTagged = 632;
localparam vpiRef = 6;
localparam vpiVirtual = 635;
localparam vpiHasActual = 636;
localparam vpiIsConstraintEnabled = 638;
localparam vpiSoft = 639;
localparam vpiClassType = 640;
localparam vpiMailboxClass = 1;
localparam vpiSemaphoreClass = 2;
localparam vpiUserDefinedClass = 3;
localparam vpiProcessClass = 4;
localparam vpiMethod = 645;
localparam vpiIsClockInferred = 649;
localparam vpiIsDeferred = 657;
localparam vpiIsFinal = 670;
localparam vpiIsCoverSequence = 659;
localparam vpiQualifier = 650;
localparam vpiNoQualifier = 0;
localparam vpiUniqueQualifier = 1;
localparam vpiPriorityQualifier = 2;
localparam vpiTaggedQualifier = 4;
localparam vpiRandQualifier = 8;
localparam vpiInsideQualifier = 16;
localparam vpiInputEdge = 651;
localparam vpiOutputEdge = 652;
localparam vpiGeneric = 653;
localparam vpiCompatibilityMode = 654;
localparam vpiMode1364v1995 = 1;
localparam vpiMode1364v2001 = 2;
localparam vpiMode1364v2005 = 3;
localparam vpiMode1800v2005 = 4;
localparam vpiMode1800v2009 = 5;
localparam vpiPackedArrayMember = 655;
localparam vpiStartLine = 661;
localparam vpiColumn = 662;
localparam vpiEndLine = 663;
localparam vpiEndColumn = 664;
localparam vpiAllocScheme = 658;
localparam vpiAutomaticScheme = 1;
localparam vpiDynamicScheme = 2;
localparam vpiOtherScheme = 3;
localparam vpiObjId = 660;
localparam vpiDPIPure = 665;
localparam vpiDPIContext = 666;
localparam vpiDPICStr = 667;
localparam vpiDPI = 1;
localparam vpiDPIC = 2;
localparam vpiDPICIdentifier = 668;
localparam vpiIsModPort = 669;
localparam vpiImplyOp = 50;
localparam vpiNonOverlapImplyOp = 51;
localparam vpiOverlapImplyOp = 52;
localparam vpiAcceptOnOp = 83;
localparam vpiRejectOnOp = 84;
localparam vpiSyncAcceptOnOp = 85;
localparam vpiSyncRejectOnOp = 86;
localparam vpiOverlapFollowedByOp = 87;
localparam vpiNonOverlapFollowedByOp = 88;
localparam vpiNexttimeOp = 89;
localparam vpiAlwaysOp = 90;
localparam vpiEventuallyOp = 91;
localparam vpiUntilOp = 92;
localparam vpiUntilWithOp = 93;
localparam vpiUnaryCycleDelayOp = 53;
localparam vpiCycleDelayOp = 54;
localparam vpiIntersectOp = 55;
localparam vpiFirstMatchOp = 56;
localparam vpiThroughoutOp = 57;
localparam vpiWithinOp = 58;
localparam vpiRepeatOp = 59;
localparam vpiConsecutiveRepeatOp = 60;
localparam vpiGotoRepeatOp = 61;
localparam vpiPostIncOp = 62;
localparam vpiPreIncOp = 63;
localparam vpiPostDecOp = 64;
localparam vpiPreDecOp = 65;
localparam vpiMatchOp = 66;
localparam vpiCastOp = 67;
localparam vpiIffOp = 68;
localparam vpiWildEqOp = 69;
localparam vpiWildNeqOp = 70;
localparam vpiStreamLROp = 71;
localparam vpiStreamRLOp = 72;
localparam vpiMatchedOp = 73;
localparam vpiTriggeredOp = 74;
localparam vpiAssignmentPatternOp = 75;
localparam vpiMultiAssignmentPatternOp = 76;
localparam vpiIfOp = 77;
localparam vpiIfElseOp = 78;
localparam vpiCompAndOp = 79;
localparam vpiCompOrOp = 80;
localparam vpiImpliesOp = 94;
localparam vpiInsideOp = 95;
localparam vpiTypeOp = 81;
localparam vpiAssignmentOp = 82;
localparam vpiOtherFunc = 6;
localparam vpiValidUnknown = 2;
localparam cbStartOfThread = 600;
localparam cbEndOfThread = 601;
localparam cbEnterThread = 602;
localparam cbStartOfFrame = 603;
localparam cbEndOfFrame = 604;
localparam cbSizeChange = 605;
localparam cbCreateObj = 700;
localparam cbReclaimObj = 701;
localparam cbEndOfObject = 702;
localparam vpiCoverageStart = 750;
localparam vpiCoverageStop = 751;
localparam vpiCoverageReset = 752;
localparam vpiCoverageCheck = 753;
localparam vpiCoverageMerge = 754;
localparam vpiCoverageSave = 755;
localparam vpiAssertCoverage = 760;
localparam vpiFsmStateCoverage = 761;
localparam vpiStatementCoverage = 762;
localparam vpiToggleCoverage = 763;
localparam vpiCovered = 765;
localparam vpiCoverMax = 766;
localparam vpiCoveredMax = 766;
localparam vpiCoveredCount = 767;
localparam vpiAssertAttemptCovered = 770;
localparam vpiAssertSuccessCovered = 771;
localparam vpiAssertFailureCovered = 772;
localparam vpiAssertVacuousSuccessCovered = 773;
localparam vpiAssertDisableCovered = 774;
localparam vpiAssertKillCovered = 777;
localparam vpiFsmStates = 775;
localparam vpiFsmStateExpression = 776;
localparam vpiFsm = 758;
localparam vpiFsmHandle = 759;
localparam cbAssertionStart = 606;
localparam cbAssertionSuccess = 607;
localparam cbAssertionFailure = 608;
localparam cbAssertionVacuousSuccess = 657;
localparam cbAssertionDisabledEvaluation = 658;
localparam cbAssertionStepSuccess = 609;
localparam cbAssertionStepFailure = 610;
localparam cbAssertionLock = 661;
localparam cbAssertionUnlock = 662;
localparam cbAssertionDisable = 611;
localparam cbAssertionEnable = 612;
localparam cbAssertionReset = 613;
localparam cbAssertionKill = 614;
localparam cbAssertionEnablePassAction = 645;
localparam cbAssertionEnableFailAction = 646;
localparam cbAssertionDisablePassAction = 647;
localparam cbAssertionDisableFailAction = 648;
localparam cbAssertionEnableNonvacuousAction = 649;
localparam cbAssertionDisableVacuousAction = 650;
localparam cbAssertionSysInitialized = 615;
localparam cbAssertionSysOn = 616;
localparam cbAssertionSysOff = 617;
localparam cbAssertionSysKill = 631;
localparam cbAssertionSysLock = 659;
localparam cbAssertionSysUnlock = 660;
localparam cbAssertionSysEnd = 618;
localparam cbAssertionSysReset = 619;
localparam cbAssertionSysEnablePassAction = 651;
localparam cbAssertionSysEnableFailAction = 652;
localparam cbAssertionSysDisablePassAction = 653;
localparam cbAssertionSysDisableFailAction = 654;
localparam cbAssertionSysEnableNonvacuousAction = 655;
localparam cbAssertionSysDisableVacuousAction = 656;
localparam vpiAssertionLock = 645;
localparam vpiAssertionUnlock = 646;
localparam vpiAssertionDisable = 620;
localparam vpiAssertionEnable = 621;
localparam vpiAssertionReset = 622;
localparam vpiAssertionKill = 623;
localparam vpiAssertionEnableStep = 624;
localparam vpiAssertionDisableStep = 625;
localparam vpiAssertionClockSteps = 626;
localparam vpiAssertionSysLock = 647;
localparam vpiAssertionSysUnlock = 648;
localparam vpiAssertionSysOn = 627;
localparam vpiAssertionSysOff = 628;
localparam vpiAssertionSysKill = 632;
localparam vpiAssertionSysEnd = 629;
localparam vpiAssertionSysReset = 630;
localparam vpiAssertionDisablePassAction = 633;
localparam vpiAssertionEnablePassAction = 634;
localparam vpiAssertionDisableFailAction = 635;
localparam vpiAssertionEnableFailAction = 636;
localparam vpiAssertionDisableVacuousAction = 637;
localparam vpiAssertionEnableNonvacuousAction = 638;
localparam vpiAssertionSysEnablePassAction = 639;
localparam vpiAssertionSysEnableFailAction = 640;
localparam vpiAssertionSysDisablePassAction = 641;
localparam vpiAssertionSysDisableFailAction = 642;
localparam vpiAssertionSysEnableNonvacuousAction = 643;
localparam vpiAssertionSysDisableVacuousAction = 644;
import "DPI-C" function vpiHandle vpi_handle_by_name(string name, vpiHandle scope);
import "DPI-C" function vpiHandle vpi_handle_by_index(string name, vpiHandle indx);
import "DPI-C" function vpiHandle vpi_handle(int arg, vpiHandle handle);
import "DPI-C" function vpiHandle vpi_iterate(int arg, vpiHandle handle);
import "DPI-C" function vpiHandle vpi_scan(vpiHandle handle);
import "DPI-C" function int vpi_get(int prop, vpiHandle obj);
import "DPI-C" function string vpi_get_str(int prop, vpiHandle obj);
import "DPI-C" function int vpi_release_handle(vpiHandle obj);

//import "DPI-C" function void vpi_get_value_4s(vpiHandle h, output reg [] value);
//import "DPI-C" function void vpi_put_value_4s(vpiHandle h, reg [] value, int flags);

endpackage
