// ****** Basic Gate Module Defination ******
module or2(out, in1, in2);
  output out;
  input in1, in2;
  wire in1, in2, out;
  assign out = in1 || in2;
endmodule

module and2(out, in1, in2);
  output out;
  input in1, in2;
  wire in1, in2, out;
  assign out = in1 && in2;
endmodule

module not1(out, in);
  output out;
  input in;
  wire in,out;
  assign out = ~in;
endmodule

module nand2(out, in1, in2);
  output out;
  input in1, in2;
  wire in1, in2, out;
  assign out = ~(in1 && in2);
endmodule
// ****** Basic Gate Module Defination End ******

// ****** Combined Logic Module Defination ******
module combLogic( w_000_000, w_000_001, w_000_002, w_000_003, w_000_004, w_000_005, w_000_006, w_000_007, w_000_008, w_000_009, w_000_010, w_000_011, w_000_012, w_000_013, w_000_014, w_000_015, w_000_016, w_000_017, w_000_018, w_000_019, w_000_020, w_000_021, w_000_022, w_000_023, w_000_024, w_000_025, w_000_026, w_000_027, w_000_028, w_000_029, w_000_030, w_000_031, w_000_032, w_000_033, w_000_034, w_000_035, w_000_036, w_000_037, w_000_038, w_000_039, w_000_040, w_000_041, w_000_042, w_000_043, w_000_044, w_000_045, w_000_046, w_000_047, w_000_048, w_000_049, w_000_050, w_000_051, w_000_052, w_000_053, w_000_054, w_000_055, w_000_056, w_000_057, w_000_058, w_000_059, w_000_060, w_000_061, w_000_062, w_000_063, w_000_064, w_000_065, w_000_066, w_000_067, w_000_068, w_000_069, w_000_070, w_000_071, w_000_072, w_000_073, w_000_074, w_000_075, w_000_076, w_000_077, w_000_078, w_000_079, w_000_080, w_000_081, w_000_082, w_000_083, w_000_084, w_000_085, w_000_086, w_000_087, w_000_088, w_000_089, w_000_090, w_000_091, w_000_092, w_000_093, w_000_094, w_000_095, w_000_096, w_000_097, w_000_098, w_000_099, w_000_100, w_000_101, w_000_102, w_000_103, w_000_104, w_000_105, w_000_106, w_000_107, w_000_108, w_000_109, w_000_110, w_000_111, w_000_112, w_000_113, w_000_114, w_000_115, w_000_116, w_000_117, w_000_118, w_000_119, w_000_120, w_000_121, w_000_122, w_000_123, w_000_124, w_000_125, w_000_126, w_000_127, w_000_128, w_000_129, w_000_130, w_000_131, w_000_132, w_000_133, w_000_134, w_000_135, w_000_136, w_000_137, w_000_138, w_000_139, w_000_140, w_000_141, w_000_142, w_000_143, w_000_144, w_000_145, w_000_146, w_000_147, w_000_148, w_000_149, w_000_150, w_000_151, w_000_152, w_000_153, w_000_154, w_000_155, w_000_156, w_000_157, w_000_158, w_000_159, w_000_160, w_000_161, w_000_162, w_000_163, w_000_164, w_000_165, w_000_166, w_000_167, w_000_168, w_000_169, w_000_170, w_000_171, w_000_172, w_000_173, w_000_174, w_000_175, w_000_176, w_000_177, w_000_178, w_000_179, w_000_180, w_000_181, w_000_182, w_000_183, w_000_184, w_000_185, w_000_186, w_000_187, w_000_188, w_000_189, w_000_190, w_000_191, w_000_192, w_000_193, w_000_194, w_000_195, w_000_196, w_000_197, w_000_198, w_000_199, w_000_200, w_000_201, w_000_202, w_000_203, w_000_204, w_000_205, w_000_206, w_000_207, w_000_208, w_000_209, w_000_210, w_000_211, w_000_212, w_000_213, w_000_214, w_000_215, w_000_216, w_000_217, w_000_218, w_000_219, w_000_220, w_000_221, w_000_222, w_000_223, w_000_224, w_000_225, w_000_226, w_000_227, w_000_228, w_000_229, w_000_230, w_000_231, w_000_232, w_000_233, w_000_234, w_000_235, w_000_236, w_000_237, w_000_238, w_000_239, w_000_240, w_000_241, w_000_242, w_000_243, w_000_244, w_000_245, w_000_246, w_000_247, w_000_248, w_000_249, w_000_250, w_000_251, w_000_252, w_000_253, w_000_254, w_000_255, w_000_256, w_000_257, w_000_258, w_000_259, w_000_260, w_000_261, w_000_262, w_000_263, w_000_264, w_000_265, w_000_266, w_000_267, w_000_268, w_000_269, w_000_270, w_000_271, w_000_272, w_000_273, w_000_274, w_000_275, w_000_276, w_000_277, w_000_278, w_000_279, w_000_280, w_000_281, w_000_282, w_000_283, w_000_284, w_000_285, w_000_286, w_000_287, w_000_288, w_000_289, w_000_290, w_000_291, w_000_292, w_000_293, w_000_294, w_000_295, w_000_296, w_000_297, w_000_298, w_000_299, w_000_300, w_000_301, w_000_302, w_000_303, w_000_304, w_000_305, w_000_306, w_000_307, w_000_308, w_000_309, w_000_310, w_000_311, w_000_312, w_000_313, w_000_314, w_000_315, w_000_316, w_000_317, w_000_318, w_000_319, w_000_320, w_000_321, w_000_322, w_000_323, w_000_324, w_000_325, w_000_326, w_000_327, w_000_328, w_000_329, w_000_330, w_000_331, w_000_332, w_000_333, w_000_334, w_000_335, w_000_336, w_000_337, w_000_338, w_000_339, w_000_340, w_000_341, w_000_342, w_000_343, w_000_344, w_000_345, w_000_346, w_000_347, w_000_348, w_000_349, w_000_350, w_000_351, w_000_352, w_000_353, w_000_354, w_000_355, w_000_356, w_000_357, w_000_358, w_000_359, w_000_360, w_000_361, w_000_362, w_000_363, w_000_364, w_000_365, w_000_366, w_000_367, w_000_368, w_000_369, w_000_370, w_000_371, w_000_372, w_000_373, w_000_374, w_000_375, w_000_376, w_000_377, w_000_378, w_000_379, w_000_380, w_000_381, w_000_382, w_000_383, w_000_384, w_000_385, w_000_386, w_000_387, w_000_388, w_000_389, w_000_390, w_000_391, w_000_392, w_000_393, w_000_394, w_000_395, w_000_396, w_000_397, w_000_398, w_000_399, w_000_400, w_000_401, w_000_402, w_000_403, w_000_404, w_000_405, w_000_406, w_000_407, w_000_408, w_000_409, w_000_410, w_000_411, w_000_412, w_000_413, w_000_414, w_000_415, w_000_416, w_000_417, w_000_418, w_000_419, w_000_420, w_000_421, w_000_422, w_000_423, w_000_424, w_000_425, w_000_426, w_000_427, w_000_428, w_000_429, w_000_430, w_000_431, w_000_432, w_000_433, w_000_434, w_000_435, w_000_436, w_000_437, w_000_438, w_000_439, w_000_440, w_000_441, w_000_442, w_000_443, w_000_444, w_000_445, w_000_446, w_000_447, w_000_448, w_000_449, w_000_450, w_000_451, w_000_452, w_000_453, w_000_454, w_000_455, w_000_456, w_000_457, w_000_458, w_000_459, w_000_460, w_000_461, w_000_462, w_000_463, w_000_464, w_000_465, w_000_466, w_000_467, w_000_468, w_000_469, w_000_470, w_000_471, w_000_472, w_000_473, w_000_474, w_000_475, w_000_476, w_000_477, w_000_478, w_000_479, w_000_480, w_000_481, w_000_482, w_000_483, w_000_484, w_000_485, w_000_486, w_000_487, w_000_488, w_000_489, w_000_490, w_000_491, w_000_492, w_000_493, w_000_494, w_000_495, w_000_496, w_000_497, w_000_498, w_000_499, w_000_500, w_000_501, w_000_502, w_000_503, w_000_504, w_000_505, w_000_506, w_000_507, w_000_508, w_000_509, w_000_510, w_000_511, w_000_512, w_000_513, w_000_514, w_000_515, w_000_516, w_000_517, w_000_518, w_000_519, w_000_520, w_000_521, w_000_522, w_000_523, w_000_524, w_000_525, w_000_526, w_000_527, w_000_528, w_000_529, w_000_530, w_000_531, w_000_532, w_000_533, w_000_534, w_000_535, w_000_536, w_000_537, w_000_538, w_000_539, w_000_540, w_000_541, w_000_542, w_000_543, w_000_544, w_000_545, w_000_546, w_000_547, w_000_548, w_000_549, w_000_550, w_000_551, w_000_552, w_000_553, w_000_554, w_000_555, w_000_556, w_000_557, w_000_558, w_000_559, w_000_560, w_000_561, w_000_562, w_000_563, w_000_564, w_000_565, w_000_566, w_000_567, w_000_568, w_000_569, w_000_570, w_000_571, w_000_572, w_000_573, w_000_574, w_000_575, w_000_576, w_000_577, w_000_578, w_000_579, w_000_580, w_000_581, w_000_582, w_000_583, w_000_584, w_000_585, w_000_586, w_000_587, w_000_588, w_000_589, w_000_590, w_000_591, w_000_592, w_000_593, w_000_594, w_000_595, w_000_596, w_000_597, w_000_598, w_000_599, w_000_600, w_000_601, w_000_602, w_000_603, w_000_604, w_000_605, w_000_606, w_000_607, w_000_608, w_000_609, w_000_610, w_000_611, w_000_612, w_000_613, w_000_614, w_000_615, w_000_616, w_000_617, w_000_618, w_000_619, w_000_620, w_000_621, w_000_622, w_000_623, w_000_624, w_000_625, w_000_626, w_000_627, w_000_628, w_000_629, w_000_630, w_000_631, w_000_632, w_000_633, w_000_634, w_000_635, w_000_636, w_000_637, w_000_638, w_000_639, w_000_640, w_000_641, w_000_642, w_000_643, w_000_644, w_000_645, w_000_646, w_000_647, w_000_648, w_000_649, w_000_650, w_000_651, w_000_652, w_000_653, w_000_654, w_000_655, w_000_656, w_000_657, w_000_658, w_000_659, w_000_660, w_000_661, w_000_662, w_000_663, w_000_664, w_000_665, w_000_666, w_000_667, w_000_668, w_000_669, w_000_670, w_000_671, w_000_672, w_000_673, w_000_674, w_000_675, w_000_676, w_000_677, w_000_678, w_000_679, w_000_680, w_000_681, w_000_682, w_000_683, w_000_684, w_000_685, w_000_686, w_000_687, w_000_688, w_000_689, w_000_690, w_000_691, w_000_692, w_000_693, w_000_694, w_000_695, w_000_696, w_000_697, w_000_698, w_000_699, w_000_700, w_000_701, w_000_702, w_000_703, w_000_704, w_000_705, w_000_706, w_000_707, w_000_708, w_000_709, w_000_710, w_000_711, w_000_712, w_000_713, w_000_714, w_000_715, w_000_716, w_000_717, w_000_718, w_000_719, w_000_720, w_000_721, w_000_722, w_000_723, w_000_724, w_000_725, w_000_726, w_000_727, w_000_728, w_000_729, w_000_730, w_000_731, w_000_732, w_000_733, w_000_734, w_000_735, w_000_736, w_000_737, w_000_738, w_000_739, w_000_740, w_000_741, w_000_742, w_000_743, w_000_744, w_000_745, w_000_746, w_000_747, w_000_748, w_000_749, w_000_750, w_000_751, w_000_752, w_000_753, w_000_754, w_000_755, w_000_756, w_000_757, w_000_758, w_000_759, w_000_760, w_000_761, w_000_762, w_000_763, w_000_764, w_000_765, w_000_766, w_000_767, w_000_768, w_000_769, w_000_770, w_000_771, w_000_772, w_000_773, w_000_774, w_000_775, w_000_776, w_000_777, w_000_778, w_000_779, w_000_780, w_000_781, w_000_782, w_000_783, w_000_784, w_000_785, w_000_786, w_000_787, w_000_788, w_000_789, w_000_790, w_000_791, w_000_792, w_000_793, w_000_794, w_000_795, w_000_796, w_000_797, w_000_798, w_000_799, w_000_800, w_000_801, w_000_802, w_000_803, w_000_804, w_000_805, w_000_806, w_000_807, w_000_808, w_000_809, w_000_810, w_000_811, w_000_812, w_000_813, w_000_814, w_000_815, w_000_816, w_000_817, w_000_818, w_000_819, w_000_820, w_000_821, w_000_822, w_000_823, w_000_824, w_000_825, w_000_826, w_000_827, w_000_828, w_000_829, w_000_830, w_000_831, w_000_832, w_000_833, w_000_834, w_000_835, w_000_836, w_000_837, w_000_838, w_000_839, w_000_840, w_000_841, w_000_842, w_000_843, w_000_844, w_000_845, w_000_846, w_000_847, w_000_848, w_000_849, w_000_850, w_000_851, w_000_852, w_000_853, w_000_854, w_000_855, w_000_856, w_000_857, w_000_858, w_000_859, w_000_860, w_000_861, w_000_862, w_000_863, w_000_864, w_000_865, w_000_866, w_000_867, w_000_868, w_000_869, w_000_870, w_000_871, w_000_872, w_000_873, w_000_874, w_000_875, w_000_876, w_000_877, w_000_878, w_000_879, w_000_880, w_000_881, w_000_882, w_000_883, w_000_884, w_000_885, w_000_886, w_000_887, w_000_888, w_000_889, w_000_890, w_000_891, w_000_892, w_000_893, w_000_894, w_000_895, w_000_896, w_000_897, w_000_898, w_000_899, w_000_900, w_000_901, w_000_902, w_000_903, w_000_904, w_000_905, w_000_906, w_000_907, w_000_908, w_000_909, w_000_910, w_000_911, w_000_912, w_000_913, w_000_914, w_000_915, w_000_916, w_000_917, w_000_918, w_000_919, w_000_920, w_000_921, w_000_922, w_000_923, w_000_924, w_000_925, w_000_926, w_000_927, w_000_928, w_000_929, w_000_930, w_000_931, w_000_932, w_000_933, w_000_934, w_000_935, w_000_936, w_000_937, w_000_938, w_000_939, w_000_940, w_000_941, w_000_942, w_000_943, w_000_944, w_000_945, w_000_946, w_000_947, w_000_948, w_000_949, w_000_950, w_000_951, w_000_952, w_000_953, w_000_954, w_000_955, w_000_956, w_000_957, w_000_958, w_000_959, w_000_960, w_000_961, w_000_962, w_000_963, w_000_964, w_000_965, w_000_966, w_000_967, w_000_968, w_000_969, w_000_970, w_000_971, w_000_972, w_000_973, w_000_974, w_000_975, w_000_976, w_000_977, w_000_978, w_000_979, w_000_980, w_000_981, w_000_982, w_000_983, w_000_984, w_000_985, w_000_986, w_000_987, w_000_988, w_000_989, w_000_990, w_000_991, w_000_992, w_000_993, w_000_994, w_000_995, w_000_996, w_000_997, w_000_998, w_000_999, w_000_1000, w_000_1001, w_000_1002, w_000_1003, w_000_1004, w_000_1005, w_000_1006, w_000_1007, w_000_1008, w_000_1009, w_000_1010, w_000_1011, w_000_1012, w_000_1013, w_000_1014, w_000_1015, w_000_1016, w_000_1017, w_000_1018, w_000_1019, w_000_1020, w_000_1021, w_000_1022, w_000_1023, w_000_1024, w_000_1025, w_000_1026, w_000_1027, w_000_1028, w_000_1029, w_000_1030, w_000_1031, w_000_1032, w_000_1033, w_000_1034, w_000_1035, w_000_1036, w_000_1037, w_000_1038, w_000_1039, w_000_1040, w_000_1041, w_000_1042, w_000_1043, w_000_1044, w_000_1045, w_000_1046, w_000_1047, w_000_1048, w_000_1049, w_000_1050, w_000_1051, w_000_1052, w_000_1053, w_000_1054, w_000_1055, w_000_1056, w_000_1057, w_000_1058, w_000_1059, w_000_1060, w_000_1061, w_000_1062, w_000_1063, w_000_1064, w_000_1065, w_000_1066, w_000_1067, w_000_1068, w_000_1069, w_000_1070, w_000_1071, w_000_1072, w_000_1073, w_000_1074, w_000_1075, w_000_1076, w_000_1077, w_000_1078, w_000_1079, w_000_1080, w_000_1081, w_000_1082, w_000_1083, w_000_1084, w_000_1085, w_000_1086, w_000_1087, w_000_1088, w_000_1089, w_000_1090, w_000_1091, w_000_1092, w_000_1093, w_000_1094, w_000_1095, w_000_1096, w_000_1097, w_000_1098, w_000_1099, w_000_1100, w_000_1101, w_000_1102, w_000_1103, w_000_1104, w_000_1105, w_000_1106, w_000_1107, w_000_1108, w_000_1109, w_000_1110, w_000_1111, w_000_1112, w_000_1113, w_000_1114, w_000_1115, w_000_1116, w_000_1117, w_000_1118, w_000_1119, w_000_1120, w_000_1121, w_000_1122, w_000_1123, w_000_1124, w_000_1125, w_000_1126, w_000_1127, w_000_1128, w_000_1129, w_000_1130, w_000_1131, w_000_1132, w_000_1133, w_000_1134, w_000_1135, w_000_1136, w_000_1137, w_000_1138, w_000_1139, w_000_1140, w_000_1141, w_000_1142, w_000_1143, w_000_1144, w_000_1145, w_000_1146, w_000_1147, w_000_1148, w_000_1149, w_000_1150, w_000_1151, w_000_1152, w_000_1153, w_000_1154, w_000_1155, w_000_1156, w_000_1157, w_000_1158, w_000_1159, w_000_1160, w_000_1161, w_000_1162, w_000_1163, w_000_1164, w_000_1165, w_000_1166, w_000_1167, w_000_1168, w_000_1169, w_000_1170, w_000_1171, w_000_1172, w_000_1173, w_000_1174, w_000_1175, w_000_1176, w_000_1177, w_000_1178, w_000_1179, w_000_1180, w_000_1181, w_000_1182, w_000_1183, w_000_1184, w_000_1185, w_000_1186, w_000_1187, w_000_1188, w_000_1189, w_000_1190, w_000_1191, w_000_1192, w_000_1193, w_000_1194, w_000_1195, w_000_1196, w_000_1197, w_000_1198, w_000_1199, w_000_1200, w_000_1201, w_000_1202, w_000_1203, w_000_1204, w_000_1205, w_000_1206, w_000_1207, w_000_1208, w_000_1209, w_000_1210, w_000_1211, w_000_1212, w_000_1213, w_000_1214, w_000_1215, w_000_1216, w_000_1217, w_000_1218, w_000_1219, w_000_1220, w_000_1221, w_000_1222, w_000_1223, w_000_1224, w_000_1225, w_000_1226, w_000_1227, w_000_1228, w_000_1229, w_000_1230, w_000_1231, w_000_1232, w_000_1233, w_000_1234, w_000_1235, w_000_1236, w_000_1237, w_000_1238, w_000_1239, w_000_1240, w_000_1241, w_000_1242, w_000_1243, w_000_1244, w_000_1245, w_000_1246, w_000_1247, w_000_1248, w_000_1249, w_000_1250, w_000_1251, w_000_1252, w_000_1253, w_000_1254, w_000_1255, w_000_1256, w_000_1257, w_000_1258, w_000_1259, w_000_1260, w_000_1261, w_000_1262, w_000_1263, w_000_1264, w_000_1265, w_000_1266, w_000_1267, w_000_1268, w_000_1269, w_000_1270, w_000_1271, w_000_1272, w_000_1273, w_000_1274, w_000_1275, w_000_1276, w_000_1277, w_000_1278, w_000_1279, w_000_1280, w_000_1281, w_000_1282, w_000_1283, w_000_1284, w_000_1285, w_000_1286, w_000_1287, w_000_1288, w_000_1289, w_000_1290, w_000_1291, w_000_1292, w_000_1293, w_000_1294, w_000_1295, w_000_1296, w_000_1297, w_000_1298, w_000_1299, w_000_1300, w_000_1301, w_000_1302, w_000_1303, w_000_1304, w_000_1305, w_000_1306, w_000_1307, w_000_1308, w_000_1309, w_000_1310, w_000_1311, w_000_1312, w_000_1313, w_000_1314, w_000_1315, w_000_1316, w_000_1317, w_000_1318, w_000_1319, w_000_1320, w_000_1321, w_000_1322, w_000_1323, w_000_1324, w_000_1325, w_000_1326, w_000_1327, w_000_1328, w_000_1329, w_000_1330, w_000_1331, w_000_1332, w_000_1333, w_000_1334, w_000_1335, w_000_1336, w_000_1337, w_000_1338, w_000_1339, w_000_1340, w_000_1341, w_000_1342, w_000_1343, w_000_1344, w_000_1345, w_000_1346, w_000_1347, w_000_1348, w_000_1349, w_000_1350, w_000_1351, w_000_1352, w_000_1353, w_000_1354, w_000_1355, w_000_1356, w_000_1357, w_000_1358, w_000_1359, w_000_1360, w_000_1361, w_000_1362, w_000_1363, w_000_1364, w_000_1365, w_000_1366, w_000_1367, w_000_1368, w_000_1369, w_000_1370, w_000_1371, w_000_1372, w_000_1373, w_000_1374, w_000_1375, w_000_1376, w_000_1377, w_000_1378, w_000_1379, w_000_1380, w_000_1381, w_000_1382, w_000_1383, w_000_1384, w_000_1385, w_000_1386, w_000_1387, w_000_1388, w_000_1389, w_000_1390, w_000_1391, w_000_1392, w_000_1393, w_000_1394, w_000_1395, w_000_1396, w_000_1397, w_000_1398, w_000_1399, w_000_1400, w_000_1401, w_000_1402, w_000_1403, w_000_1404, w_000_1405, w_000_1406, w_000_1407, w_000_1408, w_000_1409, w_000_1410, w_000_1411, w_000_1412, w_000_1413, w_000_1414, w_000_1415, w_000_1416, w_000_1417, w_000_1418, w_000_1419, w_000_1420, w_000_1421, w_000_1422, w_000_1423, w_000_1424, w_000_1425, w_000_1426, w_000_1427, w_000_1428, w_000_1429, w_000_1430, w_000_1431, w_000_1432, w_000_1433, w_000_1434, w_000_1435, w_000_1436, w_000_1437, w_000_1438, w_000_1439, w_000_1440, w_000_1441, w_000_1442, w_000_1443, w_000_1444, w_000_1445, w_000_1446, w_000_1447, w_000_1448, w_000_1449, w_000_1450, w_000_1451, w_000_1452, w_000_1453, w_000_1454, w_000_1455, w_000_1456, w_000_1457, w_000_1458, w_000_1459, w_000_1460, w_000_1461, w_000_1462, w_000_1463, w_000_1464, w_000_1465, w_000_1466, w_000_1467, w_000_1468, w_000_1469, w_000_1470, w_000_1471, w_000_1472, w_000_1473, w_000_1474, w_000_1475, w_000_1476, w_000_1477, w_000_1478, w_000_1479, w_000_1480, w_000_1481, w_000_1482, w_000_1483, w_000_1484, w_000_1485, w_000_1486, w_000_1487, w_000_1488, w_000_1489, w_000_1490, w_000_1491, w_000_1492, w_000_1493, w_000_1494, w_000_1495, w_000_1496, w_000_1497, w_000_1498, w_000_1499, w_000_1500, w_000_1501, w_000_1502, w_000_1503, w_000_1504, w_000_1505, w_000_1506, w_000_1507, w_000_1508, w_000_1509, w_000_1510, w_000_1511, w_000_1512, w_000_1513, w_000_1514, w_000_1515, w_000_1516, w_000_1517, w_000_1518, w_000_1519, w_000_1520, w_000_1521, w_000_1522, w_000_1523, w_000_1524, w_000_1525, w_000_1526, w_000_1527, w_000_1528, w_000_1529, w_000_1530, w_000_1531, w_000_1532, w_000_1533, w_000_1534, w_000_1535, w_000_1536, w_000_1537, w_000_1538, w_000_1539, w_000_1540, w_000_1541, w_000_1542, w_000_1543, w_000_1544, w_000_1545, w_000_1546, w_000_1547, w_000_1548, w_000_1549, w_000_1550, w_000_1551, w_000_1552, w_000_1553, w_000_1554, w_000_1555, w_000_1556, w_000_1557, w_000_1558, w_000_1559, w_000_1560, w_000_1561, w_000_1562, w_000_1563, w_000_1564, w_000_1565, w_000_1566, w_000_1567, w_000_1568, w_000_1569, w_000_1570, w_000_1571, w_000_1572, w_000_1573, w_000_1574, w_000_1575, w_000_1576, w_000_1577, w_000_1578, w_000_1579, w_000_1580, w_000_1581, w_000_1582, w_000_1583, w_000_1584, w_000_1585, w_000_1586, w_000_1587, w_000_1588, w_000_1589, w_000_1590, w_000_1591, w_000_1592, w_000_1593, w_000_1594, w_000_1595, w_000_1596, w_000_1597, w_000_1598, w_000_1599, w_000_1600, w_000_1601, w_000_1602, w_000_1603, w_000_1604, w_000_1605, w_000_1606, w_000_1607, w_000_1608, w_000_1609, w_000_1610, w_000_1611, w_000_1612, w_000_1613, w_000_1614, w_000_1615, w_000_1616, w_000_1617, w_000_1618, w_000_1619, w_000_1620, w_000_1621, w_000_1622, w_000_1623, w_000_1624, w_000_1625, w_000_1626, w_000_1627, w_000_1628, w_000_1629, w_000_1630, w_000_1631, w_000_1632, w_000_1633, w_000_1634, w_000_1635, w_000_1636, w_000_1637, w_000_1638, w_000_1639, w_000_1640, w_000_1641, w_000_1642, w_000_1643, w_000_1644, w_000_1645, w_000_1646, w_000_1647, w_000_1648, w_000_1649, w_000_1650, w_000_1651, w_000_1652, w_000_1653, w_000_1654, w_000_1655, w_000_1656, w_000_1657, w_000_1658, w_000_1659, w_000_1660, w_000_1661, w_000_1662, w_000_1663, w_000_1664, w_000_1665, w_000_1666, w_000_1667, w_000_1668, w_000_1669, w_000_1670, w_000_1671, w_000_1672, w_000_1673, w_000_1674, w_000_1675, w_000_1676, w_000_1677, w_000_1678, w_000_1679, w_000_1680, w_000_1681, w_000_1682, w_000_1683, w_000_1684, w_000_1685, w_000_1686, w_000_1687, w_000_1688, w_000_1689, w_000_1690, w_000_1691, w_000_1692, w_000_1693, w_000_1694, w_000_1695, w_000_1696, w_000_1697, w_000_1698, w_000_1699, w_000_1700, w_000_1701, w_000_1702, w_000_1703, w_000_1704, w_000_1705, w_000_1706, w_000_1707, w_000_1708, w_000_1709, w_000_1710, w_000_1711, w_000_1712, w_000_1713, w_000_1714, w_000_1715, w_000_1716, w_000_1717, w_000_1718, w_000_1719, w_000_1720, w_000_1721, w_000_1722, w_000_1723, w_000_1724, w_000_1725, w_000_1726, w_000_1727, w_000_1728, w_000_1729, w_000_1730, w_000_1731, w_000_1732, w_000_1733, w_000_1734, w_000_1735, w_000_1736, w_000_1737, w_000_1738, w_000_1739, w_000_1740, w_000_1741, w_000_1742, w_000_1743, w_000_1744, w_000_1745, w_000_1746, w_000_1747, w_000_1748, w_000_1749, w_000_1750, w_000_1751, w_000_1752, w_000_1753, w_000_1754, w_000_1755, w_000_1756, w_000_1757, w_000_1758, w_000_1759, w_000_1760, w_000_1761, w_000_1762, w_000_1763, w_000_1764, w_000_1765, w_000_1766, w_000_1767, w_000_1768, w_000_1769, w_000_1770, w_000_1771, w_000_1772, w_000_1773, w_000_1774, w_000_1775, w_000_1776, w_000_1777, w_000_1778, w_000_1779, w_000_1780, w_000_1781, w_000_1782, w_000_1783, w_000_1784, w_000_1785, w_000_1786, w_000_1787, w_000_1788, w_000_1789, w_000_1790, w_000_1791, w_000_1792, w_000_1793, w_000_1794, w_000_1795, w_000_1796, w_000_1797, w_000_1798, w_000_1799, w_000_1800, w_000_1801, w_000_1802, w_000_1803, w_000_1804, w_000_1805, w_000_1806, w_000_1807, w_000_1808, w_000_1809, w_000_1810, w_000_1811, w_000_1812, w_000_1813, w_000_1814, w_000_1815, w_000_1816, w_000_1817, w_000_1818, w_000_1819, w_000_1820, w_000_1821, w_000_1822, w_000_1823, w_000_1824, w_000_1825, w_000_1826, w_000_1827, w_000_1828, w_000_1829, w_000_1830, w_000_1831, w_000_1832, w_000_1833, w_000_1834, w_000_1835, w_000_1836, w_000_1837, w_000_1838, w_000_1839, w_000_1840, w_000_1841, w_000_1842, w_000_1843, w_000_1844, w_000_1845, w_000_1846, w_000_1847, w_000_1848, w_000_1849, w_000_1850, w_000_1851, w_000_1852, w_000_1853, w_000_1854, w_000_1855, w_000_1856, w_000_1857, w_000_1858, w_000_1859, w_000_1860, w_000_1861, w_000_1862, w_000_1863, w_000_1864, w_000_1865, w_000_1866, w_000_1867, w_000_1868, w_000_1869, w_000_1870, w_000_1871, w_000_1872, w_000_1873, w_000_1874, w_000_1875, w_000_1876, w_000_1877, w_000_1878, w_000_1879, w_000_1880, w_000_1881, w_000_1882, w_000_1883, w_000_1884, w_000_1885, w_000_1886, w_000_1887, w_000_1888, w_000_1889, w_000_1890, w_000_1891, w_000_1892, w_000_1893, w_000_1894, w_000_1895, w_000_1896, w_000_1897, w_000_1898, w_000_1899, w_000_1900, w_000_1901, w_000_1902, w_000_1903, w_000_1904, w_000_1905, w_000_1906, w_000_1907, w_000_1908, w_000_1909, w_000_1910, w_000_1911, w_000_1912, w_000_1913, w_000_1914, w_000_1915, w_000_1916, w_000_1917, w_000_1918, w_000_1919, w_000_1920, w_000_1921, w_000_1922, w_000_1923, w_000_1924, w_000_1925, w_000_1926, w_000_1927, w_000_1928, w_000_1929, w_000_1930, w_000_1931, w_000_1932, w_000_1933, w_000_1934, w_000_1935, w_000_1936, w_000_1937, w_000_1938, w_000_1939, w_000_1940, w_000_1941, w_000_1942, w_000_1943, w_000_1944, w_000_1945, w_000_1946, w_000_1947, w_000_1948, w_000_1949, w_000_1950, w_000_1951, w_000_1952, w_000_1953, w_000_1954, w_000_1955, w_000_1956, w_000_1957, w_000_1958, w_000_1959, w_000_1960, w_000_1961, w_000_1962, w_000_1963, w_000_1964, w_000_1965, w_000_1966, w_000_1967, w_000_1968, w_000_1969, w_000_1970, w_000_1971, w_000_1972, w_000_1973, w_000_1974, w_000_1975, w_000_1976, w_000_1977, w_000_1978, w_000_1979, w_000_1980, w_000_1981, w_000_1982, w_000_1983, w_000_1984, w_000_1985, w_000_1986, w_000_1987, w_000_1988, w_000_1989, w_000_1990, w_000_1991, w_000_1992, w_000_1993, w_000_1994, w_000_1995, w_000_1996, w_000_1997, w_000_1998, w_000_1999, w_000_2000, w_000_2001, w_000_2002, w_000_2003, w_000_2004, w_000_2005, w_000_2006, w_000_2007, w_000_2008, w_000_2009, w_000_2010, w_000_2011, w_000_2012, w_000_2013, w_000_2014, w_000_2015, w_000_2016, w_000_2017, w_000_2018, w_000_2019, w_000_2020, w_000_2021, w_000_2022, w_000_2023, w_000_2024, w_000_2025, w_000_2026, w_000_2027, w_000_2028, w_000_2029, w_000_2030, w_000_2031, w_000_2032, w_000_2033, w_000_2034, w_000_2035, w_000_2036, w_000_2037, w_000_2038, w_000_2039, w_000_2040, w_000_2041, w_000_2042, w_000_2043, w_000_2044, w_000_2045, w_000_2046, w_000_2047, w_000_2048, w_000_2049, w_000_2050, w_000_2051, w_000_2052, w_000_2053, w_000_2054, w_000_2055, w_000_2056, w_000_2057, w_000_2058, w_000_2059, w_000_2060, w_000_2061, w_000_2062, w_000_2063, w_000_2064, w_000_2065, w_000_2066, w_000_2067, w_000_2068, w_000_2069, w_000_2070, w_000_2071, w_000_2072, w_000_2073, w_000_2074, w_000_2075, w_000_2076, w_000_2077, w_000_2078, w_000_2079, w_000_2080, w_000_2081, w_000_2082, w_000_2083, w_000_2084, w_000_2085, w_000_2086, w_000_2087, w_000_2088, w_000_2089, w_000_2090, w_000_2091, w_000_2092, w_000_2093, w_000_2094, w_000_2095, w_000_2096, w_000_2097, w_000_2098, w_000_2099, w_000_2100, w_000_2101, w_000_2102, w_000_2103, w_000_2104, w_000_2105, w_000_2106, w_000_2107, w_000_2108, w_000_2109, w_000_2110, w_000_2111, w_000_2112, w_000_2113, w_000_2114, w_000_2115, w_000_2116, w_000_2117, w_000_2118, w_000_2119, w_000_2120, w_000_2121, w_000_2122, w_000_2123, w_000_2124, w_000_2125, w_000_2126, w_000_2127, w_000_2128, w_000_2129, w_000_2130, w_000_2131, w_000_2132, w_000_2133, w_000_2134, w_000_2135, w_000_2136, w_000_2137, w_000_2138, w_000_2139, w_000_2140, w_000_2141, w_000_2142, w_000_2143, w_000_2144, w_000_2145, w_000_2146, w_000_2147, w_000_2148, w_000_2149, w_000_2150, w_000_2151, w_000_2152, w_000_2153, w_000_2154, w_000_2155, w_000_2156, w_000_2157, w_000_2158, w_000_2159, w_000_2160, w_000_2161, w_000_2162, w_000_2163, w_000_2164, w_000_2165, w_000_2166, w_000_2167, w_000_2168, w_000_2169, w_000_2170, w_000_2171, w_000_2172, w_000_2173, w_000_2174, w_000_2175, w_000_2176, w_000_2177, w_000_2178, w_000_2179, w_000_2180, w_000_2181, w_000_2182, w_000_2183, w_000_2184, w_000_2185, w_000_2186, w_000_2187, w_000_2188, w_000_2189, w_000_2190, w_000_2191, w_000_2192, w_000_2193, w_000_2194, w_000_2195, w_000_2196, w_000_2197, w_000_2198, w_000_2199, w_000_2200, w_000_2201, w_000_2202, w_000_2203, w_000_2204, w_000_2205, w_000_2206, w_000_2207, w_000_2208, w_000_2209, w_000_2210, w_000_2211, w_000_2212, w_000_2213, w_000_2214, w_000_2215, w_000_2216, w_000_2217, w_000_2218, w_000_2219, w_000_2220, w_000_2221, w_000_2222, w_000_2223, w_000_2224, w_000_2225, w_000_2226, w_000_2227, w_000_2228, w_000_2229, w_000_2230, w_000_2231, w_000_2232, w_000_2233, w_000_2234, w_000_2235, w_000_2236, w_000_2237, w_000_2238, w_000_2239, w_000_2240, w_000_2241, w_000_2242, w_000_2243, w_000_2244, w_000_2245, w_000_2246, w_000_2247, w_000_2248, w_000_2249, w_000_2250, w_000_2251, w_000_2252, w_000_2253, w_000_2254, w_000_2255, w_000_2256, w_000_2257, w_000_2258, w_000_2259, w_000_2260, w_000_2261, w_000_2262, w_000_2263, w_000_2264, w_000_2265, w_000_2266, w_000_2267, w_000_2268, w_000_2269, w_000_2270, w_000_2271, w_000_2272, w_000_2273, w_000_2274, w_000_2275, w_000_2276, w_000_2277, w_000_2278, w_000_2279, w_000_2280, w_000_2281, w_000_2282, w_000_2283, w_000_2284, w_000_2285, w_000_2286, w_000_2287, w_000_2288, w_000_2289, w_000_2290, w_000_2291, w_000_2292, w_000_2293, w_000_2294, w_000_2295, w_000_2296, w_000_2297, w_000_2298, w_000_2299, w_000_2300, w_000_2301, w_000_2302, w_000_2303, w_000_2304, w_000_2305, w_000_2306, w_000_2307, w_000_2308, w_000_2309, w_000_2310, w_000_2311, w_000_2312, w_000_2313, w_000_2314, w_000_2315, w_000_2316, w_000_2317, w_000_2318, w_000_2319, w_000_2320, w_000_2321, w_000_2322, w_000_2323, w_000_2324, w_000_2325, w_000_2326, w_000_2327, w_000_2328, w_000_2329, w_000_2330, w_000_2331, w_000_2332, w_000_2333, w_000_2334, w_000_2335, w_000_2336, w_000_2337, w_000_2338, w_000_2339, w_000_2340, w_000_2341, w_000_2342, w_000_2343, w_000_2344, w_000_2345, w_000_2346, w_000_2347, w_000_2348, w_000_2349, w_000_2350, w_000_2351, w_000_2352, w_000_2353, w_000_2354, w_000_2355, w_000_2356, w_000_2357, w_000_2358, w_000_2359, w_000_2360, w_000_2361, w_000_2362, w_000_2363, w_000_2364, w_000_2365, w_000_2366, w_000_2367, w_000_2368, w_000_2369, w_000_2370, w_000_2371, w_000_2372, w_000_2373, w_000_2374, w_000_2375, w_000_2376, w_000_2377, w_000_2378, w_000_2379, w_000_2380, w_000_2381, w_000_2382, w_000_2383, w_000_2384, w_000_2385, w_000_2386, w_000_2387, w_000_2388, w_000_2389, w_000_2390, w_000_2391, w_000_2392, w_000_2393, w_000_2394, w_000_2395, w_000_2396, w_000_2397, w_000_2398, w_000_2399, w_000_2400, w_000_2401, w_000_2402, w_000_2403, w_000_2404, w_000_2405, w_000_2406, w_000_2407, w_000_2408, w_000_2409, w_000_2410, w_000_2411, w_000_2412, w_000_2413, w_000_2414, w_000_2415, w_000_2416, w_000_2417, w_000_2418, w_000_2419, w_000_2420, w_000_2421, w_000_2422, w_000_2423, w_000_2424, w_000_2425, w_000_2426, w_000_2427, w_000_2428, w_000_2429, w_000_2430, w_000_2431, w_000_2432, w_000_2433, w_000_2434, w_000_2435, w_000_2436, w_000_2437, w_000_2438, w_000_2439, w_000_2440, w_000_2441, w_000_2442, w_000_2443, w_000_2444, w_000_2445, w_000_2446, w_000_2447, w_000_2448, w_000_2449, w_000_2450, w_000_2451, w_000_2452, w_000_2453, w_000_2454, w_000_2455, w_000_2456, w_000_2457, w_000_2458, w_000_2459, w_000_2460, w_000_2461, w_000_2462, w_000_2463, w_000_2464, w_000_2465, w_000_2466, w_000_2467, w_000_2468, w_000_2469, w_000_2470, w_000_2471, w_000_2472, w_000_2473, w_000_2474, w_000_2475, w_000_2476, w_000_2477, w_000_2478, w_000_2479, w_000_2480, w_000_2481, w_000_2482, w_000_2483, w_000_2484, w_000_2485, w_000_2486, w_000_2487, w_000_2488, w_000_2489, w_000_2490, w_000_2491, w_000_2492, w_000_2493, w_000_2494, w_000_2495, w_000_2496, w_000_2497, w_000_2498, w_000_2499, w_000_2500, w_000_2501, w_000_2502, w_000_2503, w_000_2504, w_000_2505, w_000_2506, w_000_2507, w_000_2508, w_000_2509, w_000_2510, w_000_2511, w_000_2512, w_000_2513, w_000_2514, w_000_2515, w_000_2516, w_000_2517, w_000_2518, w_000_2519, w_000_2520, w_000_2521, w_000_2522, w_000_2523, w_000_2524, w_000_2525, w_000_2526, w_000_2527, w_000_2528, w_000_2529, w_000_2530, w_000_2531, w_000_2532, w_000_2533, w_000_2534, w_000_2535, w_000_2536, w_000_2537, w_000_2538, w_000_2539, w_000_2540, w_000_2541, w_000_2542, w_000_2543, w_000_2544, w_000_2545, w_000_2546, w_000_2547, w_000_2548, w_000_2549, w_000_2550, w_000_2551, w_000_2552, w_000_2553, w_000_2554, w_000_2555, w_000_2556, w_000_2557, w_000_2558, w_000_2559, w_000_2560, w_000_2561, w_000_2562, w_000_2563, w_000_2564, w_000_2565, w_000_2566, w_000_2567, w_000_2568, w_000_2569, w_000_2570, w_000_2571, w_000_2572, w_000_2573, w_000_2574, w_000_2575, w_000_2576, w_000_2577, w_000_2578, w_000_2579, w_000_2580, w_000_2581, w_000_2582, w_000_2583, w_000_2584, w_000_2585, w_000_2586, w_000_2587, w_000_2588, w_000_2589, w_000_2590, w_000_2591, w_000_2592, w_000_2593, w_000_2594, w_000_2595, w_000_2596, w_000_2597, w_000_2598, w_000_2599, w_000_2600, w_000_2601, w_000_2602, w_000_2603, w_000_2604, w_000_2605, w_000_2606, w_000_2607, w_000_2608, w_000_2609, w_000_2610, w_000_2611, w_000_2612, w_000_2613, w_000_2614, w_000_2615, w_000_2616, w_000_2617, w_000_2618, w_000_2619, w_000_2620, w_000_2621, w_000_2622, w_000_2623, w_000_2624, w_000_2625, w_000_2626, w_000_2627, w_000_2628, w_000_2629, w_000_2630, w_000_2631, w_000_2632, w_000_2633, w_000_2634, w_000_2635, w_000_2636, w_000_2637, w_000_2638, w_000_2639, w_000_2640, w_000_2641, w_000_2642, w_000_2643, w_000_2644, w_000_2645, w_000_2646, w_000_2647, w_000_2648, w_000_2649, w_000_2650, w_000_2651, w_000_2652, w_000_2653, w_000_2654, w_000_2655, w_000_2656, w_000_2657, w_000_2658, w_000_2659, w_000_2660, w_000_2661, w_000_2662, w_000_2663, w_000_2664, w_000_2665, w_000_2666, w_000_2667, w_000_2668, w_000_2669, w_000_2670, w_000_2671, w_000_2672, w_000_2673, w_000_2674, w_000_2675, w_000_2676, w_000_2677, w_000_2678, w_000_2679, w_000_2680, w_000_2681, w_000_2682, w_000_2683, w_000_2684, w_000_2685, w_000_2686, w_000_2687, w_000_2688, w_000_2689, w_000_2690, w_000_2691, w_000_2692, w_000_2693, w_000_2694, w_000_2695, w_000_2696, w_000_2697, w_000_2698, w_000_2699, w_000_2700, w_000_2701, w_000_2702, w_000_2703, w_000_2704, w_000_2705, w_000_2706, w_000_2707, w_000_2708, w_000_2709, w_000_2710, w_000_2711, w_000_2712, w_000_2713, w_000_2714, w_000_2715, w_000_2716, w_000_2717, w_000_2718, w_000_2719, w_000_2720, w_000_2721, w_000_2722, w_000_2723, w_000_2724, w_000_2725, w_000_2726, w_000_2727, w_000_2728, w_000_2729, w_000_2730, w_000_2731, w_000_2732, w_000_2733, w_000_2734, w_000_2735, w_000_2736, w_000_2737, w_000_2738, w_000_2739, w_000_2740, w_000_2741, w_000_2742, w_000_2743, w_000_2744, w_000_2745, w_000_2746, w_000_2747, w_000_2748, w_000_2749, w_000_2750, w_000_2751, w_000_2752, w_000_2753, w_000_2754, w_000_2755, w_000_2756, w_000_2757, w_000_2758, w_000_2759, w_000_2760, w_000_2761, w_000_2762, w_000_2763, w_000_2764, w_000_2765, w_000_2766, w_000_2767, w_000_2768, w_000_2769, w_000_2770, w_000_2771, w_000_2772, w_000_2773, w_000_2774, w_000_2775, w_000_2776, w_000_2777, w_000_2778, w_000_2779, w_000_2780, w_000_2781, w_000_2782, w_000_2783, w_000_2784, w_000_2785, w_000_2786, w_000_2787, w_000_2788, w_000_2789, w_000_2790, w_000_2791, w_000_2792, w_000_2793, w_000_2794, w_000_2795, w_000_2796, w_000_2797, w_000_2798, w_000_2799, w_000_2800, w_000_2801, w_000_2802, w_000_2803, w_000_2804, w_000_2805, w_000_2806, w_000_2807, w_000_2808, w_000_2809, w_000_2810, w_000_2811, w_000_2812, w_000_2813, w_000_2814, w_000_2815, w_000_2816, w_000_2817, w_000_2818, w_000_2819, w_000_2820, w_000_2821, w_000_2822, w_000_2823, w_000_2824, w_000_2825, w_000_2826, w_000_2827, w_000_2828, w_000_2829, w_000_2830, w_000_2831, w_000_2832, w_000_2833, w_000_2834, w_000_2835, w_000_2836, w_000_2837, w_000_2838, w_000_2839, w_000_2840, w_000_2841, w_000_2842, w_000_2843, w_000_2844, w_000_2845, w_000_2846, w_000_2847, w_000_2848, w_000_2849, w_000_2850, w_000_2851, w_000_2852, w_000_2853, w_000_2854, w_000_2855, w_000_2856, w_000_2857, w_000_2858, w_000_2859, w_000_2860, w_000_2861, w_000_2862, w_000_2863, w_000_2864, w_000_2865, w_000_2866, w_000_2867, w_000_2868, w_000_2869, w_000_2870, w_000_2871, w_000_2872, w_000_2873, w_000_2874, w_000_2875, w_000_2876, w_000_2877, w_000_2878, w_000_2879, w_000_2880, w_000_2881, w_000_2882, w_000_2883, w_000_2884, w_000_2885, w_000_2886, w_000_2887, w_000_2888, w_000_2889, w_000_2890, w_000_2891, w_000_2892, w_000_2893, w_000_2894, w_000_2895, w_000_2896, w_000_2897, w_000_2898, w_000_2899, w_000_2900, w_000_2901, w_000_2902, w_000_2903, w_000_2904, w_000_2905, w_000_2906, w_000_2907, w_000_2908, w_000_2909, w_000_2910, w_000_2911, w_000_2912, w_000_2913, w_000_2914, w_000_2915, w_000_2916, w_000_2917, w_000_2918, w_000_2919, w_000_2920, w_000_2921, w_000_2922, w_000_2923, w_000_2924, w_000_2925, w_000_2926, w_000_2927, w_000_2928, w_000_2929, w_000_2930, w_000_2931, w_000_2932, w_000_2933, w_000_2934, w_000_2935, w_000_2936, w_000_2937, w_000_2938, w_000_2939, w_000_2940, w_000_2941, w_000_2942, w_000_2943, w_000_2944, w_000_2945, w_000_2946, w_000_2947, w_000_2948, w_000_2949, w_000_2950, w_000_2951, w_000_2952, w_000_2953, w_000_2954, w_000_2955, w_000_2956, w_000_2957, w_000_2958, w_000_2959, w_000_2960, w_000_2961, w_000_2962, w_000_2963, w_000_2964, w_000_2965, w_000_2966, w_000_2967, w_000_2968, w_000_2969, w_000_2970, w_000_2971, w_000_2972, w_000_2973, w_000_2974, w_000_2975, w_000_2976, w_000_2977, w_000_2978, w_000_2979, w_000_2980, w_000_2981, w_000_2982, w_000_2983, w_000_2984, w_000_2985, w_000_2986, w_000_2987, w_000_2988, w_000_2989, w_000_2990, w_000_2991, w_000_2992, w_000_2993, w_000_2994, w_000_2995, w_000_2996, w_000_2997, w_000_2998, w_000_2999, w_000_3000, w_000_3001, w_000_3002, w_000_3003, w_000_3004, w_000_3005, w_000_3006, w_000_3007, w_000_3008, w_000_3009, w_000_3010, w_000_3011, w_000_3012, w_000_3013, w_000_3014, w_000_3015, w_000_3016, w_000_3017, w_000_3019, w_000_3020, w_000_3021, w_000_3022, w_000_3023, w_000_3024, w_000_3025, w_000_3026, w_000_3027, w_000_3028, w_000_3029, w_000_3030, w_000_3031, w_000_3032, w_000_3033, w_000_3034, w_000_3035, w_000_3036, w_000_3037, w_000_3038, w_000_3039, w_000_3040, w_000_3041, w_000_3042, w_000_3043, w_000_3044, w_000_3045, w_000_3046, w_000_3047, w_000_3048, w_000_3049, w_000_3050, w_000_3051, w_000_3052, w_000_3053, w_000_3054, w_000_3055, w_000_3056, w_000_3057, w_000_3058, w_000_3059, w_000_3060, w_000_3061, w_000_3062, w_000_3063, w_000_3064, w_000_3065, w_000_3066, w_000_3067, w_000_3068, w_000_3069, w_000_3070, w_000_3071, w_000_3072, w_000_3073, w_000_3074, w_000_3075, w_000_3076, w_000_3077, w_000_3078, w_000_3079, w_000_3080, w_000_3081, w_000_3082, w_000_3083, w_000_3084, w_000_3085, w_000_3086, w_000_3087, w_000_3088, w_000_3089, w_000_3090, w_000_3091, w_000_3092, w_000_3093, w_000_3094, w_000_3095, w_000_3096, w_000_3097, w_000_3098, w_000_3099, w_000_3100, w_000_3101, w_000_3102, w_000_3103, w_000_3104, w_000_3105, w_000_3106, w_000_3107, w_000_3108, w_000_3109, w_000_3110, w_000_3111, w_000_3112, w_000_3113, w_000_3114, w_000_3115, w_000_3116, w_000_3117, w_000_3118, w_000_3119, w_000_3120, w_000_3121, w_000_3122, w_000_3123, w_000_3124, w_000_3125, w_000_3126, w_000_3127, w_000_3128, w_000_3129, w_000_3130, w_000_3131, w_000_3132, w_000_3133, w_000_3134, w_000_3135, w_000_3136, w_000_3137, w_000_3138, w_000_3139, w_000_3140, w_000_3141, w_000_3142, w_000_3143, w_000_3144, w_000_3145, w_000_3146, w_000_3147, w_000_3148, w_000_3149, w_000_3150, w_000_3151, w_000_3152, w_000_3153, w_000_3154, w_000_3155, w_000_3156, w_000_3157, w_000_3158, w_000_3159, w_000_3160, w_000_3161, w_000_3162, w_000_3163, w_000_3164, w_000_3165, w_000_3166, w_000_3167, w_000_3168, w_000_3169, w_000_3170, w_000_3171, w_000_3172, w_000_3173, w_000_3174, w_000_3175, w_000_3176, w_000_3177, w_000_3178, w_000_3179, w_000_3180, w_000_3181, w_000_3182, w_000_3183, w_000_3184, w_000_3185, w_000_3186, w_000_3187, w_000_3188, w_000_3189, w_000_3190, w_000_3191, w_000_3192, w_000_3193, w_000_3194, w_000_3195, w_000_3196, w_000_3197, w_000_3198, w_000_3199, w_000_3200, w_000_3201, w_000_3202, w_000_3203, w_000_3204, w_000_3205, w_000_3206, w_000_3207, w_000_3208, w_000_3209, w_000_3210, w_000_3211, w_000_3212, w_000_3213, w_000_3214, w_000_3215, w_000_3216, w_000_3217, w_000_3218, w_000_3219, w_000_3220, w_000_3221, w_000_3222, w_000_3223, w_000_3224, w_000_3225, w_000_3226, w_000_3227, w_000_3228, w_000_3229, w_000_3230, w_000_3231, w_000_3232, w_000_3233, w_000_3234, w_000_3235, w_000_3236, w_000_3237, w_000_3238, w_000_3239, w_000_3240, w_000_3241, w_000_3242, w_000_3243, w_000_3244, w_000_3245, w_000_3246, w_000_3247, w_000_3248, w_000_3249, w_000_3250, w_000_3251, w_000_3252, w_000_3253, w_000_3254, w_000_3255, w_000_3256, w_000_3257, w_000_3258, w_000_3259, w_000_3260, w_000_3261, w_000_3262, w_000_3263, w_000_3264, w_000_3265, w_000_3266, w_000_3267, w_000_3268, w_000_3269, w_000_3270, w_000_3271, w_000_3272, w_000_3273, w_000_3274, w_000_3275, w_000_3276, w_000_3277, w_000_3278, w_000_3279, w_000_3280, w_000_3281, w_000_3282, w_000_3283, w_000_3284, w_000_3285, w_000_3286, w_000_3287, w_000_3288, w_000_3289, w_000_3290, w_000_3291, w_000_3292, w_000_3293, w_000_3294, w_000_3295, w_000_3296, w_000_3297, w_000_3298, w_000_3299, w_000_3300, w_000_3301, w_000_3302, w_000_3303, w_000_3304, w_000_3305, w_000_3306, w_000_3307, w_000_3308, w_000_3309, w_000_3310, w_000_3311, w_000_3312, w_000_3313, w_000_3314, w_000_3315, w_000_3316, w_000_3317, w_000_3318, w_000_3319, w_000_3320, w_000_3321, w_000_3322, w_000_3323, w_000_3324, w_000_3325, w_000_3326, w_000_3327, w_000_3328, w_000_3329, w_000_3330, w_000_3331, w_000_3332, w_000_3333, w_000_3334, w_000_3335, w_000_3336, w_000_3337, w_000_3338, w_000_3339, w_000_3340, w_000_3341, w_000_3342, w_000_3343, w_000_3344, w_000_3345, w_000_3346, w_000_3347, w_000_3348, w_000_3349, w_000_3350, w_000_3351, w_000_3352, w_000_3353, w_000_3354, w_000_3355, w_000_3356, w_000_3357, w_000_3358, w_000_3359, w_000_3360, w_000_3361, w_000_3362, w_000_3363, w_000_3364, w_000_3365, w_000_3366, w_000_3367, w_000_3368, w_000_3369, w_000_3370, w_000_3371, w_000_3372, w_000_3373, w_000_3374, w_000_3375, w_000_3376, w_000_3377, w_000_3378, w_000_3379, w_000_3380, w_000_3381, w_000_3382, w_000_3383, w_000_3384, w_000_3385, w_000_3386, w_000_3387, w_000_3388, w_000_3389, w_000_3390, w_000_3391, w_000_3392, w_000_3393, w_000_3394, w_000_3395, w_000_3396, w_000_3397, w_000_3398, w_000_3399, w_000_3400, w_000_3401, w_000_3402, w_000_3403, w_000_3404, w_000_3405, w_000_3406, w_000_3407, w_000_3408, w_000_3409, w_000_3410, w_000_3411, w_000_3412, w_000_3413, w_000_3414, w_000_3415, w_000_3416, w_000_3417, w_000_3418, w_000_3419, w_000_3420, w_000_3421, w_000_3422, w_000_3423, w_000_3424, w_000_3425, w_000_3426, w_000_3427, w_000_3428, w_000_3429, w_000_3430, w_000_3431, w_000_3432, w_000_3433, w_000_3434, w_000_3435, w_000_3436, w_000_3437, w_000_3438, w_000_3439, w_000_3440, w_000_3441, w_000_3442, w_000_3443, w_000_3444, w_000_3445, w_000_3446, w_000_3447, w_000_3448, w_000_3449, w_000_3450, w_000_3451, w_000_3452, w_000_3453, w_000_3454, w_000_3455, w_000_3456, w_000_3457, w_000_3458, w_000_3459, w_000_3460, w_000_3461, w_000_3462, w_000_3463, w_000_3464, w_000_3465, w_000_3466, w_000_3467, w_000_3468, w_000_3469, w_000_3470, w_000_3471, w_000_3472, w_000_3473, w_000_3474, w_000_3475, w_000_3476, w_000_3477, w_000_3478, w_000_3479, w_000_3480, w_000_3481, w_000_3482, w_000_3483, w_000_3484, w_000_3485, w_000_3486, w_000_3487, w_000_3488, w_000_3489, w_000_3490, w_000_3491, w_000_3492, w_000_3493, w_000_3494, w_000_3495, w_000_3496, w_000_3497, w_000_3498, w_000_3499, w_000_3500, w_000_3501, w_000_3502, w_000_3503, w_000_3504, w_000_3505, w_000_3506, w_000_3507, w_000_3508, w_000_3509, w_000_3510, w_000_3511, w_000_3512, w_000_3513, w_000_3514, w_000_3515, w_000_3516, w_000_3517, w_000_3518, w_000_3519, w_000_3520, w_000_3521, w_000_3522, w_000_3523, w_000_3524, w_000_3525, w_000_3526, w_000_3527, w_000_3528, w_000_3529, w_000_3530, w_000_3531, w_000_3532, w_000_3533, w_000_3534, w_000_3535, w_000_3536, w_000_3537, w_000_3538, w_000_3539, w_000_3540, w_000_3541, w_000_3542, w_000_3543, w_000_3544, w_000_3545, w_000_3546, w_000_3547, w_000_3548, w_000_3549, w_000_3550, w_000_3551, w_000_3552, w_000_3553, w_000_3554, w_000_3555, w_000_3556, w_000_3557, w_000_3558, w_000_3559, w_000_3560, w_000_3561, w_000_3562, w_000_3563, w_000_3564, w_000_3565, w_000_3566, w_000_3567, w_000_3568, w_000_3569, w_000_3570, w_000_3571, w_000_3572, w_000_3573, w_000_3574, w_000_3575, w_000_3576, w_000_3577, w_000_3578, w_000_3579, w_000_3580, w_000_3581, w_000_3582, w_000_3583, w_000_3584, w_000_3585, w_000_3586, w_000_3587, w_000_3588, w_000_3589, w_000_3590, w_000_3591, w_000_3592, w_000_3593, w_000_3594, w_000_3595, w_000_3596, w_000_3597, w_000_3598, w_000_3599, w_000_3600, w_000_3601, w_000_3602, w_000_3603, w_000_3604, w_000_3605, w_000_3606, w_000_3607, w_000_3608, w_000_3609, w_000_3610, w_000_3611, w_000_3612, w_000_3613, w_000_3614, w_000_3615, w_000_3616, w_000_3617, w_000_3618, w_000_3619, w_000_3620, w_000_3621, w_000_3622, w_000_3623, w_000_3624, w_000_3625, w_000_3626, w_000_3627, w_000_3628, w_000_3629, w_000_3630, w_000_3631, w_000_3632, w_000_3633, w_000_3634, w_000_3635, w_000_3636, w_000_3637, w_000_3638, w_000_3639, w_000_3640, w_000_3641, w_000_3642, w_000_3643, w_000_3644, w_000_3645, w_000_3646, w_000_3647, w_000_3648, w_000_3649, w_000_3650, w_000_3651, w_000_3652, w_000_3653, w_000_3654, w_000_3655, w_000_3656, w_000_3657, w_000_3658, w_000_3659, w_000_3660, w_000_3661, w_000_3662, w_000_3663, w_000_3664, w_000_3665, w_000_3666, w_000_3667, w_000_3668, w_000_3669, w_000_3670, w_000_3671, w_000_3672, w_000_3673, w_000_3674, w_000_3675, w_000_3676, w_000_3677, w_000_3678, w_000_3679, w_000_3680, w_000_3681, w_000_3682, w_000_3683, w_000_3684, w_000_3685, w_000_3686, w_000_3687, w_000_3688, w_000_3689, w_000_3690, w_000_3691, w_000_3692, w_000_3693, w_000_3694, w_000_3695, w_000_3696, w_000_3697, w_000_3698, w_000_3699, w_000_3700, w_000_3701, w_000_3702, w_000_3703, w_000_3704, w_000_3705, w_000_3706, w_000_3707, w_000_3708, w_000_3709, w_000_3710, w_000_3711, w_000_3712, w_000_3713, w_000_3714, w_000_3715, w_000_3716, w_000_3717, w_000_3718, w_000_3719, w_000_3720, w_000_3721, w_000_3722, w_000_3723, w_000_3724, w_000_3725, w_000_3726, w_000_3727, w_000_3728, w_000_3729, w_000_3730, w_000_3731, w_000_3732, w_000_3733, w_000_3734, w_000_3735, w_000_3736, w_000_3737, w_000_3738, w_000_3739, w_000_3740, w_000_3741, w_000_3742, w_000_3743, w_000_3744, w_000_3745, w_000_3746, w_000_3747, w_000_3748, w_000_3749, w_000_3750, w_000_3751, w_000_3752, w_000_3753, w_000_3754, w_000_3755, w_000_3756, w_000_3757, w_000_3758, w_000_3759, w_000_3760, w_000_3761, w_000_3762, w_000_3763, w_000_3764, w_000_3765, w_000_3766, w_000_3767, w_000_3768, w_000_3769, w_000_3770, w_000_3771, w_000_3772, w_000_3773, w_000_3774, w_000_3775, w_000_3776, w_000_3777, w_000_3778, w_000_3779, w_000_3780, w_000_3781, w_000_3782, w_000_3783, w_000_3784, w_000_3785, w_000_3786, w_000_3787, w_000_3788, w_000_3789, w_000_3790, w_000_3791, w_000_3792, w_000_3793, w_000_3794, w_000_3795, w_000_3796, w_000_3797, w_000_3798, w_000_3799, w_000_3800, w_000_3801, w_000_3802, w_000_3803, w_000_3804, w_000_3805, w_000_3806, w_000_3807, w_000_3808, w_000_3809, w_000_3810, w_000_3811, w_000_3812, w_000_3813, w_000_3814, w_000_3815, w_000_3816, w_000_3817, w_000_3818, w_000_3819, w_000_3820, w_000_3821, w_000_3822, w_000_3823, w_000_3824, w_000_3825, w_000_3826, w_000_3827, w_000_3828, w_000_3829, w_000_3830, w_000_3831, w_000_3832, w_000_3833, w_000_3834, w_000_3835, w_000_3836, w_000_3837, w_000_3838, w_000_3839, w_000_3840, w_000_3841, w_000_3842, w_000_3843, w_000_3844, w_000_3845, w_000_3846, w_000_3847, w_000_3848, w_000_3849, w_000_3850, w_000_3851, w_000_3852, w_000_3853, w_000_3854, w_000_3855, w_000_3856, w_000_3857, w_000_3858, w_000_3859, w_000_3860, w_000_3861, w_000_3862, w_000_3863, w_000_3864, w_000_3865, w_000_3866, w_000_3867, w_000_3868, w_000_3869, w_000_3870, w_000_3871, w_000_3872, w_000_3873, w_000_3874, w_000_3875, w_000_3876, w_000_3877, w_000_3878, w_000_3879, w_000_3880, w_000_3881, w_000_3882, w_000_3883, w_000_3884, w_000_3885, w_000_3886, w_000_3887, w_000_3888, w_000_3889, w_000_3890, w_000_3891, w_000_3892, w_000_3893, w_000_3894, w_000_3895, w_000_3896, w_000_3897, w_000_3898, w_000_3899, w_000_3900, w_000_3901, w_000_3902, w_000_3903, w_000_3904, w_000_3905, w_000_3906, w_000_3907, w_000_3908, w_000_3909, w_000_3910, w_000_3911, w_000_3912, w_000_3913, w_000_3914, w_000_3915, w_000_3916, w_000_3917, w_000_3918, w_000_3919, w_000_3920, w_000_3921, w_000_3922, w_000_3923, w_000_3924, w_000_3925, w_000_3926, w_000_3927, w_000_3928, w_000_3929, w_000_3930, w_000_3931, w_000_3932, w_000_3933, w_000_3934, w_000_3935, w_000_3936, w_000_3937, w_000_3938, w_000_3939, w_000_3940, w_000_3941, w_000_3942, w_000_3943, w_000_3944, w_000_3945, w_000_3946, w_000_3947, w_000_3948, w_000_3949, w_000_3950, w_000_3951, w_000_3952, w_000_3953, w_000_3954, w_000_3955, w_000_3956, w_000_3957, w_000_3958, w_000_3959, w_000_3960, w_000_3961, w_000_3962, w_000_3963, w_000_3964, w_000_3965, w_000_3966, w_000_3967, w_000_3968, w_000_3969, w_000_3970, w_000_3971, w_000_3972, w_000_3973, w_000_3974, w_000_3975, w_000_3976, w_000_3977, w_000_3978, w_000_3979, w_000_3980, w_000_3981, w_000_3982, w_000_3983, w_000_3984, w_000_3985, w_000_3986, w_000_3987, w_000_3988, w_000_3989, w_000_3990, w_000_3991, w_000_3992, w_000_3993, w_000_3994, w_000_3995, w_000_3996, w_000_3997, w_000_3998, w_000_3999, w_000_4000, w_000_4001, w_000_4002, w_000_4003, w_000_4004, w_000_4005, w_000_4006, w_000_4007, w_000_4008, w_000_4009, w_000_4010, w_000_4011, w_000_4012, w_000_4013, w_000_4014, w_000_4015, w_000_4016, w_000_4017, w_000_4018, w_000_4019, w_000_4020, w_000_4021, w_000_4022, w_000_4023, w_000_4024, w_000_4025, w_000_4026, w_000_4027, w_000_4028, w_000_4029, w_000_4030, w_000_4031, w_000_4032, w_000_4033, w_000_4034, w_000_4035, w_000_4036, w_000_4037, w_000_4038, w_000_4039, w_000_4040, w_000_4041, w_000_4042, w_000_4043, w_000_4044, w_000_4045, w_000_4046, w_000_4047, w_000_4048, w_000_4049, w_000_4050, w_000_4051, w_000_4052, w_000_4053, w_000_4054, w_000_4055, w_000_4056, w_000_4057, w_000_4058, w_000_4059, w_000_4060, w_000_4061, w_000_4062, w_000_4063, w_000_4064, w_000_4065, w_000_4066, w_000_4067, w_000_4068, w_000_4069, w_000_4070, w_000_4071, w_000_4072, w_000_4073, w_000_4074, w_000_4075, w_000_4076, w_000_4077, w_000_4078, w_000_4079, w_000_4080, w_000_4081, w_000_4082, w_000_4083, w_000_4084, w_000_4085, w_000_4086, w_000_4087, w_000_4088, w_000_4089, w_000_4090, w_000_4091, w_000_4092, w_000_4093, w_000_4094, w_000_4095, w_000_4096, w_000_4097, w_000_4098, w_000_4099, w_000_4100, w_000_4101, w_000_4102, w_000_4103, w_000_4104, w_000_4105, w_000_4106, w_000_4107, w_000_4108, w_000_4109, w_000_4110, w_000_4111, w_000_4112, w_000_4113, w_000_4114, w_000_4115, w_000_4116, w_000_4117, w_000_4118, w_000_4119, w_000_4120, w_000_4121, w_000_4122, w_000_4123, w_000_4124, w_000_4125, w_000_4126, w_000_4127, w_000_4128, w_000_4129, w_000_4130, w_000_4131, w_000_4132, w_000_4133, w_000_4134, w_000_4135, w_000_4136, w_000_4137, w_000_4138, w_000_4139, w_000_4140, w_000_4141, w_000_4142, w_000_4143, w_000_4144, w_000_4145, w_000_4146, w_000_4147, w_000_4148, w_000_4149, w_000_4150, w_000_4151, w_000_4152, w_000_4153, w_000_4154, w_000_4155, w_000_4156, w_000_4157, w_000_4158, w_000_4159, w_000_4160, w_000_4161, w_000_4162, w_000_4163, w_000_4164, w_000_4165, w_000_4166, w_000_4167, w_000_4168, w_000_4169, w_000_4170, w_000_4171, w_000_4172, w_000_4173, w_000_4174, w_000_4175, w_000_4176, w_000_4177, w_000_4178, w_000_4179, w_000_4180, w_000_4181, w_000_4182, w_000_4183, w_000_4184, w_000_4185, w_000_4186, w_000_4187, w_000_4188, w_000_4189, w_000_4190, w_000_4191, w_000_4192, w_000_4193, w_000_4194, w_000_4195, w_000_4196, w_000_4197, w_000_4198, w_000_4199, w_000_4200, w_000_4201, w_000_4202, w_000_4203, w_000_4204, w_000_4205, w_000_4206, w_000_4207, w_000_4208, w_000_4209, w_000_4210, w_000_4211, w_000_4212, w_000_4213, w_000_4215, w_000_4216, w_000_4217, w_000_4218, w_000_4219, w_000_4220, w_000_4221, w_000_4222, w_000_4223, w_000_4224, w_000_4225, w_000_4226, w_000_4227, w_000_4228, w_000_4229, w_000_4230, w_000_4231, w_000_4232, w_000_4233, w_000_4234, w_000_4235, w_000_4236, w_000_4237, w_000_4238, w_000_4239, w_000_4240, w_000_4241, w_000_4242, w_000_4243, w_000_4244, w_000_4245, w_000_4246, w_000_4247, w_000_4248, w_000_4249, w_000_4250, w_000_4251, w_000_4252, w_000_4253, w_000_4254, w_000_4255, w_000_4256, w_000_4257, w_000_4258, w_000_4259, w_000_4260, w_000_4261, w_000_4262, w_000_4263, w_000_4264, w_000_4265, w_000_4266, w_000_4267, w_000_4268, w_000_4269, w_000_4270, w_000_4271, w_000_4272, w_000_4273, w_000_4274, w_000_4275, w_000_4276, w_000_4277, w_000_4278, w_000_4279, w_000_4280, w_000_4281, w_000_4282, w_000_4283, w_000_4284, w_000_4285, w_000_4286, w_000_4287, w_000_4288, w_000_4289, w_000_4290, w_000_4291, w_000_4292, w_000_4293, w_000_4294, w_000_4295, w_000_4296, w_000_4297, w_000_4298, w_000_4299, w_000_4300, w_000_4301, w_000_4302, w_000_4303, w_000_4304, w_000_4305, w_000_4306, w_000_4307, w_000_4308, w_000_4309, w_000_4310, w_000_4311, w_000_4312, w_000_4313, w_000_4314, w_000_4315, w_000_4316, w_000_4317, w_000_4318, w_000_4319, w_000_4320, w_000_4321, w_000_4322, w_000_4323, w_000_4324, w_000_4325, w_000_4326, w_000_4327, w_000_4328, w_000_4329, w_000_4330, w_000_4331, w_000_4332, w_000_4333, w_000_4334, w_000_4335, w_000_4336, w_000_4337, w_000_4338, w_000_4339, w_000_4340, w_000_4341, w_000_4342, w_000_4343, w_000_4344, w_000_4345, w_000_4346, w_000_4347, w_000_4349, w_000_4350, w_000_4351, w_000_4352, w_000_4353, w_000_4354, w_000_4355, w_000_4356, w_000_4357, w_000_4358, w_000_4359, w_000_4360, w_000_4361, w_000_4362, w_000_4363, w_000_4364, w_000_4365, w_000_4366, w_000_4367, w_000_4368, w_000_4369, w_000_4370, w_000_4371, w_000_4372, w_000_4373, w_000_4374, w_000_4375, w_000_4376, w_000_4377, w_000_4378, w_000_4379, w_000_4380, w_000_4381, w_000_4382, w_000_4383, w_000_4384, w_000_4385, w_000_4386, w_000_4387, w_000_4388, w_000_4389, w_000_4390, w_000_4391, w_000_4392, w_000_4393, w_000_4394, w_000_4395, w_000_4396, w_000_4397, w_000_4398, w_000_4399, w_000_4400, w_000_4401, w_000_4402, w_000_4403, w_000_4404, w_000_4405, w_000_4406, w_000_4407, w_000_4408, w_000_4409, w_000_4410, w_000_4411, w_000_4412, w_000_4413, w_000_4414, w_000_4415, w_000_4416, w_000_4417, w_000_4418, w_000_4419, w_000_4420, w_000_4421, w_000_4422, w_000_4423, w_000_4424, w_000_4425, w_000_4426, w_000_4427, w_000_4428, w_000_4429, w_000_4430, w_000_4431, w_000_4432, w_000_4433, w_000_4434, w_000_4435, w_000_4436, w_000_4437, w_000_4438, w_000_4439, w_000_4440, w_000_4441, w_000_4442, w_000_4443, w_000_4444, w_000_4445, w_000_4446, w_000_4447, w_000_4448, w_000_4449, w_000_4450, w_000_4451, w_000_4452, w_000_4453, w_000_4454, w_000_4455, w_000_4456, w_000_4457, w_000_4458, w_000_4459, w_000_4460, w_000_4461, w_000_4462, w_000_4463, w_000_4464, w_000_4465, w_000_4466, w_000_4467, w_000_4468, w_000_4469, w_000_4470, w_000_4471, w_000_4472, w_000_4473, w_000_4474, w_000_4475, w_000_4476, w_000_4477, w_000_4478, w_000_4479, w_000_4480, w_000_4481, w_000_4482, w_000_4483, w_000_4484, w_000_4485, w_000_4486, w_000_4487, w_000_4488, w_000_4489, w_000_4490, w_000_4491, w_000_4492, w_000_4493, w_000_4494, w_000_4495, w_000_4496, w_000_4497, w_000_4498, w_000_4499, w_000_4500, w_000_4501, w_000_4502, w_000_4503, w_000_4504, w_000_4505, w_000_4506, w_000_4507, w_000_4508, w_000_4509, w_000_4510, w_000_4511, w_000_4512, w_000_4513, w_000_4514, w_000_4515, w_000_4516, w_000_4517, w_000_4518, w_000_4519, w_000_4520, w_000_4521, w_000_4522, w_000_4523, w_000_4524, w_000_4525, w_000_4526, w_000_4527, w_000_4528, w_000_4529, w_000_4530, w_000_4531, w_000_4532, w_000_4533, w_000_4534, w_000_4535, w_000_4536, w_000_4537, w_000_4538, w_000_4539, w_000_4540, w_000_4541, w_000_4542, w_000_4543, w_000_4544, w_000_4545, w_000_4546, w_000_4547, w_000_4548, w_000_4549, w_000_4550, w_000_4551, w_000_4552, w_000_4553, w_000_4554, w_000_4555, w_000_4556, w_000_4557, w_000_4559, w_000_4560, w_000_4561, w_000_4562, w_000_4563, w_000_4564, w_000_4565, w_000_4566, w_000_4567, w_000_4568, w_000_4569, w_000_4571, w_000_4572, w_000_4573, w_000_4574, w_000_4575, w_000_4576, w_000_4577, w_000_4578, w_000_4579, w_000_4580, w_000_4581, w_000_4582, w_000_4583, w_000_4584, w_000_4585, w_000_4586, w_000_4587, w_000_4588, w_000_4589, w_000_4590, w_000_4591, w_000_4592, w_000_4593, w_000_4594, w_000_4595, w_000_4596, w_000_4597, w_000_4598, w_000_4599, w_000_4600, w_000_4601, w_000_4602, w_000_4603, w_000_4604, w_000_4605, w_000_4606, w_000_4607, w_000_4608, w_000_4609, w_000_4610, w_000_4611, w_000_4612, w_000_4613, w_000_4614, w_000_4615, w_000_4616, w_000_4617, w_000_4618, w_000_4619, w_000_4620, w_000_4621, w_000_4622, w_000_4623, w_000_4624, w_000_4625, w_000_4626, w_000_4627, w_000_4628, w_000_4629, w_000_4630, w_000_4631, w_000_4632, w_000_4633, w_000_4634, w_000_4635, w_000_4636, w_000_4637, w_000_4638, w_000_4639, w_000_4640, w_000_4641, w_000_4642, w_000_4643, w_000_4644, w_000_4645, w_000_4646, w_000_4647, w_000_4648, w_000_4649, w_000_4650, w_000_4651, w_000_4652, w_000_4653, w_000_4654, w_000_4655, w_000_4656, w_000_4657, w_000_4658, w_000_4659, w_000_4660, w_000_4661, w_000_4662, w_000_4663, w_000_4664, w_000_4665, w_000_4666, w_000_4667, w_000_4668, w_000_4669, w_000_4670, w_000_4671, w_000_4672, w_000_4673, w_000_4674, w_000_4675, w_000_4676, w_000_4677, w_000_4678, w_000_4679, w_000_4680, w_000_4681, w_000_4682, w_000_4683, w_000_4684, w_000_4685, w_000_4686, w_000_4687, w_000_4688, w_000_4689, w_000_4690, w_000_4691, w_000_4692, w_000_4693, w_000_4694, w_000_4695, w_000_4696, w_000_4697, w_000_4698, w_000_4699, w_000_4700, w_000_4701, w_000_4702, w_000_4703, w_000_4704, w_000_4705, w_000_4706, w_000_4707, w_000_4708, w_000_4709, w_000_4710, w_000_4711, w_000_4712, w_000_4713, w_000_4714, w_000_4715, w_000_4716, w_000_4717, w_000_4718, w_000_4719, w_000_4720, w_000_4721, w_000_4722, w_000_4723, w_000_4724, w_000_4725, w_000_4726, w_000_4727, w_000_4728, w_000_4729, w_000_4730, w_000_4731, w_000_4732, w_000_4733, w_000_4734, w_000_4735, w_000_4736, w_000_4737, w_000_4738, w_000_4739, w_000_4740, w_000_4741, w_000_4742, w_000_4743, w_000_4744, w_000_4745, w_000_4746, w_000_4747, w_000_4748, w_000_4749, w_000_4750, w_000_4751, w_000_4752, w_000_4753, w_000_4754, w_000_4755, w_000_4756, w_000_4757, w_000_4758, w_000_4759, w_000_4760, w_000_4761, w_000_4762, w_000_4763, w_000_4764, w_000_4765, w_000_4766, w_000_4767, w_000_4768, w_000_4769, w_000_4770, w_000_4771, w_000_4772, w_000_4773, w_000_4774, w_000_4775, w_000_4776, w_000_4777, w_000_4778, w_000_4779, w_000_4780, w_000_4781, w_000_4782, w_000_4783, w_000_4784, w_000_4785, w_000_4786, w_000_4787, w_000_4788, w_000_4789, w_000_4790, w_000_4791, w_000_4792, w_000_4793, w_000_4794, w_000_4795, w_000_4796, w_000_4797, w_000_4798, w_000_4799, w_000_4800, w_000_4801, w_000_4803, w_000_4804, w_000_4805, w_000_4806, w_000_4807, w_000_4808, w_000_4809, w_000_4810, w_000_4811, w_000_4812, w_000_4813, w_000_4814, w_000_4815, w_000_4816, w_000_4817, w_000_4818, w_000_4819, w_000_4820, w_000_4821, w_000_4822, w_000_4823, w_000_4824, w_000_4825, w_000_4826, w_000_4827, w_000_4828, w_000_4829, w_000_4830, w_000_4831, w_000_4832, w_000_4833, w_000_4834, w_000_4835, w_000_4836, w_000_4837, w_000_4838, w_000_4839, w_000_4840, w_000_4841, w_000_4842, w_000_4843, w_000_4844, w_000_4845, w_000_4846, w_000_4847, w_000_4848, w_000_4849, w_000_4850, w_000_4851, w_000_4852, w_000_4853, w_000_4854, w_000_4855, w_000_4856, w_000_4860, w_000_4861, w_000_4862, w_000_4863, w_000_4864, w_000_4865, w_000_4866, w_000_4867, w_000_4868, w_000_4869, w_000_4870, w_000_4871, w_000_4872, w_000_4873, w_000_4874, w_000_4875, w_000_4876, w_000_4877, w_000_4878, w_000_4879, w_000_4880, w_000_4881, w_000_4882, w_000_4883, w_000_4884, w_000_4885, w_000_4886, w_000_4887, w_000_4889, w_000_4890, w_000_4891, w_000_4892, w_000_4893, w_000_4894, w_000_4895, w_000_4896, w_000_4897, w_000_4898, w_000_4900, w_000_4901, w_000_4902, w_000_4903, w_000_4905, w_000_4906, w_000_4907, w_000_4908, w_000_4909, w_000_4910, w_000_4911, w_000_4912, w_000_4914, w_000_4915, w_000_4916, w_000_4917, w_000_4918, w_000_4920, w_000_4921, w_000_4922, w_000_4923, w_000_4924, w_000_4926, w_000_4927, w_000_4928, w_000_4929, w_000_4930, w_000_4931, w_000_4932, w_000_4933, w_000_4934, w_000_4935, w_000_4936, w_000_4937, w_000_4938, w_000_4939, w_000_4941, w_000_4942, w_000_4944, w_000_4945, w_000_4946, w_000_4947, w_000_4949, w_000_4950, w_000_4952, w_000_4953, w_000_4955, w_000_4956, w_000_4957, w_000_4958, w_000_4959, w_000_4963, w_000_4964, w_000_4966, w_000_4968, w_000_4969, w_000_4970, w_000_4974, w_000_4979, w_000_4980, w_000_4984, w_000_4990, w_000_4991, w_000_4994, w_5000_000, w_5000_001, w_5000_002, w_5000_003, w_5000_004, w_5000_005, w_5000_006, w_5000_007, w_5000_008, w_5000_009, w_5000_010, w_5000_011, w_5000_012, w_5000_013, w_5000_014, w_5000_015, w_5000_016, w_5000_017, w_5000_018, w_5000_019, w_5000_020, w_5000_021, w_5000_022, w_5000_023, w_5000_024, w_5000_025, w_5000_026, w_5000_027, w_5000_028, w_5000_029, w_5000_030, w_5000_031, w_5000_032, w_5000_033, w_5000_034, w_5000_035, w_5000_036, w_5000_037, w_5000_038, w_5000_039, w_5000_040, w_5000_041, w_5000_042, w_5000_043, w_5000_044, w_5000_045, w_5000_046, w_5000_047, w_5000_048, w_5000_049, w_5000_050, w_5000_051, w_5000_052, w_5000_053, w_5000_054, w_5000_055, w_5000_056, w_5000_057, w_5000_058, w_5000_059, w_5000_060, w_5000_061, w_5000_062, w_5000_063, w_5000_064, w_5000_065, w_5000_066, w_5000_067, w_5000_068, w_5000_069, w_5000_070, w_5000_071, w_5000_072, w_5000_073, w_5000_074, w_5000_075, w_5000_076, w_5000_077, w_5000_078, w_5000_079, w_5000_080, w_5000_081, w_5000_082, w_5000_083, w_5000_084, w_5000_085, w_5000_086, w_5000_087, w_5000_088, w_5000_089, w_5000_090, w_5000_091, w_5000_092, w_5000_093, w_5000_094, w_5000_095, w_5000_096, w_5000_097, w_5000_098, w_5000_099, w_5000_100, w_5000_101, w_5000_102, w_5000_103, w_5000_104, w_5000_105, w_5000_106, w_5000_107, w_5000_108, w_5000_109, w_5000_110, w_5000_111, w_5000_112, w_5000_113, w_5000_114, w_5000_115, w_5000_116, w_5000_117, w_5000_118, w_5000_119, w_5000_120, w_5000_121, w_5000_122, w_5000_123, w_5000_124, w_5000_125, w_5000_126, w_5000_127, w_5000_128, w_5000_129, w_5000_130, w_5000_131, w_5000_132, w_5000_133, w_5000_134, w_5000_135, w_5000_136, w_5000_137, w_5000_138, w_5000_139, w_5000_140, w_5000_141, w_5000_142, w_5000_143, w_5000_144, w_5000_145, w_5000_146, w_5000_147, w_5000_148, w_5000_149, w_5000_150, w_5000_151, w_5000_152, w_5000_153, w_5000_154, w_5000_155, w_5000_156, w_5000_157, w_5000_158, w_5000_159, w_5000_160, w_5000_161, w_5000_162, w_5000_163, w_5000_164, w_5000_165, w_5000_166, w_5000_167, w_5000_168, w_5000_169, w_5000_170, w_5000_171, w_5000_172, w_5000_173, w_5000_174, w_5000_175, w_5000_176, w_5000_177, w_5000_178, w_5000_179, w_5000_180, w_5000_181, w_5000_182, w_5000_183, w_5000_184, w_5000_185, w_5000_186, w_5000_187, w_5000_188, w_5000_189, w_5000_190, w_5000_191, w_5000_192, w_5000_193, w_5000_194, w_5000_195, w_5000_196, w_5000_197, w_5000_198, w_5000_199, w_5000_200, w_5000_201, w_5000_202, w_5000_203, w_5000_204, w_5000_205, w_5000_206, w_5000_207, w_5000_208, w_5000_209, w_5000_210, w_5000_211, w_5000_212, w_5000_213, w_5000_214, w_5000_215, w_5000_216, w_5000_217, w_5000_218, w_5000_219, w_5000_220, w_5000_221, w_5000_222, w_5000_223, w_5000_224, w_5000_225, w_5000_226, w_5000_227, w_5000_228, w_5000_229, w_5000_230, w_5000_231, w_5000_232, w_5000_233, w_5000_234, w_5000_235, w_5000_236, w_5000_237, w_5000_238, w_5000_239, w_5000_240, w_5000_241, w_5000_242, w_5000_243, w_5000_244, w_5000_245, w_5000_246, w_5000_247, w_5000_248, w_5000_249, w_5000_250, w_5000_251, w_5000_252, w_5000_253, w_5000_254, w_5000_255, w_5000_256, w_5000_257, w_5000_258, w_5000_259, w_5000_260, w_5000_261, w_5000_262, w_5000_263, w_5000_264, w_5000_265, w_5000_266, w_5000_267, w_5000_268, w_5000_269, w_5000_270, w_5000_271, w_5000_272, w_5000_273, w_5000_274, w_5000_275, w_5000_276, w_5000_277, w_5000_278, w_5000_279, w_5000_280, w_5000_281, w_5000_282, w_5000_283, w_5000_284, w_5000_285, w_5000_286, w_5000_287, w_5000_288, w_5000_289, w_5000_290, w_5000_291, w_5000_292, w_5000_293, w_5000_294, w_5000_295, w_5000_296, w_5000_297, w_5000_298, w_5000_299, w_5000_300, w_5000_301, w_5000_302, w_5000_303, w_5000_304, w_5000_305, w_5000_306, w_5000_307, w_5000_308, w_5000_309, w_5000_310, w_5000_311, w_5000_312, w_5000_313, w_5000_314, w_5000_315, w_5000_316, w_5000_317, w_5000_318, w_5000_319, w_5000_320, w_5000_321, w_5000_322, w_5000_323, w_5000_324, w_5000_325, w_5000_326, w_5000_327, w_5000_328, w_5000_329, w_5000_330, w_5000_331, w_5000_332, w_5000_333, w_5000_334, w_5000_335, w_5000_336, w_5000_337, w_5000_338, w_5000_339, w_5000_340, w_5000_341, w_5000_342, w_5000_343, w_5000_344, w_5000_345, w_5000_346, w_5000_347, w_5000_348, w_5000_349, w_5000_350, w_5000_351, w_5000_352, w_5000_353, w_5000_354, w_5000_355, w_5000_356, w_5000_357, w_5000_358, w_5000_359, w_5000_360, w_5000_361, w_5000_362, w_5000_363, w_5000_364, w_5000_365, w_5000_366, w_5000_367, w_5000_368, w_5000_369, w_5000_370, w_5000_371, w_5000_372, w_5000_373, w_5000_374, w_5000_375, w_5000_376, w_5000_377, w_5000_378, w_5000_379, w_5000_380, w_5000_381, w_5000_382, w_5000_383, w_5000_384, w_5000_385, w_5000_386, w_5000_387, w_5000_388, w_5000_389, w_5000_390, w_5000_391, w_5000_392, w_5000_393, w_5000_394, w_5000_395, w_5000_396, w_5000_397, w_5000_398, w_5000_399, w_5000_400, w_5000_401, w_5000_402, w_5000_403, w_5000_404, w_5000_405, w_5000_406, w_5000_407, w_5000_408, w_5000_409, w_5000_410, w_5000_411, w_5000_412, w_5000_413, w_5000_414, w_5000_415, w_5000_416, w_5000_417, w_5000_418, w_5000_419, w_5000_420, w_5000_421, w_5000_422, w_5000_423, w_5000_424, w_5000_425, w_5000_426, w_5000_427, w_5000_428, w_5000_429, w_5000_430, w_5000_431, w_5000_432, w_5000_433, w_5000_434, w_5000_435, w_5000_436, w_5000_437, w_5000_438, w_5000_439, w_5000_440, w_5000_441, w_5000_442, w_5000_443, w_5000_444, w_5000_445, w_5000_446, w_5000_447, w_5000_448, w_5000_449, w_5000_450, w_5000_451, w_5000_452, w_5000_453, w_5000_454, w_5000_455, w_5000_456, w_5000_457, w_5000_458, w_5000_459, w_5000_460, w_5000_461, w_5000_462, w_5000_463, w_5000_464, w_5000_465, w_5000_466, w_5000_467, w_5000_468, w_5000_469, w_5000_470, w_5000_471, w_5000_472, w_5000_473, w_5000_474, w_5000_475, w_5000_476, w_5000_477, w_5000_478, w_5000_479, w_5000_480, w_5000_481, w_5000_482, w_5000_483, w_5000_484, w_5000_485, w_5000_486, w_5000_487, w_5000_488, w_5000_489, w_5000_490, w_5000_491, w_5000_492, w_5000_493, w_5000_494, w_5000_495, w_5000_496, w_5000_497, w_5000_498, w_5000_499, w_5000_500, w_5000_501, w_5000_502, w_5000_503, w_5000_504, w_5000_505, w_5000_506, w_5000_507, w_5000_508, w_5000_509, w_5000_510, w_5000_511, w_5000_512, w_5000_513, w_5000_514, w_5000_515, w_5000_516, w_5000_517, w_5000_518, w_5000_519, w_5000_520, w_5000_521, w_5000_522, w_5000_523, w_5000_524, w_5000_525, w_5000_526, w_5000_527, w_5000_528, w_5000_529, w_5000_530, w_5000_531, w_5000_532, w_5000_533, w_5000_534, w_5000_535, w_5000_536, w_5000_537, w_5000_538, w_5000_539, w_5000_540, w_5000_541, w_5000_542, w_5000_543, w_5000_544, w_5000_545, w_5000_546, w_5000_547, w_5000_548, w_5000_549, w_5000_550, w_5000_551, w_5000_552, w_5000_553, w_5000_554, w_5000_555, w_5000_556, w_5000_557, w_5000_558, w_5000_559, w_5000_560, w_5000_561, w_5000_562, w_5000_563, w_5000_564, w_5000_565, w_5000_566, w_5000_567, w_5000_568, w_5000_569, w_5000_570, w_5000_571, w_5000_572, w_5000_573, w_5000_574, w_5000_575, w_5000_576, w_5000_577, w_5000_578, w_5000_579, w_5000_580, w_5000_581, w_5000_582, w_5000_583, w_5000_584, w_5000_585, w_5000_586, w_5000_587, w_5000_588, w_5000_589, w_5000_590, w_5000_591, w_5000_592, w_5000_593, w_5000_594, w_5000_595, w_5000_596, w_5000_597, w_5000_598, w_5000_599, w_5000_600, w_5000_601, w_5000_602, w_5000_603, w_5000_604, w_5000_605, w_5000_606, w_5000_607, w_5000_608, w_5000_609, w_5000_610, w_5000_611, w_5000_612, w_5000_613, w_5000_614, w_5000_615, w_5000_616, w_5000_617, w_5000_618, w_5000_619, w_5000_620, w_5000_621, w_5000_622, w_5000_623, w_5000_624, w_5000_625, w_5000_626, w_5000_627, w_5000_628, w_5000_629, w_5000_630, w_5000_631, w_5000_632, w_5000_633, w_5000_634, w_5000_635, w_5000_636, w_5000_637, w_5000_638, w_5000_639, w_5000_640, w_5000_641, w_5000_642, w_5000_643, w_5000_644, w_5000_645, w_5000_646, w_5000_647, w_5000_648, w_5000_649, w_5000_650, w_5000_651, w_5000_652, w_5000_653, w_5000_654, w_5000_655, w_5000_656, w_5000_657, w_5000_658, w_5000_659, w_5000_660, w_5000_661, w_5000_662, w_5000_663, w_5000_664, w_5000_665, w_5000_666, w_5000_667, w_5000_668, w_5000_669, w_5000_670, w_5000_671, w_5000_672, w_5000_673, w_5000_674, w_5000_675, w_5000_676, w_5000_677, w_5000_678, w_5000_679, w_5000_680, w_5000_681, w_5000_682, w_5000_683, w_5000_684, w_5000_685, w_5000_686, w_5000_687, w_5000_688, w_5000_689, w_5000_690, w_5000_691, w_5000_692, w_5000_693, w_5000_694, w_5000_695, w_5000_696, w_5000_697, w_5000_698, w_5000_699, w_5000_700, w_5000_701, w_5000_702, w_5000_703, w_5000_704, w_5000_705, w_5000_706, w_5000_707, w_5000_708, w_5000_709, w_5000_710, w_5000_711, w_5000_712, w_5000_713, w_5000_714, w_5000_715, w_5000_716, w_5000_717, w_5000_718, w_5000_719, w_5000_720, w_5000_721, w_5000_722, w_5000_723, w_5000_724, w_5000_725, w_5000_726, w_5000_727, w_5000_728, w_5000_729, w_5000_730, w_5000_731, w_5000_732, w_5000_733, w_5000_734, w_5000_735, w_5000_736, w_5000_737, w_5000_738, w_5000_739, w_5000_740, w_5000_741, w_5000_742, w_5000_743, w_5000_744, w_5000_745, w_5000_746, w_5000_747, w_5000_748, w_5000_749, w_5000_750, w_5000_751, w_5000_752, w_5000_753, w_5000_754, w_5000_755, w_5000_756, w_5000_757, w_5000_758, w_5000_759, w_5000_760, w_5000_761, w_5000_762, w_5000_763, w_5000_764, w_5000_765, w_5000_766, w_5000_767, w_5000_768, w_5000_769, w_5000_770, w_5000_771, w_5000_772, w_5000_773, w_5000_774, w_5000_775, w_5000_776, w_5000_777, w_5000_778, w_5000_779, w_5000_780, w_5000_781, w_5000_782, w_5000_783, w_5000_784, w_5000_785, w_5000_786, w_5000_787, w_5000_788, w_5000_789, w_5000_790, w_5000_791, w_5000_792, w_5000_793, w_5000_794, w_5000_795, w_5000_796, w_5000_797, w_5000_798, w_5000_799, w_5000_800, w_5000_801, w_5000_802, w_5000_803, w_5000_804, w_5000_805, w_5000_806, w_5000_807, w_5000_808, w_5000_809, w_5000_810, w_5000_811, w_5000_812, w_5000_813, w_5000_814, w_5000_815, w_5000_816, w_5000_817, w_5000_818, w_5000_819, w_5000_820, w_5000_821, w_5000_822, w_5000_823, w_5000_824, w_5000_825, w_5000_826, w_5000_827, w_5000_828, w_5000_829, w_5000_830, w_5000_831, w_5000_832, w_5000_833, w_5000_834, w_5000_835, w_5000_836, w_5000_837, w_5000_838, w_5000_839, w_5000_840, w_5000_841, w_5000_842, w_5000_843, w_5000_844, w_5000_845, w_5000_846, w_5000_847, w_5000_848, w_5000_849, w_5000_850, w_5000_851, w_5000_852, w_5000_853, w_5000_854, w_5000_855, w_5000_856, w_5000_857, w_5000_858, w_5000_859, w_5000_860, w_5000_861, w_5000_862, w_5000_863, w_5000_864, w_5000_865, w_5000_866, w_5000_867, w_5000_868, w_5000_869, w_5000_870, w_5000_871, w_5000_872, w_5000_873, w_5000_874, w_5000_875, w_5000_876, w_5000_877, w_5000_878, w_5000_879, w_5000_880, w_5000_881, w_5000_882, w_5000_883, w_5000_884, w_5000_885, w_5000_886, w_5000_887, w_5000_888, w_5000_889, w_5000_890, w_5000_891, w_5000_892, w_5000_893, w_5000_894, w_5000_895, w_5000_896, w_5000_897, w_5000_898, w_5000_899, w_5000_900, w_5000_901, w_5000_902, w_5000_903, w_5000_904, w_5000_905, w_5000_906, w_5000_907, w_5000_908, w_5000_909, w_5000_910, w_5000_911, w_5000_912, w_5000_913, w_5000_914, w_5000_915, w_5000_916, w_5000_917, w_5000_918, w_5000_919, w_5000_920, w_5000_921, w_5000_922, w_5000_923, w_5000_924, w_5000_925, w_5000_926, w_5000_927, w_5000_928, w_5000_929, w_5000_930, w_5000_931, w_5000_932, w_5000_933, w_5000_934, w_5000_935, w_5000_936, w_5000_937, w_5000_938, w_5000_939, w_5000_940, w_5000_941, w_5000_942, w_5000_943, w_5000_944, w_5000_945, w_5000_946, w_5000_947, w_5000_948, w_5000_949, w_5000_950, w_5000_951, w_5000_952, w_5000_953, w_5000_954, w_5000_955, w_5000_956, w_5000_957, w_5000_958, w_5000_959, w_5000_960, w_5000_961, w_5000_962, w_5000_963, w_5000_964, w_5000_965, w_5000_966, w_5000_967, w_5000_968, w_5000_969, w_5000_970, w_5000_971, w_5000_972, w_5000_973, w_5000_974, w_5000_975, w_5000_976, w_5000_977, w_5000_978, w_5000_979, w_5000_980, w_5000_981, w_5000_982, w_5000_983, w_5000_984, w_5000_985, w_5000_986, w_5000_987, w_5000_988, w_5000_989, w_5000_990, w_5000_991, w_5000_992, w_5000_993, w_5000_994, w_5000_995, w_5000_996, w_5000_997, w_5000_998, w_5000_999, w_5000_1000, w_5000_1001, w_5000_1002, w_5000_1003, w_5000_1004, w_5000_1005, w_5000_1006, w_5000_1007, w_5000_1008, w_5000_1009, w_5000_1010, w_5000_1011, w_5000_1012, w_5000_1013, w_5000_1014, w_5000_1015, w_5000_1016, w_5000_1017, w_5000_1018, w_5000_1019, w_5000_1020, w_5000_1021, w_5000_1022, w_5000_1023, w_5000_1024, w_5000_1025, w_5000_1026, w_5000_1027, w_5000_1028, w_5000_1029, w_5000_1030, w_5000_1031, w_5000_1032, w_5000_1033, w_5000_1034, w_5000_1035, w_5000_1036, w_5000_1037, w_5000_1038, w_5000_1039, w_5000_1040, w_5000_1041, w_5000_1042, w_5000_1043, w_5000_1044, w_5000_1045, w_5000_1046, w_5000_1047, w_5000_1048, w_5000_1049, w_5000_1050, w_5000_1051, w_5000_1052, w_5000_1053, w_5000_1054, w_5000_1055, w_5000_1056, w_5000_1057, w_5000_1058, w_5000_1059, w_5000_1060, w_5000_1061, w_5000_1062, w_5000_1063, w_5000_1064, w_5000_1065, w_5000_1066, w_5000_1067, w_5000_1068, w_5000_1069, w_5000_1070, w_5000_1071, w_5000_1072, w_5000_1073, w_5000_1074, w_5000_1075, w_5000_1076, w_5000_1077, w_5000_1078, w_5000_1079, w_5000_1080, w_5000_1081, w_5000_1082, w_5000_1083, w_5000_1084, w_5000_1085, w_5000_1086, w_5000_1087, w_5000_1088, w_5000_1089, w_5000_1090, w_5000_1091, w_5000_1092, w_5000_1093, w_5000_1094, w_5000_1095, w_5000_1096, w_5000_1097, w_5000_1098, w_5000_1099, w_5000_1100, w_5000_1101, w_5000_1102, w_5000_1103, w_5000_1104, w_5000_1105, w_5000_1106, w_5000_1107, w_5000_1108, w_5000_1109, w_5000_1110, w_5000_1111, w_5000_1112, w_5000_1113, w_5000_1114, w_5000_1115, w_5000_1116, w_5000_1117, w_5000_1118, w_5000_1119, w_5000_1120, w_5000_1121, w_5000_1122, w_5000_1123, w_5000_1124, w_5000_1125, w_5000_1126, w_5000_1127, w_5000_1128, w_5000_1129, w_5000_1130, w_5000_1131, w_5000_1132, w_5000_1133, w_5000_1134, w_5000_1135, w_5000_1136, w_5000_1137, w_5000_1138, w_5000_1139, w_5000_1140, w_5000_1141, w_5000_1142, w_5000_1143, w_5000_1144, w_5000_1145, w_5000_1146, w_5000_1147, w_5000_1148, w_5000_1149, w_5000_1150, w_5000_1151, w_5000_1152, w_5000_1153, w_5000_1154, w_5000_1155, w_5000_1156, w_5000_1157, w_5000_1158, w_5000_1159, w_5000_1160, w_5000_1161, w_5000_1162, w_5000_1163, w_5000_1164, w_5000_1165, w_5000_1166, w_5000_1167, w_5000_1168, w_5000_1169, w_5000_1170, w_5000_1171, w_5000_1172, w_5000_1173, w_5000_1174, w_5000_1175, w_5000_1176, w_5000_1177, w_5000_1178, w_5000_1179, w_5000_1180, w_5000_1181, w_5000_1182, w_5000_1183, w_5000_1184, w_5000_1185, w_5000_1186, w_5000_1187, w_5000_1188, w_5000_1189, w_5000_1190, w_5000_1191, w_5000_1192, w_5000_1193, w_5000_1194, w_5000_1195, w_5000_1196, w_5000_1197, w_5000_1198, w_5000_1199, w_5000_1200, w_5000_1201, w_5000_1202, w_5000_1203, w_5000_1204, w_5000_1205, w_5000_1206, w_5000_1207, w_5000_1208, w_5000_1209, w_5000_1210, w_5000_1211, w_5000_1212, w_5000_1213, w_5000_1214, w_5000_1215, w_5000_1216, w_5000_1217, w_5000_1218, w_5000_1219, w_5000_1220, w_5000_1221, w_5000_1222, w_5000_1223, w_5000_1224, w_5000_1225, w_5000_1226, w_5000_1227, w_5000_1228, w_5000_1229, w_5000_1230, w_5000_1231, w_5000_1232, w_5000_1233, w_5000_1234, w_5000_1235, w_5000_1236, w_5000_1237, w_5000_1238, w_5000_1239, w_5000_1240, w_5000_1241, w_5000_1242, w_5000_1243, w_5000_1244, w_5000_1245, w_5000_1246, w_5000_1247, w_5000_1248, w_5000_1249, w_5000_1250, w_5000_1251, w_5000_1252, w_5000_1253, w_5000_1254, w_5000_1255, w_5000_1256, w_5000_1257, w_5000_1258, w_5000_1259, w_5000_1260, w_5000_1261, w_5000_1262, w_5000_1263, w_5000_1264, w_5000_1265, w_5000_1266, w_5000_1267, w_5000_1268, w_5000_1269, w_5000_1270, w_5000_1271, w_5000_1272, w_5000_1273, w_5000_1274, w_5000_1275, w_5000_1276, w_5000_1277, w_5000_1278, w_5000_1279, w_5000_1280, w_5000_1281, w_5000_1282, w_5000_1283, w_5000_1284, w_5000_1285, w_5000_1286, w_5000_1287, w_5000_1288, w_5000_1289, w_5000_1290, w_5000_1291, w_5000_1292, w_5000_1293, w_5000_1294, w_5000_1295, w_5000_1296, w_5000_1297, w_5000_1298, w_5000_1299, w_5000_1300, w_5000_1301, w_5000_1302, w_5000_1303, w_5000_1304, w_5000_1305, w_5000_1306, w_5000_1307, w_5000_1308, w_5000_1309, w_5000_1310, w_5000_1311, w_5000_1312, w_5000_1313, w_5000_1314, w_5000_1315, w_5000_1316, w_5000_1317, w_5000_1318, w_5000_1319, w_5000_1320, w_5000_1321, w_5000_1322, w_5000_1323, w_5000_1324, w_5000_1325, w_5000_1326, w_5000_1327, w_5000_1328, w_5000_1329, w_5000_1330, w_5000_1331, w_5000_1332, w_5000_1333, w_5000_1334, w_5000_1335, w_5000_1336, w_5000_1337, w_5000_1338, w_5000_1339, w_5000_1340, w_5000_1341, w_5000_1342, w_5000_1343, w_5000_1344, w_5000_1345, w_5000_1346, w_5000_1347, w_5000_1348, w_5000_1349, w_5000_1350, w_5000_1351, w_5000_1352, w_5000_1353, w_5000_1354, w_5000_1355, w_5000_1356, w_5000_1357, w_5000_1358, w_5000_1359, w_5000_1360, w_5000_1361, w_5000_1362, w_5000_1363, w_5000_1364, w_5000_1365, w_5000_1366, w_5000_1367, w_5000_1368, w_5000_1369, w_5000_1370, w_5000_1371, w_5000_1372, w_5000_1373, w_5000_1374, w_5000_1375, w_5000_1376, w_5000_1377, w_5000_1378, w_5000_1379, w_5000_1380, w_5000_1381, w_5000_1382, w_5000_1383, w_5000_1384, w_5000_1385, w_5000_1386, w_5000_1387, w_5000_1388, w_5000_1389, w_5000_1390, w_5000_1391, w_5000_1392, w_5000_1393, w_5000_1394, w_5000_1395, w_5000_1396, w_5000_1397, w_5000_1398, w_5000_1399, w_5000_1400, w_5000_1401, w_5000_1402, w_5000_1403, w_5000_1404, w_5000_1405, w_5000_1406, w_5000_1407, w_5000_1408, w_5000_1409, w_5000_1410, w_5000_1411, w_5000_1412, w_5000_1413, w_5000_1414, w_5000_1415, w_5000_1416, w_5000_1417, w_5000_1418, w_5000_1419, w_5000_1420, w_5000_1421, w_5000_1422, w_5000_1423, w_5000_1424, w_5000_1425, w_5000_1426, w_5000_1427, w_5000_1428, w_5000_1429, w_5000_1430, w_5000_1431, w_5000_1432, w_5000_1433, w_5000_1434, w_5000_1435, w_5000_1436, w_5000_1437, w_5000_1438, w_5000_1439, w_5000_1440, w_5000_1441, w_5000_1442, w_5000_1443, w_5000_1444, w_5000_1445, w_5000_1446, w_5000_1447, w_5000_1448, w_5000_1449, w_5000_1450, w_5000_1451, w_5000_1452, w_5000_1453, w_5000_1454, w_5000_1455, w_5000_1456, w_5000_1457, w_5000_1458, w_5000_1459, w_5000_1460, w_5000_1461, w_5000_1462, w_5000_1463, w_5000_1464, w_5000_1465, w_5000_1466, w_5000_1467, w_5000_1468, w_5000_1469, w_5000_1470, w_5000_1471, w_5000_1472, w_5000_1473, w_5000_1474, w_5000_1475, w_5000_1476, w_5000_1477, w_5000_1478, w_5000_1479, w_5000_1480, w_5000_1481, w_5000_1482, w_5000_1483, w_5000_1484, w_5000_1485, w_5000_1486, w_5000_1487, w_5000_1488, w_5000_1489, w_5000_1490, w_5000_1491, w_5000_1492, w_5000_1493, w_5000_1494, w_5000_1495, w_5000_1496, w_5000_1497, w_5000_1498, w_5000_1499, w_5000_1500, w_5000_1501, w_5000_1502, w_5000_1503, w_5000_1504, w_5000_1505, w_5000_1506, w_5000_1507, w_5000_1508, w_5000_1509, w_5000_1510, w_5000_1511, w_5000_1512, w_5000_1513, w_5000_1514, w_5000_1515, w_5000_1516, w_5000_1517, w_5000_1518, w_5000_1519, w_5000_1520, w_5000_1521, w_5000_1522, w_5000_1523, w_5000_1524, w_5000_1525, w_5000_1526, w_5000_1527, w_5000_1528, w_5000_1529, w_5000_1530, w_5000_1531, w_5000_1532, w_5000_1533, w_5000_1534, w_5000_1535, w_5000_1536, w_5000_1537, w_5000_1538, w_5000_1539, w_5000_1540, w_5000_1541, w_5000_1542, w_5000_1543, w_5000_1544, w_5000_1545, w_5000_1546, w_5000_1547, w_5000_1548, w_5000_1549, w_5000_1550, w_5000_1551, w_5000_1552, w_5000_1553, w_5000_1554, w_5000_1555, w_5000_1556, w_5000_1557, w_5000_1558, w_5000_1559, w_5000_1560, w_5000_1561, w_5000_1562, w_5000_1563, w_5000_1564, w_5000_1565, w_5000_1566, w_5000_1567, w_5000_1568, w_5000_1569, w_5000_1570, w_5000_1571, w_5000_1572, w_5000_1573, w_5000_1574, w_5000_1575, w_5000_1576, w_5000_1577, w_5000_1578, w_5000_1579, w_5000_1580, w_5000_1581, w_5000_1582, w_5000_1583, w_5000_1584, w_5000_1585, w_5000_1586, w_5000_1587, w_5000_1588, w_5000_1589, w_5000_1590, w_5000_1591, w_5000_1592, w_5000_1593, w_5000_1594, w_5000_1595, w_5000_1596, w_5000_1597, w_5000_1598, w_5000_1599, w_5000_1600, w_5000_1601, w_5000_1602, w_5000_1603, w_5000_1604, w_5000_1605, w_5000_1606, w_5000_1607, w_5000_1608, w_5000_1609, w_5000_1610, w_5000_1611, w_5000_1612, w_5000_1613, w_5000_1614, w_5000_1615, w_5000_1616, w_5000_1617, w_5000_1618, w_5000_1619, w_5000_1620, w_5000_1621, w_5000_1622, w_5000_1623, w_5000_1624, w_5000_1625, w_5000_1626, w_5000_1627, w_5000_1628, w_5000_1629, w_5000_1630, w_5000_1631, w_5000_1632, w_5000_1633, w_5000_1634, w_5000_1635, w_5000_1636, w_5000_1637, w_5000_1638, w_5000_1639, w_5000_1640, w_5000_1641, w_5000_1642, w_5000_1643, w_5000_1644, w_5000_1645, w_5000_1646, w_5000_1647, w_5000_1648, w_5000_1649, w_5000_1650, w_5000_1651, w_5000_1652, w_5000_1653, w_5000_1654, w_5000_1655, w_5000_1656, w_5000_1657, w_5000_1658, w_5000_1659, w_5000_1660, w_5000_1661, w_5000_1662, w_5000_1663, w_5000_1664, w_5000_1665, w_5000_1666, w_5000_1667, w_5000_1668, w_5000_1669, w_5000_1670, w_5000_1671, w_5000_1672, w_5000_1673, w_5000_1674, w_5000_1675, w_5000_1676, w_5000_1677, w_5000_1678, w_5000_1679, w_5000_1680, w_5000_1681, w_5000_1682, w_5000_1683, w_5000_1684, w_5000_1685, w_5000_1686, w_5000_1687, w_5000_1688, w_5000_1689, w_5000_1690, w_5000_1691, w_5000_1692, w_5000_1693, w_5000_1694, w_5000_1695, w_5000_1696, w_5000_1697, w_5000_1698, w_5000_1699, w_5000_1700, w_5000_1701, w_5000_1702, w_5000_1703, w_5000_1704, w_5000_1705, w_5000_1706, w_5000_1707, w_5000_1708, w_5000_1709, w_5000_1710, w_5000_1711, w_5000_1712, w_5000_1713, w_5000_1714, w_5000_1715, w_5000_1716, w_5000_1717, w_5000_1718, w_5000_1719, w_5000_1720, w_5000_1721, w_5000_1722, w_5000_1723, w_5000_1724, w_5000_1725, w_5000_1726, w_5000_1727, w_5000_1728, w_5000_1729, w_5000_1730, w_5000_1731, w_5000_1732, w_5000_1733, w_5000_1734, w_5000_1735, w_5000_1736, w_5000_1737, w_5000_1738, w_5000_1739, w_5000_1740, w_5000_1741, w_5000_1742, w_5000_1743, w_5000_1744, w_5000_1745, w_5000_1746, w_5000_1747, w_5000_1748, w_5000_1749, w_5000_1750, w_5000_1751, w_5000_1752, w_5000_1753, w_5000_1754, w_5000_1755, w_5000_1756, w_5000_1757, w_5000_1758, w_5000_1759, w_5000_1760, w_5000_1761, w_5000_1762, w_5000_1763, w_5000_1764, w_5000_1765, w_5000_1766, w_5000_1767, w_5000_1768, w_5000_1769, w_5000_1770, w_5000_1771, w_5000_1772, w_5000_1773, w_5000_1774, w_5000_1775, w_5000_1776, w_5000_1777, w_5000_1778, w_5000_1779, w_5000_1780, w_5000_1781, w_5000_1782, w_5000_1783, w_5000_1784, w_5000_1785, w_5000_1786, w_5000_1787, w_5000_1788, w_5000_1789, w_5000_1790, w_5000_1791, w_5000_1792, w_5000_1793, w_5000_1794, w_5000_1795, w_5000_1796, w_5000_1797, w_5000_1798, w_5000_1799, w_5000_1800, w_5000_1801, w_5000_1802, w_5000_1803, w_5000_1804, w_5000_1805, w_5000_1806, w_5000_1807, w_5000_1808, w_5000_1809, w_5000_1810, w_5000_1811, w_5000_1812, w_5000_1813, w_5000_1814, w_5000_1815, w_5000_1816, w_5000_1817, w_5000_1818, w_5000_1819, w_5000_1820, w_5000_1821, w_5000_1822, w_5000_1823, w_5000_1824, w_5000_1825, w_5000_1826, w_5000_1827, w_5000_1828, w_5000_1829, w_5000_1830, w_5000_1831, w_5000_1832, w_5000_1833, w_5000_1834, w_5000_1835, w_5000_1836, w_5000_1837, w_5000_1838, w_5000_1839, w_5000_1840, w_5000_1841, w_5000_1842, w_5000_1843, w_5000_1844, w_5000_1845, w_5000_1846, w_5000_1847, w_5000_1848, w_5000_1849, w_5000_1850, w_5000_1851, w_5000_1852, w_5000_1853, w_5000_1854, w_5000_1855, w_5000_1856, w_5000_1857, w_5000_1858, w_5000_1859, w_5000_1860, w_5000_1861, w_5000_1862, w_5000_1863, w_5000_1864, w_5000_1865, w_5000_1866, w_5000_1867, w_5000_1868, w_5000_1869, w_5000_1870, w_5000_1871, w_5000_1872, w_5000_1873, w_5000_1874, w_5000_1875, w_5000_1876, w_5000_1877, w_5000_1878, w_5000_1879, w_5000_1880, w_5000_1881, w_5000_1882, w_5000_1883, w_5000_1884, w_5000_1885, w_5000_1886, w_5000_1887, w_5000_1888, w_5000_1889, w_5000_1890, w_5000_1891, w_5000_1892, w_5000_1893, w_5000_1894, w_5000_1895, w_5000_1896, w_5000_1897, w_5000_1898, w_5000_1899, w_5000_1900, w_5000_1901, w_5000_1902, w_5000_1903, w_5000_1904, w_5000_1905, w_5000_1906, w_5000_1907, w_5000_1908, w_5000_1909, w_5000_1910, w_5000_1911, w_5000_1912, w_5000_1913, w_5000_1914, w_5000_1915, w_5000_1916, w_5000_1917, w_5000_1918, w_5000_1919, w_5000_1920, w_5000_1921, w_5000_1922, w_5000_1923, w_5000_1924, w_5000_1925, w_5000_1926, w_5000_1927, w_5000_1928, w_5000_1929, w_5000_1930, w_5000_1931, w_5000_1932, w_5000_1933, w_5000_1934, w_5000_1935, w_5000_1936, w_5000_1937, w_5000_1938, w_5000_1939, w_5000_1940, w_5000_1941, w_5000_1942, w_5000_1943, w_5000_1944, w_5000_1945, w_5000_1946, w_5000_1947, w_5000_1948, w_5000_1949, w_5000_1950, w_5000_1951, w_5000_1952, w_5000_1953, w_5000_1954, w_5000_1955, w_5000_1956, w_5000_1957, w_5000_1958, w_5000_1959, w_5000_1960, w_5000_1961, w_5000_1962, w_5000_1963, w_5000_1964, w_5000_1965, w_5000_1966, w_5000_1967, w_5000_1968, w_5000_1969, w_5000_1970, w_5000_1971, w_5000_1972, w_5000_1973, w_5000_1974, w_5000_1975, w_5000_1976, w_5000_1977, w_5000_1978, w_5000_1979, w_5000_1980, w_5000_1981, w_5000_1982, w_5000_1983, w_5000_1984, w_5000_1985, w_5000_1986, w_5000_1987, w_5000_1988, w_5000_1989, w_5000_1990, w_5000_1991, w_5000_1992, w_5000_1993, w_5000_1994, w_5000_1995, w_5000_1996, w_5000_1997, w_5000_1998, w_5000_1999, w_5000_2000, w_5000_2001, w_5000_2002, w_5000_2003, w_5000_2004, w_5000_2005, w_5000_2006, w_5000_2007, w_5000_2008, w_5000_2009, w_5000_2010, w_5000_2011, w_5000_2012, w_5000_2013, w_5000_2014, w_5000_2015, w_5000_2016, w_5000_2017, w_5000_2018, w_5000_2019, w_5000_2020, w_5000_2021, w_5000_2022, w_5000_2023, w_5000_2024, w_5000_2025, w_5000_2026, w_5000_2027, w_5000_2028, w_5000_2029, w_5000_2030, w_5000_2031, w_5000_2032, w_5000_2033, w_5000_2034, w_5000_2035, w_5000_2036, w_5000_2037, w_5000_2038, w_5000_2039, w_5000_2040, w_5000_2041, w_5000_2042, w_5000_2043, w_5000_2044, w_5000_2045, w_5000_2046, w_5000_2047, w_5000_2048, w_5000_2049, w_5000_2050, w_5000_2051, w_5000_2052, w_5000_2053, w_5000_2054, w_5000_2055, w_5000_2056, w_5000_2057, w_5000_2058, w_5000_2059, w_5000_2060, w_5000_2061, w_5000_2062, w_5000_2063, w_5000_2064, w_5000_2065, w_5000_2066, w_5000_2067, w_5000_2068, w_5000_2069, w_5000_2070, w_5000_2071, w_5000_2072, w_5000_2073, w_5000_2074, w_5000_2075, w_5000_2076, w_5000_2077, w_5000_2078, w_5000_2079, w_5000_2080, w_5000_2081, w_5000_2082, w_5000_2083, w_5000_2084, w_5000_2085, w_5000_2086, w_5000_2087, w_5000_2088, w_5000_2089, w_5000_2090, w_5000_2091, w_5000_2092, w_5000_2093, w_5000_2094, w_5000_2095, w_5000_2096, w_5000_2097, w_5000_2098, w_5000_2099, w_5000_2100, w_5000_2101, w_5000_2102, w_5000_2103, w_5000_2104, w_5000_2105, w_5000_2106, w_5000_2107, w_5000_2108, w_5000_2109, w_5000_2110, w_5000_2111, w_5000_2112, w_5000_2113, w_5000_2114, w_5000_2115, w_5000_2116, w_5000_2117, w_5000_2118, w_5000_2119, w_5000_2120, w_5000_2121, w_5000_2122, w_5000_2123, w_5000_2124, w_5000_2125, w_5000_2126, w_5000_2127, w_5000_2128, w_5000_2129, w_5000_2130, w_5000_2131, w_5000_2132, w_5000_2133, w_5000_2134, w_5000_2135, w_5000_2136, w_5000_2137, w_5000_2138, w_5000_2139, w_5000_2140, w_5000_2141, w_5000_2142, w_5000_2143, w_5000_2144, w_5000_2145, w_5000_2146, w_5000_2147, w_5000_2148, w_5000_2149, w_5000_2150, w_5000_2151, w_5000_2152, w_5000_2153, w_5000_2154, w_5000_2155, w_5000_2156, w_5000_2157, w_5000_2158, w_5000_2159, w_5000_2160, w_5000_2161, w_5000_2162, w_5000_2163, w_5000_2164, w_5000_2165, w_5000_2166, w_5000_2167, w_5000_2168, w_5000_2169, w_5000_2170, w_5000_2171, w_5000_2172, w_5000_2173, w_5000_2174, w_5000_2175, w_5000_2176, w_5000_2177, w_5000_2178, w_5000_2179, w_5000_2180, w_5000_2181, w_5000_2182, w_5000_2183, w_5000_2184, w_5000_2185, w_5000_2186, w_5000_2187, w_5000_2188, w_5000_2189, w_5000_2190, w_5000_2191, w_5000_2192, w_5000_2193, w_5000_2194, w_5000_2195, w_5000_2196, w_5000_2197, w_5000_2198, w_5000_2199, w_5000_2200, w_5000_2201, w_5000_2202, w_5000_2203, w_5000_2204, w_5000_2205, w_5000_2206, w_5000_2207, w_5000_2208, w_5000_2209, w_5000_2210, w_5000_2211, w_5000_2212, w_5000_2213, w_5000_2214, w_5000_2215, w_5000_2216, w_5000_2217, w_5000_2218, w_5000_2219, w_5000_2220, w_5000_2221, w_5000_2222, w_5000_2223, w_5000_2224, w_5000_2225, w_5000_2226, w_5000_2227, w_5000_2228, w_5000_2229, w_5000_2230, w_5000_2231, w_5000_2232, w_5000_2233, w_5000_2234, w_5000_2235, w_5000_2236, w_5000_2237, w_5000_2238, w_5000_2239, w_5000_2240, w_5000_2241, w_5000_2242, w_5000_2243, w_5000_2244, w_5000_2245, w_5000_2246, w_5000_2247, w_5000_2248, w_5000_2249, w_5000_2250, w_5000_2251, w_5000_2252, w_5000_2253, w_5000_2254, w_5000_2255, w_5000_2256, w_5000_2257, w_5000_2258, w_5000_2259, w_5000_2260, w_5000_2261, w_5000_2262, w_5000_2263, w_5000_2264, w_5000_2265, w_5000_2266, w_5000_2267, w_5000_2268, w_5000_2269, w_5000_2270, w_5000_2271, w_5000_2272, w_5000_2273, w_5000_2274, w_5000_2275, w_5000_2276, w_5000_2277, w_5000_2278, w_5000_2279, w_5000_2280, w_5000_2281, w_5000_2282, w_5000_2283, w_5000_2284, w_5000_2285, w_5000_2286, w_5000_2287, w_5000_2288, w_5000_2289, w_5000_2290, w_5000_2291, w_5000_2292, w_5000_2293, w_5000_2294, w_5000_2295, w_5000_2296, w_5000_2297, w_5000_2298, w_5000_2299, w_5000_2300, w_5000_2301, w_5000_2302, w_5000_2303, w_5000_2304, w_5000_2305, w_5000_2306, w_5000_2307, w_5000_2308, w_5000_2309, w_5000_2310, w_5000_2311, w_5000_2312, w_5000_2313, w_5000_2314, w_5000_2315, w_5000_2316, w_5000_2317, w_5000_2318, w_5000_2319, w_5000_2320, w_5000_2321, w_5000_2322, w_5000_2323, w_5000_2324, w_5000_2325, w_5000_2326, w_5000_2327, w_5000_2328, w_5000_2329, w_5000_2330, w_5000_2331, w_5000_2332, w_5000_2333, w_5000_2334, w_5000_2335, w_5000_2336, w_5000_2337, w_5000_2338, w_5000_2339, w_5000_2340, w_5000_2341, w_5000_2342, w_5000_2343, w_5000_2344, w_5000_2345, w_5000_2346, w_5000_2347, w_5000_2348, w_5000_2349, w_5000_2350, w_5000_2351, w_5000_2352, w_5000_2353, w_5000_2354, w_5000_2355, w_5000_2356, w_5000_2357, w_5000_2358, w_5000_2359, w_5000_2360, w_5000_2361, w_5000_2362, w_5000_2363, w_5000_2364, w_5000_2365, w_5000_2366, w_5000_2367, w_5000_2368, w_5000_2369, w_5000_2370, w_5000_2371, w_5000_2372, w_5000_2373, w_5000_2374, w_5000_2375, w_5000_2376, w_5000_2377, w_5000_2378, w_5000_2379, w_5000_2380, w_5000_2381, w_5000_2382, w_5000_2383, w_5000_2384, w_5000_2385, w_5000_2386, w_5000_2387, w_5000_2388, w_5000_2389, w_5000_2390, w_5000_2391, w_5000_2392, w_5000_2393, w_5000_2394, w_5000_2395, w_5000_2396, w_5000_2397, w_5000_2398, w_5000_2399, w_5000_2400, w_5000_2401, w_5000_2402, w_5000_2403, w_5000_2404, w_5000_2405, w_5000_2406, w_5000_2407, w_5000_2408, w_5000_2409, w_5000_2410, w_5000_2411, w_5000_2412, w_5000_2413, w_5000_2414, w_5000_2415, w_5000_2416, w_5000_2417, w_5000_2418, w_5000_2419, w_5000_2420, w_5000_2421, w_5000_2422, w_5000_2423, w_5000_2424, w_5000_2425, w_5000_2426, w_5000_2427, w_5000_2428, w_5000_2429, w_5000_2430, w_5000_2431, w_5000_2432, w_5000_2433, w_5000_2434, w_5000_2435, w_5000_2436, w_5000_2437, w_5000_2438, w_5000_2439, w_5000_2440, w_5000_2441, w_5000_2442, w_5000_2443, w_5000_2444, w_5000_2445, w_5000_2446, w_5000_2447, w_5000_2448, w_5000_2449, w_5000_2450, w_5000_2451, w_5000_2452, w_5000_2453, w_5000_2454, w_5000_2455, w_5000_2456, w_5000_2457, w_5000_2458, w_5000_2459, w_5000_2460, w_5000_2461, w_5000_2462, w_5000_2463, w_5000_2464, w_5000_2465, w_5000_2466, w_5000_2467, w_5000_2468, w_5000_2469, w_5000_2470, w_5000_2471, w_5000_2472, w_5000_2473, w_5000_2474, w_5000_2475, w_5000_2476, w_5000_2477, w_5000_2478, w_5000_2479, w_5000_2480, w_5000_2481, w_5000_2482, w_5000_2483, w_5000_2484, w_5000_2485, w_5000_2486, w_5000_2487, w_5000_2488, w_5000_2489, w_5000_2490, w_5000_2491, w_5000_2492, w_5000_2493, w_5000_2494, w_5000_2495, w_5000_2496, w_5000_2497, w_5000_2498, w_5000_2499, w_5000_2500, w_5000_2501, w_5000_2502, w_5000_2503, w_5000_2504, w_5000_2505, w_5000_2506, w_5000_2507, w_5000_2508, w_5000_2509, w_5000_2510, w_5000_2511, w_5000_2512, w_5000_2513, w_5000_2514, w_5000_2515, w_5000_2516, w_5000_2517, w_5000_2518, w_5000_2519, w_5000_2520, w_5000_2521, w_5000_2522, w_5000_2523, w_5000_2524, w_5000_2525, w_5000_2526, w_5000_2527, w_5000_2528, w_5000_2529, w_5000_2530, w_5000_2531, w_5000_2532, w_5000_2533, w_5000_2534, w_5000_2535, w_5000_2536, w_5000_2537, w_5000_2538, w_5000_2539, w_5000_2540, w_5000_2541, w_5000_2542, w_5000_2543, w_5000_2544, w_5000_2545, w_5000_2546, w_5000_2547, w_5000_2548, w_5000_2549, w_5000_2550, w_5000_2551, w_5000_2552, w_5000_2553, w_5000_2554, w_5000_2555, w_5000_2556, w_5000_2557, w_5000_2558, w_5000_2559, w_5000_2560, w_5000_2561, w_5000_2562, w_5000_2563, w_5000_2564, w_5000_2565, w_5000_2566, w_5000_2567, w_5000_2568, w_5000_2569, w_5000_2570, w_5000_2571, w_5000_2572, w_5000_2573, w_5000_2574, w_5000_2575, w_5000_2576, w_5000_2577, w_5000_2578, w_5000_2579, w_5000_2580, w_5000_2581, w_5000_2582, w_5000_2583, w_5000_2584, w_5000_2585, w_5000_2586, w_5000_2587, w_5000_2588, w_5000_2589, w_5000_2590, w_5000_2591, w_5000_2592, w_5000_2593, w_5000_2594, w_5000_2595, w_5000_2596, w_5000_2597, w_5000_2598, w_5000_2599, w_5000_2600, w_5000_2601, w_5000_2602, w_5000_2603, w_5000_2604, w_5000_2605, w_5000_2606, w_5000_2607, w_5000_2608, w_5000_2609, w_5000_2610, w_5000_2611, w_5000_2612, w_5000_2613, w_5000_2614, w_5000_2615, w_5000_2616, w_5000_2617, w_5000_2618, w_5000_2619, w_5000_2620, w_5000_2621, w_5000_2622, w_5000_2623, w_5000_2624, w_5000_2625, w_5000_2626, w_5000_2627, w_5000_2628, w_5000_2629, w_5000_2630, w_5000_2631, w_5000_2632, w_5000_2633, w_5000_2634, w_5000_2635, w_5000_2636, w_5000_2637, w_5000_2638, w_5000_2639, w_5000_2640, w_5000_2641, w_5000_2642, w_5000_2643, w_5000_2644, w_5000_2645, w_5000_2646, w_5000_2647, w_5000_2648, w_5000_2649, w_5000_2650, w_5000_2651, w_5000_2652, w_5000_2653, w_5000_2654, w_5000_2655, w_5000_2656, w_5000_2657, w_5000_2658, w_5000_2659, w_5000_2660, w_5000_2661, w_5000_2662, w_5000_2663, w_5000_2664, w_5000_2665, w_5000_2666, w_5000_2667, w_5000_2668, w_5000_2669, w_5000_2670, w_5000_2671, w_5000_2672, w_5000_2673, w_5000_2674, w_5000_2675, w_5000_2676, w_5000_2677, w_5000_2678, w_5000_2679, w_5000_2680, w_5000_2681, w_5000_2682, w_5000_2683, w_5000_2684, w_5000_2685, w_5000_2686, w_5000_2687, w_5000_2688, w_5000_2689, w_5000_2690, w_5000_2691, w_5000_2692, w_5000_2693, w_5000_2694, w_5000_2695, w_5000_2696, w_5000_2697, w_5000_2698, w_5000_2699, w_5000_2700, w_5000_2701, w_5000_2702, w_5000_2703, w_5000_2704, w_5000_2705, w_5000_2706, w_5000_2707, w_5000_2708, w_5000_2709, w_5000_2710, w_5000_2711, w_5000_2712, w_5000_2713, w_5000_2714, w_5000_2715, w_5000_2716, w_5000_2717, w_5000_2718, w_5000_2719, w_5000_2720, w_5000_2721, w_5000_2722, w_5000_2723, w_5000_2724, w_5000_2725, w_5000_2726, w_5000_2727, w_5000_2728, w_5000_2729, w_5000_2730, w_5000_2731, w_5000_2732, w_5000_2733, w_5000_2734, w_5000_2735, w_5000_2736, w_5000_2737, w_5000_2738, w_5000_2739, w_5000_2740, w_5000_2741, w_5000_2742, w_5000_2743, w_5000_2744, w_5000_2745, w_5000_2746, w_5000_2747, w_5000_2748, w_5000_2749, w_5000_2750, w_5000_2751, w_5000_2752, w_5000_2753, w_5000_2754, w_5000_2755, w_5000_2756, w_5000_2757, w_5000_2758, w_5000_2759, w_5000_2760, w_5000_2761, w_5000_2762, w_5000_2763, w_5000_2764, w_5000_2765, w_5000_2766, w_5000_2767, w_5000_2768, w_5000_2769, w_5000_2770, w_5000_2771, w_5000_2772, w_5000_2773, w_5000_2774, w_5000_2775, w_5000_2776, w_5000_2777, w_5000_2778, w_5000_2779, w_5000_2780, w_5000_2781, w_5000_2782, w_5000_2783, w_5000_2784, w_5000_2785, w_5000_2786, w_5000_2787, w_5000_2788, w_5000_2789, w_5000_2790, w_5000_2791, w_5000_2792, w_5000_2793, w_5000_2794, w_5000_2795, w_5000_2796, w_5000_2797, w_5000_2798, w_5000_2799, w_5000_2800, w_5000_2801, w_5000_2802, w_5000_2803, w_5000_2804, w_5000_2805, w_5000_2806, w_5000_2807, w_5000_2808, w_5000_2809, w_5000_2810, w_5000_2811, w_5000_2812, w_5000_2813, w_5000_2814, w_5000_2815, w_5000_2816, w_5000_2817, w_5000_2818, w_5000_2819, w_5000_2820, w_5000_2821, w_5000_2822, w_5000_2823, w_5000_2824, w_5000_2825, w_5000_2826, w_5000_2827, w_5000_2828, w_5000_2829, w_5000_2830, w_5000_2831, w_5000_2832, w_5000_2833, w_5000_2834, w_5000_2835, w_5000_2836, w_5000_2837, w_5000_2838, w_5000_2839, w_5000_2840, w_5000_2841, w_5000_2842, w_5000_2843, w_5000_2844, w_5000_2845, w_5000_2846, w_5000_2847, w_5000_2848, w_5000_2849, w_5000_2850, w_5000_2851, w_5000_2852, w_5000_2853, w_5000_2854, w_5000_2855, w_5000_2856, w_5000_2857, w_5000_2858, w_5000_2859, w_5000_2860, w_5000_2861, w_5000_2862, w_5000_2863, w_5000_2864, w_5000_2865, w_5000_2866, w_5000_2867, w_5000_2868, w_5000_2869, w_5000_2870, w_5000_2871, w_5000_2872, w_5000_2873, w_5000_2874, w_5000_2875, w_5000_2876, w_5000_2877, w_5000_2878, w_5000_2879, w_5000_2880, w_5000_2881, w_5000_2882, w_5000_2883, w_5000_2884, w_5000_2885, w_5000_2886, w_5000_2887, w_5000_2888, w_5000_2889, w_5000_2890, w_5000_2891, w_5000_2892, w_5000_2893, w_5000_2894, w_5000_2895, w_5000_2896, w_5000_2897, w_5000_2898, w_5000_2899, w_5000_2900, w_5000_2901, w_5000_2902, w_5000_2903, w_5000_2904, w_5000_2905, w_5000_2906, w_5000_2907, w_5000_2908, w_5000_2909, w_5000_2910, w_5000_2911, w_5000_2912, w_5000_2913, w_5000_2914, w_5000_2915, w_5000_2916, w_5000_2917, w_5000_2918, w_5000_2919, w_5000_2920, w_5000_2921, w_5000_2922, w_5000_2923, w_5000_2924, w_5000_2925, w_5000_2926, w_5000_2927, w_5000_2928, w_5000_2929, w_5000_2930, w_5000_2931, w_5000_2932, w_5000_2933, w_5000_2934, w_5000_2935, w_5000_2936, w_5000_2937, w_5000_2938, w_5000_2939, w_5000_2940, w_5000_2941, w_5000_2942, w_5000_2943, w_5000_2944, w_5000_2945, w_5000_2946, w_5000_2947, w_5000_2948, w_5000_2949, w_5000_2950, w_5000_2951, w_5000_2952, w_5000_2953, w_5000_2954, w_5000_2955, w_5000_2956, w_5000_2957, w_5000_2958, w_5000_2959, w_5000_2960, w_5000_2961, w_5000_2962, w_5000_2963, w_5000_2964, w_5000_2965, w_5000_2966, w_5000_2967, w_5000_2968, w_5000_2969, w_5000_2970, w_5000_2971, w_5000_2972, w_5000_2973, w_5000_2974, w_5000_2975, w_5000_2976, w_5000_2977, w_5000_2978, w_5000_2979, w_5000_2980, w_5000_2981, w_5000_2982, w_5000_2983, w_5000_2984, w_5000_2985, w_5000_2986, w_5000_2987, w_5000_2988, w_5000_2989, w_5000_2990, w_5000_2991, w_5000_2992, w_5000_2993, w_5000_2994, w_5000_2995, w_5000_2996, w_5000_2997, w_5000_2998, w_5000_2999, w_5000_3000, w_5000_3001, w_5000_3002, w_5000_3003, w_5000_3004, w_5000_3005, w_5000_3006, w_5000_3007, w_5000_3008, w_5000_3009, w_5000_3010, w_5000_3011, w_5000_3012, w_5000_3013, w_5000_3014, w_5000_3015, w_5000_3016, w_5000_3017, w_5000_3018, w_5000_3019, w_5000_3020, w_5000_3021, w_5000_3022, w_5000_3023, w_5000_3024, w_5000_3025, w_5000_3026, w_5000_3027, w_5000_3028, w_5000_3029, w_5000_3030, w_5000_3031, w_5000_3032, w_5000_3033, w_5000_3034, w_5000_3035, w_5000_3036, w_5000_3037, w_5000_3038, w_5000_3039, w_5000_3040, w_5000_3041, w_5000_3042, w_5000_3043, w_5000_3044, w_5000_3045, w_5000_3046, w_5000_3047, w_5000_3048, w_5000_3049, w_5000_3050, w_5000_3051, w_5000_3052, w_5000_3053, w_5000_3054, w_5000_3055, w_5000_3056, w_5000_3057, w_5000_3058, w_5000_3059, w_5000_3060, w_5000_3061, w_5000_3062, w_5000_3063, w_5000_3064, w_5000_3065, w_5000_3066, w_5000_3067, w_5000_3068, w_5000_3069, w_5000_3070, w_5000_3071, w_5000_3072, w_5000_3073, w_5000_3074, w_5000_3075, w_5000_3076, w_5000_3077, w_5000_3078, w_5000_3079, w_5000_3080, w_5000_3081, w_5000_3082, w_5000_3083, w_5000_3084, w_5000_3085, w_5000_3086, w_5000_3087, w_5000_3088, w_5000_3089, w_5000_3090, w_5000_3091, w_5000_3092, w_5000_3093, w_5000_3094, w_5000_3095, w_5000_3096, w_5000_3097, w_5000_3098, w_5000_3099, w_5000_3100, w_5000_3101, w_5000_3102, w_5000_3103, w_5000_3104, w_5000_3105, w_5000_3106, w_5000_3107, w_5000_3108, w_5000_3109, w_5000_3110, w_5000_3111, w_5000_3112, w_5000_3113, w_5000_3114, w_5000_3115, w_5000_3116, w_5000_3117, w_5000_3118, w_5000_3119, w_5000_3120, w_5000_3121, w_5000_3122, w_5000_3123, w_5000_3124, w_5000_3125, w_5000_3126, w_5000_3127, w_5000_3128, w_5000_3129, w_5000_3130, w_5000_3131, w_5000_3132, w_5000_3133, w_5000_3134, w_5000_3135, w_5000_3136, w_5000_3137, w_5000_3138, w_5000_3139, w_5000_3140, w_5000_3141, w_5000_3142, w_5000_3143, w_5000_3144, w_5000_3145, w_5000_3146, w_5000_3147, w_5000_3148, w_5000_3149, w_5000_3150, w_5000_3151, w_5000_3152, w_5000_3153, w_5000_3154, w_5000_3155, w_5000_3156, w_5000_3157, w_5000_3158, w_5000_3159, w_5000_3160, w_5000_3161, w_5000_3162, w_5000_3163, w_5000_3164, w_5000_3165, w_5000_3166, w_5000_3167, w_5000_3168, w_5000_3169, w_5000_3170, w_5000_3171, w_5000_3172, w_5000_3173, w_5000_3174, w_5000_3175, w_5000_3176, w_5000_3177, w_5000_3178, w_5000_3179, w_5000_3180, w_5000_3181, w_5000_3182, w_5000_3183, w_5000_3184, w_5000_3185, w_5000_3186, w_5000_3187, w_5000_3188, w_5000_3189, w_5000_3190, w_5000_3191, w_5000_3192, w_5000_3193, w_5000_3194, w_5000_3195, w_5000_3196, w_5000_3197, w_5000_3198, w_5000_3199, w_5000_3200, w_5000_3201, w_5000_3202, w_5000_3203, w_5000_3204, w_5000_3205, w_5000_3206, w_5000_3207, w_5000_3208, w_5000_3209, w_5000_3210, w_5000_3211, w_5000_3212, w_5000_3213, w_5000_3214, w_5000_3215, w_5000_3216, w_5000_3217, w_5000_3218, w_5000_3219, w_5000_3220, w_5000_3221, w_5000_3222, w_5000_3223, w_5000_3224, w_5000_3225, w_5000_3226, w_5000_3227, w_5000_3228, w_5000_3229, w_5000_3230, w_5000_3231, w_5000_3232, w_5000_3233, w_5000_3234, w_5000_3235, w_5000_3236, w_5000_3237, w_5000_3238, w_5000_3239, w_5000_3240, w_5000_3241, w_5000_3242, w_5000_3243, w_5000_3244, w_5000_3245, w_5000_3246, w_5000_3247, w_5000_3248, w_5000_3249, w_5000_3250, w_5000_3251, w_5000_3252, w_5000_3253, w_5000_3254, w_5000_3255, w_5000_3256, w_5000_3257, w_5000_3258, w_5000_3259, w_5000_3260, w_5000_3261, w_5000_3262, w_5000_3263, w_5000_3264, w_5000_3265, w_5000_3266, w_5000_3267, w_5000_3268, w_5000_3269, w_5000_3270, w_5000_3271, w_5000_3272, w_5000_3273, w_5000_3274, w_5000_3275, w_5000_3276, w_5000_3277, w_5000_3278, w_5000_3279, w_5000_3280, w_5000_3281, w_5000_3282, w_5000_3283, w_5000_3284, w_5000_3285, w_5000_3286, w_5000_3287, w_5000_3288, w_5000_3289, w_5000_3290, w_5000_3291, w_5000_3292, w_5000_3293, w_5000_3294, w_5000_3295, w_5000_3296, w_5000_3297, w_5000_3298, w_5000_3299, w_5000_3300, w_5000_3301, w_5000_3302, w_5000_3303, w_5000_3304, w_5000_3305, w_5000_3306, w_5000_3307, w_5000_3308, w_5000_3309, w_5000_3310, w_5000_3311, w_5000_3312, w_5000_3313, w_5000_3314, w_5000_3315, w_5000_3316, w_5000_3317, w_5000_3318, w_5000_3319, w_5000_3320, w_5000_3321, w_5000_3322, w_5000_3323, w_5000_3324, w_5000_3325, w_5000_3326, w_5000_3327, w_5000_3328, w_5000_3329, w_5000_3330, w_5000_3331, w_5000_3332, w_5000_3333, w_5000_3334, w_5000_3335, w_5000_3336, w_5000_3337, w_5000_3338, w_5000_3339, w_5000_3340, w_5000_3341, w_5000_3342, w_5000_3343, w_5000_3344, w_5000_3345, w_5000_3346, w_5000_3347, w_5000_3348, w_5000_3349, w_5000_3350, w_5000_3351, w_5000_3352, w_5000_3353, w_5000_3354, w_5000_3355, w_5000_3356, w_5000_3357, w_5000_3358, w_5000_3359, w_5000_3360, w_5000_3361, w_5000_3362, w_5000_3363, w_5000_3364, w_5000_3365, w_5000_3366, w_5000_3367, w_5000_3368, w_5000_3369, w_5000_3370, w_5000_3371, w_5000_3372, w_5000_3373, w_5000_3374, w_5000_3375, w_5000_3376, w_5000_3377, w_5000_3378, w_5000_3379, w_5000_3380, w_5000_3381, w_5000_3382, w_5000_3383, w_5000_3384, w_5000_3385, w_5000_3386, w_5000_3387, w_5000_3388, w_5000_3389, w_5000_3390, w_5000_3391, w_5000_3392, w_5000_3393, w_5000_3394, w_5000_3395, w_5000_3396, w_5000_3397, w_5000_3398, w_5000_3399, w_5000_3400, w_5000_3401, w_5000_3402, w_5000_3403, w_5000_3404, w_5000_3405, w_5000_3406, w_5000_3407, w_5000_3408, w_5000_3409, w_5000_3410, w_5000_3411, w_5000_3412, w_5000_3413, w_5000_3414, w_5000_3415, w_5000_3416, w_5000_3417, w_5000_3418, w_5000_3419, w_5000_3420, w_5000_3421, w_5000_3422, w_5000_3423, w_5000_3424, w_5000_3425, w_5000_3426, w_5000_3427, w_5000_3428, w_5000_3429, w_5000_3430, w_5000_3431, w_5000_3432, w_5000_3433, w_5000_3434, w_5000_3435, w_5000_3436, w_5000_3437, w_5000_3438, w_5000_3439, w_5000_3440, w_5000_3441, w_5000_3442, w_5000_3443, w_5000_3444, w_5000_3445, w_5000_3446, w_5000_3447, w_5000_3448, w_5000_3449, w_5000_3450, w_5000_3451, w_5000_3452, w_5000_3453, w_5000_3454, w_5000_3455, w_5000_3456, w_5000_3457, w_5000_3458, w_5000_3459, w_5000_3460, w_5000_3461, w_5000_3462, w_5000_3463, w_5000_3464, w_5000_3465, w_5000_3466, w_5000_3467, w_5000_3468, w_5000_3469, w_5000_3470, w_5000_3471, w_5000_3472, w_5000_3473, w_5000_3474, w_5000_3475, w_5000_3476, w_5000_3477, w_5000_3478, w_5000_3479, w_5000_3480, w_5000_3481, w_5000_3482, w_5000_3483, w_5000_3484, w_5000_3485, w_5000_3486, w_5000_3487, w_5000_3488, w_5000_3489, w_5000_3490, w_5000_3491, w_5000_3492, w_5000_3493, w_5000_3494, w_5000_3495, w_5000_3496, w_5000_3497, w_5000_3498, w_5000_3499, w_5000_3500, w_5000_3501, w_5000_3502, w_5000_3503, w_5000_3504, w_5000_3505, w_5000_3506, w_5000_3507, w_5000_3508, w_5000_3509, w_5000_3510, w_5000_3511, w_5000_3512, w_5000_3513, w_5000_3514, w_5000_3515, w_5000_3516, w_5000_3517, w_5000_3518, w_5000_3519, w_5000_3520, w_5000_3521, w_5000_3522, w_5000_3523, w_5000_3524, w_5000_3525, w_5000_3526, w_5000_3527, w_5000_3528, w_5000_3529, w_5000_3530, w_5000_3531, w_5000_3532, w_5000_3533, w_5000_3534, w_5000_3535, w_5000_3536, w_5000_3537, w_5000_3538, w_5000_3539, w_5000_3540, w_5000_3541, w_5000_3542, w_5000_3543, w_5000_3544, w_5000_3545, w_5000_3546, w_5000_3547, w_5000_3548, w_5000_3549, w_5000_3550, w_5000_3551, w_5000_3552, w_5000_3553, w_5000_3554, w_5000_3555, w_5000_3556, w_5000_3557, w_5000_3558, w_5000_3559, w_5000_3560, w_5000_3561, w_5000_3562, w_5000_3563, w_5000_3564, w_5000_3565, w_5000_3566, w_5000_3567, w_5000_3568, w_5000_3569, w_5000_3570, w_5000_3571, w_5000_3572, w_5000_3573, w_5000_3574, w_5000_3575, w_5000_3576, w_5000_3577, w_5000_3578, w_5000_3579, w_5000_3580, w_5000_3581, w_5000_3582, w_5000_3583, w_5000_3584, w_5000_3585, w_5000_3586, w_5000_3587, w_5000_3588, w_5000_3589, w_5000_3590, w_5000_3591, w_5000_3592, w_5000_3593, w_5000_3594, w_5000_3595, w_5000_3596, w_5000_3597, w_5000_3598, w_5000_3599, w_5000_3600, w_5000_3601, w_5000_3602, w_5000_3603, w_5000_3604, w_5000_3605, w_5000_3606, w_5000_3607, w_5000_3608, w_5000_3609, w_5000_3610, w_5000_3611, w_5000_3612, w_5000_3613, w_5000_3614, w_5000_3615, w_5000_3616, w_5000_3617, w_5000_3618, w_5000_3619, w_5000_3620, w_5000_3621, w_5000_3622, w_5000_3623, w_5000_3624, w_5000_3625, w_5000_3626, w_5000_3627, w_5000_3628, w_5000_3629, w_5000_3630, w_5000_3631, w_5000_3632, w_5000_3633, w_5000_3634, w_5000_3635, w_5000_3636, w_5000_3637, w_5000_3638, w_5000_3639, w_5000_3640, w_5000_3641, w_5000_3642, w_5000_3643, w_5000_3644, w_5000_3645, w_5000_3646, w_5000_3647, w_5000_3648, w_5000_3649, w_5000_3650, w_5000_3651, w_5000_3652, w_5000_3653, w_5000_3654, w_5000_3655, w_5000_3656, w_5000_3657, w_5000_3658, w_5000_3659, w_5000_3660, w_5000_3661, w_5000_3662, w_5000_3663, w_5000_3664, w_5000_3665, w_5000_3666, w_5000_3667, w_5000_3668, w_5000_3669, w_5000_3670, w_5000_3671, w_5000_3672, w_5000_3673, w_5000_3674, w_5000_3675, w_5000_3676, w_5000_3677, w_5000_3678, w_5000_3679, w_5000_3680, w_5000_3681, w_5000_3682, w_5000_3683, w_5000_3684, w_5000_3685, w_5000_3686, w_5000_3687, w_5000_3688, w_5000_3689, w_5000_3690, w_5000_3691, w_5000_3692, w_5000_3693, w_5000_3694, w_5000_3695, w_5000_3696, w_5000_3697, w_5000_3698, w_5000_3699, w_5000_3700, w_5000_3701, w_5000_3702, w_5000_3703, w_5000_3704, w_5000_3705, w_5000_3706, w_5000_3707, w_5000_3708, w_5000_3709, w_5000_3710, w_5000_3711, w_5000_3712, w_5000_3713, w_5000_3714, w_5000_3715, w_5000_3716, w_5000_3717, w_5000_3718, w_5000_3719, w_5000_3720, w_5000_3721, w_5000_3722, w_5000_3723, w_5000_3724, w_5000_3725, w_5000_3726, w_5000_3727, w_5000_3728, w_5000_3729, w_5000_3730, w_5000_3731, w_5000_3732, w_5000_3733, w_5000_3734, w_5000_3735, w_5000_3736, w_5000_3737, w_5000_3738, w_5000_3739, w_5000_3740, w_5000_3741, w_5000_3742, w_5000_3743, w_5000_3744, w_5000_3745, w_5000_3746, w_5000_3747, w_5000_3748, w_5000_3749, w_5000_3750, w_5000_3751, w_5000_3752, w_5000_3753, w_5000_3754, w_5000_3755, w_5000_3756, w_5000_3757, w_5000_3758, w_5000_3759, w_5000_3760, w_5000_3761, w_5000_3762, w_5000_3763, w_5000_3764, w_5000_3765, w_5000_3766, w_5000_3767, w_5000_3768, w_5000_3769, w_5000_3770, w_5000_3771, w_5000_3772, w_5000_3773, w_5000_3774, w_5000_3775, w_5000_3776, w_5000_3777, w_5000_3778, w_5000_3779, w_5000_3780, w_5000_3781, w_5000_3782, w_5000_3783, w_5000_3784, w_5000_3785, w_5000_3786, w_5000_3787, w_5000_3788, w_5000_3789, w_5000_3790, w_5000_3791, w_5000_3792, w_5000_3793, w_5000_3794, w_5000_3795, w_5000_3796, w_5000_3797, w_5000_3798, w_5000_3799, w_5000_3800, w_5000_3801, w_5000_3802, w_5000_3803, w_5000_3804, w_5000_3805, w_5000_3806, w_5000_3807, w_5000_3808, w_5000_3809, w_5000_3810, w_5000_3811, w_5000_3812, w_5000_3813, w_5000_3814, w_5000_3815, w_5000_3816, w_5000_3817, w_5000_3818, w_5000_3819, w_5000_3820, w_5000_3821, w_5000_3822, w_5000_3823, w_5000_3824, w_5000_3825, w_5000_3826, w_5000_3827, w_5000_3828, w_5000_3829, w_5000_3830, w_5000_3831, w_5000_3832, w_5000_3833, w_5000_3834, w_5000_3835, w_5000_3836, w_5000_3837, w_5000_3838, w_5000_3839, w_5000_3840, w_5000_3841, w_5000_3842, w_5000_3843, w_5000_3844, w_5000_3845, w_5000_3846, w_5000_3847, w_5000_3848, w_5000_3849, w_5000_3850, w_5000_3851, w_5000_3852, w_5000_3853, w_5000_3854, w_5000_3855, w_5000_3856, w_5000_3857, w_5000_3858, w_5000_3859, w_5000_3860, w_5000_3861, w_5000_3862, w_5000_3863, w_5000_3864, w_5000_3865, w_5000_3866, w_5000_3867, w_5000_3868, w_5000_3869, w_5000_3870, w_5000_3871, w_5000_3872, w_5000_3873, w_5000_3874, w_5000_3875, w_5000_3876, w_5000_3877, w_5000_3878, w_5000_3879, w_5000_3880, w_5000_3881, w_5000_3882, w_5000_3883, w_5000_3884, w_5000_3885, w_5000_3886, w_5000_3887, w_5000_3888, w_5000_3889, w_5000_3890, w_5000_3891, w_5000_3892, w_5000_3893, w_5000_3894, w_5000_3895, w_5000_3896, w_5000_3897, w_5000_3898, w_5000_3899, w_5000_3900, w_5000_3901, w_5000_3902, w_5000_3903, w_5000_3904, w_5000_3905, w_5000_3906, w_5000_3907, w_5000_3908, w_5000_3909, w_5000_3910, w_5000_3911, w_5000_3912, w_5000_3913, w_5000_3914, w_5000_3915, w_5000_3916, w_5000_3917, w_5000_3918, w_5000_3919, w_5000_3920, w_5000_3921, w_5000_3922, w_5000_3923, w_5000_3924, w_5000_3925, w_5000_3926, w_5000_3927, w_5000_3928, w_5000_3929, w_5000_3930, w_5000_3931, w_5000_3932, w_5000_3933, w_5000_3934, w_5000_3935, w_5000_3936, w_5000_3937, w_5000_3938, w_5000_3939, w_5000_3940, w_5000_3941, w_5000_3942, w_5000_3943, w_5000_3944, w_5000_3945, w_5000_3946, w_5000_3947, w_5000_3948, w_5000_3949, w_5000_3950, w_5000_3951, w_5000_3952, w_5000_3953, w_5000_3954, w_5000_3955, w_5000_3956, w_5000_3957, w_5000_3958, w_5000_3959, w_5000_3960, w_5000_3961, w_5000_3962, w_5000_3963, w_5000_3964, w_5000_3965, w_5000_3966, w_5000_3967, w_5000_3968, w_5000_3969, w_5000_3970, w_5000_3971, w_5000_3972, w_5000_3973, w_5000_3974, w_5000_3975, w_5000_3976, w_5000_3977, w_5000_3978, w_5000_3979, w_5000_3980, w_5000_3981, w_5000_3982, w_5000_3983, w_5000_3984, w_5000_3985, w_5000_3986, w_5000_3987, w_5000_3988, w_5000_3989, w_5000_3990, w_5000_3991, w_5000_3992, w_5000_3993, w_5000_3994, w_5000_3995, w_5000_3996, w_5000_3997, w_5000_3998, w_5000_3999, w_5000_4000, w_5000_4001, w_5000_4002, w_5000_4003, w_5000_4004, w_5000_4005, w_5000_4006, w_5000_4007, w_5000_4008, w_5000_4009, w_5000_4010, w_5000_4011, w_5000_4012, w_5000_4013, w_5000_4014, w_5000_4015, w_5000_4016, w_5000_4017, w_5000_4018, w_5000_4019, w_5000_4020, w_5000_4021, w_5000_4022, w_5000_4023, w_5000_4024, w_5000_4025, w_5000_4026, w_5000_4027, w_5000_4028, w_5000_4029, w_5000_4030, w_5000_4031, w_5000_4032, w_5000_4033, w_5000_4034, w_5000_4035, w_5000_4036, w_5000_4037, w_5000_4038, w_5000_4039, w_5000_4040, w_5000_4041, w_5000_4042, w_5000_4043, w_5000_4044, w_5000_4045, w_5000_4046, w_5000_4047, w_5000_4048, w_5000_4049, w_5000_4050, w_5000_4051, w_5000_4052, w_5000_4053, w_5000_4054, w_5000_4055, w_5000_4056, w_5000_4057, w_5000_4058, w_5000_4059, w_5000_4060, w_5000_4061, w_5000_4062, w_5000_4063, w_5000_4064, w_5000_4065, w_5000_4066, w_5000_4067, w_5000_4068, w_5000_4069, w_5000_4070, w_5000_4071, w_5000_4072, w_5000_4073, w_5000_4074, w_5000_4075, w_5000_4076, w_5000_4077, w_5000_4078, w_5000_4079, w_5000_4080, w_5000_4081, w_5000_4082, w_5000_4083, w_5000_4084, w_5000_4085, w_5000_4086, w_5000_4087, w_5000_4088, w_5000_4089, w_5000_4090, w_5000_4091, w_5000_4092, w_5000_4093, w_5000_4094, w_5000_4095, w_5000_4096, w_5000_4097, w_5000_4098, w_5000_4099, w_5000_4100, w_5000_4101, w_5000_4102, w_5000_4103, w_5000_4104, w_5000_4105, w_5000_4106, w_5000_4107, w_5000_4108, w_5000_4109, w_5000_4110, w_5000_4111, w_5000_4112, w_5000_4113, w_5000_4114, w_5000_4115, w_5000_4116, w_5000_4117, w_5000_4118, w_5000_4119, w_5000_4120, w_5000_4121, w_5000_4122, w_5000_4123, w_5000_4124, w_5000_4125, w_5000_4126, w_5000_4127, w_5000_4128, w_5000_4129, w_5000_4130, w_5000_4131, w_5000_4132, w_5000_4133, w_5000_4134, w_5000_4135, w_5000_4136, w_5000_4137, w_5000_4138, w_5000_4139, w_5000_4140, w_5000_4141, w_5000_4142, w_5000_4143, w_5000_4144, w_5000_4145, w_5000_4146, w_5000_4147, w_5000_4148, w_5000_4149, w_5000_4150, w_5000_4151, w_5000_4152, w_5000_4153, w_5000_4154, w_5000_4155, w_5000_4156, w_5000_4157, w_5000_4158, w_5000_4159, w_5000_4160, w_5000_4161, w_5000_4162, w_5000_4163, w_5000_4164, w_5000_4165, w_5000_4166, w_5000_4167, w_5000_4168, w_5000_4169, w_5000_4170, w_5000_4171, w_5000_4172, w_5000_4173, w_5000_4174, w_5000_4175, w_5000_4176, w_5000_4177, w_5000_4178, w_5000_4179, w_5000_4180, w_5000_4181, w_5000_4182, w_5000_4183, w_5000_4184, w_5000_4185, w_5000_4186, w_5000_4187, w_5000_4188, w_5000_4189, w_5000_4190, w_5000_4191, w_5000_4192, w_5000_4193, w_5000_4194, w_5000_4195, w_5000_4196, w_5000_4197, w_5000_4198, w_5000_4199, w_5000_4200, w_5000_4201, w_5000_4202, w_5000_4203, w_5000_4204, w_5000_4205, w_5000_4206, w_5000_4207, w_5000_4208, w_5000_4209, w_5000_4210, w_5000_4211, w_5000_4212, w_5000_4213, w_5000_4214, w_5000_4215, w_5000_4216, w_5000_4217, w_5000_4218, w_5000_4219, w_5000_4220, w_5000_4221, w_5000_4222, w_5000_4223, w_5000_4224, w_5000_4225, w_5000_4226, w_5000_4227, w_5000_4228, w_5000_4229, w_5000_4230, w_5000_4231, w_5000_4232, w_5000_4233, w_5000_4234, w_5000_4235, w_5000_4236, w_5000_4237, w_5000_4238, w_5000_4239, w_5000_4240, w_5000_4241, w_5000_4242, w_5000_4243, w_5000_4244, w_5000_4245 );
  inout w_000_000, w_000_001, w_000_002, w_000_003, w_000_004, w_000_005, w_000_006, w_000_007, w_000_008, w_000_009, w_000_010, w_000_011, w_000_012, w_000_013, w_000_014, w_000_015, w_000_016, w_000_017, w_000_018, w_000_019, w_000_020, w_000_021, w_000_022, w_000_023, w_000_024, w_000_025, w_000_026, w_000_027, w_000_028, w_000_029, w_000_030, w_000_031, w_000_032, w_000_033, w_000_034, w_000_035, w_000_036, w_000_037, w_000_038, w_000_039, w_000_040, w_000_041, w_000_042, w_000_043, w_000_044, w_000_045, w_000_046, w_000_047, w_000_048, w_000_049, w_000_050, w_000_051, w_000_052, w_000_053, w_000_054, w_000_055, w_000_056, w_000_057, w_000_058, w_000_059, w_000_060, w_000_061, w_000_062, w_000_063, w_000_064, w_000_065, w_000_066, w_000_067, w_000_068, w_000_069, w_000_070, w_000_071, w_000_072, w_000_073, w_000_074, w_000_075, w_000_076, w_000_077, w_000_078, w_000_079, w_000_080, w_000_081, w_000_082, w_000_083, w_000_084, w_000_085, w_000_086, w_000_087, w_000_088, w_000_089, w_000_090, w_000_091, w_000_092, w_000_093, w_000_094, w_000_095, w_000_096, w_000_097, w_000_098, w_000_099, w_000_100, w_000_101, w_000_102, w_000_103, w_000_104, w_000_105, w_000_106, w_000_107, w_000_108, w_000_109, w_000_110, w_000_111, w_000_112, w_000_113, w_000_114, w_000_115, w_000_116, w_000_117, w_000_118, w_000_119, w_000_120, w_000_121, w_000_122, w_000_123, w_000_124, w_000_125, w_000_126, w_000_127, w_000_128, w_000_129, w_000_130, w_000_131, w_000_132, w_000_133, w_000_134, w_000_135, w_000_136, w_000_137, w_000_138, w_000_139, w_000_140, w_000_141, w_000_142, w_000_143, w_000_144, w_000_145, w_000_146, w_000_147, w_000_148, w_000_149, w_000_150, w_000_151, w_000_152, w_000_153, w_000_154, w_000_155, w_000_156, w_000_157, w_000_158, w_000_159, w_000_160, w_000_161, w_000_162, w_000_163, w_000_164, w_000_165, w_000_166, w_000_167, w_000_168, w_000_169, w_000_170, w_000_171, w_000_172, w_000_173, w_000_174, w_000_175, w_000_176, w_000_177, w_000_178, w_000_179, w_000_180, w_000_181, w_000_182, w_000_183, w_000_184, w_000_185, w_000_186, w_000_187, w_000_188, w_000_189, w_000_190, w_000_191, w_000_192, w_000_193, w_000_194, w_000_195, w_000_196, w_000_197, w_000_198, w_000_199, w_000_200, w_000_201, w_000_202, w_000_203, w_000_204, w_000_205, w_000_206, w_000_207, w_000_208, w_000_209, w_000_210, w_000_211, w_000_212, w_000_213, w_000_214, w_000_215, w_000_216, w_000_217, w_000_218, w_000_219, w_000_220, w_000_221, w_000_222, w_000_223, w_000_224, w_000_225, w_000_226, w_000_227, w_000_228, w_000_229, w_000_230, w_000_231, w_000_232, w_000_233, w_000_234, w_000_235, w_000_236, w_000_237, w_000_238, w_000_239, w_000_240, w_000_241, w_000_242, w_000_243, w_000_244, w_000_245, w_000_246, w_000_247, w_000_248, w_000_249, w_000_250, w_000_251, w_000_252, w_000_253, w_000_254, w_000_255, w_000_256, w_000_257, w_000_258, w_000_259, w_000_260, w_000_261, w_000_262, w_000_263, w_000_264, w_000_265, w_000_266, w_000_267, w_000_268, w_000_269, w_000_270, w_000_271, w_000_272, w_000_273, w_000_274, w_000_275, w_000_276, w_000_277, w_000_278, w_000_279, w_000_280, w_000_281, w_000_282, w_000_283, w_000_284, w_000_285, w_000_286, w_000_287, w_000_288, w_000_289, w_000_290, w_000_291, w_000_292, w_000_293, w_000_294, w_000_295, w_000_296, w_000_297, w_000_298, w_000_299, w_000_300, w_000_301, w_000_302, w_000_303, w_000_304, w_000_305, w_000_306, w_000_307, w_000_308, w_000_309, w_000_310, w_000_311, w_000_312, w_000_313, w_000_314, w_000_315, w_000_316, w_000_317, w_000_318, w_000_319, w_000_320, w_000_321, w_000_322, w_000_323, w_000_324, w_000_325, w_000_326, w_000_327, w_000_328, w_000_329, w_000_330, w_000_331, w_000_332, w_000_333, w_000_334, w_000_335, w_000_336, w_000_337, w_000_338, w_000_339, w_000_340, w_000_341, w_000_342, w_000_343, w_000_344, w_000_345, w_000_346, w_000_347, w_000_348, w_000_349, w_000_350, w_000_351, w_000_352, w_000_353, w_000_354, w_000_355, w_000_356, w_000_357, w_000_358, w_000_359, w_000_360, w_000_361, w_000_362, w_000_363, w_000_364, w_000_365, w_000_366, w_000_367, w_000_368, w_000_369, w_000_370, w_000_371, w_000_372, w_000_373, w_000_374, w_000_375, w_000_376, w_000_377, w_000_378, w_000_379, w_000_380, w_000_381, w_000_382, w_000_383, w_000_384, w_000_385, w_000_386, w_000_387, w_000_388, w_000_389, w_000_390, w_000_391, w_000_392, w_000_393, w_000_394, w_000_395, w_000_396, w_000_397, w_000_398, w_000_399, w_000_400, w_000_401, w_000_402, w_000_403, w_000_404, w_000_405, w_000_406, w_000_407, w_000_408, w_000_409, w_000_410, w_000_411, w_000_412, w_000_413, w_000_414, w_000_415, w_000_416, w_000_417, w_000_418, w_000_419, w_000_420, w_000_421, w_000_422, w_000_423, w_000_424, w_000_425, w_000_426, w_000_427, w_000_428, w_000_429, w_000_430, w_000_431, w_000_432, w_000_433, w_000_434, w_000_435, w_000_436, w_000_437, w_000_438, w_000_439, w_000_440, w_000_441, w_000_442, w_000_443, w_000_444, w_000_445, w_000_446, w_000_447, w_000_448, w_000_449, w_000_450, w_000_451, w_000_452, w_000_453, w_000_454, w_000_455, w_000_456, w_000_457, w_000_458, w_000_459, w_000_460, w_000_461, w_000_462, w_000_463, w_000_464, w_000_465, w_000_466, w_000_467, w_000_468, w_000_469, w_000_470, w_000_471, w_000_472, w_000_473, w_000_474, w_000_475, w_000_476, w_000_477, w_000_478, w_000_479, w_000_480, w_000_481, w_000_482, w_000_483, w_000_484, w_000_485, w_000_486, w_000_487, w_000_488, w_000_489, w_000_490, w_000_491, w_000_492, w_000_493, w_000_494, w_000_495, w_000_496, w_000_497, w_000_498, w_000_499, w_000_500, w_000_501, w_000_502, w_000_503, w_000_504, w_000_505, w_000_506, w_000_507, w_000_508, w_000_509, w_000_510, w_000_511, w_000_512, w_000_513, w_000_514, w_000_515, w_000_516, w_000_517, w_000_518, w_000_519, w_000_520, w_000_521, w_000_522, w_000_523, w_000_524, w_000_525, w_000_526, w_000_527, w_000_528, w_000_529, w_000_530, w_000_531, w_000_532, w_000_533, w_000_534, w_000_535, w_000_536, w_000_537, w_000_538, w_000_539, w_000_540, w_000_541, w_000_542, w_000_543, w_000_544, w_000_545, w_000_546, w_000_547, w_000_548, w_000_549, w_000_550, w_000_551, w_000_552, w_000_553, w_000_554, w_000_555, w_000_556, w_000_557, w_000_558, w_000_559, w_000_560, w_000_561, w_000_562, w_000_563, w_000_564, w_000_565, w_000_566, w_000_567, w_000_568, w_000_569, w_000_570, w_000_571, w_000_572, w_000_573, w_000_574, w_000_575, w_000_576, w_000_577, w_000_578, w_000_579, w_000_580, w_000_581, w_000_582, w_000_583, w_000_584, w_000_585, w_000_586, w_000_587, w_000_588, w_000_589, w_000_590, w_000_591, w_000_592, w_000_593, w_000_594, w_000_595, w_000_596, w_000_597, w_000_598, w_000_599, w_000_600, w_000_601, w_000_602, w_000_603, w_000_604, w_000_605, w_000_606, w_000_607, w_000_608, w_000_609, w_000_610, w_000_611, w_000_612, w_000_613, w_000_614, w_000_615, w_000_616, w_000_617, w_000_618, w_000_619, w_000_620, w_000_621, w_000_622, w_000_623, w_000_624, w_000_625, w_000_626, w_000_627, w_000_628, w_000_629, w_000_630, w_000_631, w_000_632, w_000_633, w_000_634, w_000_635, w_000_636, w_000_637, w_000_638, w_000_639, w_000_640, w_000_641, w_000_642, w_000_643, w_000_644, w_000_645, w_000_646, w_000_647, w_000_648, w_000_649, w_000_650, w_000_651, w_000_652, w_000_653, w_000_654, w_000_655, w_000_656, w_000_657, w_000_658, w_000_659, w_000_660, w_000_661, w_000_662, w_000_663, w_000_664, w_000_665, w_000_666, w_000_667, w_000_668, w_000_669, w_000_670, w_000_671, w_000_672, w_000_673, w_000_674, w_000_675, w_000_676, w_000_677, w_000_678, w_000_679, w_000_680, w_000_681, w_000_682, w_000_683, w_000_684, w_000_685, w_000_686, w_000_687, w_000_688, w_000_689, w_000_690, w_000_691, w_000_692, w_000_693, w_000_694, w_000_695, w_000_696, w_000_697, w_000_698, w_000_699, w_000_700, w_000_701, w_000_702, w_000_703, w_000_704, w_000_705, w_000_706, w_000_707, w_000_708, w_000_709, w_000_710, w_000_711, w_000_712, w_000_713, w_000_714, w_000_715, w_000_716, w_000_717, w_000_718, w_000_719, w_000_720, w_000_721, w_000_722, w_000_723, w_000_724, w_000_725, w_000_726, w_000_727, w_000_728, w_000_729, w_000_730, w_000_731, w_000_732, w_000_733, w_000_734, w_000_735, w_000_736, w_000_737, w_000_738, w_000_739, w_000_740, w_000_741, w_000_742, w_000_743, w_000_744, w_000_745, w_000_746, w_000_747, w_000_748, w_000_749, w_000_750, w_000_751, w_000_752, w_000_753, w_000_754, w_000_755, w_000_756, w_000_757, w_000_758, w_000_759, w_000_760, w_000_761, w_000_762, w_000_763, w_000_764, w_000_765, w_000_766, w_000_767, w_000_768, w_000_769, w_000_770, w_000_771, w_000_772, w_000_773, w_000_774, w_000_775, w_000_776, w_000_777, w_000_778, w_000_779, w_000_780, w_000_781, w_000_782, w_000_783, w_000_784, w_000_785, w_000_786, w_000_787, w_000_788, w_000_789, w_000_790, w_000_791, w_000_792, w_000_793, w_000_794, w_000_795, w_000_796, w_000_797, w_000_798, w_000_799, w_000_800, w_000_801, w_000_802, w_000_803, w_000_804, w_000_805, w_000_806, w_000_807, w_000_808, w_000_809, w_000_810, w_000_811, w_000_812, w_000_813, w_000_814, w_000_815, w_000_816, w_000_817, w_000_818, w_000_819, w_000_820, w_000_821, w_000_822, w_000_823, w_000_824, w_000_825, w_000_826, w_000_827, w_000_828, w_000_829, w_000_830, w_000_831, w_000_832, w_000_833, w_000_834, w_000_835, w_000_836, w_000_837, w_000_838, w_000_839, w_000_840, w_000_841, w_000_842, w_000_843, w_000_844, w_000_845, w_000_846, w_000_847, w_000_848, w_000_849, w_000_850, w_000_851, w_000_852, w_000_853, w_000_854, w_000_855, w_000_856, w_000_857, w_000_858, w_000_859, w_000_860, w_000_861, w_000_862, w_000_863, w_000_864, w_000_865, w_000_866, w_000_867, w_000_868, w_000_869, w_000_870, w_000_871, w_000_872, w_000_873, w_000_874, w_000_875, w_000_876, w_000_877, w_000_878, w_000_879, w_000_880, w_000_881, w_000_882, w_000_883, w_000_884, w_000_885, w_000_886, w_000_887, w_000_888, w_000_889, w_000_890, w_000_891, w_000_892, w_000_893, w_000_894, w_000_895, w_000_896, w_000_897, w_000_898, w_000_899, w_000_900, w_000_901, w_000_902, w_000_903, w_000_904, w_000_905, w_000_906, w_000_907, w_000_908, w_000_909, w_000_910, w_000_911, w_000_912, w_000_913, w_000_914, w_000_915, w_000_916, w_000_917, w_000_918, w_000_919, w_000_920, w_000_921, w_000_922, w_000_923, w_000_924, w_000_925, w_000_926, w_000_927, w_000_928, w_000_929, w_000_930, w_000_931, w_000_932, w_000_933, w_000_934, w_000_935, w_000_936, w_000_937, w_000_938, w_000_939, w_000_940, w_000_941, w_000_942, w_000_943, w_000_944, w_000_945, w_000_946, w_000_947, w_000_948, w_000_949, w_000_950, w_000_951, w_000_952, w_000_953, w_000_954, w_000_955, w_000_956, w_000_957, w_000_958, w_000_959, w_000_960, w_000_961, w_000_962, w_000_963, w_000_964, w_000_965, w_000_966, w_000_967, w_000_968, w_000_969, w_000_970, w_000_971, w_000_972, w_000_973, w_000_974, w_000_975, w_000_976, w_000_977, w_000_978, w_000_979, w_000_980, w_000_981, w_000_982, w_000_983, w_000_984, w_000_985, w_000_986, w_000_987, w_000_988, w_000_989, w_000_990, w_000_991, w_000_992, w_000_993, w_000_994, w_000_995, w_000_996, w_000_997, w_000_998, w_000_999, w_000_1000, w_000_1001, w_000_1002, w_000_1003, w_000_1004, w_000_1005, w_000_1006, w_000_1007, w_000_1008, w_000_1009, w_000_1010, w_000_1011, w_000_1012, w_000_1013, w_000_1014, w_000_1015, w_000_1016, w_000_1017, w_000_1018, w_000_1019, w_000_1020, w_000_1021, w_000_1022, w_000_1023, w_000_1024, w_000_1025, w_000_1026, w_000_1027, w_000_1028, w_000_1029, w_000_1030, w_000_1031, w_000_1032, w_000_1033, w_000_1034, w_000_1035, w_000_1036, w_000_1037, w_000_1038, w_000_1039, w_000_1040, w_000_1041, w_000_1042, w_000_1043, w_000_1044, w_000_1045, w_000_1046, w_000_1047, w_000_1048, w_000_1049, w_000_1050, w_000_1051, w_000_1052, w_000_1053, w_000_1054, w_000_1055, w_000_1056, w_000_1057, w_000_1058, w_000_1059, w_000_1060, w_000_1061, w_000_1062, w_000_1063, w_000_1064, w_000_1065, w_000_1066, w_000_1067, w_000_1068, w_000_1069, w_000_1070, w_000_1071, w_000_1072, w_000_1073, w_000_1074, w_000_1075, w_000_1076, w_000_1077, w_000_1078, w_000_1079, w_000_1080, w_000_1081, w_000_1082, w_000_1083, w_000_1084, w_000_1085, w_000_1086, w_000_1087, w_000_1088, w_000_1089, w_000_1090, w_000_1091, w_000_1092, w_000_1093, w_000_1094, w_000_1095, w_000_1096, w_000_1097, w_000_1098, w_000_1099, w_000_1100, w_000_1101, w_000_1102, w_000_1103, w_000_1104, w_000_1105, w_000_1106, w_000_1107, w_000_1108, w_000_1109, w_000_1110, w_000_1111, w_000_1112, w_000_1113, w_000_1114, w_000_1115, w_000_1116, w_000_1117, w_000_1118, w_000_1119, w_000_1120, w_000_1121, w_000_1122, w_000_1123, w_000_1124, w_000_1125, w_000_1126, w_000_1127, w_000_1128, w_000_1129, w_000_1130, w_000_1131, w_000_1132, w_000_1133, w_000_1134, w_000_1135, w_000_1136, w_000_1137, w_000_1138, w_000_1139, w_000_1140, w_000_1141, w_000_1142, w_000_1143, w_000_1144, w_000_1145, w_000_1146, w_000_1147, w_000_1148, w_000_1149, w_000_1150, w_000_1151, w_000_1152, w_000_1153, w_000_1154, w_000_1155, w_000_1156, w_000_1157, w_000_1158, w_000_1159, w_000_1160, w_000_1161, w_000_1162, w_000_1163, w_000_1164, w_000_1165, w_000_1166, w_000_1167, w_000_1168, w_000_1169, w_000_1170, w_000_1171, w_000_1172, w_000_1173, w_000_1174, w_000_1175, w_000_1176, w_000_1177, w_000_1178, w_000_1179, w_000_1180, w_000_1181, w_000_1182, w_000_1183, w_000_1184, w_000_1185, w_000_1186, w_000_1187, w_000_1188, w_000_1189, w_000_1190, w_000_1191, w_000_1192, w_000_1193, w_000_1194, w_000_1195, w_000_1196, w_000_1197, w_000_1198, w_000_1199, w_000_1200, w_000_1201, w_000_1202, w_000_1203, w_000_1204, w_000_1205, w_000_1206, w_000_1207, w_000_1208, w_000_1209, w_000_1210, w_000_1211, w_000_1212, w_000_1213, w_000_1214, w_000_1215, w_000_1216, w_000_1217, w_000_1218, w_000_1219, w_000_1220, w_000_1221, w_000_1222, w_000_1223, w_000_1224, w_000_1225, w_000_1226, w_000_1227, w_000_1228, w_000_1229, w_000_1230, w_000_1231, w_000_1232, w_000_1233, w_000_1234, w_000_1235, w_000_1236, w_000_1237, w_000_1238, w_000_1239, w_000_1240, w_000_1241, w_000_1242, w_000_1243, w_000_1244, w_000_1245, w_000_1246, w_000_1247, w_000_1248, w_000_1249, w_000_1250, w_000_1251, w_000_1252, w_000_1253, w_000_1254, w_000_1255, w_000_1256, w_000_1257, w_000_1258, w_000_1259, w_000_1260, w_000_1261, w_000_1262, w_000_1263, w_000_1264, w_000_1265, w_000_1266, w_000_1267, w_000_1268, w_000_1269, w_000_1270, w_000_1271, w_000_1272, w_000_1273, w_000_1274, w_000_1275, w_000_1276, w_000_1277, w_000_1278, w_000_1279, w_000_1280, w_000_1281, w_000_1282, w_000_1283, w_000_1284, w_000_1285, w_000_1286, w_000_1287, w_000_1288, w_000_1289, w_000_1290, w_000_1291, w_000_1292, w_000_1293, w_000_1294, w_000_1295, w_000_1296, w_000_1297, w_000_1298, w_000_1299, w_000_1300, w_000_1301, w_000_1302, w_000_1303, w_000_1304, w_000_1305, w_000_1306, w_000_1307, w_000_1308, w_000_1309, w_000_1310, w_000_1311, w_000_1312, w_000_1313, w_000_1314, w_000_1315, w_000_1316, w_000_1317, w_000_1318, w_000_1319, w_000_1320, w_000_1321, w_000_1322, w_000_1323, w_000_1324, w_000_1325, w_000_1326, w_000_1327, w_000_1328, w_000_1329, w_000_1330, w_000_1331, w_000_1332, w_000_1333, w_000_1334, w_000_1335, w_000_1336, w_000_1337, w_000_1338, w_000_1339, w_000_1340, w_000_1341, w_000_1342, w_000_1343, w_000_1344, w_000_1345, w_000_1346, w_000_1347, w_000_1348, w_000_1349, w_000_1350, w_000_1351, w_000_1352, w_000_1353, w_000_1354, w_000_1355, w_000_1356, w_000_1357, w_000_1358, w_000_1359, w_000_1360, w_000_1361, w_000_1362, w_000_1363, w_000_1364, w_000_1365, w_000_1366, w_000_1367, w_000_1368, w_000_1369, w_000_1370, w_000_1371, w_000_1372, w_000_1373, w_000_1374, w_000_1375, w_000_1376, w_000_1377, w_000_1378, w_000_1379, w_000_1380, w_000_1381, w_000_1382, w_000_1383, w_000_1384, w_000_1385, w_000_1386, w_000_1387, w_000_1388, w_000_1389, w_000_1390, w_000_1391, w_000_1392, w_000_1393, w_000_1394, w_000_1395, w_000_1396, w_000_1397, w_000_1398, w_000_1399, w_000_1400, w_000_1401, w_000_1402, w_000_1403, w_000_1404, w_000_1405, w_000_1406, w_000_1407, w_000_1408, w_000_1409, w_000_1410, w_000_1411, w_000_1412, w_000_1413, w_000_1414, w_000_1415, w_000_1416, w_000_1417, w_000_1418, w_000_1419, w_000_1420, w_000_1421, w_000_1422, w_000_1423, w_000_1424, w_000_1425, w_000_1426, w_000_1427, w_000_1428, w_000_1429, w_000_1430, w_000_1431, w_000_1432, w_000_1433, w_000_1434, w_000_1435, w_000_1436, w_000_1437, w_000_1438, w_000_1439, w_000_1440, w_000_1441, w_000_1442, w_000_1443, w_000_1444, w_000_1445, w_000_1446, w_000_1447, w_000_1448, w_000_1449, w_000_1450, w_000_1451, w_000_1452, w_000_1453, w_000_1454, w_000_1455, w_000_1456, w_000_1457, w_000_1458, w_000_1459, w_000_1460, w_000_1461, w_000_1462, w_000_1463, w_000_1464, w_000_1465, w_000_1466, w_000_1467, w_000_1468, w_000_1469, w_000_1470, w_000_1471, w_000_1472, w_000_1473, w_000_1474, w_000_1475, w_000_1476, w_000_1477, w_000_1478, w_000_1479, w_000_1480, w_000_1481, w_000_1482, w_000_1483, w_000_1484, w_000_1485, w_000_1486, w_000_1487, w_000_1488, w_000_1489, w_000_1490, w_000_1491, w_000_1492, w_000_1493, w_000_1494, w_000_1495, w_000_1496, w_000_1497, w_000_1498, w_000_1499, w_000_1500, w_000_1501, w_000_1502, w_000_1503, w_000_1504, w_000_1505, w_000_1506, w_000_1507, w_000_1508, w_000_1509, w_000_1510, w_000_1511, w_000_1512, w_000_1513, w_000_1514, w_000_1515, w_000_1516, w_000_1517, w_000_1518, w_000_1519, w_000_1520, w_000_1521, w_000_1522, w_000_1523, w_000_1524, w_000_1525, w_000_1526, w_000_1527, w_000_1528, w_000_1529, w_000_1530, w_000_1531, w_000_1532, w_000_1533, w_000_1534, w_000_1535, w_000_1536, w_000_1537, w_000_1538, w_000_1539, w_000_1540, w_000_1541, w_000_1542, w_000_1543, w_000_1544, w_000_1545, w_000_1546, w_000_1547, w_000_1548, w_000_1549, w_000_1550, w_000_1551, w_000_1552, w_000_1553, w_000_1554, w_000_1555, w_000_1556, w_000_1557, w_000_1558, w_000_1559, w_000_1560, w_000_1561, w_000_1562, w_000_1563, w_000_1564, w_000_1565, w_000_1566, w_000_1567, w_000_1568, w_000_1569, w_000_1570, w_000_1571, w_000_1572, w_000_1573, w_000_1574, w_000_1575, w_000_1576, w_000_1577, w_000_1578, w_000_1579, w_000_1580, w_000_1581, w_000_1582, w_000_1583, w_000_1584, w_000_1585, w_000_1586, w_000_1587, w_000_1588, w_000_1589, w_000_1590, w_000_1591, w_000_1592, w_000_1593, w_000_1594, w_000_1595, w_000_1596, w_000_1597, w_000_1598, w_000_1599, w_000_1600, w_000_1601, w_000_1602, w_000_1603, w_000_1604, w_000_1605, w_000_1606, w_000_1607, w_000_1608, w_000_1609, w_000_1610, w_000_1611, w_000_1612, w_000_1613, w_000_1614, w_000_1615, w_000_1616, w_000_1617, w_000_1618, w_000_1619, w_000_1620, w_000_1621, w_000_1622, w_000_1623, w_000_1624, w_000_1625, w_000_1626, w_000_1627, w_000_1628, w_000_1629, w_000_1630, w_000_1631, w_000_1632, w_000_1633, w_000_1634, w_000_1635, w_000_1636, w_000_1637, w_000_1638, w_000_1639, w_000_1640, w_000_1641, w_000_1642, w_000_1643, w_000_1644, w_000_1645, w_000_1646, w_000_1647, w_000_1648, w_000_1649, w_000_1650, w_000_1651, w_000_1652, w_000_1653, w_000_1654, w_000_1655, w_000_1656, w_000_1657, w_000_1658, w_000_1659, w_000_1660, w_000_1661, w_000_1662, w_000_1663, w_000_1664, w_000_1665, w_000_1666, w_000_1667, w_000_1668, w_000_1669, w_000_1670, w_000_1671, w_000_1672, w_000_1673, w_000_1674, w_000_1675, w_000_1676, w_000_1677, w_000_1678, w_000_1679, w_000_1680, w_000_1681, w_000_1682, w_000_1683, w_000_1684, w_000_1685, w_000_1686, w_000_1687, w_000_1688, w_000_1689, w_000_1690, w_000_1691, w_000_1692, w_000_1693, w_000_1694, w_000_1695, w_000_1696, w_000_1697, w_000_1698, w_000_1699, w_000_1700, w_000_1701, w_000_1702, w_000_1703, w_000_1704, w_000_1705, w_000_1706, w_000_1707, w_000_1708, w_000_1709, w_000_1710, w_000_1711, w_000_1712, w_000_1713, w_000_1714, w_000_1715, w_000_1716, w_000_1717, w_000_1718, w_000_1719, w_000_1720, w_000_1721, w_000_1722, w_000_1723, w_000_1724, w_000_1725, w_000_1726, w_000_1727, w_000_1728, w_000_1729, w_000_1730, w_000_1731, w_000_1732, w_000_1733, w_000_1734, w_000_1735, w_000_1736, w_000_1737, w_000_1738, w_000_1739, w_000_1740, w_000_1741, w_000_1742, w_000_1743, w_000_1744, w_000_1745, w_000_1746, w_000_1747, w_000_1748, w_000_1749, w_000_1750, w_000_1751, w_000_1752, w_000_1753, w_000_1754, w_000_1755, w_000_1756, w_000_1757, w_000_1758, w_000_1759, w_000_1760, w_000_1761, w_000_1762, w_000_1763, w_000_1764, w_000_1765, w_000_1766, w_000_1767, w_000_1768, w_000_1769, w_000_1770, w_000_1771, w_000_1772, w_000_1773, w_000_1774, w_000_1775, w_000_1776, w_000_1777, w_000_1778, w_000_1779, w_000_1780, w_000_1781, w_000_1782, w_000_1783, w_000_1784, w_000_1785, w_000_1786, w_000_1787, w_000_1788, w_000_1789, w_000_1790, w_000_1791, w_000_1792, w_000_1793, w_000_1794, w_000_1795, w_000_1796, w_000_1797, w_000_1798, w_000_1799, w_000_1800, w_000_1801, w_000_1802, w_000_1803, w_000_1804, w_000_1805, w_000_1806, w_000_1807, w_000_1808, w_000_1809, w_000_1810, w_000_1811, w_000_1812, w_000_1813, w_000_1814, w_000_1815, w_000_1816, w_000_1817, w_000_1818, w_000_1819, w_000_1820, w_000_1821, w_000_1822, w_000_1823, w_000_1824, w_000_1825, w_000_1826, w_000_1827, w_000_1828, w_000_1829, w_000_1830, w_000_1831, w_000_1832, w_000_1833, w_000_1834, w_000_1835, w_000_1836, w_000_1837, w_000_1838, w_000_1839, w_000_1840, w_000_1841, w_000_1842, w_000_1843, w_000_1844, w_000_1845, w_000_1846, w_000_1847, w_000_1848, w_000_1849, w_000_1850, w_000_1851, w_000_1852, w_000_1853, w_000_1854, w_000_1855, w_000_1856, w_000_1857, w_000_1858, w_000_1859, w_000_1860, w_000_1861, w_000_1862, w_000_1863, w_000_1864, w_000_1865, w_000_1866, w_000_1867, w_000_1868, w_000_1869, w_000_1870, w_000_1871, w_000_1872, w_000_1873, w_000_1874, w_000_1875, w_000_1876, w_000_1877, w_000_1878, w_000_1879, w_000_1880, w_000_1881, w_000_1882, w_000_1883, w_000_1884, w_000_1885, w_000_1886, w_000_1887, w_000_1888, w_000_1889, w_000_1890, w_000_1891, w_000_1892, w_000_1893, w_000_1894, w_000_1895, w_000_1896, w_000_1897, w_000_1898, w_000_1899, w_000_1900, w_000_1901, w_000_1902, w_000_1903, w_000_1904, w_000_1905, w_000_1906, w_000_1907, w_000_1908, w_000_1909, w_000_1910, w_000_1911, w_000_1912, w_000_1913, w_000_1914, w_000_1915, w_000_1916, w_000_1917, w_000_1918, w_000_1919, w_000_1920, w_000_1921, w_000_1922, w_000_1923, w_000_1924, w_000_1925, w_000_1926, w_000_1927, w_000_1928, w_000_1929, w_000_1930, w_000_1931, w_000_1932, w_000_1933, w_000_1934, w_000_1935, w_000_1936, w_000_1937, w_000_1938, w_000_1939, w_000_1940, w_000_1941, w_000_1942, w_000_1943, w_000_1944, w_000_1945, w_000_1946, w_000_1947, w_000_1948, w_000_1949, w_000_1950, w_000_1951, w_000_1952, w_000_1953, w_000_1954, w_000_1955, w_000_1956, w_000_1957, w_000_1958, w_000_1959, w_000_1960, w_000_1961, w_000_1962, w_000_1963, w_000_1964, w_000_1965, w_000_1966, w_000_1967, w_000_1968, w_000_1969, w_000_1970, w_000_1971, w_000_1972, w_000_1973, w_000_1974, w_000_1975, w_000_1976, w_000_1977, w_000_1978, w_000_1979, w_000_1980, w_000_1981, w_000_1982, w_000_1983, w_000_1984, w_000_1985, w_000_1986, w_000_1987, w_000_1988, w_000_1989, w_000_1990, w_000_1991, w_000_1992, w_000_1993, w_000_1994, w_000_1995, w_000_1996, w_000_1997, w_000_1998, w_000_1999, w_000_2000, w_000_2001, w_000_2002, w_000_2003, w_000_2004, w_000_2005, w_000_2006, w_000_2007, w_000_2008, w_000_2009, w_000_2010, w_000_2011, w_000_2012, w_000_2013, w_000_2014, w_000_2015, w_000_2016, w_000_2017, w_000_2018, w_000_2019, w_000_2020, w_000_2021, w_000_2022, w_000_2023, w_000_2024, w_000_2025, w_000_2026, w_000_2027, w_000_2028, w_000_2029, w_000_2030, w_000_2031, w_000_2032, w_000_2033, w_000_2034, w_000_2035, w_000_2036, w_000_2037, w_000_2038, w_000_2039, w_000_2040, w_000_2041, w_000_2042, w_000_2043, w_000_2044, w_000_2045, w_000_2046, w_000_2047, w_000_2048, w_000_2049, w_000_2050, w_000_2051, w_000_2052, w_000_2053, w_000_2054, w_000_2055, w_000_2056, w_000_2057, w_000_2058, w_000_2059, w_000_2060, w_000_2061, w_000_2062, w_000_2063, w_000_2064, w_000_2065, w_000_2066, w_000_2067, w_000_2068, w_000_2069, w_000_2070, w_000_2071, w_000_2072, w_000_2073, w_000_2074, w_000_2075, w_000_2076, w_000_2077, w_000_2078, w_000_2079, w_000_2080, w_000_2081, w_000_2082, w_000_2083, w_000_2084, w_000_2085, w_000_2086, w_000_2087, w_000_2088, w_000_2089, w_000_2090, w_000_2091, w_000_2092, w_000_2093, w_000_2094, w_000_2095, w_000_2096, w_000_2097, w_000_2098, w_000_2099, w_000_2100, w_000_2101, w_000_2102, w_000_2103, w_000_2104, w_000_2105, w_000_2106, w_000_2107, w_000_2108, w_000_2109, w_000_2110, w_000_2111, w_000_2112, w_000_2113, w_000_2114, w_000_2115, w_000_2116, w_000_2117, w_000_2118, w_000_2119, w_000_2120, w_000_2121, w_000_2122, w_000_2123, w_000_2124, w_000_2125, w_000_2126, w_000_2127, w_000_2128, w_000_2129, w_000_2130, w_000_2131, w_000_2132, w_000_2133, w_000_2134, w_000_2135, w_000_2136, w_000_2137, w_000_2138, w_000_2139, w_000_2140, w_000_2141, w_000_2142, w_000_2143, w_000_2144, w_000_2145, w_000_2146, w_000_2147, w_000_2148, w_000_2149, w_000_2150, w_000_2151, w_000_2152, w_000_2153, w_000_2154, w_000_2155, w_000_2156, w_000_2157, w_000_2158, w_000_2159, w_000_2160, w_000_2161, w_000_2162, w_000_2163, w_000_2164, w_000_2165, w_000_2166, w_000_2167, w_000_2168, w_000_2169, w_000_2170, w_000_2171, w_000_2172, w_000_2173, w_000_2174, w_000_2175, w_000_2176, w_000_2177, w_000_2178, w_000_2179, w_000_2180, w_000_2181, w_000_2182, w_000_2183, w_000_2184, w_000_2185, w_000_2186, w_000_2187, w_000_2188, w_000_2189, w_000_2190, w_000_2191, w_000_2192, w_000_2193, w_000_2194, w_000_2195, w_000_2196, w_000_2197, w_000_2198, w_000_2199, w_000_2200, w_000_2201, w_000_2202, w_000_2203, w_000_2204, w_000_2205, w_000_2206, w_000_2207, w_000_2208, w_000_2209, w_000_2210, w_000_2211, w_000_2212, w_000_2213, w_000_2214, w_000_2215, w_000_2216, w_000_2217, w_000_2218, w_000_2219, w_000_2220, w_000_2221, w_000_2222, w_000_2223, w_000_2224, w_000_2225, w_000_2226, w_000_2227, w_000_2228, w_000_2229, w_000_2230, w_000_2231, w_000_2232, w_000_2233, w_000_2234, w_000_2235, w_000_2236, w_000_2237, w_000_2238, w_000_2239, w_000_2240, w_000_2241, w_000_2242, w_000_2243, w_000_2244, w_000_2245, w_000_2246, w_000_2247, w_000_2248, w_000_2249, w_000_2250, w_000_2251, w_000_2252, w_000_2253, w_000_2254, w_000_2255, w_000_2256, w_000_2257, w_000_2258, w_000_2259, w_000_2260, w_000_2261, w_000_2262, w_000_2263, w_000_2264, w_000_2265, w_000_2266, w_000_2267, w_000_2268, w_000_2269, w_000_2270, w_000_2271, w_000_2272, w_000_2273, w_000_2274, w_000_2275, w_000_2276, w_000_2277, w_000_2278, w_000_2279, w_000_2280, w_000_2281, w_000_2282, w_000_2283, w_000_2284, w_000_2285, w_000_2286, w_000_2287, w_000_2288, w_000_2289, w_000_2290, w_000_2291, w_000_2292, w_000_2293, w_000_2294, w_000_2295, w_000_2296, w_000_2297, w_000_2298, w_000_2299, w_000_2300, w_000_2301, w_000_2302, w_000_2303, w_000_2304, w_000_2305, w_000_2306, w_000_2307, w_000_2308, w_000_2309, w_000_2310, w_000_2311, w_000_2312, w_000_2313, w_000_2314, w_000_2315, w_000_2316, w_000_2317, w_000_2318, w_000_2319, w_000_2320, w_000_2321, w_000_2322, w_000_2323, w_000_2324, w_000_2325, w_000_2326, w_000_2327, w_000_2328, w_000_2329, w_000_2330, w_000_2331, w_000_2332, w_000_2333, w_000_2334, w_000_2335, w_000_2336, w_000_2337, w_000_2338, w_000_2339, w_000_2340, w_000_2341, w_000_2342, w_000_2343, w_000_2344, w_000_2345, w_000_2346, w_000_2347, w_000_2348, w_000_2349, w_000_2350, w_000_2351, w_000_2352, w_000_2353, w_000_2354, w_000_2355, w_000_2356, w_000_2357, w_000_2358, w_000_2359, w_000_2360, w_000_2361, w_000_2362, w_000_2363, w_000_2364, w_000_2365, w_000_2366, w_000_2367, w_000_2368, w_000_2369, w_000_2370, w_000_2371, w_000_2372, w_000_2373, w_000_2374, w_000_2375, w_000_2376, w_000_2377, w_000_2378, w_000_2379, w_000_2380, w_000_2381, w_000_2382, w_000_2383, w_000_2384, w_000_2385, w_000_2386, w_000_2387, w_000_2388, w_000_2389, w_000_2390, w_000_2391, w_000_2392, w_000_2393, w_000_2394, w_000_2395, w_000_2396, w_000_2397, w_000_2398, w_000_2399, w_000_2400, w_000_2401, w_000_2402, w_000_2403, w_000_2404, w_000_2405, w_000_2406, w_000_2407, w_000_2408, w_000_2409, w_000_2410, w_000_2411, w_000_2412, w_000_2413, w_000_2414, w_000_2415, w_000_2416, w_000_2417, w_000_2418, w_000_2419, w_000_2420, w_000_2421, w_000_2422, w_000_2423, w_000_2424, w_000_2425, w_000_2426, w_000_2427, w_000_2428, w_000_2429, w_000_2430, w_000_2431, w_000_2432, w_000_2433, w_000_2434, w_000_2435, w_000_2436, w_000_2437, w_000_2438, w_000_2439, w_000_2440, w_000_2441, w_000_2442, w_000_2443, w_000_2444, w_000_2445, w_000_2446, w_000_2447, w_000_2448, w_000_2449, w_000_2450, w_000_2451, w_000_2452, w_000_2453, w_000_2454, w_000_2455, w_000_2456, w_000_2457, w_000_2458, w_000_2459, w_000_2460, w_000_2461, w_000_2462, w_000_2463, w_000_2464, w_000_2465, w_000_2466, w_000_2467, w_000_2468, w_000_2469, w_000_2470, w_000_2471, w_000_2472, w_000_2473, w_000_2474, w_000_2475, w_000_2476, w_000_2477, w_000_2478, w_000_2479, w_000_2480, w_000_2481, w_000_2482, w_000_2483, w_000_2484, w_000_2485, w_000_2486, w_000_2487, w_000_2488, w_000_2489, w_000_2490, w_000_2491, w_000_2492, w_000_2493, w_000_2494, w_000_2495, w_000_2496, w_000_2497, w_000_2498, w_000_2499, w_000_2500, w_000_2501, w_000_2502, w_000_2503, w_000_2504, w_000_2505, w_000_2506, w_000_2507, w_000_2508, w_000_2509, w_000_2510, w_000_2511, w_000_2512, w_000_2513, w_000_2514, w_000_2515, w_000_2516, w_000_2517, w_000_2518, w_000_2519, w_000_2520, w_000_2521, w_000_2522, w_000_2523, w_000_2524, w_000_2525, w_000_2526, w_000_2527, w_000_2528, w_000_2529, w_000_2530, w_000_2531, w_000_2532, w_000_2533, w_000_2534, w_000_2535, w_000_2536, w_000_2537, w_000_2538, w_000_2539, w_000_2540, w_000_2541, w_000_2542, w_000_2543, w_000_2544, w_000_2545, w_000_2546, w_000_2547, w_000_2548, w_000_2549, w_000_2550, w_000_2551, w_000_2552, w_000_2553, w_000_2554, w_000_2555, w_000_2556, w_000_2557, w_000_2558, w_000_2559, w_000_2560, w_000_2561, w_000_2562, w_000_2563, w_000_2564, w_000_2565, w_000_2566, w_000_2567, w_000_2568, w_000_2569, w_000_2570, w_000_2571, w_000_2572, w_000_2573, w_000_2574, w_000_2575, w_000_2576, w_000_2577, w_000_2578, w_000_2579, w_000_2580, w_000_2581, w_000_2582, w_000_2583, w_000_2584, w_000_2585, w_000_2586, w_000_2587, w_000_2588, w_000_2589, w_000_2590, w_000_2591, w_000_2592, w_000_2593, w_000_2594, w_000_2595, w_000_2596, w_000_2597, w_000_2598, w_000_2599, w_000_2600, w_000_2601, w_000_2602, w_000_2603, w_000_2604, w_000_2605, w_000_2606, w_000_2607, w_000_2608, w_000_2609, w_000_2610, w_000_2611, w_000_2612, w_000_2613, w_000_2614, w_000_2615, w_000_2616, w_000_2617, w_000_2618, w_000_2619, w_000_2620, w_000_2621, w_000_2622, w_000_2623, w_000_2624, w_000_2625, w_000_2626, w_000_2627, w_000_2628, w_000_2629, w_000_2630, w_000_2631, w_000_2632, w_000_2633, w_000_2634, w_000_2635, w_000_2636, w_000_2637, w_000_2638, w_000_2639, w_000_2640, w_000_2641, w_000_2642, w_000_2643, w_000_2644, w_000_2645, w_000_2646, w_000_2647, w_000_2648, w_000_2649, w_000_2650, w_000_2651, w_000_2652, w_000_2653, w_000_2654, w_000_2655, w_000_2656, w_000_2657, w_000_2658, w_000_2659, w_000_2660, w_000_2661, w_000_2662, w_000_2663, w_000_2664, w_000_2665, w_000_2666, w_000_2667, w_000_2668, w_000_2669, w_000_2670, w_000_2671, w_000_2672, w_000_2673, w_000_2674, w_000_2675, w_000_2676, w_000_2677, w_000_2678, w_000_2679, w_000_2680, w_000_2681, w_000_2682, w_000_2683, w_000_2684, w_000_2685, w_000_2686, w_000_2687, w_000_2688, w_000_2689, w_000_2690, w_000_2691, w_000_2692, w_000_2693, w_000_2694, w_000_2695, w_000_2696, w_000_2697, w_000_2698, w_000_2699, w_000_2700, w_000_2701, w_000_2702, w_000_2703, w_000_2704, w_000_2705, w_000_2706, w_000_2707, w_000_2708, w_000_2709, w_000_2710, w_000_2711, w_000_2712, w_000_2713, w_000_2714, w_000_2715, w_000_2716, w_000_2717, w_000_2718, w_000_2719, w_000_2720, w_000_2721, w_000_2722, w_000_2723, w_000_2724, w_000_2725, w_000_2726, w_000_2727, w_000_2728, w_000_2729, w_000_2730, w_000_2731, w_000_2732, w_000_2733, w_000_2734, w_000_2735, w_000_2736, w_000_2737, w_000_2738, w_000_2739, w_000_2740, w_000_2741, w_000_2742, w_000_2743, w_000_2744, w_000_2745, w_000_2746, w_000_2747, w_000_2748, w_000_2749, w_000_2750, w_000_2751, w_000_2752, w_000_2753, w_000_2754, w_000_2755, w_000_2756, w_000_2757, w_000_2758, w_000_2759, w_000_2760, w_000_2761, w_000_2762, w_000_2763, w_000_2764, w_000_2765, w_000_2766, w_000_2767, w_000_2768, w_000_2769, w_000_2770, w_000_2771, w_000_2772, w_000_2773, w_000_2774, w_000_2775, w_000_2776, w_000_2777, w_000_2778, w_000_2779, w_000_2780, w_000_2781, w_000_2782, w_000_2783, w_000_2784, w_000_2785, w_000_2786, w_000_2787, w_000_2788, w_000_2789, w_000_2790, w_000_2791, w_000_2792, w_000_2793, w_000_2794, w_000_2795, w_000_2796, w_000_2797, w_000_2798, w_000_2799, w_000_2800, w_000_2801, w_000_2802, w_000_2803, w_000_2804, w_000_2805, w_000_2806, w_000_2807, w_000_2808, w_000_2809, w_000_2810, w_000_2811, w_000_2812, w_000_2813, w_000_2814, w_000_2815, w_000_2816, w_000_2817, w_000_2818, w_000_2819, w_000_2820, w_000_2821, w_000_2822, w_000_2823, w_000_2824, w_000_2825, w_000_2826, w_000_2827, w_000_2828, w_000_2829, w_000_2830, w_000_2831, w_000_2832, w_000_2833, w_000_2834, w_000_2835, w_000_2836, w_000_2837, w_000_2838, w_000_2839, w_000_2840, w_000_2841, w_000_2842, w_000_2843, w_000_2844, w_000_2845, w_000_2846, w_000_2847, w_000_2848, w_000_2849, w_000_2850, w_000_2851, w_000_2852, w_000_2853, w_000_2854, w_000_2855, w_000_2856, w_000_2857, w_000_2858, w_000_2859, w_000_2860, w_000_2861, w_000_2862, w_000_2863, w_000_2864, w_000_2865, w_000_2866, w_000_2867, w_000_2868, w_000_2869, w_000_2870, w_000_2871, w_000_2872, w_000_2873, w_000_2874, w_000_2875, w_000_2876, w_000_2877, w_000_2878, w_000_2879, w_000_2880, w_000_2881, w_000_2882, w_000_2883, w_000_2884, w_000_2885, w_000_2886, w_000_2887, w_000_2888, w_000_2889, w_000_2890, w_000_2891, w_000_2892, w_000_2893, w_000_2894, w_000_2895, w_000_2896, w_000_2897, w_000_2898, w_000_2899, w_000_2900, w_000_2901, w_000_2902, w_000_2903, w_000_2904, w_000_2905, w_000_2906, w_000_2907, w_000_2908, w_000_2909, w_000_2910, w_000_2911, w_000_2912, w_000_2913, w_000_2914, w_000_2915, w_000_2916, w_000_2917, w_000_2918, w_000_2919, w_000_2920, w_000_2921, w_000_2922, w_000_2923, w_000_2924, w_000_2925, w_000_2926, w_000_2927, w_000_2928, w_000_2929, w_000_2930, w_000_2931, w_000_2932, w_000_2933, w_000_2934, w_000_2935, w_000_2936, w_000_2937, w_000_2938, w_000_2939, w_000_2940, w_000_2941, w_000_2942, w_000_2943, w_000_2944, w_000_2945, w_000_2946, w_000_2947, w_000_2948, w_000_2949, w_000_2950, w_000_2951, w_000_2952, w_000_2953, w_000_2954, w_000_2955, w_000_2956, w_000_2957, w_000_2958, w_000_2959, w_000_2960, w_000_2961, w_000_2962, w_000_2963, w_000_2964, w_000_2965, w_000_2966, w_000_2967, w_000_2968, w_000_2969, w_000_2970, w_000_2971, w_000_2972, w_000_2973, w_000_2974, w_000_2975, w_000_2976, w_000_2977, w_000_2978, w_000_2979, w_000_2980, w_000_2981, w_000_2982, w_000_2983, w_000_2984, w_000_2985, w_000_2986, w_000_2987, w_000_2988, w_000_2989, w_000_2990, w_000_2991, w_000_2992, w_000_2993, w_000_2994, w_000_2995, w_000_2996, w_000_2997, w_000_2998, w_000_2999, w_000_3000, w_000_3001, w_000_3002, w_000_3003, w_000_3004, w_000_3005, w_000_3006, w_000_3007, w_000_3008, w_000_3009, w_000_3010, w_000_3011, w_000_3012, w_000_3013, w_000_3014, w_000_3015, w_000_3016, w_000_3017, w_000_3019, w_000_3020, w_000_3021, w_000_3022, w_000_3023, w_000_3024, w_000_3025, w_000_3026, w_000_3027, w_000_3028, w_000_3029, w_000_3030, w_000_3031, w_000_3032, w_000_3033, w_000_3034, w_000_3035, w_000_3036, w_000_3037, w_000_3038, w_000_3039, w_000_3040, w_000_3041, w_000_3042, w_000_3043, w_000_3044, w_000_3045, w_000_3046, w_000_3047, w_000_3048, w_000_3049, w_000_3050, w_000_3051, w_000_3052, w_000_3053, w_000_3054, w_000_3055, w_000_3056, w_000_3057, w_000_3058, w_000_3059, w_000_3060, w_000_3061, w_000_3062, w_000_3063, w_000_3064, w_000_3065, w_000_3066, w_000_3067, w_000_3068, w_000_3069, w_000_3070, w_000_3071, w_000_3072, w_000_3073, w_000_3074, w_000_3075, w_000_3076, w_000_3077, w_000_3078, w_000_3079, w_000_3080, w_000_3081, w_000_3082, w_000_3083, w_000_3084, w_000_3085, w_000_3086, w_000_3087, w_000_3088, w_000_3089, w_000_3090, w_000_3091, w_000_3092, w_000_3093, w_000_3094, w_000_3095, w_000_3096, w_000_3097, w_000_3098, w_000_3099, w_000_3100, w_000_3101, w_000_3102, w_000_3103, w_000_3104, w_000_3105, w_000_3106, w_000_3107, w_000_3108, w_000_3109, w_000_3110, w_000_3111, w_000_3112, w_000_3113, w_000_3114, w_000_3115, w_000_3116, w_000_3117, w_000_3118, w_000_3119, w_000_3120, w_000_3121, w_000_3122, w_000_3123, w_000_3124, w_000_3125, w_000_3126, w_000_3127, w_000_3128, w_000_3129, w_000_3130, w_000_3131, w_000_3132, w_000_3133, w_000_3134, w_000_3135, w_000_3136, w_000_3137, w_000_3138, w_000_3139, w_000_3140, w_000_3141, w_000_3142, w_000_3143, w_000_3144, w_000_3145, w_000_3146, w_000_3147, w_000_3148, w_000_3149, w_000_3150, w_000_3151, w_000_3152, w_000_3153, w_000_3154, w_000_3155, w_000_3156, w_000_3157, w_000_3158, w_000_3159, w_000_3160, w_000_3161, w_000_3162, w_000_3163, w_000_3164, w_000_3165, w_000_3166, w_000_3167, w_000_3168, w_000_3169, w_000_3170, w_000_3171, w_000_3172, w_000_3173, w_000_3174, w_000_3175, w_000_3176, w_000_3177, w_000_3178, w_000_3179, w_000_3180, w_000_3181, w_000_3182, w_000_3183, w_000_3184, w_000_3185, w_000_3186, w_000_3187, w_000_3188, w_000_3189, w_000_3190, w_000_3191, w_000_3192, w_000_3193, w_000_3194, w_000_3195, w_000_3196, w_000_3197, w_000_3198, w_000_3199, w_000_3200, w_000_3201, w_000_3202, w_000_3203, w_000_3204, w_000_3205, w_000_3206, w_000_3207, w_000_3208, w_000_3209, w_000_3210, w_000_3211, w_000_3212, w_000_3213, w_000_3214, w_000_3215, w_000_3216, w_000_3217, w_000_3218, w_000_3219, w_000_3220, w_000_3221, w_000_3222, w_000_3223, w_000_3224, w_000_3225, w_000_3226, w_000_3227, w_000_3228, w_000_3229, w_000_3230, w_000_3231, w_000_3232, w_000_3233, w_000_3234, w_000_3235, w_000_3236, w_000_3237, w_000_3238, w_000_3239, w_000_3240, w_000_3241, w_000_3242, w_000_3243, w_000_3244, w_000_3245, w_000_3246, w_000_3247, w_000_3248, w_000_3249, w_000_3250, w_000_3251, w_000_3252, w_000_3253, w_000_3254, w_000_3255, w_000_3256, w_000_3257, w_000_3258, w_000_3259, w_000_3260, w_000_3261, w_000_3262, w_000_3263, w_000_3264, w_000_3265, w_000_3266, w_000_3267, w_000_3268, w_000_3269, w_000_3270, w_000_3271, w_000_3272, w_000_3273, w_000_3274, w_000_3275, w_000_3276, w_000_3277, w_000_3278, w_000_3279, w_000_3280, w_000_3281, w_000_3282, w_000_3283, w_000_3284, w_000_3285, w_000_3286, w_000_3287, w_000_3288, w_000_3289, w_000_3290, w_000_3291, w_000_3292, w_000_3293, w_000_3294, w_000_3295, w_000_3296, w_000_3297, w_000_3298, w_000_3299, w_000_3300, w_000_3301, w_000_3302, w_000_3303, w_000_3304, w_000_3305, w_000_3306, w_000_3307, w_000_3308, w_000_3309, w_000_3310, w_000_3311, w_000_3312, w_000_3313, w_000_3314, w_000_3315, w_000_3316, w_000_3317, w_000_3318, w_000_3319, w_000_3320, w_000_3321, w_000_3322, w_000_3323, w_000_3324, w_000_3325, w_000_3326, w_000_3327, w_000_3328, w_000_3329, w_000_3330, w_000_3331, w_000_3332, w_000_3333, w_000_3334, w_000_3335, w_000_3336, w_000_3337, w_000_3338, w_000_3339, w_000_3340, w_000_3341, w_000_3342, w_000_3343, w_000_3344, w_000_3345, w_000_3346, w_000_3347, w_000_3348, w_000_3349, w_000_3350, w_000_3351, w_000_3352, w_000_3353, w_000_3354, w_000_3355, w_000_3356, w_000_3357, w_000_3358, w_000_3359, w_000_3360, w_000_3361, w_000_3362, w_000_3363, w_000_3364, w_000_3365, w_000_3366, w_000_3367, w_000_3368, w_000_3369, w_000_3370, w_000_3371, w_000_3372, w_000_3373, w_000_3374, w_000_3375, w_000_3376, w_000_3377, w_000_3378, w_000_3379, w_000_3380, w_000_3381, w_000_3382, w_000_3383, w_000_3384, w_000_3385, w_000_3386, w_000_3387, w_000_3388, w_000_3389, w_000_3390, w_000_3391, w_000_3392, w_000_3393, w_000_3394, w_000_3395, w_000_3396, w_000_3397, w_000_3398, w_000_3399, w_000_3400, w_000_3401, w_000_3402, w_000_3403, w_000_3404, w_000_3405, w_000_3406, w_000_3407, w_000_3408, w_000_3409, w_000_3410, w_000_3411, w_000_3412, w_000_3413, w_000_3414, w_000_3415, w_000_3416, w_000_3417, w_000_3418, w_000_3419, w_000_3420, w_000_3421, w_000_3422, w_000_3423, w_000_3424, w_000_3425, w_000_3426, w_000_3427, w_000_3428, w_000_3429, w_000_3430, w_000_3431, w_000_3432, w_000_3433, w_000_3434, w_000_3435, w_000_3436, w_000_3437, w_000_3438, w_000_3439, w_000_3440, w_000_3441, w_000_3442, w_000_3443, w_000_3444, w_000_3445, w_000_3446, w_000_3447, w_000_3448, w_000_3449, w_000_3450, w_000_3451, w_000_3452, w_000_3453, w_000_3454, w_000_3455, w_000_3456, w_000_3457, w_000_3458, w_000_3459, w_000_3460, w_000_3461, w_000_3462, w_000_3463, w_000_3464, w_000_3465, w_000_3466, w_000_3467, w_000_3468, w_000_3469, w_000_3470, w_000_3471, w_000_3472, w_000_3473, w_000_3474, w_000_3475, w_000_3476, w_000_3477, w_000_3478, w_000_3479, w_000_3480, w_000_3481, w_000_3482, w_000_3483, w_000_3484, w_000_3485, w_000_3486, w_000_3487, w_000_3488, w_000_3489, w_000_3490, w_000_3491, w_000_3492, w_000_3493, w_000_3494, w_000_3495, w_000_3496, w_000_3497, w_000_3498, w_000_3499, w_000_3500, w_000_3501, w_000_3502, w_000_3503, w_000_3504, w_000_3505, w_000_3506, w_000_3507, w_000_3508, w_000_3509, w_000_3510, w_000_3511, w_000_3512, w_000_3513, w_000_3514, w_000_3515, w_000_3516, w_000_3517, w_000_3518, w_000_3519, w_000_3520, w_000_3521, w_000_3522, w_000_3523, w_000_3524, w_000_3525, w_000_3526, w_000_3527, w_000_3528, w_000_3529, w_000_3530, w_000_3531, w_000_3532, w_000_3533, w_000_3534, w_000_3535, w_000_3536, w_000_3537, w_000_3538, w_000_3539, w_000_3540, w_000_3541, w_000_3542, w_000_3543, w_000_3544, w_000_3545, w_000_3546, w_000_3547, w_000_3548, w_000_3549, w_000_3550, w_000_3551, w_000_3552, w_000_3553, w_000_3554, w_000_3555, w_000_3556, w_000_3557, w_000_3558, w_000_3559, w_000_3560, w_000_3561, w_000_3562, w_000_3563, w_000_3564, w_000_3565, w_000_3566, w_000_3567, w_000_3568, w_000_3569, w_000_3570, w_000_3571, w_000_3572, w_000_3573, w_000_3574, w_000_3575, w_000_3576, w_000_3577, w_000_3578, w_000_3579, w_000_3580, w_000_3581, w_000_3582, w_000_3583, w_000_3584, w_000_3585, w_000_3586, w_000_3587, w_000_3588, w_000_3589, w_000_3590, w_000_3591, w_000_3592, w_000_3593, w_000_3594, w_000_3595, w_000_3596, w_000_3597, w_000_3598, w_000_3599, w_000_3600, w_000_3601, w_000_3602, w_000_3603, w_000_3604, w_000_3605, w_000_3606, w_000_3607, w_000_3608, w_000_3609, w_000_3610, w_000_3611, w_000_3612, w_000_3613, w_000_3614, w_000_3615, w_000_3616, w_000_3617, w_000_3618, w_000_3619, w_000_3620, w_000_3621, w_000_3622, w_000_3623, w_000_3624, w_000_3625, w_000_3626, w_000_3627, w_000_3628, w_000_3629, w_000_3630, w_000_3631, w_000_3632, w_000_3633, w_000_3634, w_000_3635, w_000_3636, w_000_3637, w_000_3638, w_000_3639, w_000_3640, w_000_3641, w_000_3642, w_000_3643, w_000_3644, w_000_3645, w_000_3646, w_000_3647, w_000_3648, w_000_3649, w_000_3650, w_000_3651, w_000_3652, w_000_3653, w_000_3654, w_000_3655, w_000_3656, w_000_3657, w_000_3658, w_000_3659, w_000_3660, w_000_3661, w_000_3662, w_000_3663, w_000_3664, w_000_3665, w_000_3666, w_000_3667, w_000_3668, w_000_3669, w_000_3670, w_000_3671, w_000_3672, w_000_3673, w_000_3674, w_000_3675, w_000_3676, w_000_3677, w_000_3678, w_000_3679, w_000_3680, w_000_3681, w_000_3682, w_000_3683, w_000_3684, w_000_3685, w_000_3686, w_000_3687, w_000_3688, w_000_3689, w_000_3690, w_000_3691, w_000_3692, w_000_3693, w_000_3694, w_000_3695, w_000_3696, w_000_3697, w_000_3698, w_000_3699, w_000_3700, w_000_3701, w_000_3702, w_000_3703, w_000_3704, w_000_3705, w_000_3706, w_000_3707, w_000_3708, w_000_3709, w_000_3710, w_000_3711, w_000_3712, w_000_3713, w_000_3714, w_000_3715, w_000_3716, w_000_3717, w_000_3718, w_000_3719, w_000_3720, w_000_3721, w_000_3722, w_000_3723, w_000_3724, w_000_3725, w_000_3726, w_000_3727, w_000_3728, w_000_3729, w_000_3730, w_000_3731, w_000_3732, w_000_3733, w_000_3734, w_000_3735, w_000_3736, w_000_3737, w_000_3738, w_000_3739, w_000_3740, w_000_3741, w_000_3742, w_000_3743, w_000_3744, w_000_3745, w_000_3746, w_000_3747, w_000_3748, w_000_3749, w_000_3750, w_000_3751, w_000_3752, w_000_3753, w_000_3754, w_000_3755, w_000_3756, w_000_3757, w_000_3758, w_000_3759, w_000_3760, w_000_3761, w_000_3762, w_000_3763, w_000_3764, w_000_3765, w_000_3766, w_000_3767, w_000_3768, w_000_3769, w_000_3770, w_000_3771, w_000_3772, w_000_3773, w_000_3774, w_000_3775, w_000_3776, w_000_3777, w_000_3778, w_000_3779, w_000_3780, w_000_3781, w_000_3782, w_000_3783, w_000_3784, w_000_3785, w_000_3786, w_000_3787, w_000_3788, w_000_3789, w_000_3790, w_000_3791, w_000_3792, w_000_3793, w_000_3794, w_000_3795, w_000_3796, w_000_3797, w_000_3798, w_000_3799, w_000_3800, w_000_3801, w_000_3802, w_000_3803, w_000_3804, w_000_3805, w_000_3806, w_000_3807, w_000_3808, w_000_3809, w_000_3810, w_000_3811, w_000_3812, w_000_3813, w_000_3814, w_000_3815, w_000_3816, w_000_3817, w_000_3818, w_000_3819, w_000_3820, w_000_3821, w_000_3822, w_000_3823, w_000_3824, w_000_3825, w_000_3826, w_000_3827, w_000_3828, w_000_3829, w_000_3830, w_000_3831, w_000_3832, w_000_3833, w_000_3834, w_000_3835, w_000_3836, w_000_3837, w_000_3838, w_000_3839, w_000_3840, w_000_3841, w_000_3842, w_000_3843, w_000_3844, w_000_3845, w_000_3846, w_000_3847, w_000_3848, w_000_3849, w_000_3850, w_000_3851, w_000_3852, w_000_3853, w_000_3854, w_000_3855, w_000_3856, w_000_3857, w_000_3858, w_000_3859, w_000_3860, w_000_3861, w_000_3862, w_000_3863, w_000_3864, w_000_3865, w_000_3866, w_000_3867, w_000_3868, w_000_3869, w_000_3870, w_000_3871, w_000_3872, w_000_3873, w_000_3874, w_000_3875, w_000_3876, w_000_3877, w_000_3878, w_000_3879, w_000_3880, w_000_3881, w_000_3882, w_000_3883, w_000_3884, w_000_3885, w_000_3886, w_000_3887, w_000_3888, w_000_3889, w_000_3890, w_000_3891, w_000_3892, w_000_3893, w_000_3894, w_000_3895, w_000_3896, w_000_3897, w_000_3898, w_000_3899, w_000_3900, w_000_3901, w_000_3902, w_000_3903, w_000_3904, w_000_3905, w_000_3906, w_000_3907, w_000_3908, w_000_3909, w_000_3910, w_000_3911, w_000_3912, w_000_3913, w_000_3914, w_000_3915, w_000_3916, w_000_3917, w_000_3918, w_000_3919, w_000_3920, w_000_3921, w_000_3922, w_000_3923, w_000_3924, w_000_3925, w_000_3926, w_000_3927, w_000_3928, w_000_3929, w_000_3930, w_000_3931, w_000_3932, w_000_3933, w_000_3934, w_000_3935, w_000_3936, w_000_3937, w_000_3938, w_000_3939, w_000_3940, w_000_3941, w_000_3942, w_000_3943, w_000_3944, w_000_3945, w_000_3946, w_000_3947, w_000_3948, w_000_3949, w_000_3950, w_000_3951, w_000_3952, w_000_3953, w_000_3954, w_000_3955, w_000_3956, w_000_3957, w_000_3958, w_000_3959, w_000_3960, w_000_3961, w_000_3962, w_000_3963, w_000_3964, w_000_3965, w_000_3966, w_000_3967, w_000_3968, w_000_3969, w_000_3970, w_000_3971, w_000_3972, w_000_3973, w_000_3974, w_000_3975, w_000_3976, w_000_3977, w_000_3978, w_000_3979, w_000_3980, w_000_3981, w_000_3982, w_000_3983, w_000_3984, w_000_3985, w_000_3986, w_000_3987, w_000_3988, w_000_3989, w_000_3990, w_000_3991, w_000_3992, w_000_3993, w_000_3994, w_000_3995, w_000_3996, w_000_3997, w_000_3998, w_000_3999, w_000_4000, w_000_4001, w_000_4002, w_000_4003, w_000_4004, w_000_4005, w_000_4006, w_000_4007, w_000_4008, w_000_4009, w_000_4010, w_000_4011, w_000_4012, w_000_4013, w_000_4014, w_000_4015, w_000_4016, w_000_4017, w_000_4018, w_000_4019, w_000_4020, w_000_4021, w_000_4022, w_000_4023, w_000_4024, w_000_4025, w_000_4026, w_000_4027, w_000_4028, w_000_4029, w_000_4030, w_000_4031, w_000_4032, w_000_4033, w_000_4034, w_000_4035, w_000_4036, w_000_4037, w_000_4038, w_000_4039, w_000_4040, w_000_4041, w_000_4042, w_000_4043, w_000_4044, w_000_4045, w_000_4046, w_000_4047, w_000_4048, w_000_4049, w_000_4050, w_000_4051, w_000_4052, w_000_4053, w_000_4054, w_000_4055, w_000_4056, w_000_4057, w_000_4058, w_000_4059, w_000_4060, w_000_4061, w_000_4062, w_000_4063, w_000_4064, w_000_4065, w_000_4066, w_000_4067, w_000_4068, w_000_4069, w_000_4070, w_000_4071, w_000_4072, w_000_4073, w_000_4074, w_000_4075, w_000_4076, w_000_4077, w_000_4078, w_000_4079, w_000_4080, w_000_4081, w_000_4082, w_000_4083, w_000_4084, w_000_4085, w_000_4086, w_000_4087, w_000_4088, w_000_4089, w_000_4090, w_000_4091, w_000_4092, w_000_4093, w_000_4094, w_000_4095, w_000_4096, w_000_4097, w_000_4098, w_000_4099, w_000_4100, w_000_4101, w_000_4102, w_000_4103, w_000_4104, w_000_4105, w_000_4106, w_000_4107, w_000_4108, w_000_4109, w_000_4110, w_000_4111, w_000_4112, w_000_4113, w_000_4114, w_000_4115, w_000_4116, w_000_4117, w_000_4118, w_000_4119, w_000_4120, w_000_4121, w_000_4122, w_000_4123, w_000_4124, w_000_4125, w_000_4126, w_000_4127, w_000_4128, w_000_4129, w_000_4130, w_000_4131, w_000_4132, w_000_4133, w_000_4134, w_000_4135, w_000_4136, w_000_4137, w_000_4138, w_000_4139, w_000_4140, w_000_4141, w_000_4142, w_000_4143, w_000_4144, w_000_4145, w_000_4146, w_000_4147, w_000_4148, w_000_4149, w_000_4150, w_000_4151, w_000_4152, w_000_4153, w_000_4154, w_000_4155, w_000_4156, w_000_4157, w_000_4158, w_000_4159, w_000_4160, w_000_4161, w_000_4162, w_000_4163, w_000_4164, w_000_4165, w_000_4166, w_000_4167, w_000_4168, w_000_4169, w_000_4170, w_000_4171, w_000_4172, w_000_4173, w_000_4174, w_000_4175, w_000_4176, w_000_4177, w_000_4178, w_000_4179, w_000_4180, w_000_4181, w_000_4182, w_000_4183, w_000_4184, w_000_4185, w_000_4186, w_000_4187, w_000_4188, w_000_4189, w_000_4190, w_000_4191, w_000_4192, w_000_4193, w_000_4194, w_000_4195, w_000_4196, w_000_4197, w_000_4198, w_000_4199, w_000_4200, w_000_4201, w_000_4202, w_000_4203, w_000_4204, w_000_4205, w_000_4206, w_000_4207, w_000_4208, w_000_4209, w_000_4210, w_000_4211, w_000_4212, w_000_4213, w_000_4215, w_000_4216, w_000_4217, w_000_4218, w_000_4219, w_000_4220, w_000_4221, w_000_4222, w_000_4223, w_000_4224, w_000_4225, w_000_4226, w_000_4227, w_000_4228, w_000_4229, w_000_4230, w_000_4231, w_000_4232, w_000_4233, w_000_4234, w_000_4235, w_000_4236, w_000_4237, w_000_4238, w_000_4239, w_000_4240, w_000_4241, w_000_4242, w_000_4243, w_000_4244, w_000_4245, w_000_4246, w_000_4247, w_000_4248, w_000_4249, w_000_4250, w_000_4251, w_000_4252, w_000_4253, w_000_4254, w_000_4255, w_000_4256, w_000_4257, w_000_4258, w_000_4259, w_000_4260, w_000_4261, w_000_4262, w_000_4263, w_000_4264, w_000_4265, w_000_4266, w_000_4267, w_000_4268, w_000_4269, w_000_4270, w_000_4271, w_000_4272, w_000_4273, w_000_4274, w_000_4275, w_000_4276, w_000_4277, w_000_4278, w_000_4279, w_000_4280, w_000_4281, w_000_4282, w_000_4283, w_000_4284, w_000_4285, w_000_4286, w_000_4287, w_000_4288, w_000_4289, w_000_4290, w_000_4291, w_000_4292, w_000_4293, w_000_4294, w_000_4295, w_000_4296, w_000_4297, w_000_4298, w_000_4299, w_000_4300, w_000_4301, w_000_4302, w_000_4303, w_000_4304, w_000_4305, w_000_4306, w_000_4307, w_000_4308, w_000_4309, w_000_4310, w_000_4311, w_000_4312, w_000_4313, w_000_4314, w_000_4315, w_000_4316, w_000_4317, w_000_4318, w_000_4319, w_000_4320, w_000_4321, w_000_4322, w_000_4323, w_000_4324, w_000_4325, w_000_4326, w_000_4327, w_000_4328, w_000_4329, w_000_4330, w_000_4331, w_000_4332, w_000_4333, w_000_4334, w_000_4335, w_000_4336, w_000_4337, w_000_4338, w_000_4339, w_000_4340, w_000_4341, w_000_4342, w_000_4343, w_000_4344, w_000_4345, w_000_4346, w_000_4347, w_000_4349, w_000_4350, w_000_4351, w_000_4352, w_000_4353, w_000_4354, w_000_4355, w_000_4356, w_000_4357, w_000_4358, w_000_4359, w_000_4360, w_000_4361, w_000_4362, w_000_4363, w_000_4364, w_000_4365, w_000_4366, w_000_4367, w_000_4368, w_000_4369, w_000_4370, w_000_4371, w_000_4372, w_000_4373, w_000_4374, w_000_4375, w_000_4376, w_000_4377, w_000_4378, w_000_4379, w_000_4380, w_000_4381, w_000_4382, w_000_4383, w_000_4384, w_000_4385, w_000_4386, w_000_4387, w_000_4388, w_000_4389, w_000_4390, w_000_4391, w_000_4392, w_000_4393, w_000_4394, w_000_4395, w_000_4396, w_000_4397, w_000_4398, w_000_4399, w_000_4400, w_000_4401, w_000_4402, w_000_4403, w_000_4404, w_000_4405, w_000_4406, w_000_4407, w_000_4408, w_000_4409, w_000_4410, w_000_4411, w_000_4412, w_000_4413, w_000_4414, w_000_4415, w_000_4416, w_000_4417, w_000_4418, w_000_4419, w_000_4420, w_000_4421, w_000_4422, w_000_4423, w_000_4424, w_000_4425, w_000_4426, w_000_4427, w_000_4428, w_000_4429, w_000_4430, w_000_4431, w_000_4432, w_000_4433, w_000_4434, w_000_4435, w_000_4436, w_000_4437, w_000_4438, w_000_4439, w_000_4440, w_000_4441, w_000_4442, w_000_4443, w_000_4444, w_000_4445, w_000_4446, w_000_4447, w_000_4448, w_000_4449, w_000_4450, w_000_4451, w_000_4452, w_000_4453, w_000_4454, w_000_4455, w_000_4456, w_000_4457, w_000_4458, w_000_4459, w_000_4460, w_000_4461, w_000_4462, w_000_4463, w_000_4464, w_000_4465, w_000_4466, w_000_4467, w_000_4468, w_000_4469, w_000_4470, w_000_4471, w_000_4472, w_000_4473, w_000_4474, w_000_4475, w_000_4476, w_000_4477, w_000_4478, w_000_4479, w_000_4480, w_000_4481, w_000_4482, w_000_4483, w_000_4484, w_000_4485, w_000_4486, w_000_4487, w_000_4488, w_000_4489, w_000_4490, w_000_4491, w_000_4492, w_000_4493, w_000_4494, w_000_4495, w_000_4496, w_000_4497, w_000_4498, w_000_4499, w_000_4500, w_000_4501, w_000_4502, w_000_4503, w_000_4504, w_000_4505, w_000_4506, w_000_4507, w_000_4508, w_000_4509, w_000_4510, w_000_4511, w_000_4512, w_000_4513, w_000_4514, w_000_4515, w_000_4516, w_000_4517, w_000_4518, w_000_4519, w_000_4520, w_000_4521, w_000_4522, w_000_4523, w_000_4524, w_000_4525, w_000_4526, w_000_4527, w_000_4528, w_000_4529, w_000_4530, w_000_4531, w_000_4532, w_000_4533, w_000_4534, w_000_4535, w_000_4536, w_000_4537, w_000_4538, w_000_4539, w_000_4540, w_000_4541, w_000_4542, w_000_4543, w_000_4544, w_000_4545, w_000_4546, w_000_4547, w_000_4548, w_000_4549, w_000_4550, w_000_4551, w_000_4552, w_000_4553, w_000_4554, w_000_4555, w_000_4556, w_000_4557, w_000_4559, w_000_4560, w_000_4561, w_000_4562, w_000_4563, w_000_4564, w_000_4565, w_000_4566, w_000_4567, w_000_4568, w_000_4569, w_000_4571, w_000_4572, w_000_4573, w_000_4574, w_000_4575, w_000_4576, w_000_4577, w_000_4578, w_000_4579, w_000_4580, w_000_4581, w_000_4582, w_000_4583, w_000_4584, w_000_4585, w_000_4586, w_000_4587, w_000_4588, w_000_4589, w_000_4590, w_000_4591, w_000_4592, w_000_4593, w_000_4594, w_000_4595, w_000_4596, w_000_4597, w_000_4598, w_000_4599, w_000_4600, w_000_4601, w_000_4602, w_000_4603, w_000_4604, w_000_4605, w_000_4606, w_000_4607, w_000_4608, w_000_4609, w_000_4610, w_000_4611, w_000_4612, w_000_4613, w_000_4614, w_000_4615, w_000_4616, w_000_4617, w_000_4618, w_000_4619, w_000_4620, w_000_4621, w_000_4622, w_000_4623, w_000_4624, w_000_4625, w_000_4626, w_000_4627, w_000_4628, w_000_4629, w_000_4630, w_000_4631, w_000_4632, w_000_4633, w_000_4634, w_000_4635, w_000_4636, w_000_4637, w_000_4638, w_000_4639, w_000_4640, w_000_4641, w_000_4642, w_000_4643, w_000_4644, w_000_4645, w_000_4646, w_000_4647, w_000_4648, w_000_4649, w_000_4650, w_000_4651, w_000_4652, w_000_4653, w_000_4654, w_000_4655, w_000_4656, w_000_4657, w_000_4658, w_000_4659, w_000_4660, w_000_4661, w_000_4662, w_000_4663, w_000_4664, w_000_4665, w_000_4666, w_000_4667, w_000_4668, w_000_4669, w_000_4670, w_000_4671, w_000_4672, w_000_4673, w_000_4674, w_000_4675, w_000_4676, w_000_4677, w_000_4678, w_000_4679, w_000_4680, w_000_4681, w_000_4682, w_000_4683, w_000_4684, w_000_4685, w_000_4686, w_000_4687, w_000_4688, w_000_4689, w_000_4690, w_000_4691, w_000_4692, w_000_4693, w_000_4694, w_000_4695, w_000_4696, w_000_4697, w_000_4698, w_000_4699, w_000_4700, w_000_4701, w_000_4702, w_000_4703, w_000_4704, w_000_4705, w_000_4706, w_000_4707, w_000_4708, w_000_4709, w_000_4710, w_000_4711, w_000_4712, w_000_4713, w_000_4714, w_000_4715, w_000_4716, w_000_4717, w_000_4718, w_000_4719, w_000_4720, w_000_4721, w_000_4722, w_000_4723, w_000_4724, w_000_4725, w_000_4726, w_000_4727, w_000_4728, w_000_4729, w_000_4730, w_000_4731, w_000_4732, w_000_4733, w_000_4734, w_000_4735, w_000_4736, w_000_4737, w_000_4738, w_000_4739, w_000_4740, w_000_4741, w_000_4742, w_000_4743, w_000_4744, w_000_4745, w_000_4746, w_000_4747, w_000_4748, w_000_4749, w_000_4750, w_000_4751, w_000_4752, w_000_4753, w_000_4754, w_000_4755, w_000_4756, w_000_4757, w_000_4758, w_000_4759, w_000_4760, w_000_4761, w_000_4762, w_000_4763, w_000_4764, w_000_4765, w_000_4766, w_000_4767, w_000_4768, w_000_4769, w_000_4770, w_000_4771, w_000_4772, w_000_4773, w_000_4774, w_000_4775, w_000_4776, w_000_4777, w_000_4778, w_000_4779, w_000_4780, w_000_4781, w_000_4782, w_000_4783, w_000_4784, w_000_4785, w_000_4786, w_000_4787, w_000_4788, w_000_4789, w_000_4790, w_000_4791, w_000_4792, w_000_4793, w_000_4794, w_000_4795, w_000_4796, w_000_4797, w_000_4798, w_000_4799, w_000_4800, w_000_4801, w_000_4803, w_000_4804, w_000_4805, w_000_4806, w_000_4807, w_000_4808, w_000_4809, w_000_4810, w_000_4811, w_000_4812, w_000_4813, w_000_4814, w_000_4815, w_000_4816, w_000_4817, w_000_4818, w_000_4819, w_000_4820, w_000_4821, w_000_4822, w_000_4823, w_000_4824, w_000_4825, w_000_4826, w_000_4827, w_000_4828, w_000_4829, w_000_4830, w_000_4831, w_000_4832, w_000_4833, w_000_4834, w_000_4835, w_000_4836, w_000_4837, w_000_4838, w_000_4839, w_000_4840, w_000_4841, w_000_4842, w_000_4843, w_000_4844, w_000_4845, w_000_4846, w_000_4847, w_000_4848, w_000_4849, w_000_4850, w_000_4851, w_000_4852, w_000_4853, w_000_4854, w_000_4855, w_000_4856, w_000_4860, w_000_4861, w_000_4862, w_000_4863, w_000_4864, w_000_4865, w_000_4866, w_000_4867, w_000_4868, w_000_4869, w_000_4870, w_000_4871, w_000_4872, w_000_4873, w_000_4874, w_000_4875, w_000_4876, w_000_4877, w_000_4878, w_000_4879, w_000_4880, w_000_4881, w_000_4882, w_000_4883, w_000_4884, w_000_4885, w_000_4886, w_000_4887, w_000_4889, w_000_4890, w_000_4891, w_000_4892, w_000_4893, w_000_4894, w_000_4895, w_000_4896, w_000_4897, w_000_4898, w_000_4900, w_000_4901, w_000_4902, w_000_4903, w_000_4905, w_000_4906, w_000_4907, w_000_4908, w_000_4909, w_000_4910, w_000_4911, w_000_4912, w_000_4914, w_000_4915, w_000_4916, w_000_4917, w_000_4918, w_000_4920, w_000_4921, w_000_4922, w_000_4923, w_000_4924, w_000_4926, w_000_4927, w_000_4928, w_000_4929, w_000_4930, w_000_4931, w_000_4932, w_000_4933, w_000_4934, w_000_4935, w_000_4936, w_000_4937, w_000_4938, w_000_4939, w_000_4941, w_000_4942, w_000_4944, w_000_4945, w_000_4946, w_000_4947, w_000_4949, w_000_4950, w_000_4952, w_000_4953, w_000_4955, w_000_4956, w_000_4957, w_000_4958, w_000_4959, w_000_4963, w_000_4964, w_000_4966, w_000_4968, w_000_4969, w_000_4970, w_000_4974, w_000_4979, w_000_4980, w_000_4984, w_000_4990, w_000_4991, w_000_4994;
  output w_5000_000, w_5000_001, w_5000_002, w_5000_003, w_5000_004, w_5000_005, w_5000_006, w_5000_007, w_5000_008, w_5000_009, w_5000_010, w_5000_011, w_5000_012, w_5000_013, w_5000_014, w_5000_015, w_5000_016, w_5000_017, w_5000_018, w_5000_019, w_5000_020, w_5000_021, w_5000_022, w_5000_023, w_5000_024, w_5000_025, w_5000_026, w_5000_027, w_5000_028, w_5000_029, w_5000_030, w_5000_031, w_5000_032, w_5000_033, w_5000_034, w_5000_035, w_5000_036, w_5000_037, w_5000_038, w_5000_039, w_5000_040, w_5000_041, w_5000_042, w_5000_043, w_5000_044, w_5000_045, w_5000_046, w_5000_047, w_5000_048, w_5000_049, w_5000_050, w_5000_051, w_5000_052, w_5000_053, w_5000_054, w_5000_055, w_5000_056, w_5000_057, w_5000_058, w_5000_059, w_5000_060, w_5000_061, w_5000_062, w_5000_063, w_5000_064, w_5000_065, w_5000_066, w_5000_067, w_5000_068, w_5000_069, w_5000_070, w_5000_071, w_5000_072, w_5000_073, w_5000_074, w_5000_075, w_5000_076, w_5000_077, w_5000_078, w_5000_079, w_5000_080, w_5000_081, w_5000_082, w_5000_083, w_5000_084, w_5000_085, w_5000_086, w_5000_087, w_5000_088, w_5000_089, w_5000_090, w_5000_091, w_5000_092, w_5000_093, w_5000_094, w_5000_095, w_5000_096, w_5000_097, w_5000_098, w_5000_099, w_5000_100, w_5000_101, w_5000_102, w_5000_103, w_5000_104, w_5000_105, w_5000_106, w_5000_107, w_5000_108, w_5000_109, w_5000_110, w_5000_111, w_5000_112, w_5000_113, w_5000_114, w_5000_115, w_5000_116, w_5000_117, w_5000_118, w_5000_119, w_5000_120, w_5000_121, w_5000_122, w_5000_123, w_5000_124, w_5000_125, w_5000_126, w_5000_127, w_5000_128, w_5000_129, w_5000_130, w_5000_131, w_5000_132, w_5000_133, w_5000_134, w_5000_135, w_5000_136, w_5000_137, w_5000_138, w_5000_139, w_5000_140, w_5000_141, w_5000_142, w_5000_143, w_5000_144, w_5000_145, w_5000_146, w_5000_147, w_5000_148, w_5000_149, w_5000_150, w_5000_151, w_5000_152, w_5000_153, w_5000_154, w_5000_155, w_5000_156, w_5000_157, w_5000_158, w_5000_159, w_5000_160, w_5000_161, w_5000_162, w_5000_163, w_5000_164, w_5000_165, w_5000_166, w_5000_167, w_5000_168, w_5000_169, w_5000_170, w_5000_171, w_5000_172, w_5000_173, w_5000_174, w_5000_175, w_5000_176, w_5000_177, w_5000_178, w_5000_179, w_5000_180, w_5000_181, w_5000_182, w_5000_183, w_5000_184, w_5000_185, w_5000_186, w_5000_187, w_5000_188, w_5000_189, w_5000_190, w_5000_191, w_5000_192, w_5000_193, w_5000_194, w_5000_195, w_5000_196, w_5000_197, w_5000_198, w_5000_199, w_5000_200, w_5000_201, w_5000_202, w_5000_203, w_5000_204, w_5000_205, w_5000_206, w_5000_207, w_5000_208, w_5000_209, w_5000_210, w_5000_211, w_5000_212, w_5000_213, w_5000_214, w_5000_215, w_5000_216, w_5000_217, w_5000_218, w_5000_219, w_5000_220, w_5000_221, w_5000_222, w_5000_223, w_5000_224, w_5000_225, w_5000_226, w_5000_227, w_5000_228, w_5000_229, w_5000_230, w_5000_231, w_5000_232, w_5000_233, w_5000_234, w_5000_235, w_5000_236, w_5000_237, w_5000_238, w_5000_239, w_5000_240, w_5000_241, w_5000_242, w_5000_243, w_5000_244, w_5000_245, w_5000_246, w_5000_247, w_5000_248, w_5000_249, w_5000_250, w_5000_251, w_5000_252, w_5000_253, w_5000_254, w_5000_255, w_5000_256, w_5000_257, w_5000_258, w_5000_259, w_5000_260, w_5000_261, w_5000_262, w_5000_263, w_5000_264, w_5000_265, w_5000_266, w_5000_267, w_5000_268, w_5000_269, w_5000_270, w_5000_271, w_5000_272, w_5000_273, w_5000_274, w_5000_275, w_5000_276, w_5000_277, w_5000_278, w_5000_279, w_5000_280, w_5000_281, w_5000_282, w_5000_283, w_5000_284, w_5000_285, w_5000_286, w_5000_287, w_5000_288, w_5000_289, w_5000_290, w_5000_291, w_5000_292, w_5000_293, w_5000_294, w_5000_295, w_5000_296, w_5000_297, w_5000_298, w_5000_299, w_5000_300, w_5000_301, w_5000_302, w_5000_303, w_5000_304, w_5000_305, w_5000_306, w_5000_307, w_5000_308, w_5000_309, w_5000_310, w_5000_311, w_5000_312, w_5000_313, w_5000_314, w_5000_315, w_5000_316, w_5000_317, w_5000_318, w_5000_319, w_5000_320, w_5000_321, w_5000_322, w_5000_323, w_5000_324, w_5000_325, w_5000_326, w_5000_327, w_5000_328, w_5000_329, w_5000_330, w_5000_331, w_5000_332, w_5000_333, w_5000_334, w_5000_335, w_5000_336, w_5000_337, w_5000_338, w_5000_339, w_5000_340, w_5000_341, w_5000_342, w_5000_343, w_5000_344, w_5000_345, w_5000_346, w_5000_347, w_5000_348, w_5000_349, w_5000_350, w_5000_351, w_5000_352, w_5000_353, w_5000_354, w_5000_355, w_5000_356, w_5000_357, w_5000_358, w_5000_359, w_5000_360, w_5000_361, w_5000_362, w_5000_363, w_5000_364, w_5000_365, w_5000_366, w_5000_367, w_5000_368, w_5000_369, w_5000_370, w_5000_371, w_5000_372, w_5000_373, w_5000_374, w_5000_375, w_5000_376, w_5000_377, w_5000_378, w_5000_379, w_5000_380, w_5000_381, w_5000_382, w_5000_383, w_5000_384, w_5000_385, w_5000_386, w_5000_387, w_5000_388, w_5000_389, w_5000_390, w_5000_391, w_5000_392, w_5000_393, w_5000_394, w_5000_395, w_5000_396, w_5000_397, w_5000_398, w_5000_399, w_5000_400, w_5000_401, w_5000_402, w_5000_403, w_5000_404, w_5000_405, w_5000_406, w_5000_407, w_5000_408, w_5000_409, w_5000_410, w_5000_411, w_5000_412, w_5000_413, w_5000_414, w_5000_415, w_5000_416, w_5000_417, w_5000_418, w_5000_419, w_5000_420, w_5000_421, w_5000_422, w_5000_423, w_5000_424, w_5000_425, w_5000_426, w_5000_427, w_5000_428, w_5000_429, w_5000_430, w_5000_431, w_5000_432, w_5000_433, w_5000_434, w_5000_435, w_5000_436, w_5000_437, w_5000_438, w_5000_439, w_5000_440, w_5000_441, w_5000_442, w_5000_443, w_5000_444, w_5000_445, w_5000_446, w_5000_447, w_5000_448, w_5000_449, w_5000_450, w_5000_451, w_5000_452, w_5000_453, w_5000_454, w_5000_455, w_5000_456, w_5000_457, w_5000_458, w_5000_459, w_5000_460, w_5000_461, w_5000_462, w_5000_463, w_5000_464, w_5000_465, w_5000_466, w_5000_467, w_5000_468, w_5000_469, w_5000_470, w_5000_471, w_5000_472, w_5000_473, w_5000_474, w_5000_475, w_5000_476, w_5000_477, w_5000_478, w_5000_479, w_5000_480, w_5000_481, w_5000_482, w_5000_483, w_5000_484, w_5000_485, w_5000_486, w_5000_487, w_5000_488, w_5000_489, w_5000_490, w_5000_491, w_5000_492, w_5000_493, w_5000_494, w_5000_495, w_5000_496, w_5000_497, w_5000_498, w_5000_499, w_5000_500, w_5000_501, w_5000_502, w_5000_503, w_5000_504, w_5000_505, w_5000_506, w_5000_507, w_5000_508, w_5000_509, w_5000_510, w_5000_511, w_5000_512, w_5000_513, w_5000_514, w_5000_515, w_5000_516, w_5000_517, w_5000_518, w_5000_519, w_5000_520, w_5000_521, w_5000_522, w_5000_523, w_5000_524, w_5000_525, w_5000_526, w_5000_527, w_5000_528, w_5000_529, w_5000_530, w_5000_531, w_5000_532, w_5000_533, w_5000_534, w_5000_535, w_5000_536, w_5000_537, w_5000_538, w_5000_539, w_5000_540, w_5000_541, w_5000_542, w_5000_543, w_5000_544, w_5000_545, w_5000_546, w_5000_547, w_5000_548, w_5000_549, w_5000_550, w_5000_551, w_5000_552, w_5000_553, w_5000_554, w_5000_555, w_5000_556, w_5000_557, w_5000_558, w_5000_559, w_5000_560, w_5000_561, w_5000_562, w_5000_563, w_5000_564, w_5000_565, w_5000_566, w_5000_567, w_5000_568, w_5000_569, w_5000_570, w_5000_571, w_5000_572, w_5000_573, w_5000_574, w_5000_575, w_5000_576, w_5000_577, w_5000_578, w_5000_579, w_5000_580, w_5000_581, w_5000_582, w_5000_583, w_5000_584, w_5000_585, w_5000_586, w_5000_587, w_5000_588, w_5000_589, w_5000_590, w_5000_591, w_5000_592, w_5000_593, w_5000_594, w_5000_595, w_5000_596, w_5000_597, w_5000_598, w_5000_599, w_5000_600, w_5000_601, w_5000_602, w_5000_603, w_5000_604, w_5000_605, w_5000_606, w_5000_607, w_5000_608, w_5000_609, w_5000_610, w_5000_611, w_5000_612, w_5000_613, w_5000_614, w_5000_615, w_5000_616, w_5000_617, w_5000_618, w_5000_619, w_5000_620, w_5000_621, w_5000_622, w_5000_623, w_5000_624, w_5000_625, w_5000_626, w_5000_627, w_5000_628, w_5000_629, w_5000_630, w_5000_631, w_5000_632, w_5000_633, w_5000_634, w_5000_635, w_5000_636, w_5000_637, w_5000_638, w_5000_639, w_5000_640, w_5000_641, w_5000_642, w_5000_643, w_5000_644, w_5000_645, w_5000_646, w_5000_647, w_5000_648, w_5000_649, w_5000_650, w_5000_651, w_5000_652, w_5000_653, w_5000_654, w_5000_655, w_5000_656, w_5000_657, w_5000_658, w_5000_659, w_5000_660, w_5000_661, w_5000_662, w_5000_663, w_5000_664, w_5000_665, w_5000_666, w_5000_667, w_5000_668, w_5000_669, w_5000_670, w_5000_671, w_5000_672, w_5000_673, w_5000_674, w_5000_675, w_5000_676, w_5000_677, w_5000_678, w_5000_679, w_5000_680, w_5000_681, w_5000_682, w_5000_683, w_5000_684, w_5000_685, w_5000_686, w_5000_687, w_5000_688, w_5000_689, w_5000_690, w_5000_691, w_5000_692, w_5000_693, w_5000_694, w_5000_695, w_5000_696, w_5000_697, w_5000_698, w_5000_699, w_5000_700, w_5000_701, w_5000_702, w_5000_703, w_5000_704, w_5000_705, w_5000_706, w_5000_707, w_5000_708, w_5000_709, w_5000_710, w_5000_711, w_5000_712, w_5000_713, w_5000_714, w_5000_715, w_5000_716, w_5000_717, w_5000_718, w_5000_719, w_5000_720, w_5000_721, w_5000_722, w_5000_723, w_5000_724, w_5000_725, w_5000_726, w_5000_727, w_5000_728, w_5000_729, w_5000_730, w_5000_731, w_5000_732, w_5000_733, w_5000_734, w_5000_735, w_5000_736, w_5000_737, w_5000_738, w_5000_739, w_5000_740, w_5000_741, w_5000_742, w_5000_743, w_5000_744, w_5000_745, w_5000_746, w_5000_747, w_5000_748, w_5000_749, w_5000_750, w_5000_751, w_5000_752, w_5000_753, w_5000_754, w_5000_755, w_5000_756, w_5000_757, w_5000_758, w_5000_759, w_5000_760, w_5000_761, w_5000_762, w_5000_763, w_5000_764, w_5000_765, w_5000_766, w_5000_767, w_5000_768, w_5000_769, w_5000_770, w_5000_771, w_5000_772, w_5000_773, w_5000_774, w_5000_775, w_5000_776, w_5000_777, w_5000_778, w_5000_779, w_5000_780, w_5000_781, w_5000_782, w_5000_783, w_5000_784, w_5000_785, w_5000_786, w_5000_787, w_5000_788, w_5000_789, w_5000_790, w_5000_791, w_5000_792, w_5000_793, w_5000_794, w_5000_795, w_5000_796, w_5000_797, w_5000_798, w_5000_799, w_5000_800, w_5000_801, w_5000_802, w_5000_803, w_5000_804, w_5000_805, w_5000_806, w_5000_807, w_5000_808, w_5000_809, w_5000_810, w_5000_811, w_5000_812, w_5000_813, w_5000_814, w_5000_815, w_5000_816, w_5000_817, w_5000_818, w_5000_819, w_5000_820, w_5000_821, w_5000_822, w_5000_823, w_5000_824, w_5000_825, w_5000_826, w_5000_827, w_5000_828, w_5000_829, w_5000_830, w_5000_831, w_5000_832, w_5000_833, w_5000_834, w_5000_835, w_5000_836, w_5000_837, w_5000_838, w_5000_839, w_5000_840, w_5000_841, w_5000_842, w_5000_843, w_5000_844, w_5000_845, w_5000_846, w_5000_847, w_5000_848, w_5000_849, w_5000_850, w_5000_851, w_5000_852, w_5000_853, w_5000_854, w_5000_855, w_5000_856, w_5000_857, w_5000_858, w_5000_859, w_5000_860, w_5000_861, w_5000_862, w_5000_863, w_5000_864, w_5000_865, w_5000_866, w_5000_867, w_5000_868, w_5000_869, w_5000_870, w_5000_871, w_5000_872, w_5000_873, w_5000_874, w_5000_875, w_5000_876, w_5000_877, w_5000_878, w_5000_879, w_5000_880, w_5000_881, w_5000_882, w_5000_883, w_5000_884, w_5000_885, w_5000_886, w_5000_887, w_5000_888, w_5000_889, w_5000_890, w_5000_891, w_5000_892, w_5000_893, w_5000_894, w_5000_895, w_5000_896, w_5000_897, w_5000_898, w_5000_899, w_5000_900, w_5000_901, w_5000_902, w_5000_903, w_5000_904, w_5000_905, w_5000_906, w_5000_907, w_5000_908, w_5000_909, w_5000_910, w_5000_911, w_5000_912, w_5000_913, w_5000_914, w_5000_915, w_5000_916, w_5000_917, w_5000_918, w_5000_919, w_5000_920, w_5000_921, w_5000_922, w_5000_923, w_5000_924, w_5000_925, w_5000_926, w_5000_927, w_5000_928, w_5000_929, w_5000_930, w_5000_931, w_5000_932, w_5000_933, w_5000_934, w_5000_935, w_5000_936, w_5000_937, w_5000_938, w_5000_939, w_5000_940, w_5000_941, w_5000_942, w_5000_943, w_5000_944, w_5000_945, w_5000_946, w_5000_947, w_5000_948, w_5000_949, w_5000_950, w_5000_951, w_5000_952, w_5000_953, w_5000_954, w_5000_955, w_5000_956, w_5000_957, w_5000_958, w_5000_959, w_5000_960, w_5000_961, w_5000_962, w_5000_963, w_5000_964, w_5000_965, w_5000_966, w_5000_967, w_5000_968, w_5000_969, w_5000_970, w_5000_971, w_5000_972, w_5000_973, w_5000_974, w_5000_975, w_5000_976, w_5000_977, w_5000_978, w_5000_979, w_5000_980, w_5000_981, w_5000_982, w_5000_983, w_5000_984, w_5000_985, w_5000_986, w_5000_987, w_5000_988, w_5000_989, w_5000_990, w_5000_991, w_5000_992, w_5000_993, w_5000_994, w_5000_995, w_5000_996, w_5000_997, w_5000_998, w_5000_999, w_5000_1000, w_5000_1001, w_5000_1002, w_5000_1003, w_5000_1004, w_5000_1005, w_5000_1006, w_5000_1007, w_5000_1008, w_5000_1009, w_5000_1010, w_5000_1011, w_5000_1012, w_5000_1013, w_5000_1014, w_5000_1015, w_5000_1016, w_5000_1017, w_5000_1018, w_5000_1019, w_5000_1020, w_5000_1021, w_5000_1022, w_5000_1023, w_5000_1024, w_5000_1025, w_5000_1026, w_5000_1027, w_5000_1028, w_5000_1029, w_5000_1030, w_5000_1031, w_5000_1032, w_5000_1033, w_5000_1034, w_5000_1035, w_5000_1036, w_5000_1037, w_5000_1038, w_5000_1039, w_5000_1040, w_5000_1041, w_5000_1042, w_5000_1043, w_5000_1044, w_5000_1045, w_5000_1046, w_5000_1047, w_5000_1048, w_5000_1049, w_5000_1050, w_5000_1051, w_5000_1052, w_5000_1053, w_5000_1054, w_5000_1055, w_5000_1056, w_5000_1057, w_5000_1058, w_5000_1059, w_5000_1060, w_5000_1061, w_5000_1062, w_5000_1063, w_5000_1064, w_5000_1065, w_5000_1066, w_5000_1067, w_5000_1068, w_5000_1069, w_5000_1070, w_5000_1071, w_5000_1072, w_5000_1073, w_5000_1074, w_5000_1075, w_5000_1076, w_5000_1077, w_5000_1078, w_5000_1079, w_5000_1080, w_5000_1081, w_5000_1082, w_5000_1083, w_5000_1084, w_5000_1085, w_5000_1086, w_5000_1087, w_5000_1088, w_5000_1089, w_5000_1090, w_5000_1091, w_5000_1092, w_5000_1093, w_5000_1094, w_5000_1095, w_5000_1096, w_5000_1097, w_5000_1098, w_5000_1099, w_5000_1100, w_5000_1101, w_5000_1102, w_5000_1103, w_5000_1104, w_5000_1105, w_5000_1106, w_5000_1107, w_5000_1108, w_5000_1109, w_5000_1110, w_5000_1111, w_5000_1112, w_5000_1113, w_5000_1114, w_5000_1115, w_5000_1116, w_5000_1117, w_5000_1118, w_5000_1119, w_5000_1120, w_5000_1121, w_5000_1122, w_5000_1123, w_5000_1124, w_5000_1125, w_5000_1126, w_5000_1127, w_5000_1128, w_5000_1129, w_5000_1130, w_5000_1131, w_5000_1132, w_5000_1133, w_5000_1134, w_5000_1135, w_5000_1136, w_5000_1137, w_5000_1138, w_5000_1139, w_5000_1140, w_5000_1141, w_5000_1142, w_5000_1143, w_5000_1144, w_5000_1145, w_5000_1146, w_5000_1147, w_5000_1148, w_5000_1149, w_5000_1150, w_5000_1151, w_5000_1152, w_5000_1153, w_5000_1154, w_5000_1155, w_5000_1156, w_5000_1157, w_5000_1158, w_5000_1159, w_5000_1160, w_5000_1161, w_5000_1162, w_5000_1163, w_5000_1164, w_5000_1165, w_5000_1166, w_5000_1167, w_5000_1168, w_5000_1169, w_5000_1170, w_5000_1171, w_5000_1172, w_5000_1173, w_5000_1174, w_5000_1175, w_5000_1176, w_5000_1177, w_5000_1178, w_5000_1179, w_5000_1180, w_5000_1181, w_5000_1182, w_5000_1183, w_5000_1184, w_5000_1185, w_5000_1186, w_5000_1187, w_5000_1188, w_5000_1189, w_5000_1190, w_5000_1191, w_5000_1192, w_5000_1193, w_5000_1194, w_5000_1195, w_5000_1196, w_5000_1197, w_5000_1198, w_5000_1199, w_5000_1200, w_5000_1201, w_5000_1202, w_5000_1203, w_5000_1204, w_5000_1205, w_5000_1206, w_5000_1207, w_5000_1208, w_5000_1209, w_5000_1210, w_5000_1211, w_5000_1212, w_5000_1213, w_5000_1214, w_5000_1215, w_5000_1216, w_5000_1217, w_5000_1218, w_5000_1219, w_5000_1220, w_5000_1221, w_5000_1222, w_5000_1223, w_5000_1224, w_5000_1225, w_5000_1226, w_5000_1227, w_5000_1228, w_5000_1229, w_5000_1230, w_5000_1231, w_5000_1232, w_5000_1233, w_5000_1234, w_5000_1235, w_5000_1236, w_5000_1237, w_5000_1238, w_5000_1239, w_5000_1240, w_5000_1241, w_5000_1242, w_5000_1243, w_5000_1244, w_5000_1245, w_5000_1246, w_5000_1247, w_5000_1248, w_5000_1249, w_5000_1250, w_5000_1251, w_5000_1252, w_5000_1253, w_5000_1254, w_5000_1255, w_5000_1256, w_5000_1257, w_5000_1258, w_5000_1259, w_5000_1260, w_5000_1261, w_5000_1262, w_5000_1263, w_5000_1264, w_5000_1265, w_5000_1266, w_5000_1267, w_5000_1268, w_5000_1269, w_5000_1270, w_5000_1271, w_5000_1272, w_5000_1273, w_5000_1274, w_5000_1275, w_5000_1276, w_5000_1277, w_5000_1278, w_5000_1279, w_5000_1280, w_5000_1281, w_5000_1282, w_5000_1283, w_5000_1284, w_5000_1285, w_5000_1286, w_5000_1287, w_5000_1288, w_5000_1289, w_5000_1290, w_5000_1291, w_5000_1292, w_5000_1293, w_5000_1294, w_5000_1295, w_5000_1296, w_5000_1297, w_5000_1298, w_5000_1299, w_5000_1300, w_5000_1301, w_5000_1302, w_5000_1303, w_5000_1304, w_5000_1305, w_5000_1306, w_5000_1307, w_5000_1308, w_5000_1309, w_5000_1310, w_5000_1311, w_5000_1312, w_5000_1313, w_5000_1314, w_5000_1315, w_5000_1316, w_5000_1317, w_5000_1318, w_5000_1319, w_5000_1320, w_5000_1321, w_5000_1322, w_5000_1323, w_5000_1324, w_5000_1325, w_5000_1326, w_5000_1327, w_5000_1328, w_5000_1329, w_5000_1330, w_5000_1331, w_5000_1332, w_5000_1333, w_5000_1334, w_5000_1335, w_5000_1336, w_5000_1337, w_5000_1338, w_5000_1339, w_5000_1340, w_5000_1341, w_5000_1342, w_5000_1343, w_5000_1344, w_5000_1345, w_5000_1346, w_5000_1347, w_5000_1348, w_5000_1349, w_5000_1350, w_5000_1351, w_5000_1352, w_5000_1353, w_5000_1354, w_5000_1355, w_5000_1356, w_5000_1357, w_5000_1358, w_5000_1359, w_5000_1360, w_5000_1361, w_5000_1362, w_5000_1363, w_5000_1364, w_5000_1365, w_5000_1366, w_5000_1367, w_5000_1368, w_5000_1369, w_5000_1370, w_5000_1371, w_5000_1372, w_5000_1373, w_5000_1374, w_5000_1375, w_5000_1376, w_5000_1377, w_5000_1378, w_5000_1379, w_5000_1380, w_5000_1381, w_5000_1382, w_5000_1383, w_5000_1384, w_5000_1385, w_5000_1386, w_5000_1387, w_5000_1388, w_5000_1389, w_5000_1390, w_5000_1391, w_5000_1392, w_5000_1393, w_5000_1394, w_5000_1395, w_5000_1396, w_5000_1397, w_5000_1398, w_5000_1399, w_5000_1400, w_5000_1401, w_5000_1402, w_5000_1403, w_5000_1404, w_5000_1405, w_5000_1406, w_5000_1407, w_5000_1408, w_5000_1409, w_5000_1410, w_5000_1411, w_5000_1412, w_5000_1413, w_5000_1414, w_5000_1415, w_5000_1416, w_5000_1417, w_5000_1418, w_5000_1419, w_5000_1420, w_5000_1421, w_5000_1422, w_5000_1423, w_5000_1424, w_5000_1425, w_5000_1426, w_5000_1427, w_5000_1428, w_5000_1429, w_5000_1430, w_5000_1431, w_5000_1432, w_5000_1433, w_5000_1434, w_5000_1435, w_5000_1436, w_5000_1437, w_5000_1438, w_5000_1439, w_5000_1440, w_5000_1441, w_5000_1442, w_5000_1443, w_5000_1444, w_5000_1445, w_5000_1446, w_5000_1447, w_5000_1448, w_5000_1449, w_5000_1450, w_5000_1451, w_5000_1452, w_5000_1453, w_5000_1454, w_5000_1455, w_5000_1456, w_5000_1457, w_5000_1458, w_5000_1459, w_5000_1460, w_5000_1461, w_5000_1462, w_5000_1463, w_5000_1464, w_5000_1465, w_5000_1466, w_5000_1467, w_5000_1468, w_5000_1469, w_5000_1470, w_5000_1471, w_5000_1472, w_5000_1473, w_5000_1474, w_5000_1475, w_5000_1476, w_5000_1477, w_5000_1478, w_5000_1479, w_5000_1480, w_5000_1481, w_5000_1482, w_5000_1483, w_5000_1484, w_5000_1485, w_5000_1486, w_5000_1487, w_5000_1488, w_5000_1489, w_5000_1490, w_5000_1491, w_5000_1492, w_5000_1493, w_5000_1494, w_5000_1495, w_5000_1496, w_5000_1497, w_5000_1498, w_5000_1499, w_5000_1500, w_5000_1501, w_5000_1502, w_5000_1503, w_5000_1504, w_5000_1505, w_5000_1506, w_5000_1507, w_5000_1508, w_5000_1509, w_5000_1510, w_5000_1511, w_5000_1512, w_5000_1513, w_5000_1514, w_5000_1515, w_5000_1516, w_5000_1517, w_5000_1518, w_5000_1519, w_5000_1520, w_5000_1521, w_5000_1522, w_5000_1523, w_5000_1524, w_5000_1525, w_5000_1526, w_5000_1527, w_5000_1528, w_5000_1529, w_5000_1530, w_5000_1531, w_5000_1532, w_5000_1533, w_5000_1534, w_5000_1535, w_5000_1536, w_5000_1537, w_5000_1538, w_5000_1539, w_5000_1540, w_5000_1541, w_5000_1542, w_5000_1543, w_5000_1544, w_5000_1545, w_5000_1546, w_5000_1547, w_5000_1548, w_5000_1549, w_5000_1550, w_5000_1551, w_5000_1552, w_5000_1553, w_5000_1554, w_5000_1555, w_5000_1556, w_5000_1557, w_5000_1558, w_5000_1559, w_5000_1560, w_5000_1561, w_5000_1562, w_5000_1563, w_5000_1564, w_5000_1565, w_5000_1566, w_5000_1567, w_5000_1568, w_5000_1569, w_5000_1570, w_5000_1571, w_5000_1572, w_5000_1573, w_5000_1574, w_5000_1575, w_5000_1576, w_5000_1577, w_5000_1578, w_5000_1579, w_5000_1580, w_5000_1581, w_5000_1582, w_5000_1583, w_5000_1584, w_5000_1585, w_5000_1586, w_5000_1587, w_5000_1588, w_5000_1589, w_5000_1590, w_5000_1591, w_5000_1592, w_5000_1593, w_5000_1594, w_5000_1595, w_5000_1596, w_5000_1597, w_5000_1598, w_5000_1599, w_5000_1600, w_5000_1601, w_5000_1602, w_5000_1603, w_5000_1604, w_5000_1605, w_5000_1606, w_5000_1607, w_5000_1608, w_5000_1609, w_5000_1610, w_5000_1611, w_5000_1612, w_5000_1613, w_5000_1614, w_5000_1615, w_5000_1616, w_5000_1617, w_5000_1618, w_5000_1619, w_5000_1620, w_5000_1621, w_5000_1622, w_5000_1623, w_5000_1624, w_5000_1625, w_5000_1626, w_5000_1627, w_5000_1628, w_5000_1629, w_5000_1630, w_5000_1631, w_5000_1632, w_5000_1633, w_5000_1634, w_5000_1635, w_5000_1636, w_5000_1637, w_5000_1638, w_5000_1639, w_5000_1640, w_5000_1641, w_5000_1642, w_5000_1643, w_5000_1644, w_5000_1645, w_5000_1646, w_5000_1647, w_5000_1648, w_5000_1649, w_5000_1650, w_5000_1651, w_5000_1652, w_5000_1653, w_5000_1654, w_5000_1655, w_5000_1656, w_5000_1657, w_5000_1658, w_5000_1659, w_5000_1660, w_5000_1661, w_5000_1662, w_5000_1663, w_5000_1664, w_5000_1665, w_5000_1666, w_5000_1667, w_5000_1668, w_5000_1669, w_5000_1670, w_5000_1671, w_5000_1672, w_5000_1673, w_5000_1674, w_5000_1675, w_5000_1676, w_5000_1677, w_5000_1678, w_5000_1679, w_5000_1680, w_5000_1681, w_5000_1682, w_5000_1683, w_5000_1684, w_5000_1685, w_5000_1686, w_5000_1687, w_5000_1688, w_5000_1689, w_5000_1690, w_5000_1691, w_5000_1692, w_5000_1693, w_5000_1694, w_5000_1695, w_5000_1696, w_5000_1697, w_5000_1698, w_5000_1699, w_5000_1700, w_5000_1701, w_5000_1702, w_5000_1703, w_5000_1704, w_5000_1705, w_5000_1706, w_5000_1707, w_5000_1708, w_5000_1709, w_5000_1710, w_5000_1711, w_5000_1712, w_5000_1713, w_5000_1714, w_5000_1715, w_5000_1716, w_5000_1717, w_5000_1718, w_5000_1719, w_5000_1720, w_5000_1721, w_5000_1722, w_5000_1723, w_5000_1724, w_5000_1725, w_5000_1726, w_5000_1727, w_5000_1728, w_5000_1729, w_5000_1730, w_5000_1731, w_5000_1732, w_5000_1733, w_5000_1734, w_5000_1735, w_5000_1736, w_5000_1737, w_5000_1738, w_5000_1739, w_5000_1740, w_5000_1741, w_5000_1742, w_5000_1743, w_5000_1744, w_5000_1745, w_5000_1746, w_5000_1747, w_5000_1748, w_5000_1749, w_5000_1750, w_5000_1751, w_5000_1752, w_5000_1753, w_5000_1754, w_5000_1755, w_5000_1756, w_5000_1757, w_5000_1758, w_5000_1759, w_5000_1760, w_5000_1761, w_5000_1762, w_5000_1763, w_5000_1764, w_5000_1765, w_5000_1766, w_5000_1767, w_5000_1768, w_5000_1769, w_5000_1770, w_5000_1771, w_5000_1772, w_5000_1773, w_5000_1774, w_5000_1775, w_5000_1776, w_5000_1777, w_5000_1778, w_5000_1779, w_5000_1780, w_5000_1781, w_5000_1782, w_5000_1783, w_5000_1784, w_5000_1785, w_5000_1786, w_5000_1787, w_5000_1788, w_5000_1789, w_5000_1790, w_5000_1791, w_5000_1792, w_5000_1793, w_5000_1794, w_5000_1795, w_5000_1796, w_5000_1797, w_5000_1798, w_5000_1799, w_5000_1800, w_5000_1801, w_5000_1802, w_5000_1803, w_5000_1804, w_5000_1805, w_5000_1806, w_5000_1807, w_5000_1808, w_5000_1809, w_5000_1810, w_5000_1811, w_5000_1812, w_5000_1813, w_5000_1814, w_5000_1815, w_5000_1816, w_5000_1817, w_5000_1818, w_5000_1819, w_5000_1820, w_5000_1821, w_5000_1822, w_5000_1823, w_5000_1824, w_5000_1825, w_5000_1826, w_5000_1827, w_5000_1828, w_5000_1829, w_5000_1830, w_5000_1831, w_5000_1832, w_5000_1833, w_5000_1834, w_5000_1835, w_5000_1836, w_5000_1837, w_5000_1838, w_5000_1839, w_5000_1840, w_5000_1841, w_5000_1842, w_5000_1843, w_5000_1844, w_5000_1845, w_5000_1846, w_5000_1847, w_5000_1848, w_5000_1849, w_5000_1850, w_5000_1851, w_5000_1852, w_5000_1853, w_5000_1854, w_5000_1855, w_5000_1856, w_5000_1857, w_5000_1858, w_5000_1859, w_5000_1860, w_5000_1861, w_5000_1862, w_5000_1863, w_5000_1864, w_5000_1865, w_5000_1866, w_5000_1867, w_5000_1868, w_5000_1869, w_5000_1870, w_5000_1871, w_5000_1872, w_5000_1873, w_5000_1874, w_5000_1875, w_5000_1876, w_5000_1877, w_5000_1878, w_5000_1879, w_5000_1880, w_5000_1881, w_5000_1882, w_5000_1883, w_5000_1884, w_5000_1885, w_5000_1886, w_5000_1887, w_5000_1888, w_5000_1889, w_5000_1890, w_5000_1891, w_5000_1892, w_5000_1893, w_5000_1894, w_5000_1895, w_5000_1896, w_5000_1897, w_5000_1898, w_5000_1899, w_5000_1900, w_5000_1901, w_5000_1902, w_5000_1903, w_5000_1904, w_5000_1905, w_5000_1906, w_5000_1907, w_5000_1908, w_5000_1909, w_5000_1910, w_5000_1911, w_5000_1912, w_5000_1913, w_5000_1914, w_5000_1915, w_5000_1916, w_5000_1917, w_5000_1918, w_5000_1919, w_5000_1920, w_5000_1921, w_5000_1922, w_5000_1923, w_5000_1924, w_5000_1925, w_5000_1926, w_5000_1927, w_5000_1928, w_5000_1929, w_5000_1930, w_5000_1931, w_5000_1932, w_5000_1933, w_5000_1934, w_5000_1935, w_5000_1936, w_5000_1937, w_5000_1938, w_5000_1939, w_5000_1940, w_5000_1941, w_5000_1942, w_5000_1943, w_5000_1944, w_5000_1945, w_5000_1946, w_5000_1947, w_5000_1948, w_5000_1949, w_5000_1950, w_5000_1951, w_5000_1952, w_5000_1953, w_5000_1954, w_5000_1955, w_5000_1956, w_5000_1957, w_5000_1958, w_5000_1959, w_5000_1960, w_5000_1961, w_5000_1962, w_5000_1963, w_5000_1964, w_5000_1965, w_5000_1966, w_5000_1967, w_5000_1968, w_5000_1969, w_5000_1970, w_5000_1971, w_5000_1972, w_5000_1973, w_5000_1974, w_5000_1975, w_5000_1976, w_5000_1977, w_5000_1978, w_5000_1979, w_5000_1980, w_5000_1981, w_5000_1982, w_5000_1983, w_5000_1984, w_5000_1985, w_5000_1986, w_5000_1987, w_5000_1988, w_5000_1989, w_5000_1990, w_5000_1991, w_5000_1992, w_5000_1993, w_5000_1994, w_5000_1995, w_5000_1996, w_5000_1997, w_5000_1998, w_5000_1999, w_5000_2000, w_5000_2001, w_5000_2002, w_5000_2003, w_5000_2004, w_5000_2005, w_5000_2006, w_5000_2007, w_5000_2008, w_5000_2009, w_5000_2010, w_5000_2011, w_5000_2012, w_5000_2013, w_5000_2014, w_5000_2015, w_5000_2016, w_5000_2017, w_5000_2018, w_5000_2019, w_5000_2020, w_5000_2021, w_5000_2022, w_5000_2023, w_5000_2024, w_5000_2025, w_5000_2026, w_5000_2027, w_5000_2028, w_5000_2029, w_5000_2030, w_5000_2031, w_5000_2032, w_5000_2033, w_5000_2034, w_5000_2035, w_5000_2036, w_5000_2037, w_5000_2038, w_5000_2039, w_5000_2040, w_5000_2041, w_5000_2042, w_5000_2043, w_5000_2044, w_5000_2045, w_5000_2046, w_5000_2047, w_5000_2048, w_5000_2049, w_5000_2050, w_5000_2051, w_5000_2052, w_5000_2053, w_5000_2054, w_5000_2055, w_5000_2056, w_5000_2057, w_5000_2058, w_5000_2059, w_5000_2060, w_5000_2061, w_5000_2062, w_5000_2063, w_5000_2064, w_5000_2065, w_5000_2066, w_5000_2067, w_5000_2068, w_5000_2069, w_5000_2070, w_5000_2071, w_5000_2072, w_5000_2073, w_5000_2074, w_5000_2075, w_5000_2076, w_5000_2077, w_5000_2078, w_5000_2079, w_5000_2080, w_5000_2081, w_5000_2082, w_5000_2083, w_5000_2084, w_5000_2085, w_5000_2086, w_5000_2087, w_5000_2088, w_5000_2089, w_5000_2090, w_5000_2091, w_5000_2092, w_5000_2093, w_5000_2094, w_5000_2095, w_5000_2096, w_5000_2097, w_5000_2098, w_5000_2099, w_5000_2100, w_5000_2101, w_5000_2102, w_5000_2103, w_5000_2104, w_5000_2105, w_5000_2106, w_5000_2107, w_5000_2108, w_5000_2109, w_5000_2110, w_5000_2111, w_5000_2112, w_5000_2113, w_5000_2114, w_5000_2115, w_5000_2116, w_5000_2117, w_5000_2118, w_5000_2119, w_5000_2120, w_5000_2121, w_5000_2122, w_5000_2123, w_5000_2124, w_5000_2125, w_5000_2126, w_5000_2127, w_5000_2128, w_5000_2129, w_5000_2130, w_5000_2131, w_5000_2132, w_5000_2133, w_5000_2134, w_5000_2135, w_5000_2136, w_5000_2137, w_5000_2138, w_5000_2139, w_5000_2140, w_5000_2141, w_5000_2142, w_5000_2143, w_5000_2144, w_5000_2145, w_5000_2146, w_5000_2147, w_5000_2148, w_5000_2149, w_5000_2150, w_5000_2151, w_5000_2152, w_5000_2153, w_5000_2154, w_5000_2155, w_5000_2156, w_5000_2157, w_5000_2158, w_5000_2159, w_5000_2160, w_5000_2161, w_5000_2162, w_5000_2163, w_5000_2164, w_5000_2165, w_5000_2166, w_5000_2167, w_5000_2168, w_5000_2169, w_5000_2170, w_5000_2171, w_5000_2172, w_5000_2173, w_5000_2174, w_5000_2175, w_5000_2176, w_5000_2177, w_5000_2178, w_5000_2179, w_5000_2180, w_5000_2181, w_5000_2182, w_5000_2183, w_5000_2184, w_5000_2185, w_5000_2186, w_5000_2187, w_5000_2188, w_5000_2189, w_5000_2190, w_5000_2191, w_5000_2192, w_5000_2193, w_5000_2194, w_5000_2195, w_5000_2196, w_5000_2197, w_5000_2198, w_5000_2199, w_5000_2200, w_5000_2201, w_5000_2202, w_5000_2203, w_5000_2204, w_5000_2205, w_5000_2206, w_5000_2207, w_5000_2208, w_5000_2209, w_5000_2210, w_5000_2211, w_5000_2212, w_5000_2213, w_5000_2214, w_5000_2215, w_5000_2216, w_5000_2217, w_5000_2218, w_5000_2219, w_5000_2220, w_5000_2221, w_5000_2222, w_5000_2223, w_5000_2224, w_5000_2225, w_5000_2226, w_5000_2227, w_5000_2228, w_5000_2229, w_5000_2230, w_5000_2231, w_5000_2232, w_5000_2233, w_5000_2234, w_5000_2235, w_5000_2236, w_5000_2237, w_5000_2238, w_5000_2239, w_5000_2240, w_5000_2241, w_5000_2242, w_5000_2243, w_5000_2244, w_5000_2245, w_5000_2246, w_5000_2247, w_5000_2248, w_5000_2249, w_5000_2250, w_5000_2251, w_5000_2252, w_5000_2253, w_5000_2254, w_5000_2255, w_5000_2256, w_5000_2257, w_5000_2258, w_5000_2259, w_5000_2260, w_5000_2261, w_5000_2262, w_5000_2263, w_5000_2264, w_5000_2265, w_5000_2266, w_5000_2267, w_5000_2268, w_5000_2269, w_5000_2270, w_5000_2271, w_5000_2272, w_5000_2273, w_5000_2274, w_5000_2275, w_5000_2276, w_5000_2277, w_5000_2278, w_5000_2279, w_5000_2280, w_5000_2281, w_5000_2282, w_5000_2283, w_5000_2284, w_5000_2285, w_5000_2286, w_5000_2287, w_5000_2288, w_5000_2289, w_5000_2290, w_5000_2291, w_5000_2292, w_5000_2293, w_5000_2294, w_5000_2295, w_5000_2296, w_5000_2297, w_5000_2298, w_5000_2299, w_5000_2300, w_5000_2301, w_5000_2302, w_5000_2303, w_5000_2304, w_5000_2305, w_5000_2306, w_5000_2307, w_5000_2308, w_5000_2309, w_5000_2310, w_5000_2311, w_5000_2312, w_5000_2313, w_5000_2314, w_5000_2315, w_5000_2316, w_5000_2317, w_5000_2318, w_5000_2319, w_5000_2320, w_5000_2321, w_5000_2322, w_5000_2323, w_5000_2324, w_5000_2325, w_5000_2326, w_5000_2327, w_5000_2328, w_5000_2329, w_5000_2330, w_5000_2331, w_5000_2332, w_5000_2333, w_5000_2334, w_5000_2335, w_5000_2336, w_5000_2337, w_5000_2338, w_5000_2339, w_5000_2340, w_5000_2341, w_5000_2342, w_5000_2343, w_5000_2344, w_5000_2345, w_5000_2346, w_5000_2347, w_5000_2348, w_5000_2349, w_5000_2350, w_5000_2351, w_5000_2352, w_5000_2353, w_5000_2354, w_5000_2355, w_5000_2356, w_5000_2357, w_5000_2358, w_5000_2359, w_5000_2360, w_5000_2361, w_5000_2362, w_5000_2363, w_5000_2364, w_5000_2365, w_5000_2366, w_5000_2367, w_5000_2368, w_5000_2369, w_5000_2370, w_5000_2371, w_5000_2372, w_5000_2373, w_5000_2374, w_5000_2375, w_5000_2376, w_5000_2377, w_5000_2378, w_5000_2379, w_5000_2380, w_5000_2381, w_5000_2382, w_5000_2383, w_5000_2384, w_5000_2385, w_5000_2386, w_5000_2387, w_5000_2388, w_5000_2389, w_5000_2390, w_5000_2391, w_5000_2392, w_5000_2393, w_5000_2394, w_5000_2395, w_5000_2396, w_5000_2397, w_5000_2398, w_5000_2399, w_5000_2400, w_5000_2401, w_5000_2402, w_5000_2403, w_5000_2404, w_5000_2405, w_5000_2406, w_5000_2407, w_5000_2408, w_5000_2409, w_5000_2410, w_5000_2411, w_5000_2412, w_5000_2413, w_5000_2414, w_5000_2415, w_5000_2416, w_5000_2417, w_5000_2418, w_5000_2419, w_5000_2420, w_5000_2421, w_5000_2422, w_5000_2423, w_5000_2424, w_5000_2425, w_5000_2426, w_5000_2427, w_5000_2428, w_5000_2429, w_5000_2430, w_5000_2431, w_5000_2432, w_5000_2433, w_5000_2434, w_5000_2435, w_5000_2436, w_5000_2437, w_5000_2438, w_5000_2439, w_5000_2440, w_5000_2441, w_5000_2442, w_5000_2443, w_5000_2444, w_5000_2445, w_5000_2446, w_5000_2447, w_5000_2448, w_5000_2449, w_5000_2450, w_5000_2451, w_5000_2452, w_5000_2453, w_5000_2454, w_5000_2455, w_5000_2456, w_5000_2457, w_5000_2458, w_5000_2459, w_5000_2460, w_5000_2461, w_5000_2462, w_5000_2463, w_5000_2464, w_5000_2465, w_5000_2466, w_5000_2467, w_5000_2468, w_5000_2469, w_5000_2470, w_5000_2471, w_5000_2472, w_5000_2473, w_5000_2474, w_5000_2475, w_5000_2476, w_5000_2477, w_5000_2478, w_5000_2479, w_5000_2480, w_5000_2481, w_5000_2482, w_5000_2483, w_5000_2484, w_5000_2485, w_5000_2486, w_5000_2487, w_5000_2488, w_5000_2489, w_5000_2490, w_5000_2491, w_5000_2492, w_5000_2493, w_5000_2494, w_5000_2495, w_5000_2496, w_5000_2497, w_5000_2498, w_5000_2499, w_5000_2500, w_5000_2501, w_5000_2502, w_5000_2503, w_5000_2504, w_5000_2505, w_5000_2506, w_5000_2507, w_5000_2508, w_5000_2509, w_5000_2510, w_5000_2511, w_5000_2512, w_5000_2513, w_5000_2514, w_5000_2515, w_5000_2516, w_5000_2517, w_5000_2518, w_5000_2519, w_5000_2520, w_5000_2521, w_5000_2522, w_5000_2523, w_5000_2524, w_5000_2525, w_5000_2526, w_5000_2527, w_5000_2528, w_5000_2529, w_5000_2530, w_5000_2531, w_5000_2532, w_5000_2533, w_5000_2534, w_5000_2535, w_5000_2536, w_5000_2537, w_5000_2538, w_5000_2539, w_5000_2540, w_5000_2541, w_5000_2542, w_5000_2543, w_5000_2544, w_5000_2545, w_5000_2546, w_5000_2547, w_5000_2548, w_5000_2549, w_5000_2550, w_5000_2551, w_5000_2552, w_5000_2553, w_5000_2554, w_5000_2555, w_5000_2556, w_5000_2557, w_5000_2558, w_5000_2559, w_5000_2560, w_5000_2561, w_5000_2562, w_5000_2563, w_5000_2564, w_5000_2565, w_5000_2566, w_5000_2567, w_5000_2568, w_5000_2569, w_5000_2570, w_5000_2571, w_5000_2572, w_5000_2573, w_5000_2574, w_5000_2575, w_5000_2576, w_5000_2577, w_5000_2578, w_5000_2579, w_5000_2580, w_5000_2581, w_5000_2582, w_5000_2583, w_5000_2584, w_5000_2585, w_5000_2586, w_5000_2587, w_5000_2588, w_5000_2589, w_5000_2590, w_5000_2591, w_5000_2592, w_5000_2593, w_5000_2594, w_5000_2595, w_5000_2596, w_5000_2597, w_5000_2598, w_5000_2599, w_5000_2600, w_5000_2601, w_5000_2602, w_5000_2603, w_5000_2604, w_5000_2605, w_5000_2606, w_5000_2607, w_5000_2608, w_5000_2609, w_5000_2610, w_5000_2611, w_5000_2612, w_5000_2613, w_5000_2614, w_5000_2615, w_5000_2616, w_5000_2617, w_5000_2618, w_5000_2619, w_5000_2620, w_5000_2621, w_5000_2622, w_5000_2623, w_5000_2624, w_5000_2625, w_5000_2626, w_5000_2627, w_5000_2628, w_5000_2629, w_5000_2630, w_5000_2631, w_5000_2632, w_5000_2633, w_5000_2634, w_5000_2635, w_5000_2636, w_5000_2637, w_5000_2638, w_5000_2639, w_5000_2640, w_5000_2641, w_5000_2642, w_5000_2643, w_5000_2644, w_5000_2645, w_5000_2646, w_5000_2647, w_5000_2648, w_5000_2649, w_5000_2650, w_5000_2651, w_5000_2652, w_5000_2653, w_5000_2654, w_5000_2655, w_5000_2656, w_5000_2657, w_5000_2658, w_5000_2659, w_5000_2660, w_5000_2661, w_5000_2662, w_5000_2663, w_5000_2664, w_5000_2665, w_5000_2666, w_5000_2667, w_5000_2668, w_5000_2669, w_5000_2670, w_5000_2671, w_5000_2672, w_5000_2673, w_5000_2674, w_5000_2675, w_5000_2676, w_5000_2677, w_5000_2678, w_5000_2679, w_5000_2680, w_5000_2681, w_5000_2682, w_5000_2683, w_5000_2684, w_5000_2685, w_5000_2686, w_5000_2687, w_5000_2688, w_5000_2689, w_5000_2690, w_5000_2691, w_5000_2692, w_5000_2693, w_5000_2694, w_5000_2695, w_5000_2696, w_5000_2697, w_5000_2698, w_5000_2699, w_5000_2700, w_5000_2701, w_5000_2702, w_5000_2703, w_5000_2704, w_5000_2705, w_5000_2706, w_5000_2707, w_5000_2708, w_5000_2709, w_5000_2710, w_5000_2711, w_5000_2712, w_5000_2713, w_5000_2714, w_5000_2715, w_5000_2716, w_5000_2717, w_5000_2718, w_5000_2719, w_5000_2720, w_5000_2721, w_5000_2722, w_5000_2723, w_5000_2724, w_5000_2725, w_5000_2726, w_5000_2727, w_5000_2728, w_5000_2729, w_5000_2730, w_5000_2731, w_5000_2732, w_5000_2733, w_5000_2734, w_5000_2735, w_5000_2736, w_5000_2737, w_5000_2738, w_5000_2739, w_5000_2740, w_5000_2741, w_5000_2742, w_5000_2743, w_5000_2744, w_5000_2745, w_5000_2746, w_5000_2747, w_5000_2748, w_5000_2749, w_5000_2750, w_5000_2751, w_5000_2752, w_5000_2753, w_5000_2754, w_5000_2755, w_5000_2756, w_5000_2757, w_5000_2758, w_5000_2759, w_5000_2760, w_5000_2761, w_5000_2762, w_5000_2763, w_5000_2764, w_5000_2765, w_5000_2766, w_5000_2767, w_5000_2768, w_5000_2769, w_5000_2770, w_5000_2771, w_5000_2772, w_5000_2773, w_5000_2774, w_5000_2775, w_5000_2776, w_5000_2777, w_5000_2778, w_5000_2779, w_5000_2780, w_5000_2781, w_5000_2782, w_5000_2783, w_5000_2784, w_5000_2785, w_5000_2786, w_5000_2787, w_5000_2788, w_5000_2789, w_5000_2790, w_5000_2791, w_5000_2792, w_5000_2793, w_5000_2794, w_5000_2795, w_5000_2796, w_5000_2797, w_5000_2798, w_5000_2799, w_5000_2800, w_5000_2801, w_5000_2802, w_5000_2803, w_5000_2804, w_5000_2805, w_5000_2806, w_5000_2807, w_5000_2808, w_5000_2809, w_5000_2810, w_5000_2811, w_5000_2812, w_5000_2813, w_5000_2814, w_5000_2815, w_5000_2816, w_5000_2817, w_5000_2818, w_5000_2819, w_5000_2820, w_5000_2821, w_5000_2822, w_5000_2823, w_5000_2824, w_5000_2825, w_5000_2826, w_5000_2827, w_5000_2828, w_5000_2829, w_5000_2830, w_5000_2831, w_5000_2832, w_5000_2833, w_5000_2834, w_5000_2835, w_5000_2836, w_5000_2837, w_5000_2838, w_5000_2839, w_5000_2840, w_5000_2841, w_5000_2842, w_5000_2843, w_5000_2844, w_5000_2845, w_5000_2846, w_5000_2847, w_5000_2848, w_5000_2849, w_5000_2850, w_5000_2851, w_5000_2852, w_5000_2853, w_5000_2854, w_5000_2855, w_5000_2856, w_5000_2857, w_5000_2858, w_5000_2859, w_5000_2860, w_5000_2861, w_5000_2862, w_5000_2863, w_5000_2864, w_5000_2865, w_5000_2866, w_5000_2867, w_5000_2868, w_5000_2869, w_5000_2870, w_5000_2871, w_5000_2872, w_5000_2873, w_5000_2874, w_5000_2875, w_5000_2876, w_5000_2877, w_5000_2878, w_5000_2879, w_5000_2880, w_5000_2881, w_5000_2882, w_5000_2883, w_5000_2884, w_5000_2885, w_5000_2886, w_5000_2887, w_5000_2888, w_5000_2889, w_5000_2890, w_5000_2891, w_5000_2892, w_5000_2893, w_5000_2894, w_5000_2895, w_5000_2896, w_5000_2897, w_5000_2898, w_5000_2899, w_5000_2900, w_5000_2901, w_5000_2902, w_5000_2903, w_5000_2904, w_5000_2905, w_5000_2906, w_5000_2907, w_5000_2908, w_5000_2909, w_5000_2910, w_5000_2911, w_5000_2912, w_5000_2913, w_5000_2914, w_5000_2915, w_5000_2916, w_5000_2917, w_5000_2918, w_5000_2919, w_5000_2920, w_5000_2921, w_5000_2922, w_5000_2923, w_5000_2924, w_5000_2925, w_5000_2926, w_5000_2927, w_5000_2928, w_5000_2929, w_5000_2930, w_5000_2931, w_5000_2932, w_5000_2933, w_5000_2934, w_5000_2935, w_5000_2936, w_5000_2937, w_5000_2938, w_5000_2939, w_5000_2940, w_5000_2941, w_5000_2942, w_5000_2943, w_5000_2944, w_5000_2945, w_5000_2946, w_5000_2947, w_5000_2948, w_5000_2949, w_5000_2950, w_5000_2951, w_5000_2952, w_5000_2953, w_5000_2954, w_5000_2955, w_5000_2956, w_5000_2957, w_5000_2958, w_5000_2959, w_5000_2960, w_5000_2961, w_5000_2962, w_5000_2963, w_5000_2964, w_5000_2965, w_5000_2966, w_5000_2967, w_5000_2968, w_5000_2969, w_5000_2970, w_5000_2971, w_5000_2972, w_5000_2973, w_5000_2974, w_5000_2975, w_5000_2976, w_5000_2977, w_5000_2978, w_5000_2979, w_5000_2980, w_5000_2981, w_5000_2982, w_5000_2983, w_5000_2984, w_5000_2985, w_5000_2986, w_5000_2987, w_5000_2988, w_5000_2989, w_5000_2990, w_5000_2991, w_5000_2992, w_5000_2993, w_5000_2994, w_5000_2995, w_5000_2996, w_5000_2997, w_5000_2998, w_5000_2999, w_5000_3000, w_5000_3001, w_5000_3002, w_5000_3003, w_5000_3004, w_5000_3005, w_5000_3006, w_5000_3007, w_5000_3008, w_5000_3009, w_5000_3010, w_5000_3011, w_5000_3012, w_5000_3013, w_5000_3014, w_5000_3015, w_5000_3016, w_5000_3017, w_5000_3018, w_5000_3019, w_5000_3020, w_5000_3021, w_5000_3022, w_5000_3023, w_5000_3024, w_5000_3025, w_5000_3026, w_5000_3027, w_5000_3028, w_5000_3029, w_5000_3030, w_5000_3031, w_5000_3032, w_5000_3033, w_5000_3034, w_5000_3035, w_5000_3036, w_5000_3037, w_5000_3038, w_5000_3039, w_5000_3040, w_5000_3041, w_5000_3042, w_5000_3043, w_5000_3044, w_5000_3045, w_5000_3046, w_5000_3047, w_5000_3048, w_5000_3049, w_5000_3050, w_5000_3051, w_5000_3052, w_5000_3053, w_5000_3054, w_5000_3055, w_5000_3056, w_5000_3057, w_5000_3058, w_5000_3059, w_5000_3060, w_5000_3061, w_5000_3062, w_5000_3063, w_5000_3064, w_5000_3065, w_5000_3066, w_5000_3067, w_5000_3068, w_5000_3069, w_5000_3070, w_5000_3071, w_5000_3072, w_5000_3073, w_5000_3074, w_5000_3075, w_5000_3076, w_5000_3077, w_5000_3078, w_5000_3079, w_5000_3080, w_5000_3081, w_5000_3082, w_5000_3083, w_5000_3084, w_5000_3085, w_5000_3086, w_5000_3087, w_5000_3088, w_5000_3089, w_5000_3090, w_5000_3091, w_5000_3092, w_5000_3093, w_5000_3094, w_5000_3095, w_5000_3096, w_5000_3097, w_5000_3098, w_5000_3099, w_5000_3100, w_5000_3101, w_5000_3102, w_5000_3103, w_5000_3104, w_5000_3105, w_5000_3106, w_5000_3107, w_5000_3108, w_5000_3109, w_5000_3110, w_5000_3111, w_5000_3112, w_5000_3113, w_5000_3114, w_5000_3115, w_5000_3116, w_5000_3117, w_5000_3118, w_5000_3119, w_5000_3120, w_5000_3121, w_5000_3122, w_5000_3123, w_5000_3124, w_5000_3125, w_5000_3126, w_5000_3127, w_5000_3128, w_5000_3129, w_5000_3130, w_5000_3131, w_5000_3132, w_5000_3133, w_5000_3134, w_5000_3135, w_5000_3136, w_5000_3137, w_5000_3138, w_5000_3139, w_5000_3140, w_5000_3141, w_5000_3142, w_5000_3143, w_5000_3144, w_5000_3145, w_5000_3146, w_5000_3147, w_5000_3148, w_5000_3149, w_5000_3150, w_5000_3151, w_5000_3152, w_5000_3153, w_5000_3154, w_5000_3155, w_5000_3156, w_5000_3157, w_5000_3158, w_5000_3159, w_5000_3160, w_5000_3161, w_5000_3162, w_5000_3163, w_5000_3164, w_5000_3165, w_5000_3166, w_5000_3167, w_5000_3168, w_5000_3169, w_5000_3170, w_5000_3171, w_5000_3172, w_5000_3173, w_5000_3174, w_5000_3175, w_5000_3176, w_5000_3177, w_5000_3178, w_5000_3179, w_5000_3180, w_5000_3181, w_5000_3182, w_5000_3183, w_5000_3184, w_5000_3185, w_5000_3186, w_5000_3187, w_5000_3188, w_5000_3189, w_5000_3190, w_5000_3191, w_5000_3192, w_5000_3193, w_5000_3194, w_5000_3195, w_5000_3196, w_5000_3197, w_5000_3198, w_5000_3199, w_5000_3200, w_5000_3201, w_5000_3202, w_5000_3203, w_5000_3204, w_5000_3205, w_5000_3206, w_5000_3207, w_5000_3208, w_5000_3209, w_5000_3210, w_5000_3211, w_5000_3212, w_5000_3213, w_5000_3214, w_5000_3215, w_5000_3216, w_5000_3217, w_5000_3218, w_5000_3219, w_5000_3220, w_5000_3221, w_5000_3222, w_5000_3223, w_5000_3224, w_5000_3225, w_5000_3226, w_5000_3227, w_5000_3228, w_5000_3229, w_5000_3230, w_5000_3231, w_5000_3232, w_5000_3233, w_5000_3234, w_5000_3235, w_5000_3236, w_5000_3237, w_5000_3238, w_5000_3239, w_5000_3240, w_5000_3241, w_5000_3242, w_5000_3243, w_5000_3244, w_5000_3245, w_5000_3246, w_5000_3247, w_5000_3248, w_5000_3249, w_5000_3250, w_5000_3251, w_5000_3252, w_5000_3253, w_5000_3254, w_5000_3255, w_5000_3256, w_5000_3257, w_5000_3258, w_5000_3259, w_5000_3260, w_5000_3261, w_5000_3262, w_5000_3263, w_5000_3264, w_5000_3265, w_5000_3266, w_5000_3267, w_5000_3268, w_5000_3269, w_5000_3270, w_5000_3271, w_5000_3272, w_5000_3273, w_5000_3274, w_5000_3275, w_5000_3276, w_5000_3277, w_5000_3278, w_5000_3279, w_5000_3280, w_5000_3281, w_5000_3282, w_5000_3283, w_5000_3284, w_5000_3285, w_5000_3286, w_5000_3287, w_5000_3288, w_5000_3289, w_5000_3290, w_5000_3291, w_5000_3292, w_5000_3293, w_5000_3294, w_5000_3295, w_5000_3296, w_5000_3297, w_5000_3298, w_5000_3299, w_5000_3300, w_5000_3301, w_5000_3302, w_5000_3303, w_5000_3304, w_5000_3305, w_5000_3306, w_5000_3307, w_5000_3308, w_5000_3309, w_5000_3310, w_5000_3311, w_5000_3312, w_5000_3313, w_5000_3314, w_5000_3315, w_5000_3316, w_5000_3317, w_5000_3318, w_5000_3319, w_5000_3320, w_5000_3321, w_5000_3322, w_5000_3323, w_5000_3324, w_5000_3325, w_5000_3326, w_5000_3327, w_5000_3328, w_5000_3329, w_5000_3330, w_5000_3331, w_5000_3332, w_5000_3333, w_5000_3334, w_5000_3335, w_5000_3336, w_5000_3337, w_5000_3338, w_5000_3339, w_5000_3340, w_5000_3341, w_5000_3342, w_5000_3343, w_5000_3344, w_5000_3345, w_5000_3346, w_5000_3347, w_5000_3348, w_5000_3349, w_5000_3350, w_5000_3351, w_5000_3352, w_5000_3353, w_5000_3354, w_5000_3355, w_5000_3356, w_5000_3357, w_5000_3358, w_5000_3359, w_5000_3360, w_5000_3361, w_5000_3362, w_5000_3363, w_5000_3364, w_5000_3365, w_5000_3366, w_5000_3367, w_5000_3368, w_5000_3369, w_5000_3370, w_5000_3371, w_5000_3372, w_5000_3373, w_5000_3374, w_5000_3375, w_5000_3376, w_5000_3377, w_5000_3378, w_5000_3379, w_5000_3380, w_5000_3381, w_5000_3382, w_5000_3383, w_5000_3384, w_5000_3385, w_5000_3386, w_5000_3387, w_5000_3388, w_5000_3389, w_5000_3390, w_5000_3391, w_5000_3392, w_5000_3393, w_5000_3394, w_5000_3395, w_5000_3396, w_5000_3397, w_5000_3398, w_5000_3399, w_5000_3400, w_5000_3401, w_5000_3402, w_5000_3403, w_5000_3404, w_5000_3405, w_5000_3406, w_5000_3407, w_5000_3408, w_5000_3409, w_5000_3410, w_5000_3411, w_5000_3412, w_5000_3413, w_5000_3414, w_5000_3415, w_5000_3416, w_5000_3417, w_5000_3418, w_5000_3419, w_5000_3420, w_5000_3421, w_5000_3422, w_5000_3423, w_5000_3424, w_5000_3425, w_5000_3426, w_5000_3427, w_5000_3428, w_5000_3429, w_5000_3430, w_5000_3431, w_5000_3432, w_5000_3433, w_5000_3434, w_5000_3435, w_5000_3436, w_5000_3437, w_5000_3438, w_5000_3439, w_5000_3440, w_5000_3441, w_5000_3442, w_5000_3443, w_5000_3444, w_5000_3445, w_5000_3446, w_5000_3447, w_5000_3448, w_5000_3449, w_5000_3450, w_5000_3451, w_5000_3452, w_5000_3453, w_5000_3454, w_5000_3455, w_5000_3456, w_5000_3457, w_5000_3458, w_5000_3459, w_5000_3460, w_5000_3461, w_5000_3462, w_5000_3463, w_5000_3464, w_5000_3465, w_5000_3466, w_5000_3467, w_5000_3468, w_5000_3469, w_5000_3470, w_5000_3471, w_5000_3472, w_5000_3473, w_5000_3474, w_5000_3475, w_5000_3476, w_5000_3477, w_5000_3478, w_5000_3479, w_5000_3480, w_5000_3481, w_5000_3482, w_5000_3483, w_5000_3484, w_5000_3485, w_5000_3486, w_5000_3487, w_5000_3488, w_5000_3489, w_5000_3490, w_5000_3491, w_5000_3492, w_5000_3493, w_5000_3494, w_5000_3495, w_5000_3496, w_5000_3497, w_5000_3498, w_5000_3499, w_5000_3500, w_5000_3501, w_5000_3502, w_5000_3503, w_5000_3504, w_5000_3505, w_5000_3506, w_5000_3507, w_5000_3508, w_5000_3509, w_5000_3510, w_5000_3511, w_5000_3512, w_5000_3513, w_5000_3514, w_5000_3515, w_5000_3516, w_5000_3517, w_5000_3518, w_5000_3519, w_5000_3520, w_5000_3521, w_5000_3522, w_5000_3523, w_5000_3524, w_5000_3525, w_5000_3526, w_5000_3527, w_5000_3528, w_5000_3529, w_5000_3530, w_5000_3531, w_5000_3532, w_5000_3533, w_5000_3534, w_5000_3535, w_5000_3536, w_5000_3537, w_5000_3538, w_5000_3539, w_5000_3540, w_5000_3541, w_5000_3542, w_5000_3543, w_5000_3544, w_5000_3545, w_5000_3546, w_5000_3547, w_5000_3548, w_5000_3549, w_5000_3550, w_5000_3551, w_5000_3552, w_5000_3553, w_5000_3554, w_5000_3555, w_5000_3556, w_5000_3557, w_5000_3558, w_5000_3559, w_5000_3560, w_5000_3561, w_5000_3562, w_5000_3563, w_5000_3564, w_5000_3565, w_5000_3566, w_5000_3567, w_5000_3568, w_5000_3569, w_5000_3570, w_5000_3571, w_5000_3572, w_5000_3573, w_5000_3574, w_5000_3575, w_5000_3576, w_5000_3577, w_5000_3578, w_5000_3579, w_5000_3580, w_5000_3581, w_5000_3582, w_5000_3583, w_5000_3584, w_5000_3585, w_5000_3586, w_5000_3587, w_5000_3588, w_5000_3589, w_5000_3590, w_5000_3591, w_5000_3592, w_5000_3593, w_5000_3594, w_5000_3595, w_5000_3596, w_5000_3597, w_5000_3598, w_5000_3599, w_5000_3600, w_5000_3601, w_5000_3602, w_5000_3603, w_5000_3604, w_5000_3605, w_5000_3606, w_5000_3607, w_5000_3608, w_5000_3609, w_5000_3610, w_5000_3611, w_5000_3612, w_5000_3613, w_5000_3614, w_5000_3615, w_5000_3616, w_5000_3617, w_5000_3618, w_5000_3619, w_5000_3620, w_5000_3621, w_5000_3622, w_5000_3623, w_5000_3624, w_5000_3625, w_5000_3626, w_5000_3627, w_5000_3628, w_5000_3629, w_5000_3630, w_5000_3631, w_5000_3632, w_5000_3633, w_5000_3634, w_5000_3635, w_5000_3636, w_5000_3637, w_5000_3638, w_5000_3639, w_5000_3640, w_5000_3641, w_5000_3642, w_5000_3643, w_5000_3644, w_5000_3645, w_5000_3646, w_5000_3647, w_5000_3648, w_5000_3649, w_5000_3650, w_5000_3651, w_5000_3652, w_5000_3653, w_5000_3654, w_5000_3655, w_5000_3656, w_5000_3657, w_5000_3658, w_5000_3659, w_5000_3660, w_5000_3661, w_5000_3662, w_5000_3663, w_5000_3664, w_5000_3665, w_5000_3666, w_5000_3667, w_5000_3668, w_5000_3669, w_5000_3670, w_5000_3671, w_5000_3672, w_5000_3673, w_5000_3674, w_5000_3675, w_5000_3676, w_5000_3677, w_5000_3678, w_5000_3679, w_5000_3680, w_5000_3681, w_5000_3682, w_5000_3683, w_5000_3684, w_5000_3685, w_5000_3686, w_5000_3687, w_5000_3688, w_5000_3689, w_5000_3690, w_5000_3691, w_5000_3692, w_5000_3693, w_5000_3694, w_5000_3695, w_5000_3696, w_5000_3697, w_5000_3698, w_5000_3699, w_5000_3700, w_5000_3701, w_5000_3702, w_5000_3703, w_5000_3704, w_5000_3705, w_5000_3706, w_5000_3707, w_5000_3708, w_5000_3709, w_5000_3710, w_5000_3711, w_5000_3712, w_5000_3713, w_5000_3714, w_5000_3715, w_5000_3716, w_5000_3717, w_5000_3718, w_5000_3719, w_5000_3720, w_5000_3721, w_5000_3722, w_5000_3723, w_5000_3724, w_5000_3725, w_5000_3726, w_5000_3727, w_5000_3728, w_5000_3729, w_5000_3730, w_5000_3731, w_5000_3732, w_5000_3733, w_5000_3734, w_5000_3735, w_5000_3736, w_5000_3737, w_5000_3738, w_5000_3739, w_5000_3740, w_5000_3741, w_5000_3742, w_5000_3743, w_5000_3744, w_5000_3745, w_5000_3746, w_5000_3747, w_5000_3748, w_5000_3749, w_5000_3750, w_5000_3751, w_5000_3752, w_5000_3753, w_5000_3754, w_5000_3755, w_5000_3756, w_5000_3757, w_5000_3758, w_5000_3759, w_5000_3760, w_5000_3761, w_5000_3762, w_5000_3763, w_5000_3764, w_5000_3765, w_5000_3766, w_5000_3767, w_5000_3768, w_5000_3769, w_5000_3770, w_5000_3771, w_5000_3772, w_5000_3773, w_5000_3774, w_5000_3775, w_5000_3776, w_5000_3777, w_5000_3778, w_5000_3779, w_5000_3780, w_5000_3781, w_5000_3782, w_5000_3783, w_5000_3784, w_5000_3785, w_5000_3786, w_5000_3787, w_5000_3788, w_5000_3789, w_5000_3790, w_5000_3791, w_5000_3792, w_5000_3793, w_5000_3794, w_5000_3795, w_5000_3796, w_5000_3797, w_5000_3798, w_5000_3799, w_5000_3800, w_5000_3801, w_5000_3802, w_5000_3803, w_5000_3804, w_5000_3805, w_5000_3806, w_5000_3807, w_5000_3808, w_5000_3809, w_5000_3810, w_5000_3811, w_5000_3812, w_5000_3813, w_5000_3814, w_5000_3815, w_5000_3816, w_5000_3817, w_5000_3818, w_5000_3819, w_5000_3820, w_5000_3821, w_5000_3822, w_5000_3823, w_5000_3824, w_5000_3825, w_5000_3826, w_5000_3827, w_5000_3828, w_5000_3829, w_5000_3830, w_5000_3831, w_5000_3832, w_5000_3833, w_5000_3834, w_5000_3835, w_5000_3836, w_5000_3837, w_5000_3838, w_5000_3839, w_5000_3840, w_5000_3841, w_5000_3842, w_5000_3843, w_5000_3844, w_5000_3845, w_5000_3846, w_5000_3847, w_5000_3848, w_5000_3849, w_5000_3850, w_5000_3851, w_5000_3852, w_5000_3853, w_5000_3854, w_5000_3855, w_5000_3856, w_5000_3857, w_5000_3858, w_5000_3859, w_5000_3860, w_5000_3861, w_5000_3862, w_5000_3863, w_5000_3864, w_5000_3865, w_5000_3866, w_5000_3867, w_5000_3868, w_5000_3869, w_5000_3870, w_5000_3871, w_5000_3872, w_5000_3873, w_5000_3874, w_5000_3875, w_5000_3876, w_5000_3877, w_5000_3878, w_5000_3879, w_5000_3880, w_5000_3881, w_5000_3882, w_5000_3883, w_5000_3884, w_5000_3885, w_5000_3886, w_5000_3887, w_5000_3888, w_5000_3889, w_5000_3890, w_5000_3891, w_5000_3892, w_5000_3893, w_5000_3894, w_5000_3895, w_5000_3896, w_5000_3897, w_5000_3898, w_5000_3899, w_5000_3900, w_5000_3901, w_5000_3902, w_5000_3903, w_5000_3904, w_5000_3905, w_5000_3906, w_5000_3907, w_5000_3908, w_5000_3909, w_5000_3910, w_5000_3911, w_5000_3912, w_5000_3913, w_5000_3914, w_5000_3915, w_5000_3916, w_5000_3917, w_5000_3918, w_5000_3919, w_5000_3920, w_5000_3921, w_5000_3922, w_5000_3923, w_5000_3924, w_5000_3925, w_5000_3926, w_5000_3927, w_5000_3928, w_5000_3929, w_5000_3930, w_5000_3931, w_5000_3932, w_5000_3933, w_5000_3934, w_5000_3935, w_5000_3936, w_5000_3937, w_5000_3938, w_5000_3939, w_5000_3940, w_5000_3941, w_5000_3942, w_5000_3943, w_5000_3944, w_5000_3945, w_5000_3946, w_5000_3947, w_5000_3948, w_5000_3949, w_5000_3950, w_5000_3951, w_5000_3952, w_5000_3953, w_5000_3954, w_5000_3955, w_5000_3956, w_5000_3957, w_5000_3958, w_5000_3959, w_5000_3960, w_5000_3961, w_5000_3962, w_5000_3963, w_5000_3964, w_5000_3965, w_5000_3966, w_5000_3967, w_5000_3968, w_5000_3969, w_5000_3970, w_5000_3971, w_5000_3972, w_5000_3973, w_5000_3974, w_5000_3975, w_5000_3976, w_5000_3977, w_5000_3978, w_5000_3979, w_5000_3980, w_5000_3981, w_5000_3982, w_5000_3983, w_5000_3984, w_5000_3985, w_5000_3986, w_5000_3987, w_5000_3988, w_5000_3989, w_5000_3990, w_5000_3991, w_5000_3992, w_5000_3993, w_5000_3994, w_5000_3995, w_5000_3996, w_5000_3997, w_5000_3998, w_5000_3999, w_5000_4000, w_5000_4001, w_5000_4002, w_5000_4003, w_5000_4004, w_5000_4005, w_5000_4006, w_5000_4007, w_5000_4008, w_5000_4009, w_5000_4010, w_5000_4011, w_5000_4012, w_5000_4013, w_5000_4014, w_5000_4015, w_5000_4016, w_5000_4017, w_5000_4018, w_5000_4019, w_5000_4020, w_5000_4021, w_5000_4022, w_5000_4023, w_5000_4024, w_5000_4025, w_5000_4026, w_5000_4027, w_5000_4028, w_5000_4029, w_5000_4030, w_5000_4031, w_5000_4032, w_5000_4033, w_5000_4034, w_5000_4035, w_5000_4036, w_5000_4037, w_5000_4038, w_5000_4039, w_5000_4040, w_5000_4041, w_5000_4042, w_5000_4043, w_5000_4044, w_5000_4045, w_5000_4046, w_5000_4047, w_5000_4048, w_5000_4049, w_5000_4050, w_5000_4051, w_5000_4052, w_5000_4053, w_5000_4054, w_5000_4055, w_5000_4056, w_5000_4057, w_5000_4058, w_5000_4059, w_5000_4060, w_5000_4061, w_5000_4062, w_5000_4063, w_5000_4064, w_5000_4065, w_5000_4066, w_5000_4067, w_5000_4068, w_5000_4069, w_5000_4070, w_5000_4071, w_5000_4072, w_5000_4073, w_5000_4074, w_5000_4075, w_5000_4076, w_5000_4077, w_5000_4078, w_5000_4079, w_5000_4080, w_5000_4081, w_5000_4082, w_5000_4083, w_5000_4084, w_5000_4085, w_5000_4086, w_5000_4087, w_5000_4088, w_5000_4089, w_5000_4090, w_5000_4091, w_5000_4092, w_5000_4093, w_5000_4094, w_5000_4095, w_5000_4096, w_5000_4097, w_5000_4098, w_5000_4099, w_5000_4100, w_5000_4101, w_5000_4102, w_5000_4103, w_5000_4104, w_5000_4105, w_5000_4106, w_5000_4107, w_5000_4108, w_5000_4109, w_5000_4110, w_5000_4111, w_5000_4112, w_5000_4113, w_5000_4114, w_5000_4115, w_5000_4116, w_5000_4117, w_5000_4118, w_5000_4119, w_5000_4120, w_5000_4121, w_5000_4122, w_5000_4123, w_5000_4124, w_5000_4125, w_5000_4126, w_5000_4127, w_5000_4128, w_5000_4129, w_5000_4130, w_5000_4131, w_5000_4132, w_5000_4133, w_5000_4134, w_5000_4135, w_5000_4136, w_5000_4137, w_5000_4138, w_5000_4139, w_5000_4140, w_5000_4141, w_5000_4142, w_5000_4143, w_5000_4144, w_5000_4145, w_5000_4146, w_5000_4147, w_5000_4148, w_5000_4149, w_5000_4150, w_5000_4151, w_5000_4152, w_5000_4153, w_5000_4154, w_5000_4155, w_5000_4156, w_5000_4157, w_5000_4158, w_5000_4159, w_5000_4160, w_5000_4161, w_5000_4162, w_5000_4163, w_5000_4164, w_5000_4165, w_5000_4166, w_5000_4167, w_5000_4168, w_5000_4169, w_5000_4170, w_5000_4171, w_5000_4172, w_5000_4173, w_5000_4174, w_5000_4175, w_5000_4176, w_5000_4177, w_5000_4178, w_5000_4179, w_5000_4180, w_5000_4181, w_5000_4182, w_5000_4183, w_5000_4184, w_5000_4185, w_5000_4186, w_5000_4187, w_5000_4188, w_5000_4189, w_5000_4190, w_5000_4191, w_5000_4192, w_5000_4193, w_5000_4194, w_5000_4195, w_5000_4196, w_5000_4197, w_5000_4198, w_5000_4199, w_5000_4200, w_5000_4201, w_5000_4202, w_5000_4203, w_5000_4204, w_5000_4205, w_5000_4206, w_5000_4207, w_5000_4208, w_5000_4209, w_5000_4210, w_5000_4211, w_5000_4212, w_5000_4213, w_5000_4214, w_5000_4215, w_5000_4216, w_5000_4217, w_5000_4218, w_5000_4219, w_5000_4220, w_5000_4221, w_5000_4222, w_5000_4223, w_5000_4224, w_5000_4225, w_5000_4226, w_5000_4227, w_5000_4228, w_5000_4229, w_5000_4230, w_5000_4231, w_5000_4232, w_5000_4233, w_5000_4234, w_5000_4235, w_5000_4236, w_5000_4237, w_5000_4238, w_5000_4239, w_5000_4240, w_5000_4241, w_5000_4242, w_5000_4243, w_5000_4244, w_5000_4245;
  wire w_000_000, w_000_001, w_000_002, w_000_003, w_000_004, w_000_005, w_000_006, w_000_007, w_000_008, w_000_009, w_000_010, w_000_011, w_000_012, w_000_013, w_000_014, w_000_015, w_000_016, w_000_017, w_000_018, w_000_019, w_000_020, w_000_021, w_000_022, w_000_023, w_000_024, w_000_025, w_000_026, w_000_027, w_000_028, w_000_029, w_000_030, w_000_031, w_000_032, w_000_033, w_000_034, w_000_035, w_000_036, w_000_037, w_000_038, w_000_039, w_000_040, w_000_041, w_000_042, w_000_043, w_000_044, w_000_045, w_000_046, w_000_047, w_000_048, w_000_049, w_000_050, w_000_051, w_000_052, w_000_053, w_000_054, w_000_055, w_000_056, w_000_057, w_000_058, w_000_059, w_000_060, w_000_061, w_000_062, w_000_063, w_000_064, w_000_065, w_000_066, w_000_067, w_000_068, w_000_069, w_000_070, w_000_071, w_000_072, w_000_073, w_000_074, w_000_075, w_000_076, w_000_077, w_000_078, w_000_079, w_000_080, w_000_081, w_000_082, w_000_083, w_000_084, w_000_085, w_000_086, w_000_087, w_000_088, w_000_089, w_000_090, w_000_091, w_000_092, w_000_093, w_000_094, w_000_095, w_000_096, w_000_097, w_000_098, w_000_099, w_000_100, w_000_101, w_000_102, w_000_103, w_000_104, w_000_105, w_000_106, w_000_107, w_000_108, w_000_109, w_000_110, w_000_111, w_000_112, w_000_113, w_000_114, w_000_115, w_000_116, w_000_117, w_000_118, w_000_119, w_000_120, w_000_121, w_000_122, w_000_123, w_000_124, w_000_125, w_000_126, w_000_127, w_000_128, w_000_129, w_000_130, w_000_131, w_000_132, w_000_133, w_000_134, w_000_135, w_000_136, w_000_137, w_000_138, w_000_139, w_000_140, w_000_141, w_000_142, w_000_143, w_000_144, w_000_145, w_000_146, w_000_147, w_000_148, w_000_149, w_000_150, w_000_151, w_000_152, w_000_153, w_000_154, w_000_155, w_000_156, w_000_157, w_000_158, w_000_159, w_000_160, w_000_161, w_000_162, w_000_163, w_000_164, w_000_165, w_000_166, w_000_167, w_000_168, w_000_169, w_000_170, w_000_171, w_000_172, w_000_173, w_000_174, w_000_175, w_000_176, w_000_177, w_000_178, w_000_179, w_000_180, w_000_181, w_000_182, w_000_183, w_000_184, w_000_185, w_000_186, w_000_187, w_000_188, w_000_189, w_000_190, w_000_191, w_000_192, w_000_193, w_000_194, w_000_195, w_000_196, w_000_197, w_000_198, w_000_199, w_000_200, w_000_201, w_000_202, w_000_203, w_000_204, w_000_205, w_000_206, w_000_207, w_000_208, w_000_209, w_000_210, w_000_211, w_000_212, w_000_213, w_000_214, w_000_215, w_000_216, w_000_217, w_000_218, w_000_219, w_000_220, w_000_221, w_000_222, w_000_223, w_000_224, w_000_225, w_000_226, w_000_227, w_000_228, w_000_229, w_000_230, w_000_231, w_000_232, w_000_233, w_000_234, w_000_235, w_000_236, w_000_237, w_000_238, w_000_239, w_000_240, w_000_241, w_000_242, w_000_243, w_000_244, w_000_245, w_000_246, w_000_247, w_000_248, w_000_249, w_000_250, w_000_251, w_000_252, w_000_253, w_000_254, w_000_255, w_000_256, w_000_257, w_000_258, w_000_259, w_000_260, w_000_261, w_000_262, w_000_263, w_000_264, w_000_265, w_000_266, w_000_267, w_000_268, w_000_269, w_000_270, w_000_271, w_000_272, w_000_273, w_000_274, w_000_275, w_000_276, w_000_277, w_000_278, w_000_279, w_000_280, w_000_281, w_000_282, w_000_283, w_000_284, w_000_285, w_000_286, w_000_287, w_000_288, w_000_289, w_000_290, w_000_291, w_000_292, w_000_293, w_000_294, w_000_295, w_000_296, w_000_297, w_000_298, w_000_299, w_000_300, w_000_301, w_000_302, w_000_303, w_000_304, w_000_305, w_000_306, w_000_307, w_000_308, w_000_309, w_000_310, w_000_311, w_000_312, w_000_313, w_000_314, w_000_315, w_000_316, w_000_317, w_000_318, w_000_319, w_000_320, w_000_321, w_000_322, w_000_323, w_000_324, w_000_325, w_000_326, w_000_327, w_000_328, w_000_329, w_000_330, w_000_331, w_000_332, w_000_333, w_000_334, w_000_335, w_000_336, w_000_337, w_000_338, w_000_339, w_000_340, w_000_341, w_000_342, w_000_343, w_000_344, w_000_345, w_000_346, w_000_347, w_000_348, w_000_349, w_000_350, w_000_351, w_000_352, w_000_353, w_000_354, w_000_355, w_000_356, w_000_357, w_000_358, w_000_359, w_000_360, w_000_361, w_000_362, w_000_363, w_000_364, w_000_365, w_000_366, w_000_367, w_000_368, w_000_369, w_000_370, w_000_371, w_000_372, w_000_373, w_000_374, w_000_375, w_000_376, w_000_377, w_000_378, w_000_379, w_000_380, w_000_381, w_000_382, w_000_383, w_000_384, w_000_385, w_000_386, w_000_387, w_000_388, w_000_389, w_000_390, w_000_391, w_000_392, w_000_393, w_000_394, w_000_395, w_000_396, w_000_397, w_000_398, w_000_399, w_000_400, w_000_401, w_000_402, w_000_403, w_000_404, w_000_405, w_000_406, w_000_407, w_000_408, w_000_409, w_000_410, w_000_411, w_000_412, w_000_413, w_000_414, w_000_415, w_000_416, w_000_417, w_000_418, w_000_419, w_000_420, w_000_421, w_000_422, w_000_423, w_000_424, w_000_425, w_000_426, w_000_427, w_000_428, w_000_429, w_000_430, w_000_431, w_000_432, w_000_433, w_000_434, w_000_435, w_000_436, w_000_437, w_000_438, w_000_439, w_000_440, w_000_441, w_000_442, w_000_443, w_000_444, w_000_445, w_000_446, w_000_447, w_000_448, w_000_449, w_000_450, w_000_451, w_000_452, w_000_453, w_000_454, w_000_455, w_000_456, w_000_457, w_000_458, w_000_459, w_000_460, w_000_461, w_000_462, w_000_463, w_000_464, w_000_465, w_000_466, w_000_467, w_000_468, w_000_469, w_000_470, w_000_471, w_000_472, w_000_473, w_000_474, w_000_475, w_000_476, w_000_477, w_000_478, w_000_479, w_000_480, w_000_481, w_000_482, w_000_483, w_000_484, w_000_485, w_000_486, w_000_487, w_000_488, w_000_489, w_000_490, w_000_491, w_000_492, w_000_493, w_000_494, w_000_495, w_000_496, w_000_497, w_000_498, w_000_499, w_000_500, w_000_501, w_000_502, w_000_503, w_000_504, w_000_505, w_000_506, w_000_507, w_000_508, w_000_509, w_000_510, w_000_511, w_000_512, w_000_513, w_000_514, w_000_515, w_000_516, w_000_517, w_000_518, w_000_519, w_000_520, w_000_521, w_000_522, w_000_523, w_000_524, w_000_525, w_000_526, w_000_527, w_000_528, w_000_529, w_000_530, w_000_531, w_000_532, w_000_533, w_000_534, w_000_535, w_000_536, w_000_537, w_000_538, w_000_539, w_000_540, w_000_541, w_000_542, w_000_543, w_000_544, w_000_545, w_000_546, w_000_547, w_000_548, w_000_549, w_000_550, w_000_551, w_000_552, w_000_553, w_000_554, w_000_555, w_000_556, w_000_557, w_000_558, w_000_559, w_000_560, w_000_561, w_000_562, w_000_563, w_000_564, w_000_565, w_000_566, w_000_567, w_000_568, w_000_569, w_000_570, w_000_571, w_000_572, w_000_573, w_000_574, w_000_575, w_000_576, w_000_577, w_000_578, w_000_579, w_000_580, w_000_581, w_000_582, w_000_583, w_000_584, w_000_585, w_000_586, w_000_587, w_000_588, w_000_589, w_000_590, w_000_591, w_000_592, w_000_593, w_000_594, w_000_595, w_000_596, w_000_597, w_000_598, w_000_599, w_000_600, w_000_601, w_000_602, w_000_603, w_000_604, w_000_605, w_000_606, w_000_607, w_000_608, w_000_609, w_000_610, w_000_611, w_000_612, w_000_613, w_000_614, w_000_615, w_000_616, w_000_617, w_000_618, w_000_619, w_000_620, w_000_621, w_000_622, w_000_623, w_000_624, w_000_625, w_000_626, w_000_627, w_000_628, w_000_629, w_000_630, w_000_631, w_000_632, w_000_633, w_000_634, w_000_635, w_000_636, w_000_637, w_000_638, w_000_639, w_000_640, w_000_641, w_000_642, w_000_643, w_000_644, w_000_645, w_000_646, w_000_647, w_000_648, w_000_649, w_000_650, w_000_651, w_000_652, w_000_653, w_000_654, w_000_655, w_000_656, w_000_657, w_000_658, w_000_659, w_000_660, w_000_661, w_000_662, w_000_663, w_000_664, w_000_665, w_000_666, w_000_667, w_000_668, w_000_669, w_000_670, w_000_671, w_000_672, w_000_673, w_000_674, w_000_675, w_000_676, w_000_677, w_000_678, w_000_679, w_000_680, w_000_681, w_000_682, w_000_683, w_000_684, w_000_685, w_000_686, w_000_687, w_000_688, w_000_689, w_000_690, w_000_691, w_000_692, w_000_693, w_000_694, w_000_695, w_000_696, w_000_697, w_000_698, w_000_699, w_000_700, w_000_701, w_000_702, w_000_703, w_000_704, w_000_705, w_000_706, w_000_707, w_000_708, w_000_709, w_000_710, w_000_711, w_000_712, w_000_713, w_000_714, w_000_715, w_000_716, w_000_717, w_000_718, w_000_719, w_000_720, w_000_721, w_000_722, w_000_723, w_000_724, w_000_725, w_000_726, w_000_727, w_000_728, w_000_729, w_000_730, w_000_731, w_000_732, w_000_733, w_000_734, w_000_735, w_000_736, w_000_737, w_000_738, w_000_739, w_000_740, w_000_741, w_000_742, w_000_743, w_000_744, w_000_745, w_000_746, w_000_747, w_000_748, w_000_749, w_000_750, w_000_751, w_000_752, w_000_753, w_000_754, w_000_755, w_000_756, w_000_757, w_000_758, w_000_759, w_000_760, w_000_761, w_000_762, w_000_763, w_000_764, w_000_765, w_000_766, w_000_767, w_000_768, w_000_769, w_000_770, w_000_771, w_000_772, w_000_773, w_000_774, w_000_775, w_000_776, w_000_777, w_000_778, w_000_779, w_000_780, w_000_781, w_000_782, w_000_783, w_000_784, w_000_785, w_000_786, w_000_787, w_000_788, w_000_789, w_000_790, w_000_791, w_000_792, w_000_793, w_000_794, w_000_795, w_000_796, w_000_797, w_000_798, w_000_799, w_000_800, w_000_801, w_000_802, w_000_803, w_000_804, w_000_805, w_000_806, w_000_807, w_000_808, w_000_809, w_000_810, w_000_811, w_000_812, w_000_813, w_000_814, w_000_815, w_000_816, w_000_817, w_000_818, w_000_819, w_000_820, w_000_821, w_000_822, w_000_823, w_000_824, w_000_825, w_000_826, w_000_827, w_000_828, w_000_829, w_000_830, w_000_831, w_000_832, w_000_833, w_000_834, w_000_835, w_000_836, w_000_837, w_000_838, w_000_839, w_000_840, w_000_841, w_000_842, w_000_843, w_000_844, w_000_845, w_000_846, w_000_847, w_000_848, w_000_849, w_000_850, w_000_851, w_000_852, w_000_853, w_000_854, w_000_855, w_000_856, w_000_857, w_000_858, w_000_859, w_000_860, w_000_861, w_000_862, w_000_863, w_000_864, w_000_865, w_000_866, w_000_867, w_000_868, w_000_869, w_000_870, w_000_871, w_000_872, w_000_873, w_000_874, w_000_875, w_000_876, w_000_877, w_000_878, w_000_879, w_000_880, w_000_881, w_000_882, w_000_883, w_000_884, w_000_885, w_000_886, w_000_887, w_000_888, w_000_889, w_000_890, w_000_891, w_000_892, w_000_893, w_000_894, w_000_895, w_000_896, w_000_897, w_000_898, w_000_899, w_000_900, w_000_901, w_000_902, w_000_903, w_000_904, w_000_905, w_000_906, w_000_907, w_000_908, w_000_909, w_000_910, w_000_911, w_000_912, w_000_913, w_000_914, w_000_915, w_000_916, w_000_917, w_000_918, w_000_919, w_000_920, w_000_921, w_000_922, w_000_923, w_000_924, w_000_925, w_000_926, w_000_927, w_000_928, w_000_929, w_000_930, w_000_931, w_000_932, w_000_933, w_000_934, w_000_935, w_000_936, w_000_937, w_000_938, w_000_939, w_000_940, w_000_941, w_000_942, w_000_943, w_000_944, w_000_945, w_000_946, w_000_947, w_000_948, w_000_949, w_000_950, w_000_951, w_000_952, w_000_953, w_000_954, w_000_955, w_000_956, w_000_957, w_000_958, w_000_959, w_000_960, w_000_961, w_000_962, w_000_963, w_000_964, w_000_965, w_000_966, w_000_967, w_000_968, w_000_969, w_000_970, w_000_971, w_000_972, w_000_973, w_000_974, w_000_975, w_000_976, w_000_977, w_000_978, w_000_979, w_000_980, w_000_981, w_000_982, w_000_983, w_000_984, w_000_985, w_000_986, w_000_987, w_000_988, w_000_989, w_000_990, w_000_991, w_000_992, w_000_993, w_000_994, w_000_995, w_000_996, w_000_997, w_000_998, w_000_999, w_000_1000, w_000_1001, w_000_1002, w_000_1003, w_000_1004, w_000_1005, w_000_1006, w_000_1007, w_000_1008, w_000_1009, w_000_1010, w_000_1011, w_000_1012, w_000_1013, w_000_1014, w_000_1015, w_000_1016, w_000_1017, w_000_1018, w_000_1019, w_000_1020, w_000_1021, w_000_1022, w_000_1023, w_000_1024, w_000_1025, w_000_1026, w_000_1027, w_000_1028, w_000_1029, w_000_1030, w_000_1031, w_000_1032, w_000_1033, w_000_1034, w_000_1035, w_000_1036, w_000_1037, w_000_1038, w_000_1039, w_000_1040, w_000_1041, w_000_1042, w_000_1043, w_000_1044, w_000_1045, w_000_1046, w_000_1047, w_000_1048, w_000_1049, w_000_1050, w_000_1051, w_000_1052, w_000_1053, w_000_1054, w_000_1055, w_000_1056, w_000_1057, w_000_1058, w_000_1059, w_000_1060, w_000_1061, w_000_1062, w_000_1063, w_000_1064, w_000_1065, w_000_1066, w_000_1067, w_000_1068, w_000_1069, w_000_1070, w_000_1071, w_000_1072, w_000_1073, w_000_1074, w_000_1075, w_000_1076, w_000_1077, w_000_1078, w_000_1079, w_000_1080, w_000_1081, w_000_1082, w_000_1083, w_000_1084, w_000_1085, w_000_1086, w_000_1087, w_000_1088, w_000_1089, w_000_1090, w_000_1091, w_000_1092, w_000_1093, w_000_1094, w_000_1095, w_000_1096, w_000_1097, w_000_1098, w_000_1099, w_000_1100, w_000_1101, w_000_1102, w_000_1103, w_000_1104, w_000_1105, w_000_1106, w_000_1107, w_000_1108, w_000_1109, w_000_1110, w_000_1111, w_000_1112, w_000_1113, w_000_1114, w_000_1115, w_000_1116, w_000_1117, w_000_1118, w_000_1119, w_000_1120, w_000_1121, w_000_1122, w_000_1123, w_000_1124, w_000_1125, w_000_1126, w_000_1127, w_000_1128, w_000_1129, w_000_1130, w_000_1131, w_000_1132, w_000_1133, w_000_1134, w_000_1135, w_000_1136, w_000_1137, w_000_1138, w_000_1139, w_000_1140, w_000_1141, w_000_1142, w_000_1143, w_000_1144, w_000_1145, w_000_1146, w_000_1147, w_000_1148, w_000_1149, w_000_1150, w_000_1151, w_000_1152, w_000_1153, w_000_1154, w_000_1155, w_000_1156, w_000_1157, w_000_1158, w_000_1159, w_000_1160, w_000_1161, w_000_1162, w_000_1163, w_000_1164, w_000_1165, w_000_1166, w_000_1167, w_000_1168, w_000_1169, w_000_1170, w_000_1171, w_000_1172, w_000_1173, w_000_1174, w_000_1175, w_000_1176, w_000_1177, w_000_1178, w_000_1179, w_000_1180, w_000_1181, w_000_1182, w_000_1183, w_000_1184, w_000_1185, w_000_1186, w_000_1187, w_000_1188, w_000_1189, w_000_1190, w_000_1191, w_000_1192, w_000_1193, w_000_1194, w_000_1195, w_000_1196, w_000_1197, w_000_1198, w_000_1199, w_000_1200, w_000_1201, w_000_1202, w_000_1203, w_000_1204, w_000_1205, w_000_1206, w_000_1207, w_000_1208, w_000_1209, w_000_1210, w_000_1211, w_000_1212, w_000_1213, w_000_1214, w_000_1215, w_000_1216, w_000_1217, w_000_1218, w_000_1219, w_000_1220, w_000_1221, w_000_1222, w_000_1223, w_000_1224, w_000_1225, w_000_1226, w_000_1227, w_000_1228, w_000_1229, w_000_1230, w_000_1231, w_000_1232, w_000_1233, w_000_1234, w_000_1235, w_000_1236, w_000_1237, w_000_1238, w_000_1239, w_000_1240, w_000_1241, w_000_1242, w_000_1243, w_000_1244, w_000_1245, w_000_1246, w_000_1247, w_000_1248, w_000_1249, w_000_1250, w_000_1251, w_000_1252, w_000_1253, w_000_1254, w_000_1255, w_000_1256, w_000_1257, w_000_1258, w_000_1259, w_000_1260, w_000_1261, w_000_1262, w_000_1263, w_000_1264, w_000_1265, w_000_1266, w_000_1267, w_000_1268, w_000_1269, w_000_1270, w_000_1271, w_000_1272, w_000_1273, w_000_1274, w_000_1275, w_000_1276, w_000_1277, w_000_1278, w_000_1279, w_000_1280, w_000_1281, w_000_1282, w_000_1283, w_000_1284, w_000_1285, w_000_1286, w_000_1287, w_000_1288, w_000_1289, w_000_1290, w_000_1291, w_000_1292, w_000_1293, w_000_1294, w_000_1295, w_000_1296, w_000_1297, w_000_1298, w_000_1299, w_000_1300, w_000_1301, w_000_1302, w_000_1303, w_000_1304, w_000_1305, w_000_1306, w_000_1307, w_000_1308, w_000_1309, w_000_1310, w_000_1311, w_000_1312, w_000_1313, w_000_1314, w_000_1315, w_000_1316, w_000_1317, w_000_1318, w_000_1319, w_000_1320, w_000_1321, w_000_1322, w_000_1323, w_000_1324, w_000_1325, w_000_1326, w_000_1327, w_000_1328, w_000_1329, w_000_1330, w_000_1331, w_000_1332, w_000_1333, w_000_1334, w_000_1335, w_000_1336, w_000_1337, w_000_1338, w_000_1339, w_000_1340, w_000_1341, w_000_1342, w_000_1343, w_000_1344, w_000_1345, w_000_1346, w_000_1347, w_000_1348, w_000_1349, w_000_1350, w_000_1351, w_000_1352, w_000_1353, w_000_1354, w_000_1355, w_000_1356, w_000_1357, w_000_1358, w_000_1359, w_000_1360, w_000_1361, w_000_1362, w_000_1363, w_000_1364, w_000_1365, w_000_1366, w_000_1367, w_000_1368, w_000_1369, w_000_1370, w_000_1371, w_000_1372, w_000_1373, w_000_1374, w_000_1375, w_000_1376, w_000_1377, w_000_1378, w_000_1379, w_000_1380, w_000_1381, w_000_1382, w_000_1383, w_000_1384, w_000_1385, w_000_1386, w_000_1387, w_000_1388, w_000_1389, w_000_1390, w_000_1391, w_000_1392, w_000_1393, w_000_1394, w_000_1395, w_000_1396, w_000_1397, w_000_1398, w_000_1399, w_000_1400, w_000_1401, w_000_1402, w_000_1403, w_000_1404, w_000_1405, w_000_1406, w_000_1407, w_000_1408, w_000_1409, w_000_1410, w_000_1411, w_000_1412, w_000_1413, w_000_1414, w_000_1415, w_000_1416, w_000_1417, w_000_1418, w_000_1419, w_000_1420, w_000_1421, w_000_1422, w_000_1423, w_000_1424, w_000_1425, w_000_1426, w_000_1427, w_000_1428, w_000_1429, w_000_1430, w_000_1431, w_000_1432, w_000_1433, w_000_1434, w_000_1435, w_000_1436, w_000_1437, w_000_1438, w_000_1439, w_000_1440, w_000_1441, w_000_1442, w_000_1443, w_000_1444, w_000_1445, w_000_1446, w_000_1447, w_000_1448, w_000_1449, w_000_1450, w_000_1451, w_000_1452, w_000_1453, w_000_1454, w_000_1455, w_000_1456, w_000_1457, w_000_1458, w_000_1459, w_000_1460, w_000_1461, w_000_1462, w_000_1463, w_000_1464, w_000_1465, w_000_1466, w_000_1467, w_000_1468, w_000_1469, w_000_1470, w_000_1471, w_000_1472, w_000_1473, w_000_1474, w_000_1475, w_000_1476, w_000_1477, w_000_1478, w_000_1479, w_000_1480, w_000_1481, w_000_1482, w_000_1483, w_000_1484, w_000_1485, w_000_1486, w_000_1487, w_000_1488, w_000_1489, w_000_1490, w_000_1491, w_000_1492, w_000_1493, w_000_1494, w_000_1495, w_000_1496, w_000_1497, w_000_1498, w_000_1499, w_000_1500, w_000_1501, w_000_1502, w_000_1503, w_000_1504, w_000_1505, w_000_1506, w_000_1507, w_000_1508, w_000_1509, w_000_1510, w_000_1511, w_000_1512, w_000_1513, w_000_1514, w_000_1515, w_000_1516, w_000_1517, w_000_1518, w_000_1519, w_000_1520, w_000_1521, w_000_1522, w_000_1523, w_000_1524, w_000_1525, w_000_1526, w_000_1527, w_000_1528, w_000_1529, w_000_1530, w_000_1531, w_000_1532, w_000_1533, w_000_1534, w_000_1535, w_000_1536, w_000_1537, w_000_1538, w_000_1539, w_000_1540, w_000_1541, w_000_1542, w_000_1543, w_000_1544, w_000_1545, w_000_1546, w_000_1547, w_000_1548, w_000_1549, w_000_1550, w_000_1551, w_000_1552, w_000_1553, w_000_1554, w_000_1555, w_000_1556, w_000_1557, w_000_1558, w_000_1559, w_000_1560, w_000_1561, w_000_1562, w_000_1563, w_000_1564, w_000_1565, w_000_1566, w_000_1567, w_000_1568, w_000_1569, w_000_1570, w_000_1571, w_000_1572, w_000_1573, w_000_1574, w_000_1575, w_000_1576, w_000_1577, w_000_1578, w_000_1579, w_000_1580, w_000_1581, w_000_1582, w_000_1583, w_000_1584, w_000_1585, w_000_1586, w_000_1587, w_000_1588, w_000_1589, w_000_1590, w_000_1591, w_000_1592, w_000_1593, w_000_1594, w_000_1595, w_000_1596, w_000_1597, w_000_1598, w_000_1599, w_000_1600, w_000_1601, w_000_1602, w_000_1603, w_000_1604, w_000_1605, w_000_1606, w_000_1607, w_000_1608, w_000_1609, w_000_1610, w_000_1611, w_000_1612, w_000_1613, w_000_1614, w_000_1615, w_000_1616, w_000_1617, w_000_1618, w_000_1619, w_000_1620, w_000_1621, w_000_1622, w_000_1623, w_000_1624, w_000_1625, w_000_1626, w_000_1627, w_000_1628, w_000_1629, w_000_1630, w_000_1631, w_000_1632, w_000_1633, w_000_1634, w_000_1635, w_000_1636, w_000_1637, w_000_1638, w_000_1639, w_000_1640, w_000_1641, w_000_1642, w_000_1643, w_000_1644, w_000_1645, w_000_1646, w_000_1647, w_000_1648, w_000_1649, w_000_1650, w_000_1651, w_000_1652, w_000_1653, w_000_1654, w_000_1655, w_000_1656, w_000_1657, w_000_1658, w_000_1659, w_000_1660, w_000_1661, w_000_1662, w_000_1663, w_000_1664, w_000_1665, w_000_1666, w_000_1667, w_000_1668, w_000_1669, w_000_1670, w_000_1671, w_000_1672, w_000_1673, w_000_1674, w_000_1675, w_000_1676, w_000_1677, w_000_1678, w_000_1679, w_000_1680, w_000_1681, w_000_1682, w_000_1683, w_000_1684, w_000_1685, w_000_1686, w_000_1687, w_000_1688, w_000_1689, w_000_1690, w_000_1691, w_000_1692, w_000_1693, w_000_1694, w_000_1695, w_000_1696, w_000_1697, w_000_1698, w_000_1699, w_000_1700, w_000_1701, w_000_1702, w_000_1703, w_000_1704, w_000_1705, w_000_1706, w_000_1707, w_000_1708, w_000_1709, w_000_1710, w_000_1711, w_000_1712, w_000_1713, w_000_1714, w_000_1715, w_000_1716, w_000_1717, w_000_1718, w_000_1719, w_000_1720, w_000_1721, w_000_1722, w_000_1723, w_000_1724, w_000_1725, w_000_1726, w_000_1727, w_000_1728, w_000_1729, w_000_1730, w_000_1731, w_000_1732, w_000_1733, w_000_1734, w_000_1735, w_000_1736, w_000_1737, w_000_1738, w_000_1739, w_000_1740, w_000_1741, w_000_1742, w_000_1743, w_000_1744, w_000_1745, w_000_1746, w_000_1747, w_000_1748, w_000_1749, w_000_1750, w_000_1751, w_000_1752, w_000_1753, w_000_1754, w_000_1755, w_000_1756, w_000_1757, w_000_1758, w_000_1759, w_000_1760, w_000_1761, w_000_1762, w_000_1763, w_000_1764, w_000_1765, w_000_1766, w_000_1767, w_000_1768, w_000_1769, w_000_1770, w_000_1771, w_000_1772, w_000_1773, w_000_1774, w_000_1775, w_000_1776, w_000_1777, w_000_1778, w_000_1779, w_000_1780, w_000_1781, w_000_1782, w_000_1783, w_000_1784, w_000_1785, w_000_1786, w_000_1787, w_000_1788, w_000_1789, w_000_1790, w_000_1791, w_000_1792, w_000_1793, w_000_1794, w_000_1795, w_000_1796, w_000_1797, w_000_1798, w_000_1799, w_000_1800, w_000_1801, w_000_1802, w_000_1803, w_000_1804, w_000_1805, w_000_1806, w_000_1807, w_000_1808, w_000_1809, w_000_1810, w_000_1811, w_000_1812, w_000_1813, w_000_1814, w_000_1815, w_000_1816, w_000_1817, w_000_1818, w_000_1819, w_000_1820, w_000_1821, w_000_1822, w_000_1823, w_000_1824, w_000_1825, w_000_1826, w_000_1827, w_000_1828, w_000_1829, w_000_1830, w_000_1831, w_000_1832, w_000_1833, w_000_1834, w_000_1835, w_000_1836, w_000_1837, w_000_1838, w_000_1839, w_000_1840, w_000_1841, w_000_1842, w_000_1843, w_000_1844, w_000_1845, w_000_1846, w_000_1847, w_000_1848, w_000_1849, w_000_1850, w_000_1851, w_000_1852, w_000_1853, w_000_1854, w_000_1855, w_000_1856, w_000_1857, w_000_1858, w_000_1859, w_000_1860, w_000_1861, w_000_1862, w_000_1863, w_000_1864, w_000_1865, w_000_1866, w_000_1867, w_000_1868, w_000_1869, w_000_1870, w_000_1871, w_000_1872, w_000_1873, w_000_1874, w_000_1875, w_000_1876, w_000_1877, w_000_1878, w_000_1879, w_000_1880, w_000_1881, w_000_1882, w_000_1883, w_000_1884, w_000_1885, w_000_1886, w_000_1887, w_000_1888, w_000_1889, w_000_1890, w_000_1891, w_000_1892, w_000_1893, w_000_1894, w_000_1895, w_000_1896, w_000_1897, w_000_1898, w_000_1899, w_000_1900, w_000_1901, w_000_1902, w_000_1903, w_000_1904, w_000_1905, w_000_1906, w_000_1907, w_000_1908, w_000_1909, w_000_1910, w_000_1911, w_000_1912, w_000_1913, w_000_1914, w_000_1915, w_000_1916, w_000_1917, w_000_1918, w_000_1919, w_000_1920, w_000_1921, w_000_1922, w_000_1923, w_000_1924, w_000_1925, w_000_1926, w_000_1927, w_000_1928, w_000_1929, w_000_1930, w_000_1931, w_000_1932, w_000_1933, w_000_1934, w_000_1935, w_000_1936, w_000_1937, w_000_1938, w_000_1939, w_000_1940, w_000_1941, w_000_1942, w_000_1943, w_000_1944, w_000_1945, w_000_1946, w_000_1947, w_000_1948, w_000_1949, w_000_1950, w_000_1951, w_000_1952, w_000_1953, w_000_1954, w_000_1955, w_000_1956, w_000_1957, w_000_1958, w_000_1959, w_000_1960, w_000_1961, w_000_1962, w_000_1963, w_000_1964, w_000_1965, w_000_1966, w_000_1967, w_000_1968, w_000_1969, w_000_1970, w_000_1971, w_000_1972, w_000_1973, w_000_1974, w_000_1975, w_000_1976, w_000_1977, w_000_1978, w_000_1979, w_000_1980, w_000_1981, w_000_1982, w_000_1983, w_000_1984, w_000_1985, w_000_1986, w_000_1987, w_000_1988, w_000_1989, w_000_1990, w_000_1991, w_000_1992, w_000_1993, w_000_1994, w_000_1995, w_000_1996, w_000_1997, w_000_1998, w_000_1999, w_000_2000, w_000_2001, w_000_2002, w_000_2003, w_000_2004, w_000_2005, w_000_2006, w_000_2007, w_000_2008, w_000_2009, w_000_2010, w_000_2011, w_000_2012, w_000_2013, w_000_2014, w_000_2015, w_000_2016, w_000_2017, w_000_2018, w_000_2019, w_000_2020, w_000_2021, w_000_2022, w_000_2023, w_000_2024, w_000_2025, w_000_2026, w_000_2027, w_000_2028, w_000_2029, w_000_2030, w_000_2031, w_000_2032, w_000_2033, w_000_2034, w_000_2035, w_000_2036, w_000_2037, w_000_2038, w_000_2039, w_000_2040, w_000_2041, w_000_2042, w_000_2043, w_000_2044, w_000_2045, w_000_2046, w_000_2047, w_000_2048, w_000_2049, w_000_2050, w_000_2051, w_000_2052, w_000_2053, w_000_2054, w_000_2055, w_000_2056, w_000_2057, w_000_2058, w_000_2059, w_000_2060, w_000_2061, w_000_2062, w_000_2063, w_000_2064, w_000_2065, w_000_2066, w_000_2067, w_000_2068, w_000_2069, w_000_2070, w_000_2071, w_000_2072, w_000_2073, w_000_2074, w_000_2075, w_000_2076, w_000_2077, w_000_2078, w_000_2079, w_000_2080, w_000_2081, w_000_2082, w_000_2083, w_000_2084, w_000_2085, w_000_2086, w_000_2087, w_000_2088, w_000_2089, w_000_2090, w_000_2091, w_000_2092, w_000_2093, w_000_2094, w_000_2095, w_000_2096, w_000_2097, w_000_2098, w_000_2099, w_000_2100, w_000_2101, w_000_2102, w_000_2103, w_000_2104, w_000_2105, w_000_2106, w_000_2107, w_000_2108, w_000_2109, w_000_2110, w_000_2111, w_000_2112, w_000_2113, w_000_2114, w_000_2115, w_000_2116, w_000_2117, w_000_2118, w_000_2119, w_000_2120, w_000_2121, w_000_2122, w_000_2123, w_000_2124, w_000_2125, w_000_2126, w_000_2127, w_000_2128, w_000_2129, w_000_2130, w_000_2131, w_000_2132, w_000_2133, w_000_2134, w_000_2135, w_000_2136, w_000_2137, w_000_2138, w_000_2139, w_000_2140, w_000_2141, w_000_2142, w_000_2143, w_000_2144, w_000_2145, w_000_2146, w_000_2147, w_000_2148, w_000_2149, w_000_2150, w_000_2151, w_000_2152, w_000_2153, w_000_2154, w_000_2155, w_000_2156, w_000_2157, w_000_2158, w_000_2159, w_000_2160, w_000_2161, w_000_2162, w_000_2163, w_000_2164, w_000_2165, w_000_2166, w_000_2167, w_000_2168, w_000_2169, w_000_2170, w_000_2171, w_000_2172, w_000_2173, w_000_2174, w_000_2175, w_000_2176, w_000_2177, w_000_2178, w_000_2179, w_000_2180, w_000_2181, w_000_2182, w_000_2183, w_000_2184, w_000_2185, w_000_2186, w_000_2187, w_000_2188, w_000_2189, w_000_2190, w_000_2191, w_000_2192, w_000_2193, w_000_2194, w_000_2195, w_000_2196, w_000_2197, w_000_2198, w_000_2199, w_000_2200, w_000_2201, w_000_2202, w_000_2203, w_000_2204, w_000_2205, w_000_2206, w_000_2207, w_000_2208, w_000_2209, w_000_2210, w_000_2211, w_000_2212, w_000_2213, w_000_2214, w_000_2215, w_000_2216, w_000_2217, w_000_2218, w_000_2219, w_000_2220, w_000_2221, w_000_2222, w_000_2223, w_000_2224, w_000_2225, w_000_2226, w_000_2227, w_000_2228, w_000_2229, w_000_2230, w_000_2231, w_000_2232, w_000_2233, w_000_2234, w_000_2235, w_000_2236, w_000_2237, w_000_2238, w_000_2239, w_000_2240, w_000_2241, w_000_2242, w_000_2243, w_000_2244, w_000_2245, w_000_2246, w_000_2247, w_000_2248, w_000_2249, w_000_2250, w_000_2251, w_000_2252, w_000_2253, w_000_2254, w_000_2255, w_000_2256, w_000_2257, w_000_2258, w_000_2259, w_000_2260, w_000_2261, w_000_2262, w_000_2263, w_000_2264, w_000_2265, w_000_2266, w_000_2267, w_000_2268, w_000_2269, w_000_2270, w_000_2271, w_000_2272, w_000_2273, w_000_2274, w_000_2275, w_000_2276, w_000_2277, w_000_2278, w_000_2279, w_000_2280, w_000_2281, w_000_2282, w_000_2283, w_000_2284, w_000_2285, w_000_2286, w_000_2287, w_000_2288, w_000_2289, w_000_2290, w_000_2291, w_000_2292, w_000_2293, w_000_2294, w_000_2295, w_000_2296, w_000_2297, w_000_2298, w_000_2299, w_000_2300, w_000_2301, w_000_2302, w_000_2303, w_000_2304, w_000_2305, w_000_2306, w_000_2307, w_000_2308, w_000_2309, w_000_2310, w_000_2311, w_000_2312, w_000_2313, w_000_2314, w_000_2315, w_000_2316, w_000_2317, w_000_2318, w_000_2319, w_000_2320, w_000_2321, w_000_2322, w_000_2323, w_000_2324, w_000_2325, w_000_2326, w_000_2327, w_000_2328, w_000_2329, w_000_2330, w_000_2331, w_000_2332, w_000_2333, w_000_2334, w_000_2335, w_000_2336, w_000_2337, w_000_2338, w_000_2339, w_000_2340, w_000_2341, w_000_2342, w_000_2343, w_000_2344, w_000_2345, w_000_2346, w_000_2347, w_000_2348, w_000_2349, w_000_2350, w_000_2351, w_000_2352, w_000_2353, w_000_2354, w_000_2355, w_000_2356, w_000_2357, w_000_2358, w_000_2359, w_000_2360, w_000_2361, w_000_2362, w_000_2363, w_000_2364, w_000_2365, w_000_2366, w_000_2367, w_000_2368, w_000_2369, w_000_2370, w_000_2371, w_000_2372, w_000_2373, w_000_2374, w_000_2375, w_000_2376, w_000_2377, w_000_2378, w_000_2379, w_000_2380, w_000_2381, w_000_2382, w_000_2383, w_000_2384, w_000_2385, w_000_2386, w_000_2387, w_000_2388, w_000_2389, w_000_2390, w_000_2391, w_000_2392, w_000_2393, w_000_2394, w_000_2395, w_000_2396, w_000_2397, w_000_2398, w_000_2399, w_000_2400, w_000_2401, w_000_2402, w_000_2403, w_000_2404, w_000_2405, w_000_2406, w_000_2407, w_000_2408, w_000_2409, w_000_2410, w_000_2411, w_000_2412, w_000_2413, w_000_2414, w_000_2415, w_000_2416, w_000_2417, w_000_2418, w_000_2419, w_000_2420, w_000_2421, w_000_2422, w_000_2423, w_000_2424, w_000_2425, w_000_2426, w_000_2427, w_000_2428, w_000_2429, w_000_2430, w_000_2431, w_000_2432, w_000_2433, w_000_2434, w_000_2435, w_000_2436, w_000_2437, w_000_2438, w_000_2439, w_000_2440, w_000_2441, w_000_2442, w_000_2443, w_000_2444, w_000_2445, w_000_2446, w_000_2447, w_000_2448, w_000_2449, w_000_2450, w_000_2451, w_000_2452, w_000_2453, w_000_2454, w_000_2455, w_000_2456, w_000_2457, w_000_2458, w_000_2459, w_000_2460, w_000_2461, w_000_2462, w_000_2463, w_000_2464, w_000_2465, w_000_2466, w_000_2467, w_000_2468, w_000_2469, w_000_2470, w_000_2471, w_000_2472, w_000_2473, w_000_2474, w_000_2475, w_000_2476, w_000_2477, w_000_2478, w_000_2479, w_000_2480, w_000_2481, w_000_2482, w_000_2483, w_000_2484, w_000_2485, w_000_2486, w_000_2487, w_000_2488, w_000_2489, w_000_2490, w_000_2491, w_000_2492, w_000_2493, w_000_2494, w_000_2495, w_000_2496, w_000_2497, w_000_2498, w_000_2499, w_000_2500, w_000_2501, w_000_2502, w_000_2503, w_000_2504, w_000_2505, w_000_2506, w_000_2507, w_000_2508, w_000_2509, w_000_2510, w_000_2511, w_000_2512, w_000_2513, w_000_2514, w_000_2515, w_000_2516, w_000_2517, w_000_2518, w_000_2519, w_000_2520, w_000_2521, w_000_2522, w_000_2523, w_000_2524, w_000_2525, w_000_2526, w_000_2527, w_000_2528, w_000_2529, w_000_2530, w_000_2531, w_000_2532, w_000_2533, w_000_2534, w_000_2535, w_000_2536, w_000_2537, w_000_2538, w_000_2539, w_000_2540, w_000_2541, w_000_2542, w_000_2543, w_000_2544, w_000_2545, w_000_2546, w_000_2547, w_000_2548, w_000_2549, w_000_2550, w_000_2551, w_000_2552, w_000_2553, w_000_2554, w_000_2555, w_000_2556, w_000_2557, w_000_2558, w_000_2559, w_000_2560, w_000_2561, w_000_2562, w_000_2563, w_000_2564, w_000_2565, w_000_2566, w_000_2567, w_000_2568, w_000_2569, w_000_2570, w_000_2571, w_000_2572, w_000_2573, w_000_2574, w_000_2575, w_000_2576, w_000_2577, w_000_2578, w_000_2579, w_000_2580, w_000_2581, w_000_2582, w_000_2583, w_000_2584, w_000_2585, w_000_2586, w_000_2587, w_000_2588, w_000_2589, w_000_2590, w_000_2591, w_000_2592, w_000_2593, w_000_2594, w_000_2595, w_000_2596, w_000_2597, w_000_2598, w_000_2599, w_000_2600, w_000_2601, w_000_2602, w_000_2603, w_000_2604, w_000_2605, w_000_2606, w_000_2607, w_000_2608, w_000_2609, w_000_2610, w_000_2611, w_000_2612, w_000_2613, w_000_2614, w_000_2615, w_000_2616, w_000_2617, w_000_2618, w_000_2619, w_000_2620, w_000_2621, w_000_2622, w_000_2623, w_000_2624, w_000_2625, w_000_2626, w_000_2627, w_000_2628, w_000_2629, w_000_2630, w_000_2631, w_000_2632, w_000_2633, w_000_2634, w_000_2635, w_000_2636, w_000_2637, w_000_2638, w_000_2639, w_000_2640, w_000_2641, w_000_2642, w_000_2643, w_000_2644, w_000_2645, w_000_2646, w_000_2647, w_000_2648, w_000_2649, w_000_2650, w_000_2651, w_000_2652, w_000_2653, w_000_2654, w_000_2655, w_000_2656, w_000_2657, w_000_2658, w_000_2659, w_000_2660, w_000_2661, w_000_2662, w_000_2663, w_000_2664, w_000_2665, w_000_2666, w_000_2667, w_000_2668, w_000_2669, w_000_2670, w_000_2671, w_000_2672, w_000_2673, w_000_2674, w_000_2675, w_000_2676, w_000_2677, w_000_2678, w_000_2679, w_000_2680, w_000_2681, w_000_2682, w_000_2683, w_000_2684, w_000_2685, w_000_2686, w_000_2687, w_000_2688, w_000_2689, w_000_2690, w_000_2691, w_000_2692, w_000_2693, w_000_2694, w_000_2695, w_000_2696, w_000_2697, w_000_2698, w_000_2699, w_000_2700, w_000_2701, w_000_2702, w_000_2703, w_000_2704, w_000_2705, w_000_2706, w_000_2707, w_000_2708, w_000_2709, w_000_2710, w_000_2711, w_000_2712, w_000_2713, w_000_2714, w_000_2715, w_000_2716, w_000_2717, w_000_2718, w_000_2719, w_000_2720, w_000_2721, w_000_2722, w_000_2723, w_000_2724, w_000_2725, w_000_2726, w_000_2727, w_000_2728, w_000_2729, w_000_2730, w_000_2731, w_000_2732, w_000_2733, w_000_2734, w_000_2735, w_000_2736, w_000_2737, w_000_2738, w_000_2739, w_000_2740, w_000_2741, w_000_2742, w_000_2743, w_000_2744, w_000_2745, w_000_2746, w_000_2747, w_000_2748, w_000_2749, w_000_2750, w_000_2751, w_000_2752, w_000_2753, w_000_2754, w_000_2755, w_000_2756, w_000_2757, w_000_2758, w_000_2759, w_000_2760, w_000_2761, w_000_2762, w_000_2763, w_000_2764, w_000_2765, w_000_2766, w_000_2767, w_000_2768, w_000_2769, w_000_2770, w_000_2771, w_000_2772, w_000_2773, w_000_2774, w_000_2775, w_000_2776, w_000_2777, w_000_2778, w_000_2779, w_000_2780, w_000_2781, w_000_2782, w_000_2783, w_000_2784, w_000_2785, w_000_2786, w_000_2787, w_000_2788, w_000_2789, w_000_2790, w_000_2791, w_000_2792, w_000_2793, w_000_2794, w_000_2795, w_000_2796, w_000_2797, w_000_2798, w_000_2799, w_000_2800, w_000_2801, w_000_2802, w_000_2803, w_000_2804, w_000_2805, w_000_2806, w_000_2807, w_000_2808, w_000_2809, w_000_2810, w_000_2811, w_000_2812, w_000_2813, w_000_2814, w_000_2815, w_000_2816, w_000_2817, w_000_2818, w_000_2819, w_000_2820, w_000_2821, w_000_2822, w_000_2823, w_000_2824, w_000_2825, w_000_2826, w_000_2827, w_000_2828, w_000_2829, w_000_2830, w_000_2831, w_000_2832, w_000_2833, w_000_2834, w_000_2835, w_000_2836, w_000_2837, w_000_2838, w_000_2839, w_000_2840, w_000_2841, w_000_2842, w_000_2843, w_000_2844, w_000_2845, w_000_2846, w_000_2847, w_000_2848, w_000_2849, w_000_2850, w_000_2851, w_000_2852, w_000_2853, w_000_2854, w_000_2855, w_000_2856, w_000_2857, w_000_2858, w_000_2859, w_000_2860, w_000_2861, w_000_2862, w_000_2863, w_000_2864, w_000_2865, w_000_2866, w_000_2867, w_000_2868, w_000_2869, w_000_2870, w_000_2871, w_000_2872, w_000_2873, w_000_2874, w_000_2875, w_000_2876, w_000_2877, w_000_2878, w_000_2879, w_000_2880, w_000_2881, w_000_2882, w_000_2883, w_000_2884, w_000_2885, w_000_2886, w_000_2887, w_000_2888, w_000_2889, w_000_2890, w_000_2891, w_000_2892, w_000_2893, w_000_2894, w_000_2895, w_000_2896, w_000_2897, w_000_2898, w_000_2899, w_000_2900, w_000_2901, w_000_2902, w_000_2903, w_000_2904, w_000_2905, w_000_2906, w_000_2907, w_000_2908, w_000_2909, w_000_2910, w_000_2911, w_000_2912, w_000_2913, w_000_2914, w_000_2915, w_000_2916, w_000_2917, w_000_2918, w_000_2919, w_000_2920, w_000_2921, w_000_2922, w_000_2923, w_000_2924, w_000_2925, w_000_2926, w_000_2927, w_000_2928, w_000_2929, w_000_2930, w_000_2931, w_000_2932, w_000_2933, w_000_2934, w_000_2935, w_000_2936, w_000_2937, w_000_2938, w_000_2939, w_000_2940, w_000_2941, w_000_2942, w_000_2943, w_000_2944, w_000_2945, w_000_2946, w_000_2947, w_000_2948, w_000_2949, w_000_2950, w_000_2951, w_000_2952, w_000_2953, w_000_2954, w_000_2955, w_000_2956, w_000_2957, w_000_2958, w_000_2959, w_000_2960, w_000_2961, w_000_2962, w_000_2963, w_000_2964, w_000_2965, w_000_2966, w_000_2967, w_000_2968, w_000_2969, w_000_2970, w_000_2971, w_000_2972, w_000_2973, w_000_2974, w_000_2975, w_000_2976, w_000_2977, w_000_2978, w_000_2979, w_000_2980, w_000_2981, w_000_2982, w_000_2983, w_000_2984, w_000_2985, w_000_2986, w_000_2987, w_000_2988, w_000_2989, w_000_2990, w_000_2991, w_000_2992, w_000_2993, w_000_2994, w_000_2995, w_000_2996, w_000_2997, w_000_2998, w_000_2999, w_000_3000, w_000_3001, w_000_3002, w_000_3003, w_000_3004, w_000_3005, w_000_3006, w_000_3007, w_000_3008, w_000_3009, w_000_3010, w_000_3011, w_000_3012, w_000_3013, w_000_3014, w_000_3015, w_000_3016, w_000_3017, w_000_3019, w_000_3020, w_000_3021, w_000_3022, w_000_3023, w_000_3024, w_000_3025, w_000_3026, w_000_3027, w_000_3028, w_000_3029, w_000_3030, w_000_3031, w_000_3032, w_000_3033, w_000_3034, w_000_3035, w_000_3036, w_000_3037, w_000_3038, w_000_3039, w_000_3040, w_000_3041, w_000_3042, w_000_3043, w_000_3044, w_000_3045, w_000_3046, w_000_3047, w_000_3048, w_000_3049, w_000_3050, w_000_3051, w_000_3052, w_000_3053, w_000_3054, w_000_3055, w_000_3056, w_000_3057, w_000_3058, w_000_3059, w_000_3060, w_000_3061, w_000_3062, w_000_3063, w_000_3064, w_000_3065, w_000_3066, w_000_3067, w_000_3068, w_000_3069, w_000_3070, w_000_3071, w_000_3072, w_000_3073, w_000_3074, w_000_3075, w_000_3076, w_000_3077, w_000_3078, w_000_3079, w_000_3080, w_000_3081, w_000_3082, w_000_3083, w_000_3084, w_000_3085, w_000_3086, w_000_3087, w_000_3088, w_000_3089, w_000_3090, w_000_3091, w_000_3092, w_000_3093, w_000_3094, w_000_3095, w_000_3096, w_000_3097, w_000_3098, w_000_3099, w_000_3100, w_000_3101, w_000_3102, w_000_3103, w_000_3104, w_000_3105, w_000_3106, w_000_3107, w_000_3108, w_000_3109, w_000_3110, w_000_3111, w_000_3112, w_000_3113, w_000_3114, w_000_3115, w_000_3116, w_000_3117, w_000_3118, w_000_3119, w_000_3120, w_000_3121, w_000_3122, w_000_3123, w_000_3124, w_000_3125, w_000_3126, w_000_3127, w_000_3128, w_000_3129, w_000_3130, w_000_3131, w_000_3132, w_000_3133, w_000_3134, w_000_3135, w_000_3136, w_000_3137, w_000_3138, w_000_3139, w_000_3140, w_000_3141, w_000_3142, w_000_3143, w_000_3144, w_000_3145, w_000_3146, w_000_3147, w_000_3148, w_000_3149, w_000_3150, w_000_3151, w_000_3152, w_000_3153, w_000_3154, w_000_3155, w_000_3156, w_000_3157, w_000_3158, w_000_3159, w_000_3160, w_000_3161, w_000_3162, w_000_3163, w_000_3164, w_000_3165, w_000_3166, w_000_3167, w_000_3168, w_000_3169, w_000_3170, w_000_3171, w_000_3172, w_000_3173, w_000_3174, w_000_3175, w_000_3176, w_000_3177, w_000_3178, w_000_3179, w_000_3180, w_000_3181, w_000_3182, w_000_3183, w_000_3184, w_000_3185, w_000_3186, w_000_3187, w_000_3188, w_000_3189, w_000_3190, w_000_3191, w_000_3192, w_000_3193, w_000_3194, w_000_3195, w_000_3196, w_000_3197, w_000_3198, w_000_3199, w_000_3200, w_000_3201, w_000_3202, w_000_3203, w_000_3204, w_000_3205, w_000_3206, w_000_3207, w_000_3208, w_000_3209, w_000_3210, w_000_3211, w_000_3212, w_000_3213, w_000_3214, w_000_3215, w_000_3216, w_000_3217, w_000_3218, w_000_3219, w_000_3220, w_000_3221, w_000_3222, w_000_3223, w_000_3224, w_000_3225, w_000_3226, w_000_3227, w_000_3228, w_000_3229, w_000_3230, w_000_3231, w_000_3232, w_000_3233, w_000_3234, w_000_3235, w_000_3236, w_000_3237, w_000_3238, w_000_3239, w_000_3240, w_000_3241, w_000_3242, w_000_3243, w_000_3244, w_000_3245, w_000_3246, w_000_3247, w_000_3248, w_000_3249, w_000_3250, w_000_3251, w_000_3252, w_000_3253, w_000_3254, w_000_3255, w_000_3256, w_000_3257, w_000_3258, w_000_3259, w_000_3260, w_000_3261, w_000_3262, w_000_3263, w_000_3264, w_000_3265, w_000_3266, w_000_3267, w_000_3268, w_000_3269, w_000_3270, w_000_3271, w_000_3272, w_000_3273, w_000_3274, w_000_3275, w_000_3276, w_000_3277, w_000_3278, w_000_3279, w_000_3280, w_000_3281, w_000_3282, w_000_3283, w_000_3284, w_000_3285, w_000_3286, w_000_3287, w_000_3288, w_000_3289, w_000_3290, w_000_3291, w_000_3292, w_000_3293, w_000_3294, w_000_3295, w_000_3296, w_000_3297, w_000_3298, w_000_3299, w_000_3300, w_000_3301, w_000_3302, w_000_3303, w_000_3304, w_000_3305, w_000_3306, w_000_3307, w_000_3308, w_000_3309, w_000_3310, w_000_3311, w_000_3312, w_000_3313, w_000_3314, w_000_3315, w_000_3316, w_000_3317, w_000_3318, w_000_3319, w_000_3320, w_000_3321, w_000_3322, w_000_3323, w_000_3324, w_000_3325, w_000_3326, w_000_3327, w_000_3328, w_000_3329, w_000_3330, w_000_3331, w_000_3332, w_000_3333, w_000_3334, w_000_3335, w_000_3336, w_000_3337, w_000_3338, w_000_3339, w_000_3340, w_000_3341, w_000_3342, w_000_3343, w_000_3344, w_000_3345, w_000_3346, w_000_3347, w_000_3348, w_000_3349, w_000_3350, w_000_3351, w_000_3352, w_000_3353, w_000_3354, w_000_3355, w_000_3356, w_000_3357, w_000_3358, w_000_3359, w_000_3360, w_000_3361, w_000_3362, w_000_3363, w_000_3364, w_000_3365, w_000_3366, w_000_3367, w_000_3368, w_000_3369, w_000_3370, w_000_3371, w_000_3372, w_000_3373, w_000_3374, w_000_3375, w_000_3376, w_000_3377, w_000_3378, w_000_3379, w_000_3380, w_000_3381, w_000_3382, w_000_3383, w_000_3384, w_000_3385, w_000_3386, w_000_3387, w_000_3388, w_000_3389, w_000_3390, w_000_3391, w_000_3392, w_000_3393, w_000_3394, w_000_3395, w_000_3396, w_000_3397, w_000_3398, w_000_3399, w_000_3400, w_000_3401, w_000_3402, w_000_3403, w_000_3404, w_000_3405, w_000_3406, w_000_3407, w_000_3408, w_000_3409, w_000_3410, w_000_3411, w_000_3412, w_000_3413, w_000_3414, w_000_3415, w_000_3416, w_000_3417, w_000_3418, w_000_3419, w_000_3420, w_000_3421, w_000_3422, w_000_3423, w_000_3424, w_000_3425, w_000_3426, w_000_3427, w_000_3428, w_000_3429, w_000_3430, w_000_3431, w_000_3432, w_000_3433, w_000_3434, w_000_3435, w_000_3436, w_000_3437, w_000_3438, w_000_3439, w_000_3440, w_000_3441, w_000_3442, w_000_3443, w_000_3444, w_000_3445, w_000_3446, w_000_3447, w_000_3448, w_000_3449, w_000_3450, w_000_3451, w_000_3452, w_000_3453, w_000_3454, w_000_3455, w_000_3456, w_000_3457, w_000_3458, w_000_3459, w_000_3460, w_000_3461, w_000_3462, w_000_3463, w_000_3464, w_000_3465, w_000_3466, w_000_3467, w_000_3468, w_000_3469, w_000_3470, w_000_3471, w_000_3472, w_000_3473, w_000_3474, w_000_3475, w_000_3476, w_000_3477, w_000_3478, w_000_3479, w_000_3480, w_000_3481, w_000_3482, w_000_3483, w_000_3484, w_000_3485, w_000_3486, w_000_3487, w_000_3488, w_000_3489, w_000_3490, w_000_3491, w_000_3492, w_000_3493, w_000_3494, w_000_3495, w_000_3496, w_000_3497, w_000_3498, w_000_3499, w_000_3500, w_000_3501, w_000_3502, w_000_3503, w_000_3504, w_000_3505, w_000_3506, w_000_3507, w_000_3508, w_000_3509, w_000_3510, w_000_3511, w_000_3512, w_000_3513, w_000_3514, w_000_3515, w_000_3516, w_000_3517, w_000_3518, w_000_3519, w_000_3520, w_000_3521, w_000_3522, w_000_3523, w_000_3524, w_000_3525, w_000_3526, w_000_3527, w_000_3528, w_000_3529, w_000_3530, w_000_3531, w_000_3532, w_000_3533, w_000_3534, w_000_3535, w_000_3536, w_000_3537, w_000_3538, w_000_3539, w_000_3540, w_000_3541, w_000_3542, w_000_3543, w_000_3544, w_000_3545, w_000_3546, w_000_3547, w_000_3548, w_000_3549, w_000_3550, w_000_3551, w_000_3552, w_000_3553, w_000_3554, w_000_3555, w_000_3556, w_000_3557, w_000_3558, w_000_3559, w_000_3560, w_000_3561, w_000_3562, w_000_3563, w_000_3564, w_000_3565, w_000_3566, w_000_3567, w_000_3568, w_000_3569, w_000_3570, w_000_3571, w_000_3572, w_000_3573, w_000_3574, w_000_3575, w_000_3576, w_000_3577, w_000_3578, w_000_3579, w_000_3580, w_000_3581, w_000_3582, w_000_3583, w_000_3584, w_000_3585, w_000_3586, w_000_3587, w_000_3588, w_000_3589, w_000_3590, w_000_3591, w_000_3592, w_000_3593, w_000_3594, w_000_3595, w_000_3596, w_000_3597, w_000_3598, w_000_3599, w_000_3600, w_000_3601, w_000_3602, w_000_3603, w_000_3604, w_000_3605, w_000_3606, w_000_3607, w_000_3608, w_000_3609, w_000_3610, w_000_3611, w_000_3612, w_000_3613, w_000_3614, w_000_3615, w_000_3616, w_000_3617, w_000_3618, w_000_3619, w_000_3620, w_000_3621, w_000_3622, w_000_3623, w_000_3624, w_000_3625, w_000_3626, w_000_3627, w_000_3628, w_000_3629, w_000_3630, w_000_3631, w_000_3632, w_000_3633, w_000_3634, w_000_3635, w_000_3636, w_000_3637, w_000_3638, w_000_3639, w_000_3640, w_000_3641, w_000_3642, w_000_3643, w_000_3644, w_000_3645, w_000_3646, w_000_3647, w_000_3648, w_000_3649, w_000_3650, w_000_3651, w_000_3652, w_000_3653, w_000_3654, w_000_3655, w_000_3656, w_000_3657, w_000_3658, w_000_3659, w_000_3660, w_000_3661, w_000_3662, w_000_3663, w_000_3664, w_000_3665, w_000_3666, w_000_3667, w_000_3668, w_000_3669, w_000_3670, w_000_3671, w_000_3672, w_000_3673, w_000_3674, w_000_3675, w_000_3676, w_000_3677, w_000_3678, w_000_3679, w_000_3680, w_000_3681, w_000_3682, w_000_3683, w_000_3684, w_000_3685, w_000_3686, w_000_3687, w_000_3688, w_000_3689, w_000_3690, w_000_3691, w_000_3692, w_000_3693, w_000_3694, w_000_3695, w_000_3696, w_000_3697, w_000_3698, w_000_3699, w_000_3700, w_000_3701, w_000_3702, w_000_3703, w_000_3704, w_000_3705, w_000_3706, w_000_3707, w_000_3708, w_000_3709, w_000_3710, w_000_3711, w_000_3712, w_000_3713, w_000_3714, w_000_3715, w_000_3716, w_000_3717, w_000_3718, w_000_3719, w_000_3720, w_000_3721, w_000_3722, w_000_3723, w_000_3724, w_000_3725, w_000_3726, w_000_3727, w_000_3728, w_000_3729, w_000_3730, w_000_3731, w_000_3732, w_000_3733, w_000_3734, w_000_3735, w_000_3736, w_000_3737, w_000_3738, w_000_3739, w_000_3740, w_000_3741, w_000_3742, w_000_3743, w_000_3744, w_000_3745, w_000_3746, w_000_3747, w_000_3748, w_000_3749, w_000_3750, w_000_3751, w_000_3752, w_000_3753, w_000_3754, w_000_3755, w_000_3756, w_000_3757, w_000_3758, w_000_3759, w_000_3760, w_000_3761, w_000_3762, w_000_3763, w_000_3764, w_000_3765, w_000_3766, w_000_3767, w_000_3768, w_000_3769, w_000_3770, w_000_3771, w_000_3772, w_000_3773, w_000_3774, w_000_3775, w_000_3776, w_000_3777, w_000_3778, w_000_3779, w_000_3780, w_000_3781, w_000_3782, w_000_3783, w_000_3784, w_000_3785, w_000_3786, w_000_3787, w_000_3788, w_000_3789, w_000_3790, w_000_3791, w_000_3792, w_000_3793, w_000_3794, w_000_3795, w_000_3796, w_000_3797, w_000_3798, w_000_3799, w_000_3800, w_000_3801, w_000_3802, w_000_3803, w_000_3804, w_000_3805, w_000_3806, w_000_3807, w_000_3808, w_000_3809, w_000_3810, w_000_3811, w_000_3812, w_000_3813, w_000_3814, w_000_3815, w_000_3816, w_000_3817, w_000_3818, w_000_3819, w_000_3820, w_000_3821, w_000_3822, w_000_3823, w_000_3824, w_000_3825, w_000_3826, w_000_3827, w_000_3828, w_000_3829, w_000_3830, w_000_3831, w_000_3832, w_000_3833, w_000_3834, w_000_3835, w_000_3836, w_000_3837, w_000_3838, w_000_3839, w_000_3840, w_000_3841, w_000_3842, w_000_3843, w_000_3844, w_000_3845, w_000_3846, w_000_3847, w_000_3848, w_000_3849, w_000_3850, w_000_3851, w_000_3852, w_000_3853, w_000_3854, w_000_3855, w_000_3856, w_000_3857, w_000_3858, w_000_3859, w_000_3860, w_000_3861, w_000_3862, w_000_3863, w_000_3864, w_000_3865, w_000_3866, w_000_3867, w_000_3868, w_000_3869, w_000_3870, w_000_3871, w_000_3872, w_000_3873, w_000_3874, w_000_3875, w_000_3876, w_000_3877, w_000_3878, w_000_3879, w_000_3880, w_000_3881, w_000_3882, w_000_3883, w_000_3884, w_000_3885, w_000_3886, w_000_3887, w_000_3888, w_000_3889, w_000_3890, w_000_3891, w_000_3892, w_000_3893, w_000_3894, w_000_3895, w_000_3896, w_000_3897, w_000_3898, w_000_3899, w_000_3900, w_000_3901, w_000_3902, w_000_3903, w_000_3904, w_000_3905, w_000_3906, w_000_3907, w_000_3908, w_000_3909, w_000_3910, w_000_3911, w_000_3912, w_000_3913, w_000_3914, w_000_3915, w_000_3916, w_000_3917, w_000_3918, w_000_3919, w_000_3920, w_000_3921, w_000_3922, w_000_3923, w_000_3924, w_000_3925, w_000_3926, w_000_3927, w_000_3928, w_000_3929, w_000_3930, w_000_3931, w_000_3932, w_000_3933, w_000_3934, w_000_3935, w_000_3936, w_000_3937, w_000_3938, w_000_3939, w_000_3940, w_000_3941, w_000_3942, w_000_3943, w_000_3944, w_000_3945, w_000_3946, w_000_3947, w_000_3948, w_000_3949, w_000_3950, w_000_3951, w_000_3952, w_000_3953, w_000_3954, w_000_3955, w_000_3956, w_000_3957, w_000_3958, w_000_3959, w_000_3960, w_000_3961, w_000_3962, w_000_3963, w_000_3964, w_000_3965, w_000_3966, w_000_3967, w_000_3968, w_000_3969, w_000_3970, w_000_3971, w_000_3972, w_000_3973, w_000_3974, w_000_3975, w_000_3976, w_000_3977, w_000_3978, w_000_3979, w_000_3980, w_000_3981, w_000_3982, w_000_3983, w_000_3984, w_000_3985, w_000_3986, w_000_3987, w_000_3988, w_000_3989, w_000_3990, w_000_3991, w_000_3992, w_000_3993, w_000_3994, w_000_3995, w_000_3996, w_000_3997, w_000_3998, w_000_3999, w_000_4000, w_000_4001, w_000_4002, w_000_4003, w_000_4004, w_000_4005, w_000_4006, w_000_4007, w_000_4008, w_000_4009, w_000_4010, w_000_4011, w_000_4012, w_000_4013, w_000_4014, w_000_4015, w_000_4016, w_000_4017, w_000_4018, w_000_4019, w_000_4020, w_000_4021, w_000_4022, w_000_4023, w_000_4024, w_000_4025, w_000_4026, w_000_4027, w_000_4028, w_000_4029, w_000_4030, w_000_4031, w_000_4032, w_000_4033, w_000_4034, w_000_4035, w_000_4036, w_000_4037, w_000_4038, w_000_4039, w_000_4040, w_000_4041, w_000_4042, w_000_4043, w_000_4044, w_000_4045, w_000_4046, w_000_4047, w_000_4048, w_000_4049, w_000_4050, w_000_4051, w_000_4052, w_000_4053, w_000_4054, w_000_4055, w_000_4056, w_000_4057, w_000_4058, w_000_4059, w_000_4060, w_000_4061, w_000_4062, w_000_4063, w_000_4064, w_000_4065, w_000_4066, w_000_4067, w_000_4068, w_000_4069, w_000_4070, w_000_4071, w_000_4072, w_000_4073, w_000_4074, w_000_4075, w_000_4076, w_000_4077, w_000_4078, w_000_4079, w_000_4080, w_000_4081, w_000_4082, w_000_4083, w_000_4084, w_000_4085, w_000_4086, w_000_4087, w_000_4088, w_000_4089, w_000_4090, w_000_4091, w_000_4092, w_000_4093, w_000_4094, w_000_4095, w_000_4096, w_000_4097, w_000_4098, w_000_4099, w_000_4100, w_000_4101, w_000_4102, w_000_4103, w_000_4104, w_000_4105, w_000_4106, w_000_4107, w_000_4108, w_000_4109, w_000_4110, w_000_4111, w_000_4112, w_000_4113, w_000_4114, w_000_4115, w_000_4116, w_000_4117, w_000_4118, w_000_4119, w_000_4120, w_000_4121, w_000_4122, w_000_4123, w_000_4124, w_000_4125, w_000_4126, w_000_4127, w_000_4128, w_000_4129, w_000_4130, w_000_4131, w_000_4132, w_000_4133, w_000_4134, w_000_4135, w_000_4136, w_000_4137, w_000_4138, w_000_4139, w_000_4140, w_000_4141, w_000_4142, w_000_4143, w_000_4144, w_000_4145, w_000_4146, w_000_4147, w_000_4148, w_000_4149, w_000_4150, w_000_4151, w_000_4152, w_000_4153, w_000_4154, w_000_4155, w_000_4156, w_000_4157, w_000_4158, w_000_4159, w_000_4160, w_000_4161, w_000_4162, w_000_4163, w_000_4164, w_000_4165, w_000_4166, w_000_4167, w_000_4168, w_000_4169, w_000_4170, w_000_4171, w_000_4172, w_000_4173, w_000_4174, w_000_4175, w_000_4176, w_000_4177, w_000_4178, w_000_4179, w_000_4180, w_000_4181, w_000_4182, w_000_4183, w_000_4184, w_000_4185, w_000_4186, w_000_4187, w_000_4188, w_000_4189, w_000_4190, w_000_4191, w_000_4192, w_000_4193, w_000_4194, w_000_4195, w_000_4196, w_000_4197, w_000_4198, w_000_4199, w_000_4200, w_000_4201, w_000_4202, w_000_4203, w_000_4204, w_000_4205, w_000_4206, w_000_4207, w_000_4208, w_000_4209, w_000_4210, w_000_4211, w_000_4212, w_000_4213, w_000_4215, w_000_4216, w_000_4217, w_000_4218, w_000_4219, w_000_4220, w_000_4221, w_000_4222, w_000_4223, w_000_4224, w_000_4225, w_000_4226, w_000_4227, w_000_4228, w_000_4229, w_000_4230, w_000_4231, w_000_4232, w_000_4233, w_000_4234, w_000_4235, w_000_4236, w_000_4237, w_000_4238, w_000_4239, w_000_4240, w_000_4241, w_000_4242, w_000_4243, w_000_4244, w_000_4245, w_000_4246, w_000_4247, w_000_4248, w_000_4249, w_000_4250, w_000_4251, w_000_4252, w_000_4253, w_000_4254, w_000_4255, w_000_4256, w_000_4257, w_000_4258, w_000_4259, w_000_4260, w_000_4261, w_000_4262, w_000_4263, w_000_4264, w_000_4265, w_000_4266, w_000_4267, w_000_4268, w_000_4269, w_000_4270, w_000_4271, w_000_4272, w_000_4273, w_000_4274, w_000_4275, w_000_4276, w_000_4277, w_000_4278, w_000_4279, w_000_4280, w_000_4281, w_000_4282, w_000_4283, w_000_4284, w_000_4285, w_000_4286, w_000_4287, w_000_4288, w_000_4289, w_000_4290, w_000_4291, w_000_4292, w_000_4293, w_000_4294, w_000_4295, w_000_4296, w_000_4297, w_000_4298, w_000_4299, w_000_4300, w_000_4301, w_000_4302, w_000_4303, w_000_4304, w_000_4305, w_000_4306, w_000_4307, w_000_4308, w_000_4309, w_000_4310, w_000_4311, w_000_4312, w_000_4313, w_000_4314, w_000_4315, w_000_4316, w_000_4317, w_000_4318, w_000_4319, w_000_4320, w_000_4321, w_000_4322, w_000_4323, w_000_4324, w_000_4325, w_000_4326, w_000_4327, w_000_4328, w_000_4329, w_000_4330, w_000_4331, w_000_4332, w_000_4333, w_000_4334, w_000_4335, w_000_4336, w_000_4337, w_000_4338, w_000_4339, w_000_4340, w_000_4341, w_000_4342, w_000_4343, w_000_4344, w_000_4345, w_000_4346, w_000_4347, w_000_4349, w_000_4350, w_000_4351, w_000_4352, w_000_4353, w_000_4354, w_000_4355, w_000_4356, w_000_4357, w_000_4358, w_000_4359, w_000_4360, w_000_4361, w_000_4362, w_000_4363, w_000_4364, w_000_4365, w_000_4366, w_000_4367, w_000_4368, w_000_4369, w_000_4370, w_000_4371, w_000_4372, w_000_4373, w_000_4374, w_000_4375, w_000_4376, w_000_4377, w_000_4378, w_000_4379, w_000_4380, w_000_4381, w_000_4382, w_000_4383, w_000_4384, w_000_4385, w_000_4386, w_000_4387, w_000_4388, w_000_4389, w_000_4390, w_000_4391, w_000_4392, w_000_4393, w_000_4394, w_000_4395, w_000_4396, w_000_4397, w_000_4398, w_000_4399, w_000_4400, w_000_4401, w_000_4402, w_000_4403, w_000_4404, w_000_4405, w_000_4406, w_000_4407, w_000_4408, w_000_4409, w_000_4410, w_000_4411, w_000_4412, w_000_4413, w_000_4414, w_000_4415, w_000_4416, w_000_4417, w_000_4418, w_000_4419, w_000_4420, w_000_4421, w_000_4422, w_000_4423, w_000_4424, w_000_4425, w_000_4426, w_000_4427, w_000_4428, w_000_4429, w_000_4430, w_000_4431, w_000_4432, w_000_4433, w_000_4434, w_000_4435, w_000_4436, w_000_4437, w_000_4438, w_000_4439, w_000_4440, w_000_4441, w_000_4442, w_000_4443, w_000_4444, w_000_4445, w_000_4446, w_000_4447, w_000_4448, w_000_4449, w_000_4450, w_000_4451, w_000_4452, w_000_4453, w_000_4454, w_000_4455, w_000_4456, w_000_4457, w_000_4458, w_000_4459, w_000_4460, w_000_4461, w_000_4462, w_000_4463, w_000_4464, w_000_4465, w_000_4466, w_000_4467, w_000_4468, w_000_4469, w_000_4470, w_000_4471, w_000_4472, w_000_4473, w_000_4474, w_000_4475, w_000_4476, w_000_4477, w_000_4478, w_000_4479, w_000_4480, w_000_4481, w_000_4482, w_000_4483, w_000_4484, w_000_4485, w_000_4486, w_000_4487, w_000_4488, w_000_4489, w_000_4490, w_000_4491, w_000_4492, w_000_4493, w_000_4494, w_000_4495, w_000_4496, w_000_4497, w_000_4498, w_000_4499, w_000_4500, w_000_4501, w_000_4502, w_000_4503, w_000_4504, w_000_4505, w_000_4506, w_000_4507, w_000_4508, w_000_4509, w_000_4510, w_000_4511, w_000_4512, w_000_4513, w_000_4514, w_000_4515, w_000_4516, w_000_4517, w_000_4518, w_000_4519, w_000_4520, w_000_4521, w_000_4522, w_000_4523, w_000_4524, w_000_4525, w_000_4526, w_000_4527, w_000_4528, w_000_4529, w_000_4530, w_000_4531, w_000_4532, w_000_4533, w_000_4534, w_000_4535, w_000_4536, w_000_4537, w_000_4538, w_000_4539, w_000_4540, w_000_4541, w_000_4542, w_000_4543, w_000_4544, w_000_4545, w_000_4546, w_000_4547, w_000_4548, w_000_4549, w_000_4550, w_000_4551, w_000_4552, w_000_4553, w_000_4554, w_000_4555, w_000_4556, w_000_4557, w_000_4559, w_000_4560, w_000_4561, w_000_4562, w_000_4563, w_000_4564, w_000_4565, w_000_4566, w_000_4567, w_000_4568, w_000_4569, w_000_4571, w_000_4572, w_000_4573, w_000_4574, w_000_4575, w_000_4576, w_000_4577, w_000_4578, w_000_4579, w_000_4580, w_000_4581, w_000_4582, w_000_4583, w_000_4584, w_000_4585, w_000_4586, w_000_4587, w_000_4588, w_000_4589, w_000_4590, w_000_4591, w_000_4592, w_000_4593, w_000_4594, w_000_4595, w_000_4596, w_000_4597, w_000_4598, w_000_4599, w_000_4600, w_000_4601, w_000_4602, w_000_4603, w_000_4604, w_000_4605, w_000_4606, w_000_4607, w_000_4608, w_000_4609, w_000_4610, w_000_4611, w_000_4612, w_000_4613, w_000_4614, w_000_4615, w_000_4616, w_000_4617, w_000_4618, w_000_4619, w_000_4620, w_000_4621, w_000_4622, w_000_4623, w_000_4624, w_000_4625, w_000_4626, w_000_4627, w_000_4628, w_000_4629, w_000_4630, w_000_4631, w_000_4632, w_000_4633, w_000_4634, w_000_4635, w_000_4636, w_000_4637, w_000_4638, w_000_4639, w_000_4640, w_000_4641, w_000_4642, w_000_4643, w_000_4644, w_000_4645, w_000_4646, w_000_4647, w_000_4648, w_000_4649, w_000_4650, w_000_4651, w_000_4652, w_000_4653, w_000_4654, w_000_4655, w_000_4656, w_000_4657, w_000_4658, w_000_4659, w_000_4660, w_000_4661, w_000_4662, w_000_4663, w_000_4664, w_000_4665, w_000_4666, w_000_4667, w_000_4668, w_000_4669, w_000_4670, w_000_4671, w_000_4672, w_000_4673, w_000_4674, w_000_4675, w_000_4676, w_000_4677, w_000_4678, w_000_4679, w_000_4680, w_000_4681, w_000_4682, w_000_4683, w_000_4684, w_000_4685, w_000_4686, w_000_4687, w_000_4688, w_000_4689, w_000_4690, w_000_4691, w_000_4692, w_000_4693, w_000_4694, w_000_4695, w_000_4696, w_000_4697, w_000_4698, w_000_4699, w_000_4700, w_000_4701, w_000_4702, w_000_4703, w_000_4704, w_000_4705, w_000_4706, w_000_4707, w_000_4708, w_000_4709, w_000_4710, w_000_4711, w_000_4712, w_000_4713, w_000_4714, w_000_4715, w_000_4716, w_000_4717, w_000_4718, w_000_4719, w_000_4720, w_000_4721, w_000_4722, w_000_4723, w_000_4724, w_000_4725, w_000_4726, w_000_4727, w_000_4728, w_000_4729, w_000_4730, w_000_4731, w_000_4732, w_000_4733, w_000_4734, w_000_4735, w_000_4736, w_000_4737, w_000_4738, w_000_4739, w_000_4740, w_000_4741, w_000_4742, w_000_4743, w_000_4744, w_000_4745, w_000_4746, w_000_4747, w_000_4748, w_000_4749, w_000_4750, w_000_4751, w_000_4752, w_000_4753, w_000_4754, w_000_4755, w_000_4756, w_000_4757, w_000_4758, w_000_4759, w_000_4760, w_000_4761, w_000_4762, w_000_4763, w_000_4764, w_000_4765, w_000_4766, w_000_4767, w_000_4768, w_000_4769, w_000_4770, w_000_4771, w_000_4772, w_000_4773, w_000_4774, w_000_4775, w_000_4776, w_000_4777, w_000_4778, w_000_4779, w_000_4780, w_000_4781, w_000_4782, w_000_4783, w_000_4784, w_000_4785, w_000_4786, w_000_4787, w_000_4788, w_000_4789, w_000_4790, w_000_4791, w_000_4792, w_000_4793, w_000_4794, w_000_4795, w_000_4796, w_000_4797, w_000_4798, w_000_4799, w_000_4800, w_000_4801, w_000_4803, w_000_4804, w_000_4805, w_000_4806, w_000_4807, w_000_4808, w_000_4809, w_000_4810, w_000_4811, w_000_4812, w_000_4813, w_000_4814, w_000_4815, w_000_4816, w_000_4817, w_000_4818, w_000_4819, w_000_4820, w_000_4821, w_000_4822, w_000_4823, w_000_4824, w_000_4825, w_000_4826, w_000_4827, w_000_4828, w_000_4829, w_000_4830, w_000_4831, w_000_4832, w_000_4833, w_000_4834, w_000_4835, w_000_4836, w_000_4837, w_000_4838, w_000_4839, w_000_4840, w_000_4841, w_000_4842, w_000_4843, w_000_4844, w_000_4845, w_000_4846, w_000_4847, w_000_4848, w_000_4849, w_000_4850, w_000_4851, w_000_4852, w_000_4853, w_000_4854, w_000_4855, w_000_4856, w_000_4860, w_000_4861, w_000_4862, w_000_4863, w_000_4864, w_000_4865, w_000_4866, w_000_4867, w_000_4868, w_000_4869, w_000_4870, w_000_4871, w_000_4872, w_000_4873, w_000_4874, w_000_4875, w_000_4876, w_000_4877, w_000_4878, w_000_4879, w_000_4880, w_000_4881, w_000_4882, w_000_4883, w_000_4884, w_000_4885, w_000_4886, w_000_4887, w_000_4889, w_000_4890, w_000_4891, w_000_4892, w_000_4893, w_000_4894, w_000_4895, w_000_4896, w_000_4897, w_000_4898, w_000_4900, w_000_4901, w_000_4902, w_000_4903, w_000_4905, w_000_4906, w_000_4907, w_000_4908, w_000_4909, w_000_4910, w_000_4911, w_000_4912, w_000_4914, w_000_4915, w_000_4916, w_000_4917, w_000_4918, w_000_4920, w_000_4921, w_000_4922, w_000_4923, w_000_4924, w_000_4926, w_000_4927, w_000_4928, w_000_4929, w_000_4930, w_000_4931, w_000_4932, w_000_4933, w_000_4934, w_000_4935, w_000_4936, w_000_4937, w_000_4938, w_000_4939, w_000_4941, w_000_4942, w_000_4944, w_000_4945, w_000_4946, w_000_4947, w_000_4949, w_000_4950, w_000_4952, w_000_4953, w_000_4955, w_000_4956, w_000_4957, w_000_4958, w_000_4959, w_000_4963, w_000_4964, w_000_4966, w_000_4968, w_000_4969, w_000_4970, w_000_4974, w_000_4979, w_000_4980, w_000_4984, w_000_4990, w_000_4991, w_000_4994;
  wire w_001_000, w_001_001, w_001_002, w_001_003, w_001_004, w_001_005, w_001_006, w_001_007, w_001_008, w_001_009, w_001_010, w_001_011, w_001_012, w_001_013, w_001_014, w_001_015, w_001_016, w_001_017, w_001_018, w_001_019, w_001_020, w_001_021, w_001_022, w_001_023, w_001_024, w_001_025, w_001_026, w_001_027, w_001_028, w_001_029, w_001_030, w_001_031, w_001_032, w_001_033, w_001_034, w_001_035, w_001_036, w_001_037, w_001_038, w_001_039, w_001_040, w_001_041, w_001_042, w_001_043, w_001_044, w_001_045, w_001_046, w_001_047, w_001_048, w_001_049, w_001_050, w_001_051, w_001_052, w_001_053, w_001_054, w_001_055, w_001_056, w_001_057, w_001_058, w_001_059, w_001_060, w_001_061, w_001_062, w_001_063, w_001_064, w_001_065, w_001_066, w_001_067, w_001_068, w_001_069, w_001_070, w_001_071, w_001_072, w_001_073, w_001_074, w_001_075, w_001_076, w_001_077, w_001_078, w_001_079, w_001_080, w_001_081, w_001_082, w_001_083, w_001_084, w_001_085, w_001_086, w_001_087, w_001_088, w_001_089, w_001_090, w_001_091, w_001_092, w_001_093, w_001_094, w_001_095, w_001_096, w_001_097, w_001_098, w_001_099, w_001_100, w_001_101, w_001_102, w_001_103, w_001_104, w_001_105, w_001_106, w_001_107, w_001_108, w_001_109, w_001_110, w_001_111, w_001_112, w_001_113, w_001_114, w_001_115, w_001_116, w_001_117, w_001_118, w_001_119, w_001_120, w_001_121, w_001_122, w_001_123, w_001_124, w_001_125, w_001_126, w_001_127, w_001_128, w_001_129, w_001_130, w_001_131, w_001_132, w_001_133, w_001_134, w_001_135, w_001_136, w_001_137, w_001_138, w_001_139, w_001_140, w_001_141, w_001_142, w_001_143, w_001_144, w_001_145, w_001_146, w_001_147, w_001_148, w_001_149, w_001_150, w_001_151, w_001_152, w_001_153, w_001_154, w_001_155, w_001_156, w_001_157, w_001_158, w_001_159, w_001_160, w_001_161, w_001_162, w_001_163, w_001_164, w_001_165, w_001_166, w_001_167, w_001_168, w_001_169, w_001_170, w_001_171, w_001_172, w_001_173, w_001_174, w_001_175, w_001_176, w_001_177, w_001_178, w_001_179, w_001_180, w_001_181, w_001_182, w_001_183, w_001_184, w_001_185, w_001_186, w_001_187, w_001_188, w_001_189, w_001_190, w_001_191, w_001_192, w_001_193, w_001_194, w_001_195, w_001_196, w_001_197, w_001_198, w_001_199, w_001_200, w_001_201, w_001_202, w_001_203, w_001_204, w_001_205, w_001_206, w_001_207, w_001_208, w_001_209, w_001_210, w_001_211, w_001_212, w_001_213, w_001_214, w_001_215, w_001_216, w_001_217, w_001_218, w_001_219, w_001_220, w_001_221, w_001_222, w_001_223, w_001_224, w_001_225, w_001_226, w_001_227, w_001_228, w_001_229, w_001_230, w_001_231, w_001_232, w_001_233, w_001_234, w_001_235, w_001_236, w_001_237, w_001_238, w_001_239, w_001_240, w_001_241, w_001_242, w_001_243, w_001_244, w_001_245, w_001_246, w_001_247, w_001_248, w_001_249, w_001_250, w_001_251, w_001_252, w_001_253, w_001_254, w_001_255, w_001_256, w_001_257, w_001_258, w_001_259, w_001_260, w_001_261, w_001_262, w_001_263, w_001_264, w_001_265, w_001_266, w_001_267, w_001_268, w_001_269, w_001_270, w_001_271, w_001_272, w_001_273, w_001_274, w_001_275, w_001_276, w_001_277, w_001_278, w_001_279, w_001_280, w_001_281, w_001_282, w_001_283, w_001_284, w_001_285, w_001_286, w_001_287, w_001_288, w_001_289, w_001_290, w_001_291, w_001_292, w_001_293, w_001_294, w_001_295, w_001_296, w_001_297, w_001_298, w_001_299, w_001_300, w_001_301, w_001_302, w_001_303, w_001_304, w_001_305, w_001_306, w_001_307, w_001_308, w_001_309, w_001_310, w_001_311, w_001_312, w_001_313, w_001_314, w_001_315, w_001_316, w_001_317, w_001_318, w_001_319, w_001_320, w_001_321, w_001_322, w_001_323, w_001_324, w_001_325, w_001_326, w_001_327, w_001_328, w_001_329, w_001_330, w_001_331, w_001_332, w_001_333, w_001_334, w_001_335, w_001_336, w_001_337, w_001_338, w_001_339, w_001_340, w_001_341, w_001_342, w_001_343, w_001_344, w_001_345, w_001_346, w_001_347, w_001_348, w_001_349, w_001_350, w_001_351, w_001_352, w_001_353, w_001_354, w_001_355, w_001_356, w_001_357, w_001_358, w_001_359, w_001_360, w_001_361, w_001_362, w_001_363, w_001_364, w_001_365, w_001_366, w_001_367, w_001_368, w_001_369, w_001_370, w_001_371, w_001_372, w_001_373, w_001_374, w_001_375, w_001_376, w_001_377, w_001_378, w_001_379, w_001_380, w_001_381, w_001_382, w_001_383, w_001_384, w_001_385, w_001_386, w_001_387, w_001_388, w_001_389, w_001_390, w_001_391, w_001_392, w_001_393, w_001_394, w_001_395, w_001_396, w_001_397, w_001_398, w_001_399, w_001_400, w_001_401, w_001_402, w_001_403, w_001_404, w_001_405, w_001_406, w_001_407, w_001_408, w_001_409, w_001_410, w_001_411, w_001_412, w_001_413, w_001_414, w_001_415, w_001_416, w_001_417, w_001_418, w_001_419, w_001_420, w_001_421, w_001_422, w_001_423, w_001_424, w_001_425, w_001_426, w_001_427, w_001_428, w_001_429, w_001_430, w_001_431, w_001_432, w_001_433, w_001_434, w_001_435, w_001_436, w_001_437, w_001_438, w_001_439, w_001_440, w_001_441, w_001_442, w_001_443, w_001_444, w_001_445, w_001_446, w_001_447, w_001_448, w_001_449, w_001_450, w_001_451, w_001_453, w_001_454, w_001_455, w_001_456, w_001_457, w_001_458, w_001_459, w_001_460, w_001_461, w_001_462, w_001_463, w_001_464, w_001_465, w_001_466, w_001_467, w_001_468, w_001_469, w_001_470, w_001_471, w_001_472, w_001_473, w_001_474, w_001_475, w_001_476, w_001_477, w_001_478, w_001_479, w_001_480, w_001_481, w_001_482, w_001_483, w_001_484, w_001_485, w_001_486, w_001_487, w_001_488, w_001_489, w_001_490, w_001_491, w_001_492, w_001_493, w_001_494, w_001_495, w_001_496, w_001_497, w_001_498, w_001_499, w_001_500, w_001_501, w_001_502, w_001_503, w_001_504, w_001_505, w_001_506, w_001_507, w_001_508, w_001_509, w_001_510, w_001_511, w_001_512, w_001_513, w_001_514, w_001_515, w_001_516, w_001_517, w_001_518, w_001_519, w_001_520, w_001_521, w_001_522, w_001_523, w_001_524, w_001_525, w_001_526, w_001_527, w_001_528, w_001_529, w_001_530, w_001_531, w_001_532, w_001_533, w_001_534, w_001_535, w_001_536, w_001_537, w_001_538, w_001_539, w_001_540, w_001_541, w_001_542, w_001_543, w_001_544, w_001_545, w_001_546, w_001_547, w_001_548, w_001_549, w_001_550, w_001_551, w_001_552, w_001_553, w_001_554, w_001_555, w_001_556, w_001_557, w_001_558, w_001_559, w_001_560, w_001_561, w_001_562, w_001_563, w_001_564, w_001_565, w_001_566, w_001_567, w_001_568, w_001_569, w_001_570, w_001_571, w_001_572, w_001_573, w_001_574, w_001_575, w_001_576, w_001_577, w_001_578, w_001_579, w_001_580, w_001_581, w_001_582, w_001_583, w_001_584, w_001_585, w_001_586, w_001_587, w_001_588, w_001_589, w_001_590, w_001_591, w_001_592, w_001_593, w_001_594, w_001_595, w_001_596, w_001_597, w_001_598, w_001_599, w_001_600, w_001_601, w_001_602, w_001_603, w_001_604, w_001_605, w_001_606, w_001_607, w_001_608, w_001_609, w_001_610, w_001_611, w_001_612, w_001_613, w_001_614, w_001_615, w_001_616, w_001_617, w_001_618, w_001_619, w_001_620, w_001_621, w_001_622, w_001_623, w_001_624, w_001_625, w_001_626, w_001_627, w_001_628, w_001_629, w_001_630, w_001_631, w_001_632, w_001_633, w_001_634, w_001_635, w_001_636, w_001_637, w_001_638, w_001_639, w_001_640, w_001_641, w_001_642, w_001_643, w_001_644, w_001_645, w_001_646, w_001_647, w_001_648, w_001_649, w_001_650, w_001_651, w_001_652, w_001_653, w_001_654, w_001_655, w_001_656, w_001_657, w_001_658, w_001_659, w_001_660, w_001_661, w_001_662, w_001_663, w_001_664, w_001_665, w_001_666, w_001_667, w_001_668, w_001_669, w_001_670, w_001_671, w_001_672, w_001_673, w_001_674, w_001_675, w_001_676, w_001_677, w_001_678, w_001_679, w_001_680, w_001_681, w_001_682, w_001_683, w_001_684, w_001_685, w_001_686, w_001_687, w_001_688, w_001_689, w_001_690, w_001_691, w_001_692, w_001_693, w_001_694, w_001_695, w_001_696, w_001_697, w_001_698, w_001_699, w_001_700, w_001_701, w_001_702, w_001_703, w_001_704, w_001_705, w_001_706, w_001_707, w_001_708, w_001_709, w_001_710, w_001_711, w_001_712, w_001_713, w_001_714, w_001_715, w_001_716, w_001_717, w_001_718, w_001_719, w_001_720, w_001_721, w_001_722, w_001_723, w_001_724, w_001_725, w_001_726, w_001_727, w_001_728, w_001_729, w_001_730, w_001_731, w_001_732, w_001_733, w_001_734, w_001_735, w_001_736, w_001_737, w_001_738, w_001_739, w_001_740, w_001_741, w_001_742, w_001_743, w_001_744, w_001_745, w_001_746, w_001_747, w_001_748, w_001_749, w_001_750, w_001_751, w_001_752, w_001_753, w_001_754, w_001_755, w_001_756, w_001_757, w_001_758, w_001_759, w_001_760, w_001_761, w_001_762, w_001_763, w_001_764, w_001_765, w_001_766, w_001_767, w_001_768, w_001_769, w_001_770, w_001_771, w_001_772, w_001_773, w_001_774, w_001_775, w_001_776, w_001_777, w_001_778, w_001_779, w_001_780, w_001_781, w_001_782, w_001_783, w_001_784, w_001_785, w_001_786, w_001_787, w_001_788, w_001_789, w_001_790, w_001_791, w_001_792, w_001_793, w_001_794, w_001_795, w_001_796, w_001_797, w_001_798, w_001_799, w_001_800, w_001_801, w_001_802, w_001_803, w_001_804, w_001_805, w_001_806, w_001_807, w_001_808, w_001_809, w_001_810, w_001_811, w_001_812, w_001_813, w_001_814, w_001_815, w_001_816, w_001_817, w_001_818, w_001_819, w_001_820, w_001_821, w_001_822, w_001_823, w_001_824, w_001_825, w_001_826, w_001_827, w_001_828, w_001_829, w_001_830, w_001_831, w_001_832, w_001_833, w_001_834, w_001_835, w_001_836, w_001_837, w_001_838, w_001_839, w_001_840, w_001_841, w_001_842, w_001_843, w_001_844, w_001_845, w_001_846, w_001_847, w_001_848, w_001_849, w_001_850, w_001_851, w_001_852, w_001_853, w_001_854, w_001_855, w_001_856, w_001_857, w_001_858, w_001_859, w_001_860, w_001_861, w_001_862, w_001_863, w_001_864, w_001_865, w_001_866, w_001_867, w_001_868, w_001_869, w_001_870, w_001_871, w_001_872, w_001_873, w_001_874, w_001_875, w_001_876, w_001_877, w_001_878, w_001_879, w_001_880, w_001_881, w_001_882, w_001_883, w_001_884, w_001_885, w_001_886, w_001_887, w_001_888, w_001_889, w_001_890, w_001_891, w_001_892, w_001_893, w_001_894, w_001_895, w_001_896, w_001_897, w_001_898, w_001_899, w_001_900, w_001_901, w_001_902, w_001_903, w_001_904, w_001_905, w_001_906, w_001_907, w_001_908, w_001_909, w_001_910, w_001_911, w_001_912, w_001_913, w_001_914, w_001_915, w_001_916, w_001_917, w_001_918, w_001_919, w_001_920, w_001_921, w_001_922, w_001_923, w_001_924, w_001_925, w_001_926, w_001_927, w_001_928, w_001_929, w_001_930, w_001_931, w_001_932, w_001_933, w_001_934, w_001_935, w_001_936, w_001_937, w_001_938, w_001_939, w_001_940, w_001_941, w_001_942, w_001_943, w_001_944, w_001_945, w_001_946, w_001_947, w_001_948, w_001_949, w_001_950, w_001_951, w_001_952, w_001_953, w_001_954, w_001_955, w_001_956, w_001_957, w_001_958, w_001_959, w_001_960, w_001_961, w_001_962, w_001_963, w_001_964, w_001_965, w_001_966, w_001_967, w_001_968, w_001_969, w_001_970, w_001_971, w_001_972, w_001_973, w_001_974, w_001_975, w_001_976, w_001_977, w_001_978, w_001_979, w_001_980, w_001_981, w_001_982, w_001_983, w_001_984, w_001_985, w_001_986, w_001_987, w_001_988, w_001_989, w_001_990, w_001_991, w_001_992, w_001_993, w_001_994, w_001_995, w_001_996, w_001_997, w_001_998, w_001_999, w_001_1000, w_001_1001, w_001_1002, w_001_1003, w_001_1004, w_001_1005, w_001_1006, w_001_1007, w_001_1008, w_001_1009, w_001_1010, w_001_1011, w_001_1012, w_001_1013, w_001_1014, w_001_1015, w_001_1016, w_001_1017, w_001_1018, w_001_1019, w_001_1020, w_001_1021, w_001_1022, w_001_1023, w_001_1024, w_001_1025, w_001_1026, w_001_1027, w_001_1028, w_001_1029, w_001_1030, w_001_1031, w_001_1032, w_001_1033, w_001_1034, w_001_1035, w_001_1036, w_001_1037, w_001_1038, w_001_1039, w_001_1040, w_001_1041, w_001_1042, w_001_1043, w_001_1044, w_001_1045, w_001_1046, w_001_1047, w_001_1048, w_001_1049, w_001_1050, w_001_1051, w_001_1052, w_001_1053, w_001_1054, w_001_1055, w_001_1056, w_001_1057, w_001_1058, w_001_1059, w_001_1060, w_001_1061, w_001_1062, w_001_1063, w_001_1064, w_001_1065, w_001_1066, w_001_1067, w_001_1068, w_001_1069, w_001_1070, w_001_1071, w_001_1072, w_001_1073, w_001_1074, w_001_1075, w_001_1076, w_001_1077, w_001_1078, w_001_1079, w_001_1080, w_001_1081, w_001_1082, w_001_1083, w_001_1084, w_001_1085, w_001_1086, w_001_1087, w_001_1088, w_001_1089, w_001_1090, w_001_1091, w_001_1092, w_001_1093, w_001_1094, w_001_1095, w_001_1096, w_001_1097, w_001_1098, w_001_1099, w_001_1100, w_001_1101, w_001_1102, w_001_1103, w_001_1104, w_001_1105, w_001_1106, w_001_1107, w_001_1108, w_001_1109, w_001_1110, w_001_1111, w_001_1112, w_001_1113, w_001_1114, w_001_1115, w_001_1116, w_001_1117, w_001_1118, w_001_1119, w_001_1120, w_001_1121, w_001_1122, w_001_1123, w_001_1124, w_001_1125, w_001_1126, w_001_1127, w_001_1128, w_001_1129, w_001_1130, w_001_1131, w_001_1132, w_001_1133, w_001_1134, w_001_1135, w_001_1136, w_001_1137, w_001_1138, w_001_1139, w_001_1140, w_001_1141, w_001_1142, w_001_1143, w_001_1144, w_001_1145, w_001_1146, w_001_1147, w_001_1148, w_001_1149, w_001_1150, w_001_1151, w_001_1152, w_001_1153, w_001_1154, w_001_1155, w_001_1156, w_001_1157, w_001_1158, w_001_1159, w_001_1160, w_001_1161, w_001_1162, w_001_1163, w_001_1164, w_001_1165, w_001_1166, w_001_1167, w_001_1168, w_001_1169, w_001_1170, w_001_1171, w_001_1172, w_001_1173, w_001_1174, w_001_1175, w_001_1176, w_001_1177, w_001_1178, w_001_1179, w_001_1180, w_001_1181, w_001_1182, w_001_1183, w_001_1184, w_001_1185, w_001_1186, w_001_1187, w_001_1188, w_001_1189, w_001_1190, w_001_1191, w_001_1192, w_001_1193, w_001_1194, w_001_1195, w_001_1196, w_001_1197, w_001_1198, w_001_1199, w_001_1200, w_001_1201, w_001_1202, w_001_1203, w_001_1204, w_001_1205, w_001_1206, w_001_1207, w_001_1208, w_001_1209, w_001_1210, w_001_1211, w_001_1212, w_001_1213, w_001_1214, w_001_1215, w_001_1216, w_001_1217, w_001_1218, w_001_1219, w_001_1220, w_001_1221, w_001_1222, w_001_1224, w_001_1225, w_001_1226, w_001_1227, w_001_1228, w_001_1229, w_001_1230, w_001_1231, w_001_1232, w_001_1233, w_001_1234, w_001_1235, w_001_1236, w_001_1237, w_001_1238, w_001_1239, w_001_1240, w_001_1241, w_001_1242, w_001_1243, w_001_1244, w_001_1245, w_001_1246, w_001_1247, w_001_1248, w_001_1249, w_001_1250, w_001_1251, w_001_1252, w_001_1253, w_001_1254, w_001_1255, w_001_1256, w_001_1257, w_001_1258, w_001_1259, w_001_1260, w_001_1261, w_001_1262, w_001_1263, w_001_1264, w_001_1265, w_001_1266, w_001_1267, w_001_1268, w_001_1269, w_001_1270, w_001_1271, w_001_1272, w_001_1273, w_001_1274, w_001_1275, w_001_1276, w_001_1277, w_001_1278, w_001_1279, w_001_1280, w_001_1281, w_001_1282, w_001_1283, w_001_1284, w_001_1285, w_001_1286, w_001_1287, w_001_1288, w_001_1289, w_001_1290, w_001_1291, w_001_1292, w_001_1293, w_001_1294, w_001_1295, w_001_1296, w_001_1297, w_001_1298, w_001_1299, w_001_1300, w_001_1301, w_001_1302, w_001_1303, w_001_1304, w_001_1305, w_001_1306, w_001_1307, w_001_1308, w_001_1309, w_001_1310, w_001_1311, w_001_1312, w_001_1313, w_001_1314, w_001_1315, w_001_1316, w_001_1317, w_001_1318, w_001_1319, w_001_1320, w_001_1321, w_001_1322, w_001_1323, w_001_1324, w_001_1325, w_001_1326, w_001_1327, w_001_1328, w_001_1329, w_001_1330, w_001_1331, w_001_1332, w_001_1333, w_001_1334, w_001_1335, w_001_1336, w_001_1337, w_001_1338, w_001_1339, w_001_1340, w_001_1341, w_001_1342, w_001_1343, w_001_1344, w_001_1345, w_001_1346, w_001_1347, w_001_1348, w_001_1349, w_001_1350, w_001_1351, w_001_1352, w_001_1353, w_001_1354, w_001_1355, w_001_1356, w_001_1357, w_001_1358, w_001_1359, w_001_1360, w_001_1361, w_001_1362, w_001_1363, w_001_1364, w_001_1365, w_001_1366, w_001_1367, w_001_1368, w_001_1369, w_001_1370, w_001_1371, w_001_1372, w_001_1373, w_001_1374, w_001_1375, w_001_1376, w_001_1377, w_001_1378, w_001_1379, w_001_1380, w_001_1381, w_001_1382, w_001_1383, w_001_1384, w_001_1385, w_001_1386, w_001_1387, w_001_1388, w_001_1389, w_001_1390, w_001_1391, w_001_1392, w_001_1393, w_001_1394, w_001_1395, w_001_1396, w_001_1397, w_001_1398, w_001_1399, w_001_1400, w_001_1401, w_001_1402, w_001_1403, w_001_1404, w_001_1405, w_001_1406, w_001_1407, w_001_1408, w_001_1409, w_001_1410, w_001_1411, w_001_1412, w_001_1413, w_001_1414, w_001_1415, w_001_1416, w_001_1417, w_001_1418, w_001_1419, w_001_1420, w_001_1422, w_001_1423, w_001_1424, w_001_1425, w_001_1426, w_001_1427, w_001_1428, w_001_1429, w_001_1431, w_001_1432, w_001_1433, w_001_1434, w_001_1436, w_001_1437, w_001_1438, w_001_1439, w_001_1440, w_001_1441, w_001_1442, w_001_1443, w_001_1444, w_001_1445, w_001_1446, w_001_1447, w_001_1448, w_001_1449, w_001_1450, w_001_1451, w_001_1452, w_001_1453, w_001_1454, w_001_1455, w_001_1456, w_001_1457, w_001_1458, w_001_1459, w_001_1460, w_001_1461, w_001_1462, w_001_1463, w_001_1464, w_001_1465, w_001_1466, w_001_1467, w_001_1468, w_001_1469, w_001_1470, w_001_1471, w_001_1472, w_001_1473, w_001_1474, w_001_1475, w_001_1476, w_001_1477, w_001_1478, w_001_1479, w_001_1480, w_001_1481, w_001_1482, w_001_1483, w_001_1485, w_001_1486, w_001_1487, w_001_1488, w_001_1489, w_001_1490, w_001_1491, w_001_1492, w_001_1493, w_001_1494, w_001_1495, w_001_1496, w_001_1497, w_001_1498, w_001_1499, w_001_1500, w_001_1501, w_001_1502, w_001_1503, w_001_1504, w_001_1505, w_001_1506, w_001_1507, w_001_1508, w_001_1509, w_001_1510, w_001_1511, w_001_1512, w_001_1513, w_001_1514, w_001_1515, w_001_1516, w_001_1517, w_001_1518, w_001_1519, w_001_1520, w_001_1521, w_001_1522, w_001_1523, w_001_1524, w_001_1525, w_001_1526, w_001_1527, w_001_1528, w_001_1529, w_001_1530, w_001_1531, w_001_1532, w_001_1533, w_001_1534, w_001_1535, w_001_1536, w_001_1537, w_001_1538, w_001_1539, w_001_1540, w_001_1541, w_001_1542, w_001_1543, w_001_1544, w_001_1545, w_001_1546, w_001_1547, w_001_1548, w_001_1549, w_001_1550, w_001_1552, w_001_1553, w_001_1554, w_001_1555, w_001_1556, w_001_1557, w_001_1558, w_001_1559, w_001_1560, w_001_1561, w_001_1562, w_001_1563, w_001_1564, w_001_1565, w_001_1566, w_001_1567, w_001_1568, w_001_1569, w_001_1570, w_001_1571, w_001_1572, w_001_1574, w_001_1575, w_001_1576, w_001_1577, w_001_1578, w_001_1579, w_001_1580, w_001_1581, w_001_1582, w_001_1583, w_001_1584, w_001_1585, w_001_1586, w_001_1587, w_001_1588, w_001_1589, w_001_1590, w_001_1591, w_001_1592, w_001_1593, w_001_1594, w_001_1595, w_001_1597, w_001_1598, w_001_1599, w_001_1600, w_001_1601, w_001_1602, w_001_1603, w_001_1604, w_001_1605, w_001_1606, w_001_1607, w_001_1608, w_001_1609, w_001_1610, w_001_1611, w_001_1612, w_001_1613, w_001_1614, w_001_1616, w_001_1617, w_001_1618, w_001_1619, w_001_1621, w_001_1622, w_001_1623, w_001_1624, w_001_1625, w_001_1626, w_001_1627, w_001_1628, w_001_1629, w_001_1630, w_001_1631, w_001_1632, w_001_1633, w_001_1634, w_001_1635, w_001_1637, w_001_1638, w_001_1639, w_001_1640, w_001_1641, w_001_1642, w_001_1643, w_001_1644, w_001_1645, w_001_1646, w_001_1647, w_001_1648, w_001_1649, w_001_1650, w_001_1652, w_001_1653, w_001_1654, w_001_1655, w_001_1656, w_001_1657, w_001_1658, w_001_1659, w_001_1660, w_001_1661, w_001_1662, w_001_1663, w_001_1664, w_001_1665, w_001_1666, w_001_1667, w_001_1668, w_001_1669, w_001_1670, w_001_1671, w_001_1672, w_001_1674, w_001_1675, w_001_1676, w_001_1677, w_001_1678, w_001_1679, w_001_1680, w_001_1681, w_001_1682, w_001_1683, w_001_1684, w_001_1685, w_001_1686, w_001_1687, w_001_1688, w_001_1689, w_001_1690, w_001_1691, w_001_1692, w_001_1693, w_001_1694, w_001_1696, w_001_1697, w_001_1699, w_001_1700, w_001_1701, w_001_1702, w_001_1703, w_001_1704, w_001_1705, w_001_1706, w_001_1707, w_001_1708, w_001_1709, w_001_1710, w_001_1711, w_001_1712, w_001_1713, w_001_1715, w_001_1716, w_001_1717, w_001_1718, w_001_1719, w_001_1720, w_001_1721, w_001_1722, w_001_1723, w_001_1725, w_001_1726, w_001_1727, w_001_1728, w_001_1729, w_001_1730, w_001_1731, w_001_1732, w_001_1733, w_001_1734, w_001_1735, w_001_1736, w_001_1737, w_001_1738, w_001_1739, w_001_1740, w_001_1741, w_001_1742, w_001_1743, w_001_1744, w_001_1745, w_001_1746, w_001_1747, w_001_1748, w_001_1749, w_001_1750, w_001_1751, w_001_1752, w_001_1753, w_001_1754, w_001_1755, w_001_1756, w_001_1757, w_001_1758, w_001_1759, w_001_1760, w_001_1761, w_001_1763, w_001_1764, w_001_1765, w_001_1766, w_001_1767, w_001_1768, w_001_1769, w_001_1770, w_001_1771, w_001_1772, w_001_1773, w_001_1774, w_001_1775, w_001_1776, w_001_1777, w_001_1778, w_001_1779, w_001_1781, w_001_1782, w_001_1783, w_001_1784, w_001_1785, w_001_1786, w_001_1787, w_001_1788, w_001_1789, w_001_1790, w_001_1791, w_001_1792, w_001_1793, w_001_1794, w_001_1795, w_001_1796, w_001_1797, w_001_1798, w_001_1799, w_001_1800, w_001_1801, w_001_1802, w_001_1805, w_001_1806, w_001_1807, w_001_1808, w_001_1809, w_001_1810, w_001_1811, w_001_1812, w_001_1813, w_001_1814, w_001_1815, w_001_1816, w_001_1817, w_001_1818, w_001_1819, w_001_1820, w_001_1821, w_001_1822, w_001_1823, w_001_1824, w_001_1825, w_001_1826, w_001_1827, w_001_1828, w_001_1829, w_001_1830, w_001_1831, w_001_1832, w_001_1833, w_001_1834, w_001_1835, w_001_1836, w_001_1837, w_001_1838, w_001_1839, w_001_1840, w_001_1841, w_001_1842, w_001_1843, w_001_1844, w_001_1845, w_001_1846, w_001_1847, w_001_1848, w_001_1849, w_001_1850, w_001_1851, w_001_1852, w_001_1853, w_001_1854, w_001_1855, w_001_1856, w_001_1857, w_001_1858, w_001_1859, w_001_1860, w_001_1861, w_001_1862, w_001_1863, w_001_1864, w_001_1865, w_001_1866, w_001_1867, w_001_1868, w_001_1869, w_001_1870, w_001_1871, w_001_1872, w_001_1873, w_001_1874, w_001_1875, w_001_1876, w_001_1877, w_001_1878, w_001_1879, w_001_1880, w_001_1881, w_001_1882, w_001_1884, w_001_1885, w_001_1886, w_001_1887, w_001_1888, w_001_1889, w_001_1890, w_001_1891, w_001_1892, w_001_1893, w_001_1894, w_001_1895, w_001_1896, w_001_1897, w_001_1898, w_001_1899, w_001_1900, w_001_1901, w_001_1903, w_001_1904, w_001_1905, w_001_1906, w_001_1907, w_001_1909, w_001_1910, w_001_1911, w_001_1913, w_001_1914, w_001_1915, w_001_1916, w_001_1917, w_001_1918, w_001_1919, w_001_1920, w_001_1921, w_001_1922, w_001_1923, w_001_1924, w_001_1925, w_001_1926, w_001_1927, w_001_1928, w_001_1929, w_001_1930, w_001_1931, w_001_1932, w_001_1933, w_001_1934, w_001_1935, w_001_1936, w_001_1937, w_001_1938, w_001_1939, w_001_1941, w_001_1942, w_001_1943, w_001_1944, w_001_1945, w_001_1946, w_001_1947, w_001_1948, w_001_1949, w_001_1950, w_001_1951, w_001_1952, w_001_1953, w_001_1954, w_001_1955, w_001_1956, w_001_1957, w_001_1958, w_001_1959, w_001_1960, w_001_1961, w_001_1962, w_001_1963, w_001_1964, w_001_1965, w_001_1966, w_001_1967, w_001_1968, w_001_1969, w_001_1970, w_001_1971, w_001_1972, w_001_1973, w_001_1974, w_001_1975, w_001_1976, w_001_1977, w_001_1978, w_001_1979, w_001_1980, w_001_1981, w_001_1982, w_001_1984, w_001_1985, w_001_1986, w_001_1987, w_001_1988, w_001_1989, w_001_1990, w_001_1991, w_001_1992, w_001_1993, w_001_1994, w_001_1995, w_001_1996, w_001_1997, w_001_1999, w_001_2000, w_001_2001, w_001_2002, w_001_2003, w_001_2004, w_001_2005, w_001_2006, w_001_2007, w_001_2008, w_001_2009, w_001_2010, w_001_2011, w_001_2012, w_001_2013, w_001_2014, w_001_2015, w_001_2016, w_001_2017, w_001_2018, w_001_2019, w_001_2020, w_001_2021, w_001_2022, w_001_2023, w_001_2024, w_001_2025, w_001_2026, w_001_2027, w_001_2028, w_001_2029, w_001_2030, w_001_2031, w_001_2032, w_001_2033, w_001_2034, w_001_2035, w_001_2036, w_001_2037, w_001_2038, w_001_2039, w_001_2040, w_001_2041, w_001_2042, w_001_2043, w_001_2044, w_001_2045, w_001_2046, w_001_2047, w_001_2048, w_001_2049, w_001_2050, w_001_2051, w_001_2052, w_001_2054, w_001_2055, w_001_2056, w_001_2057, w_001_2058, w_001_2059, w_001_2060, w_001_2061, w_001_2062, w_001_2063, w_001_2064, w_001_2065, w_001_2066, w_001_2067, w_001_2068, w_001_2069, w_001_2070, w_001_2071, w_001_2072, w_001_2073, w_001_2074, w_001_2075, w_001_2076, w_001_2077, w_001_2078, w_001_2079, w_001_2080, w_001_2081, w_001_2082, w_001_2083, w_001_2084, w_001_2085, w_001_2086, w_001_2087, w_001_2088, w_001_2089, w_001_2090, w_001_2091, w_001_2092, w_001_2093, w_001_2094, w_001_2095, w_001_2096, w_001_2097, w_001_2098, w_001_2099, w_001_2100, w_001_2101, w_001_2102, w_001_2103, w_001_2105, w_001_2106, w_001_2107, w_001_2108, w_001_2109, w_001_2111, w_001_2112, w_001_2113, w_001_2114, w_001_2115, w_001_2116, w_001_2117, w_001_2118, w_001_2119, w_001_2120, w_001_2122, w_001_2123, w_001_2124, w_001_2125, w_001_2126, w_001_2127, w_001_2128, w_001_2129, w_001_2130, w_001_2131, w_001_2132, w_001_2133, w_001_2134, w_001_2135, w_001_2138, w_001_2139, w_001_2140, w_001_2141, w_001_2142, w_001_2143, w_001_2144, w_001_2145, w_001_2146, w_001_2147, w_001_2148, w_001_2149, w_001_2150, w_001_2151, w_001_2152, w_001_2153, w_001_2154, w_001_2155, w_001_2156, w_001_2157, w_001_2158, w_001_2159, w_001_2160, w_001_2161, w_001_2162, w_001_2163, w_001_2164, w_001_2165, w_001_2166, w_001_2167, w_001_2168, w_001_2169, w_001_2170, w_001_2171, w_001_2172, w_001_2173, w_001_2174, w_001_2175, w_001_2177, w_001_2178, w_001_2180, w_001_2181, w_001_2182, w_001_2183, w_001_2184, w_001_2185, w_001_2186, w_001_2187, w_001_2188, w_001_2189, w_001_2190, w_001_2191, w_001_2192, w_001_2193, w_001_2194, w_001_2195, w_001_2196, w_001_2197, w_001_2198, w_001_2199, w_001_2200, w_001_2201, w_001_2202, w_001_2203, w_001_2204, w_001_2205, w_001_2206, w_001_2207, w_001_2208, w_001_2209, w_001_2210, w_001_2211, w_001_2212, w_001_2213, w_001_2214, w_001_2215, w_001_2216, w_001_2217, w_001_2218, w_001_2219, w_001_2220, w_001_2221, w_001_2222, w_001_2223, w_001_2224, w_001_2225, w_001_2226, w_001_2227, w_001_2228, w_001_2229, w_001_2230, w_001_2232, w_001_2233, w_001_2234, w_001_2235, w_001_2236, w_001_2237, w_001_2238, w_001_2239, w_001_2240, w_001_2241, w_001_2242, w_001_2243, w_001_2244, w_001_2245, w_001_2246, w_001_2247, w_001_2248, w_001_2250, w_001_2252, w_001_2253, w_001_2254, w_001_2255, w_001_2256, w_001_2258, w_001_2259, w_001_2260, w_001_2261, w_001_2262, w_001_2263, w_001_2264, w_001_2265, w_001_2266, w_001_2267, w_001_2268, w_001_2270, w_001_2271, w_001_2272, w_001_2273, w_001_2274, w_001_2275, w_001_2276, w_001_2277, w_001_2279, w_001_2280, w_001_2281, w_001_2282, w_001_2283, w_001_2284, w_001_2285, w_001_2287, w_001_2288, w_001_2289, w_001_2290, w_001_2291, w_001_2292, w_001_2293, w_001_2294, w_001_2295, w_001_2296, w_001_2297, w_001_2298, w_001_2299, w_001_2300, w_001_2301, w_001_2302, w_001_2303, w_001_2304, w_001_2305, w_001_2306, w_001_2307, w_001_2308, w_001_2309, w_001_2310, w_001_2311, w_001_2312, w_001_2313, w_001_2315, w_001_2316, w_001_2317, w_001_2318, w_001_2319, w_001_2320, w_001_2321, w_001_2322, w_001_2323, w_001_2324, w_001_2325, w_001_2326, w_001_2327, w_001_2328, w_001_2329, w_001_2330, w_001_2331, w_001_2332, w_001_2333, w_001_2334, w_001_2335, w_001_2336, w_001_2337, w_001_2338, w_001_2339, w_001_2340, w_001_2341, w_001_2342, w_001_2343, w_001_2344, w_001_2345, w_001_2346, w_001_2347, w_001_2348, w_001_2349, w_001_2350, w_001_2351, w_001_2352, w_001_2353, w_001_2355, w_001_2356, w_001_2357, w_001_2358, w_001_2359, w_001_2360, w_001_2361, w_001_2362, w_001_2363, w_001_2364, w_001_2365, w_001_2366, w_001_2367, w_001_2369, w_001_2370, w_001_2371, w_001_2372, w_001_2373, w_001_2374, w_001_2377, w_001_2378, w_001_2379, w_001_2380, w_001_2381, w_001_2382, w_001_2383, w_001_2384, w_001_2385, w_001_2386, w_001_2387, w_001_2388, w_001_2389, w_001_2390, w_001_2391, w_001_2392, w_001_2393, w_001_2394, w_001_2395, w_001_2396, w_001_2397, w_001_2398, w_001_2399, w_001_2400, w_001_2401, w_001_2402, w_001_2403, w_001_2404, w_001_2405, w_001_2406, w_001_2407, w_001_2408, w_001_2409, w_001_2410, w_001_2411, w_001_2412, w_001_2413, w_001_2414, w_001_2415, w_001_2416, w_001_2417, w_001_2418, w_001_2419, w_001_2420, w_001_2421, w_001_2422, w_001_2423, w_001_2424, w_001_2425, w_001_2426, w_001_2427, w_001_2428, w_001_2429, w_001_2430, w_001_2431, w_001_2432, w_001_2433, w_001_2434, w_001_2435, w_001_2436, w_001_2437, w_001_2438, w_001_2439, w_001_2440, w_001_2441, w_001_2442, w_001_2443, w_001_2444, w_001_2445, w_001_2446, w_001_2447, w_001_2448, w_001_2449, w_001_2450, w_001_2451, w_001_2452, w_001_2453, w_001_2454, w_001_2455, w_001_2456, w_001_2457, w_001_2458, w_001_2459, w_001_2460, w_001_2461, w_001_2462, w_001_2463, w_001_2464, w_001_2465, w_001_2466, w_001_2467, w_001_2468, w_001_2469, w_001_2470, w_001_2471, w_001_2472, w_001_2473, w_001_2474, w_001_2475, w_001_2476, w_001_2477, w_001_2478, w_001_2479, w_001_2480, w_001_2481, w_001_2482, w_001_2483, w_001_2484, w_001_2485, w_001_2486, w_001_2487, w_001_2488, w_001_2489, w_001_2490, w_001_2491, w_001_2492, w_001_2493, w_001_2494, w_001_2495, w_001_2496, w_001_2497, w_001_2498, w_001_2499, w_001_2500, w_001_2501, w_001_2502, w_001_2503, w_001_2504, w_001_2505, w_001_2506, w_001_2507, w_001_2508, w_001_2509, w_001_2510, w_001_2511, w_001_2512, w_001_2513, w_001_2514, w_001_2515, w_001_2516, w_001_2517, w_001_2518, w_001_2519, w_001_2520, w_001_2521, w_001_2522, w_001_2523, w_001_2524, w_001_2525, w_001_2526, w_001_2527, w_001_2528, w_001_2529, w_001_2530, w_001_2531, w_001_2532, w_001_2533, w_001_2534, w_001_2535, w_001_2536, w_001_2537, w_001_2538, w_001_2539, w_001_2540, w_001_2541, w_001_2542, w_001_2543, w_001_2544, w_001_2545, w_001_2546, w_001_2547, w_001_2548, w_001_2549, w_001_2550, w_001_2551, w_001_2552, w_001_2553, w_001_2554, w_001_2555, w_001_2556, w_001_2557, w_001_2558, w_001_2559, w_001_2560, w_001_2561, w_001_2562, w_001_2563, w_001_2564, w_001_2565, w_001_2566, w_001_2567, w_001_2568, w_001_2569, w_001_2571, w_001_2572, w_001_2573, w_001_2574, w_001_2575, w_001_2576, w_001_2577, w_001_2579, w_001_2580, w_001_2581, w_001_2584, w_001_2585, w_001_2586, w_001_2587, w_001_2588, w_001_2589, w_001_2590, w_001_2591, w_001_2592, w_001_2593, w_001_2594, w_001_2595, w_001_2596, w_001_2597, w_001_2598, w_001_2599, w_001_2600, w_001_2601, w_001_2602, w_001_2603, w_001_2604, w_001_2605, w_001_2606, w_001_2608, w_001_2609, w_001_2610, w_001_2611, w_001_2612, w_001_2613, w_001_2614, w_001_2615, w_001_2616, w_001_2617, w_001_2618, w_001_2619, w_001_2620, w_001_2621, w_001_2622, w_001_2623, w_001_2624, w_001_2625, w_001_2626, w_001_2627, w_001_2628, w_001_2629, w_001_2630, w_001_2631, w_001_2632, w_001_2633, w_001_2634, w_001_2635, w_001_2636, w_001_2637, w_001_2638, w_001_2639, w_001_2640, w_001_2641, w_001_2642, w_001_2643, w_001_2644, w_001_2645, w_001_2646, w_001_2647, w_001_2648, w_001_2649, w_001_2650, w_001_2651, w_001_2652, w_001_2653, w_001_2654, w_001_2655, w_001_2656, w_001_2657, w_001_2658, w_001_2659, w_001_2660, w_001_2661, w_001_2662, w_001_2663, w_001_2664, w_001_2665, w_001_2666, w_001_2667, w_001_2668, w_001_2669, w_001_2670, w_001_2671, w_001_2672, w_001_2673, w_001_2674, w_001_2675, w_001_2676, w_001_2677, w_001_2678, w_001_2679, w_001_2681, w_001_2682, w_001_2683, w_001_2684, w_001_2685, w_001_2686, w_001_2687, w_001_2688, w_001_2689, w_001_2690, w_001_2691, w_001_2692, w_001_2693, w_001_2694, w_001_2695, w_001_2696, w_001_2697, w_001_2698, w_001_2699, w_001_2700, w_001_2701, w_001_2702, w_001_2703, w_001_2704, w_001_2705, w_001_2706, w_001_2707, w_001_2708, w_001_2709, w_001_2710, w_001_2711, w_001_2712, w_001_2713, w_001_2715, w_001_2716, w_001_2717, w_001_2718, w_001_2719, w_001_2720, w_001_2721, w_001_2722, w_001_2723, w_001_2724, w_001_2725, w_001_2727, w_001_2728, w_001_2729, w_001_2730, w_001_2731, w_001_2732, w_001_2733, w_001_2734, w_001_2735, w_001_2736, w_001_2737, w_001_2738, w_001_2739, w_001_2740, w_001_2741, w_001_2742, w_001_2743, w_001_2744, w_001_2745, w_001_2746, w_001_2747, w_001_2748, w_001_2749, w_001_2750, w_001_2751, w_001_2752, w_001_2754, w_001_2755, w_001_2756, w_001_2757, w_001_2758, w_001_2759, w_001_2760, w_001_2761, w_001_2762, w_001_2763, w_001_2764, w_001_2765, w_001_2766, w_001_2767, w_001_2768, w_001_2769, w_001_2770, w_001_2771, w_001_2772, w_001_2773, w_001_2774, w_001_2775, w_001_2776, w_001_2777, w_001_2778, w_001_2779, w_001_2780, w_001_2781, w_001_2782, w_001_2783, w_001_2784, w_001_2785, w_001_2786, w_001_2787, w_001_2788, w_001_2789, w_001_2790, w_001_2791, w_001_2792, w_001_2793, w_001_2794, w_001_2795, w_001_2796, w_001_2797, w_001_2798, w_001_2799, w_001_2800, w_001_2801, w_001_2802, w_001_2804, w_001_2805, w_001_2806, w_001_2807, w_001_2808, w_001_2809, w_001_2810, w_001_2811, w_001_2812, w_001_2813, w_001_2814, w_001_2815, w_001_2816, w_001_2817, w_001_2818, w_001_2819, w_001_2820, w_001_2821, w_001_2822, w_001_2823, w_001_2824, w_001_2825, w_001_2826, w_001_2827, w_001_2828, w_001_2829, w_001_2830, w_001_2831, w_001_2832, w_001_2833, w_001_2834, w_001_2835, w_001_2836, w_001_2837, w_001_2838, w_001_2839, w_001_2840, w_001_2841, w_001_2842, w_001_2843, w_001_2845, w_001_2846, w_001_2847, w_001_2848, w_001_2849, w_001_2850, w_001_2851, w_001_2852, w_001_2853, w_001_2854, w_001_2855, w_001_2856, w_001_2857, w_001_2858, w_001_2859, w_001_2860, w_001_2861, w_001_2862, w_001_2863, w_001_2864, w_001_2865, w_001_2866, w_001_2867, w_001_2868, w_001_2869, w_001_2870, w_001_2871, w_001_2872, w_001_2873, w_001_2874, w_001_2875, w_001_2877, w_001_2878, w_001_2879, w_001_2880, w_001_2881, w_001_2882, w_001_2883, w_001_2884, w_001_2885, w_001_2886, w_001_2887, w_001_2888, w_001_2889, w_001_2890, w_001_2891, w_001_2892, w_001_2894, w_001_2895, w_001_2896, w_001_2897, w_001_2898, w_001_2899, w_001_2900, w_001_2901, w_001_2902, w_001_2903, w_001_2904, w_001_2905, w_001_2906, w_001_2907, w_001_2908, w_001_2909, w_001_2910, w_001_2911, w_001_2912, w_001_2913, w_001_2914, w_001_2915, w_001_2916, w_001_2917, w_001_2918, w_001_2919, w_001_2920, w_001_2921, w_001_2922, w_001_2923, w_001_2924, w_001_2925, w_001_2926, w_001_2927, w_001_2928, w_001_2929, w_001_2930, w_001_2931, w_001_2932, w_001_2933, w_001_2934, w_001_2935, w_001_2936, w_001_2937, w_001_2938, w_001_2939, w_001_2940, w_001_2941, w_001_2942, w_001_2943, w_001_2944, w_001_2945, w_001_2946, w_001_2947, w_001_2948, w_001_2949, w_001_2950, w_001_2951, w_001_2952, w_001_2953, w_001_2954, w_001_2955, w_001_2956, w_001_2957, w_001_2958, w_001_2959, w_001_2960, w_001_2962, w_001_2963, w_001_2964, w_001_2965, w_001_2966, w_001_2967, w_001_2968, w_001_2969, w_001_2970, w_001_2971, w_001_2972, w_001_2973, w_001_2974, w_001_2975, w_001_2976, w_001_2977, w_001_2978, w_001_2979, w_001_2981, w_001_2982, w_001_2983, w_001_2984, w_001_2985, w_001_2986, w_001_2987, w_001_2988, w_001_2989, w_001_2990, w_001_2991, w_001_2992, w_001_2993, w_001_2994, w_001_2995, w_001_2996, w_001_2997, w_001_2998, w_001_2999, w_001_3000, w_001_3001, w_001_3002, w_001_3003, w_001_3004, w_001_3005, w_001_3006, w_001_3007, w_001_3008, w_001_3009, w_001_3010, w_001_3011, w_001_3012, w_001_3013, w_001_3014, w_001_3015, w_001_3016, w_001_3017, w_001_3018, w_001_3019, w_001_3020, w_001_3021, w_001_3022, w_001_3023, w_001_3024, w_001_3026, w_001_3027, w_001_3028, w_001_3029, w_001_3030, w_001_3031, w_001_3032, w_001_3033, w_001_3034, w_001_3035, w_001_3036, w_001_3037, w_001_3038, w_001_3039, w_001_3040, w_001_3041, w_001_3042, w_001_3043, w_001_3044, w_001_3045, w_001_3046, w_001_3047, w_001_3048, w_001_3049, w_001_3050, w_001_3051, w_001_3052, w_001_3053, w_001_3054, w_001_3055, w_001_3056, w_001_3057, w_001_3059, w_001_3060, w_001_3061, w_001_3062, w_001_3063, w_001_3064, w_001_3065, w_001_3066, w_001_3067, w_001_3068, w_001_3069, w_001_3071, w_001_3072, w_001_3073, w_001_3074, w_001_3075, w_001_3076, w_001_3077, w_001_3079, w_001_3080, w_001_3082, w_001_3083, w_001_3084, w_001_3085, w_001_3086, w_001_3087, w_001_3088, w_001_3089, w_001_3090, w_001_3091, w_001_3092, w_001_3093, w_001_3094, w_001_3095, w_001_3096, w_001_3097, w_001_3098, w_001_3099, w_001_3100, w_001_3101, w_001_3102, w_001_3103, w_001_3104, w_001_3105, w_001_3106, w_001_3107, w_001_3108, w_001_3109, w_001_3110, w_001_3111, w_001_3112, w_001_3113, w_001_3114, w_001_3115, w_001_3116, w_001_3117, w_001_3118, w_001_3119, w_001_3120, w_001_3121, w_001_3122, w_001_3123, w_001_3124, w_001_3125, w_001_3126, w_001_3127, w_001_3128, w_001_3129, w_001_3130, w_001_3131, w_001_3132, w_001_3133, w_001_3134, w_001_3135, w_001_3136, w_001_3137, w_001_3138, w_001_3139, w_001_3140, w_001_3141, w_001_3142, w_001_3143, w_001_3144, w_001_3145, w_001_3146, w_001_3147, w_001_3148, w_001_3149, w_001_3150, w_001_3151, w_001_3152, w_001_3153, w_001_3154, w_001_3155, w_001_3156, w_001_3157, w_001_3158, w_001_3159, w_001_3160, w_001_3161, w_001_3162, w_001_3163, w_001_3164, w_001_3165, w_001_3166, w_001_3167, w_001_3168, w_001_3169, w_001_3170, w_001_3171, w_001_3172, w_001_3173, w_001_3174, w_001_3175, w_001_3176, w_001_3177, w_001_3178, w_001_3179, w_001_3180, w_001_3181, w_001_3182, w_001_3183, w_001_3184, w_001_3185, w_001_3186, w_001_3187, w_001_3188, w_001_3189, w_001_3190, w_001_3191, w_001_3192, w_001_3193, w_001_3194, w_001_3195, w_001_3196, w_001_3197, w_001_3198, w_001_3199, w_001_3200, w_001_3201, w_001_3202, w_001_3203, w_001_3204, w_001_3205, w_001_3206, w_001_3207, w_001_3208, w_001_3209, w_001_3210, w_001_3211, w_001_3212, w_001_3213, w_001_3214, w_001_3215, w_001_3216, w_001_3217, w_001_3218, w_001_3219, w_001_3220, w_001_3221, w_001_3222, w_001_3223, w_001_3224, w_001_3225, w_001_3226, w_001_3228, w_001_3229, w_001_3230, w_001_3231, w_001_3232, w_001_3233, w_001_3234, w_001_3235, w_001_3236, w_001_3237, w_001_3238, w_001_3239, w_001_3240, w_001_3241, w_001_3242, w_001_3243, w_001_3244, w_001_3245, w_001_3246, w_001_3247, w_001_3248, w_001_3249, w_001_3250, w_001_3251, w_001_3252, w_001_3253, w_001_3254, w_001_3255, w_001_3256, w_001_3257, w_001_3258, w_001_3259, w_001_3260, w_001_3261, w_001_3262, w_001_3263, w_001_3264, w_001_3265, w_001_3266, w_001_3267, w_001_3268, w_001_3269, w_001_3270, w_001_3271, w_001_3272, w_001_3273, w_001_3274, w_001_3275, w_001_3276, w_001_3277, w_001_3278, w_001_3280, w_001_3281, w_001_3282, w_001_3283, w_001_3284, w_001_3285, w_001_3286, w_001_3287, w_001_3288, w_001_3289, w_001_3290, w_001_3291, w_001_3292, w_001_3294, w_001_3295, w_001_3296, w_001_3297, w_001_3298, w_001_3299, w_001_3300, w_001_3301, w_001_3302, w_001_3303, w_001_3304, w_001_3305, w_001_3307, w_001_3308, w_001_3309, w_001_3310, w_001_3311, w_001_3312, w_001_3313, w_001_3314, w_001_3315, w_001_3316, w_001_3317, w_001_3318, w_001_3319, w_001_3320, w_001_3321, w_001_3322, w_001_3323, w_001_3324, w_001_3325, w_001_3326, w_001_3327, w_001_3328, w_001_3329, w_001_3330, w_001_3332, w_001_3333, w_001_3334, w_001_3335, w_001_3336, w_001_3337, w_001_3338, w_001_3339, w_001_3340, w_001_3341, w_001_3342, w_001_3343, w_001_3344, w_001_3345, w_001_3346, w_001_3347, w_001_3348, w_001_3349, w_001_3350, w_001_3351, w_001_3352, w_001_3353, w_001_3354, w_001_3355, w_001_3356, w_001_3357, w_001_3358, w_001_3359, w_001_3360, w_001_3361, w_001_3362, w_001_3363, w_001_3364, w_001_3365, w_001_3366, w_001_3367, w_001_3368, w_001_3370, w_001_3371, w_001_3372, w_001_3373, w_001_3374, w_001_3375, w_001_3376, w_001_3377, w_001_3378, w_001_3379, w_001_3380, w_001_3381, w_001_3382, w_001_3383, w_001_3384, w_001_3385, w_001_3386, w_001_3387, w_001_3388, w_001_3389, w_001_3390, w_001_3391, w_001_3392, w_001_3393, w_001_3394, w_001_3395, w_001_3396, w_001_3397, w_001_3398, w_001_3399, w_001_3400, w_001_3401, w_001_3402, w_001_3403, w_001_3404, w_001_3405, w_001_3406, w_001_3407, w_001_3408, w_001_3409, w_001_3410, w_001_3411, w_001_3412, w_001_3413, w_001_3414, w_001_3415, w_001_3416, w_001_3417, w_001_3418, w_001_3419, w_001_3420, w_001_3422, w_001_3423, w_001_3424, w_001_3425, w_001_3426, w_001_3427, w_001_3428, w_001_3429, w_001_3430, w_001_3431, w_001_3432, w_001_3433, w_001_3434, w_001_3435, w_001_3436, w_001_3437, w_001_3438, w_001_3439, w_001_3440, w_001_3441, w_001_3442, w_001_3443, w_001_3444, w_001_3445, w_001_3446, w_001_3447, w_001_3448, w_001_3449, w_001_3450, w_001_3451, w_001_3452, w_001_3453, w_001_3454, w_001_3455, w_001_3456, w_001_3457, w_001_3458, w_001_3459, w_001_3460, w_001_3461, w_001_3462, w_001_3463, w_001_3464, w_001_3465, w_001_3466, w_001_3467, w_001_3468, w_001_3469, w_001_3470, w_001_3471, w_001_3472, w_001_3473, w_001_3474, w_001_3475, w_001_3476, w_001_3477, w_001_3478, w_001_3479, w_001_3480, w_001_3481, w_001_3482, w_001_3483, w_001_3484, w_001_3485, w_001_3486, w_001_3487, w_001_3488, w_001_3489, w_001_3490, w_001_3491, w_001_3492, w_001_3493, w_001_3494, w_001_3495, w_001_3496, w_001_3497, w_001_3498, w_001_3499, w_001_3500, w_001_3501, w_001_3502, w_001_3503, w_001_3504, w_001_3505, w_001_3506, w_001_3507, w_001_3508, w_001_3509, w_001_3510, w_001_3511, w_001_3513, w_001_3514, w_001_3515, w_001_3516, w_001_3517, w_001_3518, w_001_3519, w_001_3520, w_001_3521, w_001_3522, w_001_3523, w_001_3524, w_001_3525, w_001_3526, w_001_3528, w_001_3529, w_001_3530, w_001_3531, w_001_3532, w_001_3533, w_001_3534, w_001_3535, w_001_3536, w_001_3537, w_001_3539, w_001_3540, w_001_3541, w_001_3542, w_001_3543, w_001_3544, w_001_3545, w_001_3546, w_001_3547, w_001_3548, w_001_3550, w_001_3551, w_001_3552, w_001_3553, w_001_3554, w_001_3555, w_001_3556, w_001_3557, w_001_3559, w_001_3560, w_001_3562, w_001_3563, w_001_3564, w_001_3565, w_001_3566, w_001_3567, w_001_3568, w_001_3569, w_001_3570, w_001_3571, w_001_3572, w_001_3573, w_001_3574, w_001_3575, w_001_3576, w_001_3577, w_001_3578, w_001_3579, w_001_3580, w_001_3581, w_001_3582, w_001_3583, w_001_3584, w_001_3585, w_001_3586, w_001_3587, w_001_3588, w_001_3589, w_001_3590, w_001_3591, w_001_3592, w_001_3594, w_001_3595, w_001_3596, w_001_3597;
  wire w_002_000, w_002_001, w_002_002, w_002_003, w_002_004, w_002_005, w_002_006, w_002_007, w_002_008, w_002_009, w_002_010, w_002_011, w_002_012, w_002_013, w_002_014, w_002_015, w_002_016, w_002_017, w_002_018, w_002_019, w_002_020, w_002_021, w_002_022, w_002_023, w_002_024, w_002_025, w_002_026, w_002_027, w_002_028, w_002_029, w_002_030, w_002_031, w_002_032, w_002_033, w_002_034, w_002_035, w_002_036, w_002_037, w_002_038, w_002_039, w_002_040, w_002_041, w_002_042, w_002_043, w_002_044, w_002_045, w_002_046, w_002_047, w_002_048, w_002_049, w_002_050, w_002_051, w_002_052, w_002_053, w_002_054, w_002_055, w_002_056, w_002_057, w_002_058, w_002_059, w_002_060, w_002_061, w_002_062, w_002_063, w_002_064, w_002_065, w_002_066, w_002_067, w_002_068, w_002_069, w_002_070, w_002_071, w_002_072, w_002_073, w_002_074, w_002_075, w_002_076, w_002_077, w_002_078, w_002_079, w_002_080, w_002_081, w_002_082, w_002_083, w_002_084, w_002_085, w_002_086, w_002_087, w_002_088, w_002_089, w_002_090, w_002_091, w_002_092, w_002_093, w_002_094, w_002_095, w_002_096, w_002_097, w_002_098, w_002_099, w_002_100, w_002_101, w_002_102, w_002_103, w_002_104, w_002_105, w_002_106, w_002_107, w_002_108, w_002_109, w_002_110, w_002_111, w_002_112, w_002_113, w_002_114, w_002_115, w_002_116, w_002_117, w_002_118, w_002_119, w_002_120, w_002_121, w_002_122, w_002_123, w_002_124, w_002_125, w_002_126, w_002_127, w_002_128, w_002_129, w_002_130, w_002_131, w_002_132, w_002_133, w_002_134, w_002_135, w_002_136, w_002_137, w_002_138, w_002_139, w_002_140, w_002_141, w_002_142, w_002_143, w_002_144, w_002_145, w_002_146, w_002_147, w_002_148, w_002_149, w_002_150, w_002_151, w_002_152, w_002_153, w_002_154, w_002_155, w_002_156, w_002_157, w_002_158, w_002_159, w_002_160, w_002_161, w_002_162, w_002_163, w_002_164, w_002_165, w_002_166, w_002_167, w_002_168, w_002_169, w_002_170, w_002_171, w_002_172, w_002_173, w_002_174, w_002_175, w_002_176, w_002_177, w_002_178, w_002_179, w_002_180, w_002_181, w_002_182, w_002_183, w_002_184, w_002_185, w_002_186, w_002_187, w_002_188, w_002_189, w_002_190, w_002_191, w_002_192, w_002_193, w_002_194, w_002_195, w_002_196, w_002_197, w_002_198, w_002_199, w_002_200, w_002_201, w_002_202, w_002_203, w_002_204, w_002_205, w_002_206, w_002_207, w_002_208, w_002_209, w_002_210, w_002_211, w_002_212, w_002_213, w_002_214, w_002_215, w_002_216, w_002_217, w_002_218, w_002_219, w_002_220, w_002_221, w_002_222, w_002_223, w_002_224, w_002_225, w_002_226, w_002_227, w_002_228, w_002_229, w_002_230, w_002_231, w_002_232, w_002_233, w_002_234, w_002_235, w_002_236, w_002_237, w_002_238, w_002_239, w_002_240, w_002_241, w_002_242, w_002_243, w_002_244, w_002_245, w_002_246, w_002_247, w_002_248, w_002_249, w_002_250, w_002_251, w_002_252, w_002_253, w_002_254, w_002_255, w_002_256, w_002_257, w_002_258, w_002_259, w_002_260, w_002_261, w_002_262, w_002_263, w_002_264, w_002_265, w_002_266, w_002_267, w_002_268, w_002_269, w_002_270, w_002_271, w_002_272, w_002_273, w_002_274, w_002_275, w_002_276, w_002_277, w_002_278, w_002_279, w_002_280, w_002_281, w_002_282, w_002_283, w_002_284, w_002_285, w_002_286, w_002_287, w_002_288, w_002_289, w_002_290, w_002_291, w_002_292, w_002_293, w_002_294, w_002_295, w_002_296, w_002_297, w_002_298, w_002_299, w_002_300, w_002_301, w_002_302, w_002_303, w_002_304, w_002_305, w_002_306, w_002_307, w_002_308, w_002_309, w_002_310, w_002_311, w_002_312, w_002_313, w_002_314, w_002_315, w_002_316, w_002_317, w_002_318, w_002_319, w_002_320, w_002_321, w_002_322, w_002_323, w_002_324, w_002_325, w_002_326, w_002_327, w_002_328, w_002_329, w_002_330, w_002_331, w_002_332, w_002_333, w_002_334, w_002_335, w_002_336, w_002_337, w_002_338, w_002_339, w_002_340, w_002_341, w_002_342, w_002_343, w_002_344, w_002_345, w_002_346, w_002_347, w_002_348, w_002_349, w_002_350, w_002_351, w_002_352, w_002_353, w_002_354, w_002_355, w_002_356, w_002_357, w_002_358, w_002_359, w_002_360, w_002_361, w_002_362, w_002_363, w_002_364, w_002_365, w_002_366, w_002_367, w_002_368, w_002_369, w_002_370, w_002_371, w_002_372, w_002_373, w_002_374, w_002_375, w_002_376, w_002_377, w_002_378, w_002_379, w_002_380, w_002_381, w_002_382, w_002_383, w_002_384, w_002_385, w_002_386, w_002_387, w_002_388, w_002_389, w_002_390, w_002_391, w_002_392, w_002_393, w_002_394, w_002_395, w_002_396, w_002_397, w_002_398, w_002_399, w_002_400, w_002_401, w_002_402, w_002_403, w_002_404, w_002_405, w_002_406, w_002_407, w_002_408, w_002_409, w_002_410, w_002_411, w_002_412, w_002_413, w_002_414, w_002_415, w_002_416, w_002_417, w_002_418, w_002_419, w_002_420, w_002_421, w_002_422, w_002_423, w_002_424, w_002_425, w_002_426, w_002_427, w_002_428, w_002_429, w_002_430, w_002_431, w_002_432, w_002_433, w_002_434, w_002_435, w_002_436, w_002_437, w_002_438, w_002_439, w_002_440, w_002_441, w_002_442, w_002_443, w_002_444, w_002_445, w_002_446, w_002_447, w_002_448, w_002_449, w_002_450, w_002_451, w_002_452, w_002_453, w_002_454, w_002_455, w_002_456, w_002_457, w_002_458, w_002_459, w_002_460, w_002_461, w_002_462, w_002_463, w_002_464, w_002_465, w_002_466, w_002_467, w_002_468, w_002_469, w_002_470, w_002_471, w_002_472, w_002_473, w_002_474, w_002_475, w_002_476, w_002_477, w_002_478, w_002_479, w_002_480, w_002_481, w_002_482, w_002_483, w_002_484, w_002_485, w_002_486, w_002_487, w_002_488, w_002_489, w_002_490, w_002_491, w_002_492, w_002_493, w_002_494, w_002_495, w_002_496, w_002_497, w_002_498, w_002_499, w_002_500, w_002_501, w_002_502, w_002_503, w_002_504, w_002_505, w_002_506, w_002_507, w_002_508, w_002_509, w_002_510, w_002_511, w_002_512, w_002_513, w_002_514, w_002_515, w_002_516, w_002_517, w_002_518, w_002_519, w_002_520, w_002_521, w_002_522, w_002_523, w_002_524, w_002_525, w_002_526, w_002_527, w_002_528, w_002_529, w_002_530, w_002_531, w_002_532, w_002_533, w_002_534, w_002_535, w_002_536, w_002_537, w_002_538, w_002_539, w_002_540, w_002_541, w_002_542, w_002_543, w_002_544, w_002_545, w_002_546, w_002_547, w_002_548, w_002_549, w_002_550, w_002_551, w_002_552, w_002_553, w_002_554, w_002_555, w_002_556, w_002_557, w_002_558, w_002_559, w_002_560, w_002_561, w_002_562, w_002_563, w_002_564, w_002_565, w_002_566, w_002_567, w_002_568, w_002_569, w_002_570, w_002_571, w_002_572, w_002_573, w_002_574, w_002_575, w_002_576, w_002_577, w_002_578, w_002_579, w_002_580, w_002_581, w_002_582, w_002_583, w_002_584, w_002_585, w_002_586, w_002_587, w_002_588, w_002_589, w_002_590, w_002_591, w_002_592, w_002_593, w_002_594, w_002_595, w_002_596, w_002_597, w_002_598, w_002_599, w_002_600, w_002_601, w_002_602, w_002_603, w_002_604, w_002_605, w_002_606, w_002_607, w_002_608, w_002_609, w_002_610, w_002_611, w_002_612, w_002_613, w_002_614, w_002_615, w_002_616, w_002_617, w_002_618, w_002_619, w_002_620, w_002_621, w_002_622, w_002_623, w_002_624, w_002_625, w_002_626, w_002_627, w_002_628, w_002_629, w_002_630, w_002_631, w_002_632, w_002_633, w_002_634, w_002_635, w_002_636, w_002_637, w_002_638, w_002_639, w_002_640, w_002_641, w_002_642, w_002_643, w_002_644, w_002_645, w_002_646, w_002_647, w_002_648, w_002_649, w_002_650, w_002_651, w_002_652, w_002_653, w_002_654, w_002_655, w_002_656, w_002_657, w_002_658, w_002_659, w_002_660, w_002_661, w_002_662, w_002_663, w_002_664, w_002_665, w_002_666, w_002_667, w_002_668, w_002_669, w_002_670, w_002_671, w_002_672, w_002_673, w_002_674, w_002_675, w_002_676, w_002_677, w_002_678, w_002_679, w_002_680, w_002_681, w_002_682, w_002_683, w_002_684, w_002_685, w_002_686, w_002_687, w_002_688, w_002_689, w_002_690, w_002_691, w_002_692, w_002_693, w_002_694, w_002_695, w_002_696, w_002_697, w_002_698, w_002_699, w_002_700, w_002_701, w_002_702, w_002_703, w_002_704, w_002_705, w_002_706, w_002_707, w_002_708, w_002_709, w_002_710, w_002_711, w_002_712, w_002_713, w_002_714, w_002_715, w_002_716, w_002_717, w_002_718, w_002_719, w_002_720, w_002_721, w_002_722, w_002_723, w_002_724, w_002_725, w_002_726, w_002_727, w_002_728, w_002_729, w_002_730, w_002_731, w_002_732, w_002_733, w_002_734, w_002_735, w_002_736, w_002_737, w_002_738, w_002_739, w_002_740, w_002_741, w_002_742, w_002_743, w_002_744, w_002_745, w_002_746, w_002_747, w_002_748, w_002_749, w_002_750, w_002_751, w_002_752, w_002_753, w_002_754, w_002_755, w_002_756, w_002_757, w_002_758, w_002_759, w_002_760, w_002_761, w_002_762, w_002_763, w_002_764, w_002_765, w_002_766, w_002_767, w_002_768, w_002_769, w_002_770, w_002_771, w_002_772, w_002_773, w_002_774, w_002_775, w_002_776, w_002_777, w_002_778, w_002_779, w_002_780, w_002_781, w_002_782, w_002_783, w_002_784, w_002_785, w_002_786, w_002_787, w_002_788, w_002_789, w_002_790, w_002_791, w_002_792, w_002_793, w_002_794, w_002_795, w_002_796, w_002_797, w_002_798, w_002_799, w_002_800, w_002_801, w_002_802, w_002_803, w_002_804, w_002_805, w_002_806, w_002_807, w_002_808, w_002_809, w_002_810, w_002_811, w_002_812, w_002_813, w_002_814, w_002_815, w_002_816, w_002_817, w_002_818, w_002_819, w_002_820, w_002_821, w_002_822, w_002_823, w_002_824, w_002_825, w_002_826, w_002_827, w_002_828, w_002_829, w_002_830, w_002_831, w_002_832, w_002_833, w_002_834, w_002_835, w_002_836, w_002_837, w_002_838, w_002_839, w_002_840, w_002_841, w_002_842, w_002_843, w_002_844, w_002_845, w_002_846, w_002_847, w_002_848, w_002_849, w_002_850, w_002_851, w_002_852, w_002_853, w_002_854, w_002_855, w_002_856, w_002_857, w_002_858, w_002_859, w_002_860, w_002_861, w_002_862, w_002_863, w_002_864, w_002_865, w_002_866, w_002_867, w_002_868, w_002_869, w_002_870, w_002_871, w_002_872;
  wire w_003_000, w_003_001, w_003_002, w_003_003, w_003_004, w_003_005, w_003_006, w_003_007, w_003_008, w_003_009, w_003_010, w_003_011, w_003_012, w_003_013, w_003_014, w_003_015, w_003_016, w_003_017, w_003_018, w_003_019, w_003_020, w_003_021, w_003_022, w_003_023, w_003_024, w_003_025, w_003_026, w_003_027, w_003_028, w_003_029, w_003_030, w_003_031, w_003_032, w_003_033, w_003_034, w_003_035, w_003_036, w_003_037, w_003_038, w_003_039, w_003_040, w_003_041, w_003_042, w_003_043, w_003_044, w_003_045, w_003_046, w_003_047, w_003_048, w_003_049, w_003_050, w_003_051, w_003_052, w_003_053, w_003_054, w_003_055, w_003_056, w_003_057, w_003_058, w_003_059, w_003_060, w_003_061, w_003_062, w_003_063, w_003_064, w_003_065, w_003_066, w_003_067, w_003_068, w_003_069, w_003_070, w_003_071, w_003_072, w_003_073, w_003_074, w_003_075, w_003_076, w_003_077, w_003_078, w_003_079, w_003_080, w_003_081, w_003_082, w_003_083, w_003_084, w_003_085, w_003_086, w_003_087, w_003_088, w_003_089, w_003_090, w_003_091, w_003_092, w_003_093, w_003_094, w_003_095, w_003_096, w_003_097, w_003_098, w_003_099, w_003_100, w_003_101, w_003_102, w_003_103, w_003_104, w_003_105, w_003_106, w_003_107, w_003_108, w_003_109, w_003_110, w_003_111, w_003_112, w_003_113, w_003_114, w_003_115, w_003_116, w_003_117, w_003_118, w_003_119, w_003_120, w_003_121, w_003_122, w_003_123, w_003_124, w_003_125, w_003_126, w_003_127, w_003_128, w_003_129, w_003_130, w_003_131, w_003_132, w_003_133, w_003_134, w_003_135, w_003_136, w_003_137, w_003_138, w_003_139, w_003_140, w_003_141, w_003_142, w_003_143, w_003_144, w_003_145, w_003_146, w_003_147, w_003_148, w_003_149, w_003_150, w_003_151, w_003_152, w_003_153, w_003_154, w_003_155, w_003_156, w_003_157, w_003_158, w_003_159, w_003_160, w_003_161, w_003_162, w_003_163, w_003_164, w_003_165, w_003_166, w_003_167, w_003_168, w_003_169, w_003_170, w_003_171, w_003_172, w_003_173, w_003_174, w_003_175, w_003_176, w_003_177, w_003_178, w_003_179, w_003_180, w_003_181, w_003_182, w_003_183, w_003_184, w_003_185, w_003_186, w_003_187, w_003_188, w_003_189, w_003_190, w_003_191, w_003_192, w_003_193, w_003_194, w_003_195, w_003_196, w_003_197, w_003_198, w_003_199, w_003_200, w_003_201, w_003_202, w_003_203, w_003_204, w_003_205, w_003_206, w_003_207, w_003_208, w_003_209, w_003_210, w_003_211, w_003_212, w_003_213, w_003_214, w_003_215, w_003_216, w_003_217, w_003_218, w_003_219, w_003_220, w_003_221, w_003_222, w_003_223, w_003_224, w_003_225, w_003_226, w_003_227, w_003_228, w_003_229, w_003_230, w_003_231, w_003_232, w_003_233, w_003_234, w_003_235, w_003_236, w_003_237, w_003_238, w_003_239, w_003_240, w_003_241, w_003_242, w_003_243, w_003_244, w_003_245, w_003_246, w_003_247, w_003_248, w_003_249, w_003_250, w_003_251, w_003_252, w_003_253, w_003_254, w_003_255, w_003_256, w_003_257, w_003_258, w_003_259, w_003_260, w_003_261, w_003_262, w_003_263, w_003_264, w_003_265, w_003_266, w_003_267, w_003_268, w_003_269, w_003_270, w_003_271, w_003_272, w_003_273, w_003_274, w_003_275, w_003_276, w_003_277, w_003_278, w_003_279, w_003_280, w_003_281, w_003_282, w_003_283, w_003_284, w_003_285, w_003_286, w_003_287, w_003_288, w_003_289, w_003_290, w_003_291, w_003_292, w_003_293, w_003_294, w_003_295, w_003_296, w_003_297, w_003_298, w_003_299, w_003_300, w_003_301, w_003_302, w_003_303, w_003_304, w_003_305, w_003_306, w_003_307, w_003_308, w_003_309, w_003_310, w_003_311, w_003_312, w_003_313, w_003_314, w_003_315, w_003_316, w_003_317, w_003_318, w_003_319, w_003_320, w_003_321, w_003_322, w_003_323, w_003_324, w_003_325, w_003_326, w_003_327, w_003_328, w_003_329, w_003_330, w_003_331, w_003_332, w_003_333, w_003_334, w_003_335, w_003_336, w_003_337, w_003_338, w_003_339, w_003_340, w_003_341, w_003_342, w_003_343, w_003_344, w_003_345, w_003_346, w_003_347, w_003_348, w_003_349, w_003_350, w_003_351, w_003_352, w_003_353, w_003_354, w_003_355, w_003_356, w_003_357, w_003_358, w_003_359, w_003_360, w_003_361, w_003_362, w_003_363, w_003_364, w_003_365, w_003_366, w_003_367, w_003_368, w_003_369, w_003_370, w_003_371, w_003_372, w_003_373, w_003_374, w_003_375, w_003_376, w_003_377, w_003_378, w_003_379, w_003_380, w_003_381, w_003_382, w_003_383, w_003_384, w_003_385, w_003_386, w_003_387, w_003_388, w_003_389, w_003_390, w_003_391, w_003_392, w_003_393, w_003_394, w_003_395, w_003_396, w_003_397, w_003_398, w_003_399, w_003_400, w_003_401, w_003_402, w_003_403, w_003_404, w_003_405, w_003_406, w_003_407, w_003_408, w_003_409, w_003_410, w_003_411, w_003_412, w_003_413, w_003_414, w_003_415, w_003_416, w_003_417, w_003_418, w_003_419, w_003_420, w_003_421, w_003_422, w_003_423, w_003_424, w_003_425, w_003_426, w_003_427, w_003_428, w_003_429, w_003_430, w_003_431, w_003_432, w_003_433, w_003_434, w_003_435, w_003_436, w_003_437, w_003_438, w_003_439, w_003_440, w_003_441, w_003_442, w_003_443, w_003_444, w_003_445, w_003_446, w_003_447, w_003_448, w_003_449, w_003_450, w_003_451, w_003_452, w_003_453, w_003_454, w_003_455, w_003_456, w_003_457, w_003_458, w_003_459, w_003_460, w_003_461, w_003_462, w_003_463, w_003_464, w_003_465, w_003_466, w_003_467, w_003_468, w_003_469, w_003_470, w_003_471, w_003_472, w_003_473, w_003_474, w_003_475, w_003_476, w_003_477, w_003_478, w_003_479, w_003_480, w_003_481, w_003_482, w_003_483, w_003_484, w_003_485, w_003_486, w_003_487, w_003_488, w_003_489, w_003_490, w_003_491, w_003_492, w_003_493, w_003_494, w_003_495, w_003_496, w_003_497, w_003_498, w_003_499, w_003_500, w_003_501, w_003_502, w_003_503, w_003_504, w_003_505, w_003_506, w_003_507, w_003_508, w_003_509, w_003_510, w_003_511, w_003_512, w_003_513, w_003_514, w_003_515, w_003_516, w_003_517, w_003_518, w_003_519, w_003_520, w_003_521, w_003_522, w_003_523, w_003_524, w_003_525, w_003_526, w_003_527, w_003_528, w_003_529, w_003_530, w_003_531, w_003_532, w_003_533, w_003_534, w_003_535, w_003_536, w_003_537, w_003_538, w_003_539, w_003_540, w_003_541, w_003_542, w_003_543, w_003_544, w_003_545, w_003_546, w_003_547, w_003_548, w_003_549, w_003_550, w_003_551, w_003_552, w_003_553, w_003_554, w_003_555, w_003_556, w_003_557, w_003_558, w_003_559, w_003_560, w_003_561, w_003_562, w_003_563, w_003_564, w_003_566, w_003_567, w_003_568, w_003_569, w_003_570, w_003_571, w_003_572, w_003_573, w_003_574, w_003_575, w_003_576, w_003_577, w_003_578, w_003_579, w_003_580, w_003_581, w_003_582, w_003_583, w_003_584, w_003_585, w_003_586, w_003_587, w_003_588, w_003_589, w_003_590, w_003_591, w_003_592, w_003_593, w_003_594, w_003_595, w_003_596, w_003_597, w_003_598, w_003_599, w_003_600, w_003_601, w_003_602, w_003_603, w_003_604, w_003_605, w_003_606, w_003_607, w_003_608, w_003_609, w_003_610, w_003_611, w_003_612, w_003_613, w_003_614, w_003_615, w_003_616, w_003_617, w_003_618, w_003_619, w_003_620, w_003_621, w_003_622, w_003_623, w_003_624, w_003_625, w_003_626, w_003_627, w_003_628, w_003_629, w_003_630, w_003_631, w_003_632, w_003_633, w_003_634, w_003_635, w_003_636, w_003_637, w_003_638, w_003_639, w_003_640, w_003_641, w_003_642, w_003_643, w_003_644, w_003_645, w_003_646, w_003_647, w_003_648, w_003_649, w_003_650, w_003_651, w_003_652, w_003_653, w_003_654, w_003_655, w_003_656, w_003_657, w_003_658, w_003_659, w_003_660, w_003_661, w_003_662, w_003_663, w_003_664, w_003_665, w_003_666, w_003_667, w_003_668, w_003_669, w_003_670, w_003_671, w_003_672, w_003_673, w_003_674, w_003_675, w_003_676, w_003_677, w_003_678, w_003_679, w_003_680, w_003_681, w_003_682, w_003_683, w_003_684, w_003_685, w_003_686, w_003_687, w_003_688, w_003_689, w_003_690, w_003_691, w_003_692, w_003_693, w_003_694, w_003_695, w_003_696, w_003_697, w_003_698, w_003_699, w_003_700, w_003_701, w_003_702, w_003_703, w_003_704, w_003_705, w_003_706, w_003_707, w_003_708, w_003_709, w_003_710, w_003_711, w_003_712, w_003_713, w_003_714, w_003_715, w_003_716, w_003_717, w_003_718, w_003_719, w_003_720, w_003_721, w_003_722, w_003_723, w_003_724, w_003_725, w_003_726, w_003_727, w_003_728, w_003_729, w_003_730, w_003_731, w_003_732, w_003_733, w_003_734, w_003_735, w_003_736, w_003_737, w_003_738, w_003_739, w_003_740, w_003_741, w_003_742, w_003_743, w_003_744, w_003_745, w_003_746, w_003_747, w_003_748, w_003_749, w_003_750, w_003_751, w_003_752, w_003_753, w_003_754, w_003_755, w_003_756, w_003_757, w_003_758, w_003_759, w_003_760, w_003_761, w_003_762, w_003_763, w_003_764, w_003_765, w_003_766, w_003_767, w_003_768, w_003_769, w_003_770, w_003_771, w_003_772, w_003_773, w_003_774, w_003_775, w_003_776, w_003_777, w_003_778, w_003_779, w_003_780, w_003_781, w_003_782, w_003_783, w_003_784, w_003_785, w_003_786, w_003_787, w_003_788, w_003_789, w_003_790, w_003_791, w_003_792, w_003_793, w_003_794, w_003_795, w_003_796, w_003_797, w_003_798, w_003_799, w_003_800, w_003_801, w_003_802, w_003_803, w_003_804, w_003_805, w_003_806, w_003_807, w_003_808, w_003_809, w_003_810, w_003_811, w_003_812, w_003_813, w_003_814, w_003_815, w_003_816, w_003_817, w_003_818, w_003_819, w_003_820, w_003_821, w_003_822, w_003_823, w_003_824, w_003_825, w_003_826, w_003_827, w_003_828, w_003_829, w_003_830, w_003_831, w_003_832, w_003_833, w_003_834, w_003_835, w_003_836, w_003_837, w_003_838, w_003_839, w_003_840, w_003_841, w_003_842, w_003_843, w_003_844, w_003_845, w_003_846, w_003_847, w_003_848, w_003_849, w_003_850, w_003_851, w_003_852, w_003_853, w_003_854, w_003_855, w_003_856, w_003_857, w_003_858, w_003_859, w_003_860, w_003_861, w_003_862, w_003_863, w_003_864, w_003_865, w_003_866, w_003_867, w_003_868, w_003_869, w_003_870, w_003_871, w_003_872, w_003_873, w_003_874, w_003_875, w_003_876, w_003_877, w_003_878, w_003_879, w_003_880, w_003_881, w_003_882, w_003_883, w_003_884, w_003_885, w_003_886, w_003_887, w_003_888, w_003_889, w_003_890, w_003_891, w_003_892, w_003_893, w_003_894, w_003_895, w_003_896, w_003_897, w_003_898, w_003_899, w_003_900, w_003_901, w_003_902, w_003_903, w_003_904, w_003_905, w_003_906, w_003_907, w_003_908, w_003_909, w_003_910, w_003_911, w_003_912, w_003_913, w_003_914, w_003_915, w_003_916, w_003_917, w_003_918, w_003_919, w_003_920, w_003_921, w_003_922, w_003_923, w_003_924, w_003_925, w_003_926, w_003_927, w_003_928, w_003_929, w_003_930, w_003_931, w_003_932, w_003_933, w_003_934, w_003_935, w_003_936, w_003_937, w_003_938, w_003_939, w_003_940, w_003_941, w_003_942, w_003_943, w_003_944, w_003_945, w_003_946, w_003_947, w_003_948, w_003_949, w_003_950, w_003_951, w_003_952, w_003_953, w_003_954, w_003_955, w_003_956, w_003_957, w_003_958, w_003_959, w_003_960, w_003_961, w_003_963, w_003_964, w_003_965, w_003_966, w_003_967, w_003_968, w_003_969, w_003_970, w_003_971, w_003_972, w_003_973, w_003_974, w_003_975, w_003_976, w_003_977, w_003_978, w_003_979, w_003_980, w_003_981, w_003_982, w_003_983, w_003_984, w_003_985, w_003_986, w_003_987, w_003_988, w_003_989, w_003_990, w_003_991, w_003_992, w_003_993, w_003_994, w_003_995, w_003_996, w_003_997, w_003_998, w_003_999, w_003_1000, w_003_1001, w_003_1002, w_003_1003, w_003_1004, w_003_1005, w_003_1006, w_003_1007, w_003_1008, w_003_1009, w_003_1010, w_003_1011, w_003_1012, w_003_1013, w_003_1014, w_003_1015, w_003_1016, w_003_1017, w_003_1018, w_003_1019, w_003_1020, w_003_1021, w_003_1022, w_003_1023, w_003_1024, w_003_1025, w_003_1026, w_003_1027, w_003_1028, w_003_1029, w_003_1030, w_003_1031, w_003_1032, w_003_1033, w_003_1034, w_003_1035, w_003_1036, w_003_1037, w_003_1038, w_003_1039, w_003_1040, w_003_1041, w_003_1042, w_003_1043, w_003_1044, w_003_1045, w_003_1046, w_003_1047, w_003_1048, w_003_1049, w_003_1050, w_003_1051, w_003_1052, w_003_1053, w_003_1054, w_003_1055, w_003_1056, w_003_1057, w_003_1058, w_003_1059, w_003_1060, w_003_1061, w_003_1062, w_003_1063, w_003_1064, w_003_1065, w_003_1066, w_003_1067, w_003_1068, w_003_1069, w_003_1070, w_003_1071, w_003_1072, w_003_1073, w_003_1074, w_003_1075, w_003_1076, w_003_1077, w_003_1078, w_003_1079, w_003_1080, w_003_1081, w_003_1082, w_003_1083, w_003_1085, w_003_1086, w_003_1087, w_003_1088, w_003_1089, w_003_1090, w_003_1091, w_003_1092, w_003_1093, w_003_1095, w_003_1096, w_003_1097, w_003_1098, w_003_1099, w_003_1100, w_003_1101, w_003_1102, w_003_1103, w_003_1104, w_003_1105, w_003_1106, w_003_1107, w_003_1108, w_003_1109, w_003_1110, w_003_1111, w_003_1112, w_003_1113, w_003_1114, w_003_1115, w_003_1116, w_003_1117, w_003_1118, w_003_1119, w_003_1120, w_003_1121, w_003_1122, w_003_1123, w_003_1124, w_003_1125, w_003_1126, w_003_1127, w_003_1128, w_003_1129, w_003_1130, w_003_1131, w_003_1132, w_003_1133, w_003_1134, w_003_1135, w_003_1136, w_003_1137, w_003_1138, w_003_1139, w_003_1140, w_003_1141, w_003_1142, w_003_1143, w_003_1144, w_003_1145, w_003_1146, w_003_1147, w_003_1148, w_003_1149, w_003_1150, w_003_1151, w_003_1152, w_003_1153, w_003_1154, w_003_1155, w_003_1156, w_003_1157, w_003_1158, w_003_1159, w_003_1160, w_003_1161, w_003_1162, w_003_1163, w_003_1164, w_003_1165, w_003_1166, w_003_1167, w_003_1168, w_003_1169, w_003_1170, w_003_1171, w_003_1172, w_003_1173, w_003_1174, w_003_1175, w_003_1176, w_003_1177, w_003_1178, w_003_1179, w_003_1180, w_003_1181, w_003_1182, w_003_1183, w_003_1184, w_003_1185, w_003_1186, w_003_1187, w_003_1188, w_003_1189, w_003_1190, w_003_1191, w_003_1192, w_003_1193, w_003_1194, w_003_1195, w_003_1196, w_003_1197, w_003_1198, w_003_1199, w_003_1200, w_003_1201, w_003_1202, w_003_1203, w_003_1204, w_003_1205, w_003_1206, w_003_1207, w_003_1208, w_003_1209, w_003_1210, w_003_1211, w_003_1212, w_003_1213, w_003_1214, w_003_1215, w_003_1216, w_003_1217, w_003_1218, w_003_1219, w_003_1220, w_003_1221, w_003_1222, w_003_1223, w_003_1224, w_003_1225, w_003_1226, w_003_1227, w_003_1228, w_003_1229, w_003_1230, w_003_1231, w_003_1232, w_003_1233, w_003_1234, w_003_1235, w_003_1236, w_003_1237, w_003_1238, w_003_1239, w_003_1240, w_003_1241, w_003_1243, w_003_1244, w_003_1245, w_003_1246, w_003_1247, w_003_1248, w_003_1249, w_003_1250, w_003_1251, w_003_1252, w_003_1253, w_003_1254, w_003_1255, w_003_1256, w_003_1257, w_003_1258, w_003_1259, w_003_1260, w_003_1261, w_003_1262, w_003_1263, w_003_1264, w_003_1265, w_003_1266, w_003_1267, w_003_1268, w_003_1269, w_003_1270, w_003_1271, w_003_1272, w_003_1273, w_003_1274, w_003_1275, w_003_1276, w_003_1277, w_003_1278, w_003_1279, w_003_1280, w_003_1281, w_003_1282, w_003_1283, w_003_1284, w_003_1285, w_003_1286, w_003_1287, w_003_1288, w_003_1289, w_003_1290, w_003_1291, w_003_1292, w_003_1293, w_003_1294, w_003_1295, w_003_1296, w_003_1297, w_003_1298, w_003_1299, w_003_1300, w_003_1301, w_003_1302, w_003_1303, w_003_1304, w_003_1305, w_003_1306, w_003_1307, w_003_1308, w_003_1309, w_003_1310, w_003_1311, w_003_1312, w_003_1313, w_003_1314, w_003_1315, w_003_1316, w_003_1317, w_003_1318, w_003_1319, w_003_1320, w_003_1321, w_003_1322, w_003_1323, w_003_1324, w_003_1325, w_003_1326, w_003_1328, w_003_1329, w_003_1330, w_003_1331, w_003_1332, w_003_1333, w_003_1334, w_003_1335, w_003_1336, w_003_1337, w_003_1338, w_003_1339, w_003_1340, w_003_1341, w_003_1342, w_003_1343, w_003_1344, w_003_1345, w_003_1346, w_003_1347, w_003_1348, w_003_1349, w_003_1350, w_003_1351, w_003_1352, w_003_1353, w_003_1354, w_003_1355, w_003_1356, w_003_1357, w_003_1358, w_003_1359, w_003_1360, w_003_1361, w_003_1362, w_003_1363, w_003_1364, w_003_1365, w_003_1366, w_003_1367, w_003_1368, w_003_1369, w_003_1370, w_003_1371, w_003_1372, w_003_1373, w_003_1374, w_003_1375, w_003_1376, w_003_1377, w_003_1378, w_003_1379, w_003_1380, w_003_1381, w_003_1382, w_003_1383, w_003_1384, w_003_1385, w_003_1386, w_003_1387, w_003_1388, w_003_1389, w_003_1390, w_003_1391, w_003_1392, w_003_1393, w_003_1394, w_003_1395, w_003_1396, w_003_1397, w_003_1398, w_003_1399, w_003_1400, w_003_1401, w_003_1402, w_003_1403, w_003_1404, w_003_1405, w_003_1406, w_003_1407, w_003_1408, w_003_1409, w_003_1410, w_003_1411, w_003_1412, w_003_1413, w_003_1414, w_003_1415, w_003_1416, w_003_1417, w_003_1418, w_003_1419, w_003_1420, w_003_1421, w_003_1422, w_003_1423, w_003_1424, w_003_1425, w_003_1426, w_003_1427, w_003_1428, w_003_1429, w_003_1430, w_003_1431, w_003_1432, w_003_1433, w_003_1434, w_003_1435, w_003_1436, w_003_1437, w_003_1438, w_003_1439, w_003_1440, w_003_1441, w_003_1442, w_003_1443, w_003_1444, w_003_1445, w_003_1446, w_003_1447, w_003_1448, w_003_1449, w_003_1450, w_003_1451, w_003_1452, w_003_1453, w_003_1454, w_003_1455, w_003_1456, w_003_1457, w_003_1458, w_003_1459, w_003_1460, w_003_1461, w_003_1462, w_003_1463, w_003_1464, w_003_1465, w_003_1466, w_003_1467, w_003_1468, w_003_1469, w_003_1470, w_003_1471, w_003_1472, w_003_1473, w_003_1474, w_003_1475, w_003_1476, w_003_1477, w_003_1478, w_003_1479, w_003_1480, w_003_1481, w_003_1482, w_003_1483, w_003_1484, w_003_1485, w_003_1486, w_003_1487, w_003_1488, w_003_1489, w_003_1490, w_003_1491, w_003_1492, w_003_1493, w_003_1494, w_003_1495, w_003_1496, w_003_1497, w_003_1498, w_003_1499, w_003_1500, w_003_1501, w_003_1502, w_003_1503, w_003_1504, w_003_1505, w_003_1506, w_003_1507, w_003_1508, w_003_1509, w_003_1510, w_003_1511, w_003_1512, w_003_1513, w_003_1514, w_003_1515, w_003_1516, w_003_1517, w_003_1518, w_003_1519, w_003_1520, w_003_1521, w_003_1522, w_003_1523, w_003_1524, w_003_1525, w_003_1526, w_003_1527, w_003_1528, w_003_1529, w_003_1530, w_003_1531, w_003_1532, w_003_1533, w_003_1534, w_003_1535, w_003_1536, w_003_1537, w_003_1538, w_003_1539, w_003_1540, w_003_1541, w_003_1542, w_003_1543, w_003_1544, w_003_1545, w_003_1546, w_003_1547, w_003_1548, w_003_1549, w_003_1550, w_003_1551, w_003_1552, w_003_1553, w_003_1554, w_003_1555, w_003_1556, w_003_1557, w_003_1558, w_003_1559, w_003_1560, w_003_1561, w_003_1562, w_003_1563, w_003_1564, w_003_1565, w_003_1566, w_003_1567, w_003_1568, w_003_1569, w_003_1570, w_003_1571, w_003_1572, w_003_1573, w_003_1574, w_003_1575, w_003_1576, w_003_1577, w_003_1578, w_003_1579, w_003_1580, w_003_1581, w_003_1582, w_003_1583, w_003_1584, w_003_1585, w_003_1586, w_003_1587, w_003_1588, w_003_1589, w_003_1590, w_003_1591, w_003_1592, w_003_1593, w_003_1594, w_003_1595, w_003_1596, w_003_1597, w_003_1598, w_003_1599, w_003_1600, w_003_1601, w_003_1602, w_003_1603, w_003_1604, w_003_1605, w_003_1606, w_003_1607, w_003_1608, w_003_1609, w_003_1610, w_003_1611, w_003_1612, w_003_1613, w_003_1614, w_003_1615, w_003_1616, w_003_1617, w_003_1618, w_003_1619, w_003_1620, w_003_1621, w_003_1622, w_003_1623, w_003_1624, w_003_1625, w_003_1626, w_003_1627, w_003_1628, w_003_1629, w_003_1630, w_003_1631, w_003_1632, w_003_1633, w_003_1634, w_003_1635, w_003_1636, w_003_1637, w_003_1638, w_003_1639, w_003_1640, w_003_1641, w_003_1642, w_003_1643, w_003_1644, w_003_1645, w_003_1646, w_003_1647, w_003_1648, w_003_1649, w_003_1650, w_003_1651, w_003_1652, w_003_1653, w_003_1654, w_003_1655, w_003_1656, w_003_1657, w_003_1658, w_003_1659, w_003_1660, w_003_1661, w_003_1662, w_003_1663, w_003_1664, w_003_1665, w_003_1666, w_003_1667, w_003_1668, w_003_1669, w_003_1670, w_003_1671, w_003_1672, w_003_1673, w_003_1674, w_003_1675, w_003_1676, w_003_1678, w_003_1679, w_003_1680, w_003_1681, w_003_1682, w_003_1683, w_003_1684, w_003_1685, w_003_1686, w_003_1687, w_003_1689, w_003_1690, w_003_1691, w_003_1693, w_003_1694, w_003_1695, w_003_1696, w_003_1697, w_003_1698, w_003_1699, w_003_1700, w_003_1701, w_003_1702, w_003_1703, w_003_1704, w_003_1705, w_003_1706, w_003_1707, w_003_1708, w_003_1709, w_003_1710, w_003_1711, w_003_1712, w_003_1713, w_003_1714, w_003_1715, w_003_1716, w_003_1717, w_003_1718, w_003_1719, w_003_1720, w_003_1721, w_003_1722, w_003_1723, w_003_1724, w_003_1725, w_003_1726, w_003_1727, w_003_1728, w_003_1729, w_003_1731, w_003_1732, w_003_1733, w_003_1734, w_003_1735, w_003_1736, w_003_1737, w_003_1738, w_003_1739, w_003_1740, w_003_1741, w_003_1742, w_003_1743, w_003_1744, w_003_1745, w_003_1746, w_003_1747, w_003_1748, w_003_1750, w_003_1751, w_003_1752, w_003_1753, w_003_1754, w_003_1755, w_003_1756, w_003_1757, w_003_1758, w_003_1759, w_003_1761, w_003_1762, w_003_1763, w_003_1764, w_003_1765, w_003_1767, w_003_1768, w_003_1769, w_003_1770, w_003_1771, w_003_1774, w_003_1775, w_003_1776, w_003_1777, w_003_1778, w_003_1779, w_003_1780, w_003_1781, w_003_1782, w_003_1783, w_003_1784, w_003_1785, w_003_1786, w_003_1787, w_003_1788, w_003_1789, w_003_1790, w_003_1791, w_003_1792, w_003_1793, w_003_1794, w_003_1795, w_003_1796, w_003_1797, w_003_1798, w_003_1799, w_003_1800, w_003_1801, w_003_1802, w_003_1803, w_003_1804, w_003_1805, w_003_1807, w_003_1808, w_003_1809, w_003_1811, w_003_1812, w_003_1813, w_003_1814, w_003_1815, w_003_1817, w_003_1818, w_003_1819, w_003_1820, w_003_1821, w_003_1822, w_003_1823, w_003_1824, w_003_1825, w_003_1826, w_003_1827, w_003_1828, w_003_1829, w_003_1830, w_003_1831, w_003_1832, w_003_1833, w_003_1834, w_003_1835, w_003_1836, w_003_1837, w_003_1838, w_003_1839, w_003_1841, w_003_1842, w_003_1843, w_003_1844, w_003_1845, w_003_1846, w_003_1847, w_003_1848, w_003_1849, w_003_1850, w_003_1851, w_003_1852, w_003_1854, w_003_1855, w_003_1856, w_003_1857, w_003_1858, w_003_1859, w_003_1860, w_003_1861, w_003_1862, w_003_1863, w_003_1864, w_003_1865, w_003_1866, w_003_1867, w_003_1868, w_003_1869, w_003_1870, w_003_1871, w_003_1872, w_003_1873, w_003_1874, w_003_1875, w_003_1876, w_003_1877, w_003_1878, w_003_1879, w_003_1880, w_003_1881, w_003_1882, w_003_1883, w_003_1884, w_003_1885, w_003_1886, w_003_1887, w_003_1888, w_003_1889, w_003_1890, w_003_1891, w_003_1892, w_003_1893, w_003_1894, w_003_1895, w_003_1897, w_003_1898, w_003_1899, w_003_1900, w_003_1901, w_003_1902, w_003_1904, w_003_1905, w_003_1906, w_003_1907, w_003_1908, w_003_1910, w_003_1911, w_003_1912, w_003_1913, w_003_1914, w_003_1915, w_003_1916, w_003_1917, w_003_1918, w_003_1919, w_003_1920, w_003_1921, w_003_1922, w_003_1923, w_003_1924, w_003_1925, w_003_1926, w_003_1927, w_003_1928, w_003_1929, w_003_1930, w_003_1931, w_003_1932, w_003_1933, w_003_1934, w_003_1935, w_003_1936, w_003_1937, w_003_1938, w_003_1939, w_003_1940, w_003_1942, w_003_1944, w_003_1946, w_003_1947, w_003_1948, w_003_1949, w_003_1950, w_003_1951, w_003_1952, w_003_1953, w_003_1954, w_003_1955, w_003_1956, w_003_1958, w_003_1959, w_003_1960, w_003_1961, w_003_1962, w_003_1963, w_003_1964, w_003_1966, w_003_1967, w_003_1968, w_003_1969, w_003_1970, w_003_1971, w_003_1972, w_003_1973, w_003_1974, w_003_1975, w_003_1976, w_003_1977, w_003_1978, w_003_1979, w_003_1980, w_003_1981, w_003_1982, w_003_1983, w_003_1985, w_003_1986, w_003_1987, w_003_1988, w_003_1990, w_003_1991, w_003_1992, w_003_1993, w_003_1994, w_003_1995, w_003_1996, w_003_1997, w_003_1998, w_003_1999, w_003_2000, w_003_2001, w_003_2002, w_003_2003, w_003_2004, w_003_2005, w_003_2006, w_003_2008, w_003_2009, w_003_2010, w_003_2011, w_003_2012, w_003_2013, w_003_2014, w_003_2015, w_003_2016, w_003_2017, w_003_2019, w_003_2020, w_003_2021, w_003_2022, w_003_2023, w_003_2024, w_003_2025, w_003_2026, w_003_2027, w_003_2030, w_003_2031, w_003_2033, w_003_2035, w_003_2036, w_003_2037, w_003_2038, w_003_2039, w_003_2040, w_003_2041, w_003_2042, w_003_2043, w_003_2044, w_003_2045, w_003_2046, w_003_2047, w_003_2048, w_003_2049, w_003_2050, w_003_2051, w_003_2052, w_003_2053, w_003_2054, w_003_2055, w_003_2056, w_003_2057, w_003_2058, w_003_2059, w_003_2060, w_003_2062, w_003_2063, w_003_2064, w_003_2065, w_003_2066, w_003_2067, w_003_2068, w_003_2069, w_003_2070, w_003_2071, w_003_2072, w_003_2074, w_003_2075, w_003_2076, w_003_2077, w_003_2078, w_003_2079, w_003_2080, w_003_2081, w_003_2082, w_003_2083, w_003_2084, w_003_2085, w_003_2086, w_003_2088, w_003_2089, w_003_2090, w_003_2091, w_003_2092, w_003_2093, w_003_2094, w_003_2095, w_003_2096, w_003_2097, w_003_2098, w_003_2101, w_003_2102, w_003_2103, w_003_2104, w_003_2105, w_003_2106, w_003_2107, w_003_2108, w_003_2109, w_003_2110, w_003_2111, w_003_2112, w_003_2113, w_003_2114, w_003_2115, w_003_2116, w_003_2117, w_003_2118, w_003_2119, w_003_2120, w_003_2121, w_003_2122, w_003_2123, w_003_2124, w_003_2125, w_003_2126, w_003_2127, w_003_2128, w_003_2129, w_003_2130, w_003_2131, w_003_2132, w_003_2133, w_003_2134, w_003_2135, w_003_2136, w_003_2137, w_003_2138, w_003_2139, w_003_2140, w_003_2141, w_003_2142, w_003_2143, w_003_2144, w_003_2145, w_003_2146, w_003_2147, w_003_2148, w_003_2149, w_003_2150, w_003_2151, w_003_2152, w_003_2153, w_003_2154, w_003_2155, w_003_2156, w_003_2157, w_003_2158, w_003_2160, w_003_2161, w_003_2162, w_003_2163, w_003_2165, w_003_2166, w_003_2168, w_003_2170, w_003_2171, w_003_2172, w_003_2173, w_003_2174, w_003_2175, w_003_2176, w_003_2177, w_003_2178, w_003_2179, w_003_2180, w_003_2181, w_003_2182, w_003_2183, w_003_2184, w_003_2186, w_003_2187, w_003_2188, w_003_2189, w_003_2190, w_003_2191, w_003_2192, w_003_2193, w_003_2194, w_003_2195, w_003_2196, w_003_2197, w_003_2198, w_003_2199, w_003_2200, w_003_2201, w_003_2202, w_003_2203, w_003_2204, w_003_2205, w_003_2206, w_003_2208, w_003_2209, w_003_2210, w_003_2211, w_003_2212, w_003_2213, w_003_2214, w_003_2215, w_003_2216, w_003_2217, w_003_2219, w_003_2220, w_003_2221, w_003_2223, w_003_2224, w_003_2225, w_003_2226, w_003_2227, w_003_2228, w_003_2229, w_003_2230, w_003_2232, w_003_2233, w_003_2234, w_003_2235, w_003_2236, w_003_2237, w_003_2238, w_003_2239, w_003_2240, w_003_2241, w_003_2242, w_003_2243, w_003_2244, w_003_2246, w_003_2247, w_003_2248, w_003_2249, w_003_2250, w_003_2251, w_003_2252, w_003_2253, w_003_2254, w_003_2255, w_003_2256, w_003_2257, w_003_2258, w_003_2259, w_003_2260, w_003_2261, w_003_2262, w_003_2263, w_003_2264, w_003_2265, w_003_2266, w_003_2267, w_003_2268, w_003_2269, w_003_2270, w_003_2271, w_003_2272, w_003_2273, w_003_2274, w_003_2275, w_003_2276, w_003_2277, w_003_2278, w_003_2279, w_003_2280, w_003_2281, w_003_2282, w_003_2283, w_003_2284, w_003_2285, w_003_2286, w_003_2288, w_003_2289, w_003_2290, w_003_2291, w_003_2292, w_003_2293, w_003_2294, w_003_2295, w_003_2296, w_003_2297, w_003_2298, w_003_2299, w_003_2300, w_003_2301, w_003_2302, w_003_2303, w_003_2304, w_003_2305, w_003_2306, w_003_2307, w_003_2308, w_003_2309, w_003_2310, w_003_2311, w_003_2312, w_003_2313, w_003_2314, w_003_2315, w_003_2316, w_003_2317, w_003_2318, w_003_2319, w_003_2320, w_003_2321, w_003_2322, w_003_2323, w_003_2324, w_003_2326, w_003_2327, w_003_2328, w_003_2329, w_003_2330, w_003_2331, w_003_2332, w_003_2333, w_003_2334, w_003_2335, w_003_2337, w_003_2338, w_003_2339, w_003_2340, w_003_2341, w_003_2342, w_003_2343, w_003_2344, w_003_2345, w_003_2346, w_003_2347, w_003_2348, w_003_2349, w_003_2350, w_003_2351, w_003_2352, w_003_2354, w_003_2355, w_003_2356, w_003_2357, w_003_2358, w_003_2359, w_003_2360, w_003_2361, w_003_2362, w_003_2363, w_003_2364, w_003_2365, w_003_2366, w_003_2367, w_003_2368, w_003_2369, w_003_2370, w_003_2371, w_003_2372, w_003_2373, w_003_2374, w_003_2375, w_003_2376, w_003_2378, w_003_2379, w_003_2380, w_003_2382, w_003_2383, w_003_2384, w_003_2385, w_003_2387, w_003_2388, w_003_2389, w_003_2390, w_003_2391, w_003_2392, w_003_2393, w_003_2394, w_003_2395, w_003_2396, w_003_2397, w_003_2398, w_003_2399, w_003_2400, w_003_2401, w_003_2402, w_003_2403, w_003_2404, w_003_2405, w_003_2406, w_003_2407, w_003_2408, w_003_2409, w_003_2410, w_003_2411, w_003_2412, w_003_2413, w_003_2414, w_003_2415, w_003_2416, w_003_2417, w_003_2418, w_003_2419, w_003_2420, w_003_2421, w_003_2422, w_003_2423, w_003_2424, w_003_2425, w_003_2426, w_003_2427, w_003_2428, w_003_2429, w_003_2430, w_003_2431, w_003_2433, w_003_2434, w_003_2435, w_003_2436, w_003_2437, w_003_2438, w_003_2439, w_003_2440, w_003_2441, w_003_2442, w_003_2443, w_003_2444, w_003_2445, w_003_2446, w_003_2448, w_003_2449, w_003_2450, w_003_2451, w_003_2452, w_003_2453, w_003_2454, w_003_2455, w_003_2456, w_003_2457, w_003_2458, w_003_2460, w_003_2461, w_003_2463, w_003_2464, w_003_2465, w_003_2466, w_003_2467, w_003_2468, w_003_2469, w_003_2470, w_003_2471, w_003_2472, w_003_2473, w_003_2474, w_003_2475, w_003_2476, w_003_2477, w_003_2478, w_003_2479, w_003_2480, w_003_2481, w_003_2482, w_003_2483, w_003_2484, w_003_2485, w_003_2486, w_003_2487, w_003_2488, w_003_2489, w_003_2490, w_003_2491, w_003_2492, w_003_2493, w_003_2494, w_003_2495, w_003_2496, w_003_2497, w_003_2498, w_003_2499, w_003_2500, w_003_2501, w_003_2502, w_003_2503, w_003_2504, w_003_2505, w_003_2506, w_003_2507, w_003_2508, w_003_2509, w_003_2510, w_003_2511, w_003_2512, w_003_2513, w_003_2515, w_003_2516, w_003_2517, w_003_2518, w_003_2519, w_003_2520, w_003_2522, w_003_2523, w_003_2524, w_003_2525, w_003_2526, w_003_2527, w_003_2528, w_003_2529, w_003_2530, w_003_2531, w_003_2532, w_003_2533, w_003_2535, w_003_2536, w_003_2537, w_003_2538, w_003_2539, w_003_2540, w_003_2541, w_003_2542, w_003_2543, w_003_2544, w_003_2545, w_003_2546, w_003_2547, w_003_2549, w_003_2550, w_003_2551, w_003_2552, w_003_2553, w_003_2554, w_003_2555, w_003_2556, w_003_2557, w_003_2558, w_003_2559, w_003_2560, w_003_2561, w_003_2562, w_003_2563, w_003_2564, w_003_2565, w_003_2566, w_003_2567, w_003_2568, w_003_2569, w_003_2570, w_003_2571, w_003_2572, w_003_2574, w_003_2575, w_003_2576, w_003_2577, w_003_2578, w_003_2579, w_003_2580, w_003_2581, w_003_2582, w_003_2583, w_003_2584, w_003_2585, w_003_2586, w_003_2587, w_003_2588, w_003_2589, w_003_2590, w_003_2591, w_003_2592, w_003_2593, w_003_2594, w_003_2595, w_003_2596, w_003_2597, w_003_2598, w_003_2599, w_003_2600, w_003_2602, w_003_2603, w_003_2606, w_003_2607, w_003_2608, w_003_2609, w_003_2610, w_003_2611, w_003_2612, w_003_2614, w_003_2615, w_003_2616, w_003_2617, w_003_2618, w_003_2619, w_003_2620, w_003_2621, w_003_2622, w_003_2623, w_003_2624, w_003_2625, w_003_2626, w_003_2627, w_003_2628, w_003_2629, w_003_2630, w_003_2631, w_003_2632, w_003_2634, w_003_2635, w_003_2636, w_003_2637, w_003_2639, w_003_2640, w_003_2641, w_003_2642, w_003_2643, w_003_2644, w_003_2645, w_003_2648, w_003_2649, w_003_2650, w_003_2651, w_003_2652, w_003_2653, w_003_2654, w_003_2655, w_003_2656, w_003_2657, w_003_2658, w_003_2659, w_003_2660, w_003_2661, w_003_2662, w_003_2663, w_003_2664, w_003_2665, w_003_2666, w_003_2667, w_003_2668, w_003_2669, w_003_2670, w_003_2671, w_003_2672, w_003_2673, w_003_2674, w_003_2675, w_003_2676, w_003_2677, w_003_2678, w_003_2679, w_003_2680, w_003_2681, w_003_2682, w_003_2683, w_003_2684, w_003_2685, w_003_2686, w_003_2687, w_003_2688, w_003_2689, w_003_2690, w_003_2691, w_003_2692, w_003_2693, w_003_2694, w_003_2696, w_003_2697, w_003_2698, w_003_2699, w_003_2700, w_003_2701, w_003_2702, w_003_2703, w_003_2704, w_003_2705, w_003_2706, w_003_2707, w_003_2708, w_003_2709, w_003_2710, w_003_2711, w_003_2712, w_003_2713, w_003_2714, w_003_2715, w_003_2716, w_003_2717, w_003_2718, w_003_2719, w_003_2720, w_003_2721, w_003_2722, w_003_2723, w_003_2724, w_003_2725, w_003_2726, w_003_2727, w_003_2728, w_003_2729, w_003_2730, w_003_2731, w_003_2732, w_003_2733, w_003_2734, w_003_2735, w_003_2736, w_003_2737, w_003_2738, w_003_2739, w_003_2740, w_003_2741, w_003_2742, w_003_2743, w_003_2744, w_003_2745, w_003_2747, w_003_2748, w_003_2749, w_003_2750, w_003_2751, w_003_2752, w_003_2753, w_003_2754, w_003_2755, w_003_2756, w_003_2758, w_003_2759, w_003_2760, w_003_2761, w_003_2762, w_003_2763, w_003_2764, w_003_2765, w_003_2766, w_003_2767, w_003_2768, w_003_2769, w_003_2770, w_003_2771, w_003_2772, w_003_2773, w_003_2774, w_003_2775, w_003_2776, w_003_2777, w_003_2778, w_003_2779, w_003_2780, w_003_2781, w_003_2782, w_003_2784, w_003_2785, w_003_2786, w_003_2787, w_003_2788, w_003_2789, w_003_2790, w_003_2791, w_003_2792, w_003_2793, w_003_2794, w_003_2795, w_003_2796, w_003_2797, w_003_2798, w_003_2799, w_003_2800, w_003_2801, w_003_2802, w_003_2803, w_003_2804, w_003_2805, w_003_2806, w_003_2807, w_003_2808, w_003_2809, w_003_2810, w_003_2811, w_003_2812, w_003_2814, w_003_2815, w_003_2816, w_003_2817, w_003_2818, w_003_2819, w_003_2820, w_003_2821, w_003_2822, w_003_2823, w_003_2824, w_003_2825, w_003_2826, w_003_2827, w_003_2828, w_003_2829, w_003_2830, w_003_2832, w_003_2833, w_003_2834, w_003_2835, w_003_2836, w_003_2837, w_003_2838, w_003_2839, w_003_2840, w_003_2841, w_003_2842, w_003_2843, w_003_2844, w_003_2846, w_003_2847, w_003_2848, w_003_2849, w_003_2850, w_003_2851, w_003_2852, w_003_2853, w_003_2854, w_003_2855, w_003_2856, w_003_2857, w_003_2858, w_003_2859, w_003_2860, w_003_2861, w_003_2862, w_003_2863, w_003_2864, w_003_2865, w_003_2866, w_003_2868, w_003_2869, w_003_2870, w_003_2871, w_003_2872, w_003_2873, w_003_2874, w_003_2876, w_003_2877, w_003_2878, w_003_2879, w_003_2880, w_003_2881, w_003_2882, w_003_2883, w_003_2884, w_003_2885, w_003_2886, w_003_2887, w_003_2888, w_003_2889, w_003_2890, w_003_2892, w_003_2893, w_003_2894, w_003_2895, w_003_2896, w_003_2897, w_003_2898, w_003_2899, w_003_2900, w_003_2901, w_003_2902, w_003_2903, w_003_2904, w_003_2905, w_003_2906, w_003_2907, w_003_2908, w_003_2910, w_003_2911, w_003_2912, w_003_2913, w_003_2914, w_003_2917, w_003_2918, w_003_2919, w_003_2920, w_003_2921, w_003_2922, w_003_2923, w_003_2924, w_003_2925, w_003_2926, w_003_2927, w_003_2928, w_003_2929, w_003_2930, w_003_2931, w_003_2932, w_003_2933, w_003_2934, w_003_2935, w_003_2936, w_003_2937, w_003_2938, w_003_2939, w_003_2940, w_003_2941, w_003_2942, w_003_2943, w_003_2944, w_003_2945, w_003_2946, w_003_2947, w_003_2948, w_003_2949, w_003_2950, w_003_2951, w_003_2952, w_003_2953, w_003_2954, w_003_2955, w_003_2956, w_003_2957, w_003_2958, w_003_2959, w_003_2960, w_003_2962, w_003_2963, w_003_2964, w_003_2965, w_003_2966, w_003_2967, w_003_2968, w_003_2970, w_003_2972, w_003_2973, w_003_2974, w_003_2975, w_003_2976, w_003_2977, w_003_2978, w_003_2979, w_003_2980, w_003_2981, w_003_2982, w_003_2983, w_003_2984, w_003_2985, w_003_2986, w_003_2987, w_003_2988, w_003_2989, w_003_2990, w_003_2991, w_003_2992, w_003_2993, w_003_2994, w_003_2995, w_003_2997, w_003_2998, w_003_2999, w_003_3000, w_003_3001, w_003_3002, w_003_3003, w_003_3004, w_003_3005, w_003_3006, w_003_3007, w_003_3008, w_003_3010, w_003_3011, w_003_3012, w_003_3013, w_003_3014, w_003_3015, w_003_3016, w_003_3017, w_003_3018, w_003_3019, w_003_3020, w_003_3021, w_003_3022, w_003_3023, w_003_3024, w_003_3025, w_003_3026, w_003_3027, w_003_3028, w_003_3029, w_003_3030, w_003_3031, w_003_3033, w_003_3034, w_003_3035, w_003_3036, w_003_3037, w_003_3038, w_003_3039, w_003_3040, w_003_3041, w_003_3042, w_003_3043, w_003_3044, w_003_3045, w_003_3046, w_003_3047, w_003_3048, w_003_3049, w_003_3050, w_003_3051, w_003_3052, w_003_3053, w_003_3054, w_003_3055, w_003_3056, w_003_3057, w_003_3058, w_003_3059, w_003_3060, w_003_3061, w_003_3062, w_003_3063, w_003_3064, w_003_3065, w_003_3067, w_003_3068, w_003_3069, w_003_3070, w_003_3071, w_003_3072, w_003_3073, w_003_3074, w_003_3075, w_003_3076, w_003_3077, w_003_3078, w_003_3079, w_003_3080, w_003_3081, w_003_3082, w_003_3083, w_003_3084, w_003_3085, w_003_3086, w_003_3087, w_003_3088, w_003_3089, w_003_3090, w_003_3091, w_003_3092, w_003_3093, w_003_3094, w_003_3095, w_003_3096, w_003_3097, w_003_3098, w_003_3099, w_003_3100, w_003_3101, w_003_3102, w_003_3103, w_003_3105, w_003_3106, w_003_3107, w_003_3108, w_003_3109, w_003_3111, w_003_3112, w_003_3113, w_003_3114, w_003_3115, w_003_3116, w_003_3117, w_003_3118, w_003_3119, w_003_3120, w_003_3121, w_003_3122, w_003_3123, w_003_3124, w_003_3125, w_003_3126, w_003_3127, w_003_3128, w_003_3129, w_003_3130, w_003_3131, w_003_3132, w_003_3133, w_003_3134, w_003_3135, w_003_3136, w_003_3137, w_003_3138, w_003_3139, w_003_3140, w_003_3141, w_003_3142, w_003_3143, w_003_3144, w_003_3145, w_003_3146, w_003_3147, w_003_3148, w_003_3149, w_003_3150, w_003_3151, w_003_3152, w_003_3153, w_003_3155, w_003_3156, w_003_3157, w_003_3158, w_003_3159, w_003_3160, w_003_3161, w_003_3162, w_003_3163, w_003_3164, w_003_3165, w_003_3166, w_003_3168, w_003_3169, w_003_3171, w_003_3172, w_003_3173, w_003_3174, w_003_3175, w_003_3176, w_003_3177, w_003_3178, w_003_3179, w_003_3180, w_003_3181, w_003_3182, w_003_3183, w_003_3184, w_003_3185, w_003_3186, w_003_3187, w_003_3188, w_003_3189, w_003_3190, w_003_3191, w_003_3192, w_003_3193, w_003_3194, w_003_3195, w_003_3197, w_003_3198, w_003_3199, w_003_3200, w_003_3201, w_003_3202, w_003_3203, w_003_3205, w_003_3206, w_003_3207, w_003_3208, w_003_3209, w_003_3210, w_003_3211, w_003_3212, w_003_3213, w_003_3214, w_003_3215, w_003_3216, w_003_3217, w_003_3220, w_003_3221, w_003_3222, w_003_3223, w_003_3224, w_003_3225, w_003_3226, w_003_3227, w_003_3228, w_003_3229, w_003_3230, w_003_3231, w_003_3232, w_003_3233, w_003_3234, w_003_3235, w_003_3236, w_003_3237, w_003_3238, w_003_3239, w_003_3240, w_003_3241, w_003_3242, w_003_3243, w_003_3244, w_003_3246, w_003_3247, w_003_3248, w_003_3250, w_003_3251, w_003_3252, w_003_3253, w_003_3254, w_003_3255, w_003_3256, w_003_3257, w_003_3258, w_003_3259, w_003_3260, w_003_3261, w_003_3262, w_003_3263, w_003_3264, w_003_3265, w_003_3266, w_003_3267, w_003_3268, w_003_3269, w_003_3271, w_003_3272, w_003_3274, w_003_3275, w_003_3276, w_003_3277, w_003_3278, w_003_3279, w_003_3280, w_003_3281, w_003_3283, w_003_3284, w_003_3285, w_003_3286, w_003_3287, w_003_3288, w_003_3289, w_003_3290, w_003_3294, w_003_3295, w_003_3296, w_003_3298, w_003_3299, w_003_3300, w_003_3301, w_003_3302, w_003_3303, w_003_3305, w_003_3306, w_003_3307, w_003_3308, w_003_3309, w_003_3311, w_003_3312, w_003_3313, w_003_3314, w_003_3315, w_003_3316, w_003_3317, w_003_3318, w_003_3319, w_003_3320, w_003_3321, w_003_3322, w_003_3323;
  wire w_004_000, w_004_002, w_004_003, w_004_004, w_004_005, w_004_006, w_004_007, w_004_008, w_004_009, w_004_010, w_004_011, w_004_012, w_004_013, w_004_014, w_004_015, w_004_016, w_004_017, w_004_018, w_004_019, w_004_020, w_004_021, w_004_022, w_004_023, w_004_024, w_004_025, w_004_026, w_004_027, w_004_028, w_004_029, w_004_030, w_004_031, w_004_032, w_004_033, w_004_034, w_004_035, w_004_036, w_004_037, w_004_038, w_004_039, w_004_040, w_004_041, w_004_042, w_004_043, w_004_044, w_004_045, w_004_046, w_004_047, w_004_048, w_004_049, w_004_050, w_004_051, w_004_052, w_004_053, w_004_054, w_004_055, w_004_056, w_004_057, w_004_058, w_004_059, w_004_060, w_004_061, w_004_062, w_004_063, w_004_064, w_004_065, w_004_066, w_004_067, w_004_068, w_004_069, w_004_070, w_004_071, w_004_072, w_004_073, w_004_074, w_004_075, w_004_076, w_004_077, w_004_078, w_004_079, w_004_080, w_004_081, w_004_082, w_004_083, w_004_084, w_004_085, w_004_086, w_004_087, w_004_088, w_004_089, w_004_090, w_004_091, w_004_092, w_004_093, w_004_094, w_004_095, w_004_096, w_004_097, w_004_098, w_004_099, w_004_100, w_004_101, w_004_102, w_004_103, w_004_104, w_004_105, w_004_106, w_004_107, w_004_108, w_004_109, w_004_110, w_004_111, w_004_112, w_004_113, w_004_115, w_004_116, w_004_117, w_004_118, w_004_119, w_004_120, w_004_121, w_004_122, w_004_123, w_004_124, w_004_125, w_004_126, w_004_127, w_004_128, w_004_129, w_004_130, w_004_131, w_004_132, w_004_133, w_004_135, w_004_136, w_004_137, w_004_138, w_004_139, w_004_140, w_004_141, w_004_142, w_004_143, w_004_144, w_004_145, w_004_146, w_004_147, w_004_148, w_004_149, w_004_150, w_004_151, w_004_152, w_004_153, w_004_154, w_004_155, w_004_156, w_004_157, w_004_158, w_004_159, w_004_160, w_004_161, w_004_162, w_004_163, w_004_164, w_004_165, w_004_166, w_004_167, w_004_168, w_004_169, w_004_170, w_004_171, w_004_172, w_004_173, w_004_174, w_004_175, w_004_176, w_004_177, w_004_178, w_004_179, w_004_180, w_004_181, w_004_182, w_004_183, w_004_184, w_004_185, w_004_186, w_004_187, w_004_188, w_004_189, w_004_190, w_004_191, w_004_192, w_004_193, w_004_194, w_004_195, w_004_196, w_004_197, w_004_198, w_004_199, w_004_200, w_004_201, w_004_202, w_004_203, w_004_204, w_004_205, w_004_206, w_004_207, w_004_208, w_004_209, w_004_210, w_004_211, w_004_212, w_004_213, w_004_214, w_004_215, w_004_216, w_004_217, w_004_218, w_004_219, w_004_220, w_004_221, w_004_222, w_004_223, w_004_224, w_004_225, w_004_226, w_004_227, w_004_228, w_004_229, w_004_230, w_004_231, w_004_232, w_004_233, w_004_234, w_004_235, w_004_236, w_004_237, w_004_238, w_004_239, w_004_240, w_004_241, w_004_242, w_004_243, w_004_244, w_004_245, w_004_246, w_004_247, w_004_248, w_004_249, w_004_250, w_004_251, w_004_252, w_004_253, w_004_254, w_004_255, w_004_256, w_004_257, w_004_259, w_004_260, w_004_261, w_004_262, w_004_265, w_004_266, w_004_267, w_004_268, w_004_269, w_004_270, w_004_272, w_004_273, w_004_274, w_004_275, w_004_277, w_004_278, w_004_279, w_004_280, w_004_281, w_004_282, w_004_284, w_004_285, w_004_287, w_004_288, w_004_289, w_004_290, w_004_291, w_004_292, w_004_293, w_004_294, w_004_295, w_004_296, w_004_297, w_004_299, w_004_300, w_004_303, w_004_304, w_004_305, w_004_306, w_004_307, w_004_308, w_004_309, w_004_310, w_004_311, w_004_312, w_004_313, w_004_314, w_004_315, w_004_316, w_004_317, w_004_318, w_004_319, w_004_320, w_004_321, w_004_322, w_004_323, w_004_324, w_004_326, w_004_327, w_004_328, w_004_329, w_004_331, w_004_332, w_004_334, w_004_335, w_004_336, w_004_337, w_004_338, w_004_339, w_004_340, w_004_341, w_004_343, w_004_344, w_004_345, w_004_346, w_004_347, w_004_348, w_004_349, w_004_351, w_004_353, w_004_354, w_004_356, w_004_357, w_004_358, w_004_359, w_004_360, w_004_361, w_004_362, w_004_363, w_004_364, w_004_365, w_004_366, w_004_367, w_004_368, w_004_369, w_004_370, w_004_371, w_004_372, w_004_373, w_004_374, w_004_375, w_004_376, w_004_378, w_004_379, w_004_381, w_004_382, w_004_383, w_004_385, w_004_386, w_004_387, w_004_389, w_004_390, w_004_391, w_004_392, w_004_396, w_004_397, w_004_398, w_004_399, w_004_400, w_004_401, w_004_403, w_004_404, w_004_405, w_004_406, w_004_407, w_004_408, w_004_409, w_004_410, w_004_411, w_004_412, w_004_413, w_004_414, w_004_415, w_004_416, w_004_417, w_004_418, w_004_419, w_004_420, w_004_421, w_004_422, w_004_423, w_004_424, w_004_425, w_004_427, w_004_428, w_004_430, w_004_431, w_004_433, w_004_434, w_004_435, w_004_436, w_004_437, w_004_438, w_004_439, w_004_442, w_004_443, w_004_444, w_004_445, w_004_446, w_004_447, w_004_448, w_004_449, w_004_450, w_004_451, w_004_452, w_004_453, w_004_454, w_004_455, w_004_456, w_004_459, w_004_460, w_004_461, w_004_462, w_004_463, w_004_464, w_004_465, w_004_466, w_004_467, w_004_469, w_004_471, w_004_472, w_004_474, w_004_475, w_004_476, w_004_477, w_004_478, w_004_479, w_004_481, w_004_482, w_004_483, w_004_484, w_004_485, w_004_486, w_004_487, w_004_489, w_004_490, w_004_491, w_004_492, w_004_493, w_004_494, w_004_495, w_004_497, w_004_499, w_004_500, w_004_501, w_004_502, w_004_503, w_004_504, w_004_505, w_004_506, w_004_507, w_004_508, w_004_509, w_004_510, w_004_511, w_004_512, w_004_513, w_004_514, w_004_515, w_004_516, w_004_517, w_004_518, w_004_519, w_004_520, w_004_521, w_004_522, w_004_523, w_004_524, w_004_526, w_004_527, w_004_528, w_004_529, w_004_530, w_004_531, w_004_532, w_004_533, w_004_534, w_004_535, w_004_536, w_004_537, w_004_538, w_004_539, w_004_540, w_004_541, w_004_542, w_004_543, w_004_544, w_004_546, w_004_547, w_004_548, w_004_550, w_004_551, w_004_552, w_004_553, w_004_554, w_004_555, w_004_556, w_004_558, w_004_559, w_004_560, w_004_561, w_004_563, w_004_564, w_004_565, w_004_566, w_004_567, w_004_568, w_004_569, w_004_570, w_004_571, w_004_572, w_004_573, w_004_574, w_004_575, w_004_576, w_004_577, w_004_578, w_004_579, w_004_580, w_004_581, w_004_582, w_004_583, w_004_584, w_004_585, w_004_586, w_004_587, w_004_588, w_004_589, w_004_590, w_004_591, w_004_592, w_004_593, w_004_594, w_004_595, w_004_596, w_004_597, w_004_598, w_004_600, w_004_601, w_004_602, w_004_603, w_004_604, w_004_605, w_004_606, w_004_607, w_004_608, w_004_609, w_004_610, w_004_611, w_004_612, w_004_614, w_004_615, w_004_616, w_004_617, w_004_618, w_004_619, w_004_621, w_004_622, w_004_623, w_004_624, w_004_625, w_004_626, w_004_627, w_004_628, w_004_629, w_004_630, w_004_631, w_004_632, w_004_633, w_004_634, w_004_635, w_004_636, w_004_637, w_004_639, w_004_640, w_004_641, w_004_642, w_004_643, w_004_645, w_004_646, w_004_647, w_004_648, w_004_649, w_004_650, w_004_651, w_004_652, w_004_653, w_004_654, w_004_655, w_004_656, w_004_657, w_004_658, w_004_659, w_004_660, w_004_661, w_004_662, w_004_663, w_004_664, w_004_665, w_004_666, w_004_667, w_004_668, w_004_669, w_004_670, w_004_671, w_004_673, w_004_674, w_004_675, w_004_678, w_004_679, w_004_680, w_004_681, w_004_682, w_004_683, w_004_684, w_004_685, w_004_686, w_004_687, w_004_688, w_004_689, w_004_690, w_004_691, w_004_692, w_004_693, w_004_694, w_004_695, w_004_696, w_004_697, w_004_698, w_004_700, w_004_701, w_004_702, w_004_703, w_004_704, w_004_705, w_004_706, w_004_707, w_004_708, w_004_709, w_004_710, w_004_711, w_004_713, w_004_714, w_004_715, w_004_716, w_004_717, w_004_718, w_004_719, w_004_720, w_004_722, w_004_724, w_004_725, w_004_726, w_004_727, w_004_728, w_004_729, w_004_730, w_004_731, w_004_732, w_004_733, w_004_734, w_004_735, w_004_736, w_004_737, w_004_738, w_004_739, w_004_740, w_004_741, w_004_743, w_004_744, w_004_745, w_004_746, w_004_747, w_004_748, w_004_749, w_004_750, w_004_751, w_004_752, w_004_754, w_004_755, w_004_756, w_004_757, w_004_758, w_004_759, w_004_760, w_004_761, w_004_762, w_004_763, w_004_764, w_004_765, w_004_766, w_004_767, w_004_768, w_004_769, w_004_770, w_004_771, w_004_772, w_004_773, w_004_774, w_004_775, w_004_776, w_004_777, w_004_779, w_004_780, w_004_781, w_004_782, w_004_783, w_004_784, w_004_786, w_004_787, w_004_788, w_004_789, w_004_790, w_004_791, w_004_792, w_004_793, w_004_794, w_004_795, w_004_796, w_004_797, w_004_798, w_004_799, w_004_800, w_004_802, w_004_805, w_004_806, w_004_807, w_004_808, w_004_809, w_004_810, w_004_811, w_004_812, w_004_813, w_004_814, w_004_815, w_004_816, w_004_817, w_004_818, w_004_819, w_004_821, w_004_823, w_004_824, w_004_825, w_004_826, w_004_827, w_004_828, w_004_829, w_004_830, w_004_831, w_004_832, w_004_833, w_004_834, w_004_835, w_004_837, w_004_839, w_004_840, w_004_841, w_004_842, w_004_843, w_004_845, w_004_846, w_004_847, w_004_848, w_004_849, w_004_850, w_004_851, w_004_852, w_004_853, w_004_854, w_004_856, w_004_857, w_004_858, w_004_860, w_004_861, w_004_862, w_004_863, w_004_864, w_004_865, w_004_866, w_004_867, w_004_868, w_004_869, w_004_870, w_004_871, w_004_872, w_004_873, w_004_874, w_004_876, w_004_877, w_004_878, w_004_879, w_004_880, w_004_881, w_004_882, w_004_883, w_004_884, w_004_885, w_004_886, w_004_887, w_004_888, w_004_889, w_004_890, w_004_891, w_004_892, w_004_893, w_004_894, w_004_895, w_004_896, w_004_897, w_004_898, w_004_899, w_004_900, w_004_901, w_004_902, w_004_903, w_004_904, w_004_905, w_004_906, w_004_907, w_004_908, w_004_909, w_004_910, w_004_911, w_004_912, w_004_913, w_004_914, w_004_915, w_004_916, w_004_917, w_004_918, w_004_919, w_004_920, w_004_921, w_004_922, w_004_923, w_004_925, w_004_926, w_004_927, w_004_929, w_004_930, w_004_931, w_004_932, w_004_933, w_004_934, w_004_935, w_004_936, w_004_937, w_004_939, w_004_940, w_004_941, w_004_942, w_004_943, w_004_944, w_004_945, w_004_946, w_004_947, w_004_949, w_004_950, w_004_951, w_004_952, w_004_953, w_004_954, w_004_956, w_004_957, w_004_958, w_004_959, w_004_960, w_004_961, w_004_962, w_004_963, w_004_964, w_004_966, w_004_967, w_004_970, w_004_971, w_004_972, w_004_973, w_004_974, w_004_975, w_004_976, w_004_977, w_004_978, w_004_979, w_004_980, w_004_981, w_004_983, w_004_984, w_004_985, w_004_986, w_004_987, w_004_988, w_004_989, w_004_990, w_004_991, w_004_992, w_004_993, w_004_994, w_004_995, w_004_996, w_004_997, w_004_998, w_004_999, w_004_1000, w_004_1001, w_004_1002, w_004_1003, w_004_1004, w_004_1006, w_004_1007, w_004_1008, w_004_1009, w_004_1010, w_004_1011, w_004_1012, w_004_1013, w_004_1014, w_004_1015, w_004_1016, w_004_1018, w_004_1020, w_004_1021, w_004_1022, w_004_1023, w_004_1025, w_004_1026, w_004_1027, w_004_1028, w_004_1029, w_004_1030, w_004_1032, w_004_1033, w_004_1034, w_004_1035, w_004_1036, w_004_1037, w_004_1038, w_004_1039, w_004_1040, w_004_1041, w_004_1042, w_004_1043, w_004_1044, w_004_1045, w_004_1046, w_004_1047, w_004_1048, w_004_1050, w_004_1051, w_004_1052, w_004_1053, w_004_1055, w_004_1056, w_004_1057, w_004_1058, w_004_1059, w_004_1060, w_004_1061, w_004_1062, w_004_1064, w_004_1065, w_004_1066, w_004_1067, w_004_1068, w_004_1069, w_004_1070, w_004_1071, w_004_1072, w_004_1073, w_004_1074, w_004_1076, w_004_1077, w_004_1078, w_004_1079, w_004_1080, w_004_1081, w_004_1082, w_004_1083, w_004_1084, w_004_1085, w_004_1086, w_004_1087, w_004_1091, w_004_1092, w_004_1093, w_004_1095, w_004_1096, w_004_1097, w_004_1098, w_004_1099, w_004_1100, w_004_1101, w_004_1103, w_004_1104, w_004_1105, w_004_1106, w_004_1108, w_004_1109, w_004_1110, w_004_1111, w_004_1112, w_004_1113, w_004_1114, w_004_1116, w_004_1117, w_004_1118, w_004_1119, w_004_1120, w_004_1121, w_004_1122, w_004_1123, w_004_1124, w_004_1125, w_004_1126, w_004_1127, w_004_1128, w_004_1129, w_004_1130, w_004_1131, w_004_1132, w_004_1134, w_004_1135, w_004_1136, w_004_1137, w_004_1138, w_004_1140, w_004_1141, w_004_1142, w_004_1143, w_004_1144, w_004_1146, w_004_1147, w_004_1148, w_004_1149, w_004_1150, w_004_1151, w_004_1152, w_004_1153, w_004_1154, w_004_1156, w_004_1157, w_004_1158, w_004_1159, w_004_1160, w_004_1161, w_004_1162, w_004_1163, w_004_1164, w_004_1166, w_004_1168, w_004_1169, w_004_1170, w_004_1171, w_004_1172, w_004_1173, w_004_1174, w_004_1175, w_004_1176, w_004_1177, w_004_1178, w_004_1179, w_004_1180, w_004_1181, w_004_1182, w_004_1183, w_004_1184, w_004_1185, w_004_1186, w_004_1187, w_004_1188, w_004_1189, w_004_1190, w_004_1191, w_004_1193, w_004_1195, w_004_1196, w_004_1197, w_004_1198, w_004_1199, w_004_1201, w_004_1202, w_004_1203, w_004_1204, w_004_1205, w_004_1206, w_004_1207, w_004_1208, w_004_1209, w_004_1210, w_004_1211, w_004_1212, w_004_1213, w_004_1214, w_004_1215, w_004_1216, w_004_1217, w_004_1218, w_004_1219, w_004_1220, w_004_1222, w_004_1223, w_004_1224, w_004_1225, w_004_1227, w_004_1229, w_004_1230, w_004_1231, w_004_1232, w_004_1234, w_004_1235, w_004_1237, w_004_1238, w_004_1239, w_004_1240, w_004_1241, w_004_1242, w_004_1243, w_004_1244, w_004_1245, w_004_1246, w_004_1247, w_004_1248, w_004_1249, w_004_1250, w_004_1251, w_004_1252, w_004_1253, w_004_1254, w_004_1255, w_004_1256, w_004_1257, w_004_1258, w_004_1259, w_004_1260, w_004_1261, w_004_1262, w_004_1264, w_004_1266, w_004_1267, w_004_1269, w_004_1270, w_004_1271, w_004_1273, w_004_1274, w_004_1275, w_004_1276, w_004_1279, w_004_1280, w_004_1281, w_004_1282, w_004_1283, w_004_1284, w_004_1285, w_004_1286, w_004_1287, w_004_1288, w_004_1289, w_004_1290, w_004_1291, w_004_1292, w_004_1293, w_004_1294, w_004_1295, w_004_1296, w_004_1297, w_004_1298, w_004_1300, w_004_1301, w_004_1302, w_004_1304, w_004_1305, w_004_1306, w_004_1307, w_004_1309, w_004_1310, w_004_1311, w_004_1312, w_004_1313, w_004_1314, w_004_1315, w_004_1316, w_004_1317, w_004_1318, w_004_1319, w_004_1320, w_004_1321, w_004_1322, w_004_1324, w_004_1325, w_004_1326, w_004_1327, w_004_1328, w_004_1329, w_004_1330, w_004_1331, w_004_1332, w_004_1333, w_004_1334, w_004_1335, w_004_1336, w_004_1337, w_004_1338, w_004_1339, w_004_1340, w_004_1342, w_004_1343, w_004_1344, w_004_1345, w_004_1347, w_004_1348, w_004_1349, w_004_1350, w_004_1351, w_004_1352, w_004_1353, w_004_1354, w_004_1355, w_004_1356, w_004_1357, w_004_1358, w_004_1360, w_004_1361, w_004_1362, w_004_1363, w_004_1364, w_004_1366, w_004_1367, w_004_1368, w_004_1369, w_004_1371, w_004_1372, w_004_1373, w_004_1374, w_004_1375, w_004_1376, w_004_1377, w_004_1379, w_004_1380, w_004_1381, w_004_1382, w_004_1383, w_004_1386, w_004_1387, w_004_1388, w_004_1389, w_004_1390, w_004_1391, w_004_1392, w_004_1393, w_004_1394, w_004_1395, w_004_1396, w_004_1397, w_004_1398, w_004_1399, w_004_1401, w_004_1402, w_004_1403, w_004_1404, w_004_1405, w_004_1406, w_004_1407, w_004_1408, w_004_1410, w_004_1411, w_004_1412, w_004_1413, w_004_1414, w_004_1415, w_004_1416, w_004_1417, w_004_1418, w_004_1419, w_004_1420, w_004_1421, w_004_1422, w_004_1423, w_004_1424, w_004_1425, w_004_1426, w_004_1427, w_004_1428, w_004_1429, w_004_1430, w_004_1431, w_004_1432, w_004_1433, w_004_1434, w_004_1435, w_004_1436, w_004_1437, w_004_1438, w_004_1439, w_004_1440, w_004_1442, w_004_1443, w_004_1444, w_004_1445, w_004_1446, w_004_1447, w_004_1448, w_004_1449, w_004_1450, w_004_1451, w_004_1452, w_004_1453, w_004_1454, w_004_1455, w_004_1457, w_004_1458, w_004_1459, w_004_1460, w_004_1461, w_004_1462, w_004_1464, w_004_1465, w_004_1467, w_004_1468, w_004_1469, w_004_1471, w_004_1472, w_004_1474, w_004_1475, w_004_1476, w_004_1477, w_004_1478, w_004_1479, w_004_1480, w_004_1482, w_004_1483, w_004_1484, w_004_1485, w_004_1487, w_004_1488, w_004_1489, w_004_1491, w_004_1492, w_004_1493, w_004_1494, w_004_1496, w_004_1497, w_004_1498, w_004_1499, w_004_1500, w_004_1501, w_004_1502, w_004_1504, w_004_1505, w_004_1506, w_004_1508, w_004_1509, w_004_1510, w_004_1511, w_004_1513, w_004_1514, w_004_1515, w_004_1516, w_004_1517, w_004_1518, w_004_1519, w_004_1520, w_004_1522, w_004_1524, w_004_1525, w_004_1526, w_004_1528, w_004_1529, w_004_1531, w_004_1532, w_004_1533, w_004_1534, w_004_1535, w_004_1536, w_004_1538, w_004_1539, w_004_1540, w_004_1541, w_004_1542, w_004_1543, w_004_1545, w_004_1546, w_004_1547, w_004_1548, w_004_1549, w_004_1550, w_004_1551, w_004_1552, w_004_1553, w_004_1554, w_004_1555, w_004_1556, w_004_1557, w_004_1558, w_004_1559, w_004_1560, w_004_1561, w_004_1562, w_004_1563, w_004_1564, w_004_1565, w_004_1566, w_004_1567, w_004_1568, w_004_1569, w_004_1570, w_004_1571, w_004_1573, w_004_1574, w_004_1575, w_004_1576, w_004_1577, w_004_1578, w_004_1579, w_004_1580, w_004_1581, w_004_1582, w_004_1583, w_004_1584, w_004_1585, w_004_1586, w_004_1587, w_004_1588, w_004_1589, w_004_1590, w_004_1591, w_004_1592, w_004_1593, w_004_1594, w_004_1595, w_004_1596, w_004_1597, w_004_1599, w_004_1600, w_004_1601, w_004_1602, w_004_1603, w_004_1604, w_004_1605, w_004_1606, w_004_1607, w_004_1608, w_004_1611, w_004_1612, w_004_1613, w_004_1614, w_004_1615, w_004_1616, w_004_1618, w_004_1619, w_004_1620, w_004_1621, w_004_1622, w_004_1623, w_004_1624, w_004_1625, w_004_1626, w_004_1627, w_004_1628, w_004_1630, w_004_1631, w_004_1632, w_004_1633, w_004_1634, w_004_1635, w_004_1636, w_004_1637, w_004_1638, w_004_1639, w_004_1640, w_004_1641, w_004_1642, w_004_1643, w_004_1644, w_004_1645, w_004_1646, w_004_1647, w_004_1648, w_004_1649, w_004_1651, w_004_1652, w_004_1653, w_004_1654, w_004_1655, w_004_1657, w_004_1658, w_004_1659, w_004_1660, w_004_1661, w_004_1662, w_004_1663, w_004_1664, w_004_1665, w_004_1666, w_004_1667, w_004_1668, w_004_1669, w_004_1670, w_004_1671, w_004_1672, w_004_1673, w_004_1674, w_004_1675, w_004_1676, w_004_1677, w_004_1678, w_004_1679, w_004_1680, w_004_1681, w_004_1682, w_004_1683, w_004_1684, w_004_1686, w_004_1687, w_004_1688, w_004_1689, w_004_1690, w_004_1691, w_004_1692, w_004_1693, w_004_1694, w_004_1695, w_004_1696, w_004_1697, w_004_1698, w_004_1699, w_004_1700, w_004_1701, w_004_1702, w_004_1703, w_004_1704, w_004_1705, w_004_1706, w_004_1709, w_004_1710, w_004_1713, w_004_1714, w_004_1715, w_004_1716, w_004_1717, w_004_1718, w_004_1719, w_004_1720, w_004_1722, w_004_1723, w_004_1724, w_004_1726, w_004_1727, w_004_1728, w_004_1729, w_004_1730, w_004_1731, w_004_1732, w_004_1733, w_004_1734, w_004_1736, w_004_1737, w_004_1738, w_004_1739, w_004_1740, w_004_1741, w_004_1742, w_004_1743, w_004_1744, w_004_1745, w_004_1746, w_004_1747, w_004_1748, w_004_1749, w_004_1750, w_004_1751, w_004_1752, w_004_1753, w_004_1754, w_004_1755, w_004_1756, w_004_1757, w_004_1758, w_004_1759, w_004_1760, w_004_1761, w_004_1762, w_004_1763, w_004_1764, w_004_1765, w_004_1766, w_004_1767, w_004_1768, w_004_1769, w_004_1770, w_004_1772, w_004_1773, w_004_1774, w_004_1775, w_004_1776, w_004_1777, w_004_1778, w_004_1779, w_004_1780, w_004_1781, w_004_1782, w_004_1783, w_004_1784, w_004_1785, w_004_1787, w_004_1788, w_004_1789, w_004_1790, w_004_1791, w_004_1793, w_004_1794, w_004_1795, w_004_1796, w_004_1797, w_004_1798, w_004_1799, w_004_1800, w_004_1801, w_004_1802, w_004_1803, w_004_1804, w_004_1806, w_004_1807, w_004_1808, w_004_1809, w_004_1811, w_004_1812, w_004_1813, w_004_1814, w_004_1816, w_004_1817, w_004_1818, w_004_1819, w_004_1820, w_004_1821, w_004_1822, w_004_1825, w_004_1826, w_004_1827, w_004_1828, w_004_1829, w_004_1831, w_004_1832, w_004_1834, w_004_1835, w_004_1836, w_004_1837, w_004_1838, w_004_1839, w_004_1840, w_004_1842, w_004_1843, w_004_1844, w_004_1845, w_004_1847, w_004_1848, w_004_1849, w_004_1850, w_004_1851, w_004_1853, w_004_1855, w_004_1856, w_004_1857, w_004_1858, w_004_1859, w_004_1860, w_004_1861, w_004_1862, w_004_1863, w_004_1864, w_004_1866, w_004_1867, w_004_1868, w_004_1869, w_004_1870, w_004_1871, w_004_1872, w_004_1873, w_004_1874, w_004_1875, w_004_1876, w_004_1877, w_004_1878, w_004_1879, w_004_1880, w_004_1881, w_004_1882, w_004_1883, w_004_1884, w_004_1885, w_004_1886, w_004_1887, w_004_1888, w_004_1889, w_004_1890, w_004_1891, w_004_1892, w_004_1893, w_004_1894, w_004_1895, w_004_1896, w_004_1897, w_004_1898, w_004_1899, w_004_1900, w_004_1901, w_004_1902, w_004_1903, w_004_1904, w_004_1905, w_004_1906, w_004_1907, w_004_1909, w_004_1910, w_004_1911, w_004_1912, w_004_1913, w_004_1914, w_004_1915, w_004_1916, w_004_1918, w_004_1919, w_004_1920, w_004_1922, w_004_1923, w_004_1924, w_004_1927, w_004_1928, w_004_1929, w_004_1930, w_004_1931, w_004_1932, w_004_1933, w_004_1934, w_004_1935, w_004_1936, w_004_1937, w_004_1938, w_004_1939, w_004_1940, w_004_1941, w_004_1942, w_004_1943, w_004_1944, w_004_1945, w_004_1946, w_004_1947, w_004_1948, w_004_1949, w_004_1951, w_004_1952, w_004_1953, w_004_1955, w_004_1956, w_004_1957, w_004_1958, w_004_1959, w_004_1960, w_004_1961, w_004_1962, w_004_1964, w_004_1965, w_004_1966, w_004_1967, w_004_1968, w_004_1969, w_004_1970, w_004_1971, w_004_1972, w_004_1973, w_004_1974, w_004_1975, w_004_1976, w_004_1977, w_004_1978, w_004_1979, w_004_1980, w_004_1981, w_004_1982, w_004_1983, w_004_1984, w_004_1985, w_004_1986, w_004_1987, w_004_1988, w_004_1989, w_004_1990, w_004_1992, w_004_1993, w_004_1994, w_004_1995, w_004_1996, w_004_1997, w_004_1998, w_004_1999, w_004_2000, w_004_2001, w_004_2002, w_004_2003, w_004_2004, w_004_2005, w_004_2006, w_004_2007, w_004_2008, w_004_2009, w_004_2010, w_004_2011, w_004_2012, w_004_2013, w_004_2014, w_004_2015, w_004_2016, w_004_2017, w_004_2019, w_004_2020, w_004_2021, w_004_2022, w_004_2023, w_004_2024, w_004_2025, w_004_2026, w_004_2027, w_004_2028, w_004_2029, w_004_2030, w_004_2031, w_004_2032, w_004_2033, w_004_2034, w_004_2035, w_004_2036, w_004_2037, w_004_2038, w_004_2039, w_004_2040, w_004_2041, w_004_2042, w_004_2043, w_004_2044, w_004_2046, w_004_2047, w_004_2048, w_004_2049, w_004_2050, w_004_2051, w_004_2052, w_004_2053, w_004_2054, w_004_2055, w_004_2056, w_004_2057, w_004_2058, w_004_2060, w_004_2061, w_004_2062, w_004_2063, w_004_2064, w_004_2065, w_004_2066, w_004_2067, w_004_2069, w_004_2070, w_004_2071, w_004_2072, w_004_2074, w_004_2075, w_004_2076, w_004_2077, w_004_2078, w_004_2079, w_004_2080, w_004_2081, w_004_2082, w_004_2083, w_004_2084, w_004_2085, w_004_2086, w_004_2088, w_004_2089, w_004_2090, w_004_2091, w_004_2092, w_004_2093, w_004_2094, w_004_2095, w_004_2096, w_004_2097, w_004_2098, w_004_2099, w_004_2100, w_004_2101, w_004_2102, w_004_2103, w_004_2104, w_004_2105, w_004_2106, w_004_2108, w_004_2109, w_004_2110, w_004_2111, w_004_2112, w_004_2113, w_004_2114, w_004_2115, w_004_2117, w_004_2118, w_004_2119, w_004_2120, w_004_2121, w_004_2122, w_004_2123, w_004_2124, w_004_2125, w_004_2126, w_004_2127, w_004_2128, w_004_2129, w_004_2130, w_004_2131, w_004_2132, w_004_2133, w_004_2134, w_004_2136, w_004_2138, w_004_2140, w_004_2141, w_004_2142, w_004_2143, w_004_2144, w_004_2145, w_004_2146, w_004_2147, w_004_2148, w_004_2149, w_004_2150, w_004_2151, w_004_2152, w_004_2155, w_004_2157, w_004_2159, w_004_2160, w_004_2161, w_004_2162, w_004_2163, w_004_2164, w_004_2165, w_004_2166, w_004_2168, w_004_2169, w_004_2170, w_004_2171, w_004_2172, w_004_2173, w_004_2174, w_004_2175, w_004_2176, w_004_2177, w_004_2178, w_004_2179, w_004_2180, w_004_2181, w_004_2182, w_004_2183, w_004_2184, w_004_2185, w_004_2186, w_004_2187, w_004_2188, w_004_2189, w_004_2190, w_004_2191, w_004_2192, w_004_2194, w_004_2195, w_004_2196, w_004_2197, w_004_2198, w_004_2200, w_004_2201, w_004_2202, w_004_2203, w_004_2204, w_004_2205, w_004_2206, w_004_2207, w_004_2208, w_004_2209, w_004_2210, w_004_2211, w_004_2212, w_004_2213, w_004_2214, w_004_2215, w_004_2216, w_004_2217, w_004_2218, w_004_2219, w_004_2220, w_004_2221, w_004_2222, w_004_2223, w_004_2224, w_004_2225, w_004_2226, w_004_2228, w_004_2229, w_004_2230, w_004_2231, w_004_2232, w_004_2233, w_004_2234, w_004_2235, w_004_2236, w_004_2237, w_004_2238, w_004_2239, w_004_2240, w_004_2241, w_004_2242, w_004_2243, w_004_2244, w_004_2245, w_004_2246, w_004_2247, w_004_2248, w_004_2249, w_004_2250, w_004_2251, w_004_2252, w_004_2253, w_004_2254, w_004_2255, w_004_2256, w_004_2257, w_004_2258, w_004_2259, w_004_2260, w_004_2261, w_004_2262, w_004_2263, w_004_2264, w_004_2265, w_004_2266, w_004_2267, w_004_2268, w_004_2269, w_004_2270, w_004_2271, w_004_2272, w_004_2273, w_004_2275, w_004_2276, w_004_2277, w_004_2278, w_004_2279, w_004_2280, w_004_2281, w_004_2284, w_004_2286, w_004_2288, w_004_2289, w_004_2290, w_004_2292, w_004_2293, w_004_2294, w_004_2295, w_004_2296, w_004_2297, w_004_2298, w_004_2299, w_004_2300, w_004_2302, w_004_2304, w_004_2305, w_004_2306, w_004_2307, w_004_2308, w_004_2309, w_004_2310, w_004_2311, w_004_2312, w_004_2313, w_004_2314, w_004_2315, w_004_2316, w_004_2319, w_004_2320, w_004_2321, w_004_2322, w_004_2323, w_004_2324, w_004_2325, w_004_2326, w_004_2327, w_004_2328, w_004_2329, w_004_2330, w_004_2331, w_004_2332, w_004_2333, w_004_2334, w_004_2335, w_004_2336, w_004_2337, w_004_2338, w_004_2339, w_004_2340, w_004_2341, w_004_2342, w_004_2343, w_004_2344, w_004_2345, w_004_2346, w_004_2347, w_004_2348, w_004_2349, w_004_2350, w_004_2351, w_004_2353, w_004_2354, w_004_2355, w_004_2356, w_004_2357, w_004_2358, w_004_2359, w_004_2360, w_004_2361, w_004_2362, w_004_2363, w_004_2366, w_004_2368, w_004_2369, w_004_2370, w_004_2371, w_004_2372, w_004_2374, w_004_2375, w_004_2376, w_004_2378, w_004_2379, w_004_2380, w_004_2381, w_004_2382, w_004_2383, w_004_2384, w_004_2385, w_004_2386, w_004_2387, w_004_2389, w_004_2390, w_004_2391, w_004_2392, w_004_2393, w_004_2394, w_004_2395, w_004_2396, w_004_2397, w_004_2398, w_004_2399, w_004_2400, w_004_2402, w_004_2403, w_004_2404, w_004_2405, w_004_2406, w_004_2407, w_004_2409, w_004_2410, w_004_2412, w_004_2413, w_004_2414, w_004_2415, w_004_2416, w_004_2417, w_004_2418, w_004_2420, w_004_2421, w_004_2422, w_004_2423, w_004_2424, w_004_2425, w_004_2426, w_004_2427, w_004_2428, w_004_2429, w_004_2430, w_004_2431, w_004_2432, w_004_2433, w_004_2434, w_004_2435, w_004_2436, w_004_2437, w_004_2439, w_004_2440, w_004_2441, w_004_2442, w_004_2443, w_004_2444, w_004_2445, w_004_2446, w_004_2447, w_004_2448, w_004_2452, w_004_2453, w_004_2454, w_004_2456, w_004_2457, w_004_2458, w_004_2459, w_004_2460, w_004_2461, w_004_2462, w_004_2463, w_004_2464, w_004_2465, w_004_2466, w_004_2467, w_004_2469, w_004_2470, w_004_2471, w_004_2472, w_004_2474, w_004_2475, w_004_2476, w_004_2477, w_004_2478, w_004_2479, w_004_2480, w_004_2481, w_004_2482, w_004_2483, w_004_2484, w_004_2485, w_004_2486, w_004_2487, w_004_2488, w_004_2489, w_004_2490, w_004_2492, w_004_2493, w_004_2494, w_004_2495, w_004_2496, w_004_2498, w_004_2499, w_004_2500, w_004_2501, w_004_2502, w_004_2506, w_004_2507, w_004_2508, w_004_2509, w_004_2512, w_004_2513, w_004_2514, w_004_2515, w_004_2516, w_004_2517, w_004_2518, w_004_2519, w_004_2520, w_004_2521, w_004_2522, w_004_2523, w_004_2524, w_004_2525, w_004_2526, w_004_2527, w_004_2528, w_004_2530, w_004_2531, w_004_2532, w_004_2533, w_004_2535, w_004_2536, w_004_2537, w_004_2538, w_004_2539, w_004_2540, w_004_2541, w_004_2542, w_004_2543, w_004_2544, w_004_2545, w_004_2546, w_004_2547, w_004_2548, w_004_2549, w_004_2550, w_004_2551, w_004_2553, w_004_2554, w_004_2555, w_004_2556, w_004_2557, w_004_2558, w_004_2559, w_004_2560, w_004_2562, w_004_2563, w_004_2564, w_004_2565, w_004_2566, w_004_2567, w_004_2568, w_004_2569, w_004_2571, w_004_2572, w_004_2574, w_004_2575, w_004_2576, w_004_2577, w_004_2578, w_004_2579, w_004_2580, w_004_2581, w_004_2582, w_004_2583, w_004_2584, w_004_2585, w_004_2586, w_004_2587, w_004_2588, w_004_2589, w_004_2590, w_004_2591, w_004_2593, w_004_2594, w_004_2595, w_004_2596, w_004_2597, w_004_2598, w_004_2599, w_004_2600, w_004_2601, w_004_2602, w_004_2603, w_004_2604, w_004_2605, w_004_2606, w_004_2607, w_004_2608, w_004_2609, w_004_2610, w_004_2611, w_004_2612, w_004_2613, w_004_2614, w_004_2615, w_004_2616, w_004_2617, w_004_2618, w_004_2619, w_004_2620, w_004_2621, w_004_2622, w_004_2623, w_004_2624, w_004_2625, w_004_2626, w_004_2627, w_004_2628, w_004_2629, w_004_2630, w_004_2631, w_004_2632, w_004_2633, w_004_2634, w_004_2635, w_004_2636, w_004_2637, w_004_2638, w_004_2639, w_004_2640, w_004_2641, w_004_2642, w_004_2643, w_004_2644, w_004_2645, w_004_2646, w_004_2647, w_004_2648, w_004_2649, w_004_2650, w_004_2651, w_004_2652, w_004_2653, w_004_2654, w_004_2655, w_004_2657, w_004_2658, w_004_2659, w_004_2660, w_004_2661, w_004_2662, w_004_2663, w_004_2664, w_004_2665, w_004_2666, w_004_2667, w_004_2668, w_004_2670, w_004_2671, w_004_2673, w_004_2675, w_004_2676, w_004_2677, w_004_2678, w_004_2680, w_004_2681, w_004_2682, w_004_2683, w_004_2684, w_004_2687, w_004_2688, w_004_2689, w_004_2690, w_004_2691, w_004_2692, w_004_2693, w_004_2694, w_004_2695, w_004_2697, w_004_2698, w_004_2699, w_004_2701, w_004_2702, w_004_2703, w_004_2704, w_004_2705, w_004_2706, w_004_2707, w_004_2708, w_004_2709, w_004_2711, w_004_2712, w_004_2713, w_004_2714, w_004_2715, w_004_2716, w_004_2717, w_004_2718, w_004_2719, w_004_2720, w_004_2721, w_004_2722, w_004_2723, w_004_2724, w_004_2725, w_004_2726, w_004_2727, w_004_2728, w_004_2729, w_004_2731, w_004_2732, w_004_2734, w_004_2735, w_004_2736, w_004_2737, w_004_2738, w_004_2739, w_004_2740, w_004_2741, w_004_2742, w_004_2743, w_004_2744, w_004_2745, w_004_2746, w_004_2747, w_004_2748, w_004_2750, w_004_2751, w_004_2752, w_004_2753, w_004_2754, w_004_2755, w_004_2756, w_004_2757, w_004_2758, w_004_2759, w_004_2760, w_004_2762, w_004_2763, w_004_2764, w_004_2765, w_004_2766, w_004_2767, w_004_2768, w_004_2769, w_004_2770, w_004_2771, w_004_2772, w_004_2773, w_004_2774, w_004_2775, w_004_2776, w_004_2777, w_004_2778, w_004_2779, w_004_2780, w_004_2781, w_004_2782, w_004_2783, w_004_2784, w_004_2785, w_004_2786, w_004_2787, w_004_2788, w_004_2789, w_004_2790, w_004_2792, w_004_2793, w_004_2794, w_004_2796, w_004_2797, w_004_2798, w_004_2799, w_004_2800, w_004_2801, w_004_2802, w_004_2803, w_004_2804, w_004_2805, w_004_2806, w_004_2807, w_004_2808, w_004_2809, w_004_2810, w_004_2811, w_004_2812, w_004_2813, w_004_2814, w_004_2815, w_004_2816, w_004_2817, w_004_2819, w_004_2820, w_004_2822, w_004_2823, w_004_2824, w_004_2825, w_004_2826, w_004_2827, w_004_2828, w_004_2830, w_004_2831, w_004_2832, w_004_2833, w_004_2834, w_004_2835, w_004_2836, w_004_2837, w_004_2838, w_004_2839, w_004_2840, w_004_2841, w_004_2842, w_004_2843, w_004_2844, w_004_2845, w_004_2846, w_004_2847, w_004_2848, w_004_2849, w_004_2850, w_004_2851, w_004_2852, w_004_2853, w_004_2854, w_004_2855, w_004_2856, w_004_2857, w_004_2858, w_004_2860, w_004_2863, w_004_2864, w_004_2865, w_004_2866, w_004_2867, w_004_2868, w_004_2869, w_004_2870, w_004_2871, w_004_2872, w_004_2873, w_004_2874, w_004_2875, w_004_2876, w_004_2878, w_004_2879, w_004_2880, w_004_2881, w_004_2882, w_004_2883, w_004_2884, w_004_2885, w_004_2886, w_004_2887, w_004_2888, w_004_2890, w_004_2891, w_004_2892, w_004_2893, w_004_2894, w_004_2895, w_004_2896, w_004_2897, w_004_2898, w_004_2899, w_004_2900, w_004_2901, w_004_2902, w_004_2903, w_004_2905, w_004_2906, w_004_2907, w_004_2908, w_004_2911, w_004_2912, w_004_2913, w_004_2914, w_004_2915, w_004_2916, w_004_2918, w_004_2919, w_004_2920, w_004_2922, w_004_2923, w_004_2924, w_004_2925, w_004_2926, w_004_2927, w_004_2928, w_004_2929, w_004_2930, w_004_2931, w_004_2933, w_004_2934, w_004_2935, w_004_2937, w_004_2938, w_004_2939, w_004_2940, w_004_2941, w_004_2942, w_004_2943, w_004_2944, w_004_2945, w_004_2946, w_004_2947, w_004_2948, w_004_2949, w_004_2950, w_004_2951, w_004_2952, w_004_2953, w_004_2954, w_004_2955, w_004_2956, w_004_2957, w_004_2958, w_004_2959, w_004_2960, w_004_2961, w_004_2963, w_004_2964, w_004_2965, w_004_2966, w_004_2967, w_004_2968, w_004_2969, w_004_2970, w_004_2971, w_004_2972, w_004_2973, w_004_2974, w_004_2975, w_004_2976, w_004_2977, w_004_2978, w_004_2979, w_004_2980, w_004_2981, w_004_2982, w_004_2983, w_004_2984, w_004_2985, w_004_2986, w_004_2987, w_004_2988, w_004_2989, w_004_2990, w_004_2991, w_004_2993, w_004_2994, w_004_2995, w_004_2996, w_004_2997, w_004_2998, w_004_2999, w_004_3000, w_004_3001, w_004_3002, w_004_3003, w_004_3004, w_004_3005, w_004_3006, w_004_3007, w_004_3008, w_004_3009, w_004_3010, w_004_3011, w_004_3012, w_004_3013, w_004_3014, w_004_3015, w_004_3016, w_004_3017, w_004_3018, w_004_3019, w_004_3020, w_004_3021, w_004_3022, w_004_3023, w_004_3024, w_004_3025, w_004_3026, w_004_3027, w_004_3028, w_004_3029, w_004_3030, w_004_3031, w_004_3032, w_004_3033, w_004_3034, w_004_3035, w_004_3036, w_004_3037, w_004_3038, w_004_3039, w_004_3040, w_004_3041, w_004_3042, w_004_3043, w_004_3044, w_004_3045, w_004_3046, w_004_3047, w_004_3048, w_004_3049, w_004_3050, w_004_3051, w_004_3052, w_004_3054, w_004_3055, w_004_3057, w_004_3058, w_004_3059, w_004_3060, w_004_3061, w_004_3062, w_004_3063, w_004_3064, w_004_3065, w_004_3066, w_004_3068, w_004_3069, w_004_3071, w_004_3072, w_004_3073, w_004_3074, w_004_3075, w_004_3076, w_004_3077, w_004_3078, w_004_3079, w_004_3080, w_004_3081, w_004_3082, w_004_3083, w_004_3084, w_004_3085, w_004_3086, w_004_3087, w_004_3088, w_004_3089, w_004_3090, w_004_3091, w_004_3092, w_004_3093, w_004_3094, w_004_3095, w_004_3096, w_004_3097, w_004_3098, w_004_3099, w_004_3100, w_004_3101, w_004_3102, w_004_3103, w_004_3104, w_004_3105, w_004_3106, w_004_3108, w_004_3109, w_004_3111, w_004_3112, w_004_3113, w_004_3114, w_004_3115, w_004_3116, w_004_3117, w_004_3118, w_004_3119, w_004_3120, w_004_3121, w_004_3122, w_004_3124, w_004_3126, w_004_3127, w_004_3128, w_004_3129, w_004_3132, w_004_3133, w_004_3135, w_004_3136, w_004_3137, w_004_3138, w_004_3139, w_004_3140, w_004_3141, w_004_3142, w_004_3144, w_004_3145, w_004_3146, w_004_3147, w_004_3148, w_004_3149, w_004_3150, w_004_3151, w_004_3153, w_004_3154, w_004_3155, w_004_3156, w_004_3157, w_004_3158, w_004_3159, w_004_3160, w_004_3161, w_004_3162, w_004_3163, w_004_3164, w_004_3166, w_004_3167, w_004_3168, w_004_3169, w_004_3171, w_004_3172, w_004_3174, w_004_3175, w_004_3176, w_004_3177, w_004_3178, w_004_3179, w_004_3180, w_004_3181, w_004_3182, w_004_3183, w_004_3184, w_004_3185, w_004_3186, w_004_3187, w_004_3188, w_004_3189, w_004_3190, w_004_3192, w_004_3193, w_004_3194, w_004_3195, w_004_3197, w_004_3198, w_004_3199, w_004_3200, w_004_3201, w_004_3202, w_004_3203, w_004_3205, w_004_3206, w_004_3207, w_004_3209, w_004_3211, w_004_3212, w_004_3214, w_004_3215, w_004_3216, w_004_3218, w_004_3219, w_004_3220, w_004_3222, w_004_3223, w_004_3224, w_004_3225, w_004_3226, w_004_3228, w_004_3230, w_004_3231, w_004_3232, w_004_3233, w_004_3234, w_004_3235, w_004_3236, w_004_3237, w_004_3238, w_004_3239, w_004_3240, w_004_3241, w_004_3242, w_004_3243, w_004_3244, w_004_3245, w_004_3246, w_004_3247, w_004_3248, w_004_3251, w_004_3252, w_004_3254, w_004_3255, w_004_3257, w_004_3258, w_004_3260, w_004_3262, w_004_3263, w_004_3264, w_004_3265, w_004_3266, w_004_3267, w_004_3268, w_004_3269, w_004_3271, w_004_3272, w_004_3273, w_004_3274, w_004_3275, w_004_3276, w_004_3278, w_004_3279, w_004_3280, w_004_3281, w_004_3282, w_004_3283, w_004_3284, w_004_3285, w_004_3286, w_004_3287, w_004_3288, w_004_3289, w_004_3290, w_004_3291, w_004_3292, w_004_3293, w_004_3294, w_004_3295, w_004_3296, w_004_3298, w_004_3299, w_004_3300, w_004_3301, w_004_3302, w_004_3303, w_004_3304, w_004_3305, w_004_3306, w_004_3307, w_004_3308, w_004_3309, w_004_3310, w_004_3311, w_004_3312, w_004_3313, w_004_3314, w_004_3315, w_004_3316, w_004_3318, w_004_3319, w_004_3320, w_004_3321, w_004_3322, w_004_3323, w_004_3324, w_004_3325, w_004_3327, w_004_3328, w_004_3329, w_004_3330, w_004_3331, w_004_3332, w_004_3333, w_004_3334, w_004_3335, w_004_3336, w_004_3337, w_004_3338, w_004_3339, w_004_3340, w_004_3341, w_004_3342, w_004_3343, w_004_3344, w_004_3345, w_004_3346, w_004_3347, w_004_3348, w_004_3349, w_004_3350, w_004_3351, w_004_3353, w_004_3354, w_004_3355, w_004_3356, w_004_3357, w_004_3358, w_004_3359, w_004_3360, w_004_3361, w_004_3362, w_004_3363, w_004_3364, w_004_3365, w_004_3366, w_004_3367, w_004_3368, w_004_3369, w_004_3370, w_004_3371, w_004_3372, w_004_3373, w_004_3374, w_004_3375, w_004_3376, w_004_3377, w_004_3378, w_004_3379, w_004_3380, w_004_3381, w_004_3382, w_004_3383, w_004_3384, w_004_3385, w_004_3386, w_004_3387, w_004_3388, w_004_3389, w_004_3390, w_004_3391, w_004_3393, w_004_3394, w_004_3395, w_004_3396, w_004_3397, w_004_3398, w_004_3400, w_004_3401, w_004_3402, w_004_3403, w_004_3404, w_004_3405, w_004_3406, w_004_3407, w_004_3408, w_004_3409, w_004_3410, w_004_3411, w_004_3412, w_004_3413, w_004_3414, w_004_3415, w_004_3416, w_004_3418, w_004_3419, w_004_3420, w_004_3422, w_004_3423, w_004_3424, w_004_3425, w_004_3426, w_004_3427, w_004_3428, w_004_3429, w_004_3430, w_004_3431, w_004_3432, w_004_3433, w_004_3434, w_004_3435, w_004_3436, w_004_3437, w_004_3438, w_004_3439, w_004_3440, w_004_3441, w_004_3442, w_004_3443, w_004_3445, w_004_3446, w_004_3447, w_004_3448, w_004_3449, w_004_3451, w_004_3452, w_004_3453, w_004_3454, w_004_3455, w_004_3456, w_004_3457, w_004_3458, w_004_3459, w_004_3460, w_004_3461, w_004_3463, w_004_3464, w_004_3465, w_004_3467, w_004_3468, w_004_3469, w_004_3470, w_004_3471, w_004_3472, w_004_3473, w_004_3474, w_004_3476, w_004_3477, w_004_3478, w_004_3479, w_004_3480, w_004_3481, w_004_3482, w_004_3483, w_004_3484, w_004_3485, w_004_3486, w_004_3487, w_004_3488, w_004_3489, w_004_3490, w_004_3491, w_004_3492, w_004_3493, w_004_3494, w_004_3495, w_004_3497, w_004_3498, w_004_3499, w_004_3500, w_004_3501, w_004_3502, w_004_3503, w_004_3504, w_004_3505, w_004_3506, w_004_3507, w_004_3508, w_004_3509, w_004_3510, w_004_3511, w_004_3512, w_004_3514, w_004_3515, w_004_3517, w_004_3518, w_004_3519, w_004_3520, w_004_3521, w_004_3522, w_004_3523, w_004_3524, w_004_3525, w_004_3526, w_004_3527, w_004_3528, w_004_3529, w_004_3530, w_004_3531, w_004_3532, w_004_3533, w_004_3534, w_004_3536, w_004_3537, w_004_3539, w_004_3540, w_004_3541, w_004_3542, w_004_3543, w_004_3544, w_004_3546, w_004_3547, w_004_3548, w_004_3549, w_004_3550, w_004_3551, w_004_3552, w_004_3553, w_004_3554, w_004_3556, w_004_3557, w_004_3558, w_004_3559, w_004_3560, w_004_3561, w_004_3562, w_004_3563, w_004_3564, w_004_3565, w_004_3566, w_004_3567, w_004_3568, w_004_3569, w_004_3570, w_004_3573, w_004_3574, w_004_3575, w_004_3576, w_004_3577, w_004_3578, w_004_3581, w_004_3582, w_004_3583, w_004_3584, w_004_3586, w_004_3587, w_004_3588, w_004_3589, w_004_3590, w_004_3591, w_004_3592, w_004_3593, w_004_3594, w_004_3595, w_004_3596, w_004_3597, w_004_3598, w_004_3599, w_004_3600, w_004_3601, w_004_3602, w_004_3603, w_004_3604, w_004_3605, w_004_3606, w_004_3607, w_004_3608, w_004_3609, w_004_3611, w_004_3612, w_004_3613, w_004_3615, w_004_3616, w_004_3617, w_004_3618, w_004_3619, w_004_3620, w_004_3621, w_004_3622, w_004_3623, w_004_3624, w_004_3625, w_004_3626, w_004_3627, w_004_3628, w_004_3629, w_004_3630, w_004_3631, w_004_3632, w_004_3633, w_004_3634, w_004_3635, w_004_3636, w_004_3637, w_004_3638, w_004_3639, w_004_3640, w_004_3641, w_004_3642, w_004_3643, w_004_3644, w_004_3645, w_004_3647, w_004_3648, w_004_3649, w_004_3650, w_004_3651, w_004_3652, w_004_3653, w_004_3654, w_004_3655, w_004_3657, w_004_3658, w_004_3659, w_004_3660, w_004_3661, w_004_3662, w_004_3663, w_004_3664, w_004_3665, w_004_3666, w_004_3667, w_004_3668, w_004_3669, w_004_3670, w_004_3672, w_004_3673, w_004_3674, w_004_3676, w_004_3677, w_004_3678, w_004_3679, w_004_3680, w_004_3682, w_004_3683, w_004_3684, w_004_3685, w_004_3686, w_004_3687, w_004_3689, w_004_3690, w_004_3691, w_004_3692, w_004_3693, w_004_3696, w_004_3697, w_004_3698, w_004_3700, w_004_3701, w_004_3702, w_004_3703, w_004_3704, w_004_3705, w_004_3706, w_004_3707, w_004_3708, w_004_3709, w_004_3710, w_004_3711, w_004_3712, w_004_3713, w_004_3715, w_004_3716, w_004_3717, w_004_3718, w_004_3719, w_004_3720, w_004_3721, w_004_3722, w_004_3723, w_004_3724, w_004_3725, w_004_3727, w_004_3728, w_004_3729, w_004_3730, w_004_3731, w_004_3734, w_004_3735, w_004_3736, w_004_3737, w_004_3738, w_004_3739, w_004_3741, w_004_3742, w_004_3743, w_004_3744, w_004_3745, w_004_3746, w_004_3747, w_004_3748, w_004_3749, w_004_3750, w_004_3751, w_004_3752, w_004_3753, w_004_3754, w_004_3755, w_004_3756, w_004_3757, w_004_3758, w_004_3759, w_004_3760, w_004_3761, w_004_3762, w_004_3763, w_004_3764, w_004_3765, w_004_3766, w_004_3767, w_004_3768, w_004_3769, w_004_3770, w_004_3771, w_004_3772, w_004_3773, w_004_3774, w_004_3775, w_004_3777, w_004_3778, w_004_3779, w_004_3780, w_004_3781, w_004_3783, w_004_3784, w_004_3785, w_004_3786, w_004_3787, w_004_3788, w_004_3789, w_004_3790, w_004_3791, w_004_3792, w_004_3793, w_004_3794, w_004_3795, w_004_3796, w_004_3797, w_004_3798, w_004_3799, w_004_3800, w_004_3801, w_004_3802, w_004_3803, w_004_3804, w_004_3805, w_004_3806, w_004_3807, w_004_3808, w_004_3809, w_004_3810, w_004_3811, w_004_3813, w_004_3814, w_004_3815, w_004_3816, w_004_3817, w_004_3818, w_004_3819, w_004_3820, w_004_3822, w_004_3823, w_004_3824, w_004_3825, w_004_3826, w_004_3827, w_004_3828, w_004_3829, w_004_3830, w_004_3831, w_004_3832, w_004_3833, w_004_3834, w_004_3835, w_004_3836, w_004_3837, w_004_3838, w_004_3839, w_004_3840, w_004_3841, w_004_3842, w_004_3843, w_004_3844, w_004_3845, w_004_3846, w_004_3847, w_004_3848, w_004_3849, w_004_3850, w_004_3851, w_004_3853, w_004_3854, w_004_3855, w_004_3856, w_004_3857, w_004_3858, w_004_3859, w_004_3860, w_004_3861, w_004_3862, w_004_3863, w_004_3864, w_004_3866, w_004_3867, w_004_3868, w_004_3869, w_004_3870, w_004_3871, w_004_3872, w_004_3874, w_004_3875, w_004_3876, w_004_3877, w_004_3878, w_004_3879, w_004_3880, w_004_3881, w_004_3882, w_004_3883, w_004_3884, w_004_3885, w_004_3886, w_004_3887, w_004_3888, w_004_3889, w_004_3891, w_004_3892, w_004_3894, w_004_3895, w_004_3896, w_004_3897, w_004_3898, w_004_3899, w_004_3900, w_004_3902, w_004_3903, w_004_3904, w_004_3905, w_004_3906, w_004_3907, w_004_3908, w_004_3909, w_004_3910, w_004_3912, w_004_3913, w_004_3914, w_004_3915, w_004_3916, w_004_3917, w_004_3920, w_004_3921, w_004_3922, w_004_3924, w_004_3925, w_004_3927, w_004_3928, w_004_3929, w_004_3930, w_004_3931, w_004_3932, w_004_3933, w_004_3934, w_004_3935, w_004_3936, w_004_3938, w_004_3939, w_004_3941, w_004_3942, w_004_3943, w_004_3944, w_004_3945, w_004_3946, w_004_3947, w_004_3948, w_004_3949, w_004_3950, w_004_3951, w_004_3952, w_004_3953, w_004_3954, w_004_3955, w_004_3956, w_004_3957, w_004_3958, w_004_3959, w_004_3960, w_004_3961, w_004_3962, w_004_3963, w_004_3964, w_004_3965, w_004_3966, w_004_3967, w_004_3968, w_004_3969, w_004_3970, w_004_3971, w_004_3972, w_004_3973, w_004_3974, w_004_3976, w_004_3977, w_004_3978, w_004_3979, w_004_3980, w_004_3981, w_004_3982, w_004_3983, w_004_3984, w_004_3986, w_004_3987, w_004_3988, w_004_3989, w_004_3990, w_004_3991, w_004_3992, w_004_3993, w_004_3994, w_004_3995, w_004_3996, w_004_3998, w_004_3999, w_004_4000, w_004_4001, w_004_4002, w_004_4003, w_004_4004, w_004_4005, w_004_4006, w_004_4007, w_004_4010, w_004_4011, w_004_4012, w_004_4013, w_004_4014, w_004_4016, w_004_4017, w_004_4018, w_004_4019, w_004_4020, w_004_4021, w_004_4023, w_004_4024, w_004_4025, w_004_4027, w_004_4028, w_004_4029, w_004_4030, w_004_4031, w_004_4032, w_004_4033, w_004_4034, w_004_4035, w_004_4036, w_004_4037, w_004_4038, w_004_4039, w_004_4040, w_004_4041, w_004_4042, w_004_4043, w_004_4044, w_004_4045, w_004_4046, w_004_4047, w_004_4048, w_004_4049, w_004_4050, w_004_4051, w_004_4052, w_004_4053, w_004_4054, w_004_4055, w_004_4056, w_004_4058, w_004_4059, w_004_4060, w_004_4063, w_004_4064, w_004_4065, w_004_4066, w_004_4067, w_004_4068, w_004_4069, w_004_4070, w_004_4071, w_004_4072, w_004_4073, w_004_4074, w_004_4076, w_004_4077, w_004_4078, w_004_4079, w_004_4080, w_004_4081, w_004_4082, w_004_4083, w_004_4084, w_004_4085, w_004_4086, w_004_4087, w_004_4089, w_004_4090, w_004_4091, w_004_4092, w_004_4093, w_004_4094, w_004_4095, w_004_4096, w_004_4097, w_004_4098, w_004_4099, w_004_4100, w_004_4101, w_004_4102, w_004_4103, w_004_4104, w_004_4105, w_004_4106, w_004_4107, w_004_4109, w_004_4110, w_004_4111, w_004_4112, w_004_4113, w_004_4114, w_004_4115, w_004_4116, w_004_4117, w_004_4118, w_004_4119, w_004_4121, w_004_4122, w_004_4123, w_004_4124, w_004_4125, w_004_4126, w_004_4127, w_004_4128, w_004_4129, w_004_4130, w_004_4131, w_004_4132, w_004_4134, w_004_4135, w_004_4136, w_004_4137, w_004_4138, w_004_4139, w_004_4140, w_004_4141, w_004_4142, w_004_4143, w_004_4144, w_004_4145, w_004_4146, w_004_4147, w_004_4148, w_004_4149, w_004_4150, w_004_4151, w_004_4152, w_004_4153, w_004_4154, w_004_4155, w_004_4156, w_004_4157, w_004_4158, w_004_4159, w_004_4160, w_004_4161, w_004_4162, w_004_4163, w_004_4164, w_004_4165, w_004_4166, w_004_4168, w_004_4169, w_004_4170, w_004_4171, w_004_4172, w_004_4173, w_004_4174, w_004_4175, w_004_4176, w_004_4177, w_004_4180, w_004_4182, w_004_4184, w_004_4185, w_004_4186, w_004_4187, w_004_4188, w_004_4189, w_004_4190, w_004_4191, w_004_4192, w_004_4193, w_004_4194, w_004_4195, w_004_4196, w_004_4197, w_004_4198, w_004_4200, w_004_4201, w_004_4202, w_004_4203, w_004_4204, w_004_4205, w_004_4206, w_004_4207, w_004_4208, w_004_4209, w_004_4210, w_004_4211, w_004_4212, w_004_4213, w_004_4214, w_004_4215, w_004_4216, w_004_4217, w_004_4218, w_004_4219, w_004_4220, w_004_4222, w_004_4224, w_004_4225, w_004_4226, w_004_4227, w_004_4228, w_004_4229, w_004_4230, w_004_4231, w_004_4233, w_004_4234, w_004_4235, w_004_4236, w_004_4237, w_004_4238, w_004_4239, w_004_4240, w_004_4241, w_004_4243, w_004_4244, w_004_4245, w_004_4246, w_004_4247, w_004_4248, w_004_4249, w_004_4250, w_004_4251, w_004_4252, w_004_4253, w_004_4256, w_004_4257, w_004_4258, w_004_4259, w_004_4260, w_004_4261, w_004_4262, w_004_4263, w_004_4264, w_004_4265, w_004_4266, w_004_4267, w_004_4268, w_004_4269, w_004_4270, w_004_4271, w_004_4272, w_004_4273, w_004_4275, w_004_4276, w_004_4277, w_004_4278, w_004_4279, w_004_4280, w_004_4281, w_004_4282, w_004_4283, w_004_4284, w_004_4285, w_004_4286, w_004_4288, w_004_4289, w_004_4290, w_004_4291, w_004_4292, w_004_4293, w_004_4294, w_004_4295, w_004_4296, w_004_4298, w_004_4299, w_004_4300, w_004_4301, w_004_4302, w_004_4303, w_004_4304, w_004_4305, w_004_4306, w_004_4307, w_004_4308, w_004_4310, w_004_4312, w_004_4313, w_004_4314, w_004_4315, w_004_4316, w_004_4317, w_004_4318, w_004_4319, w_004_4320, w_004_4321, w_004_4322, w_004_4323, w_004_4324, w_004_4325, w_004_4326, w_004_4327, w_004_4328, w_004_4329, w_004_4330, w_004_4331, w_004_4332, w_004_4333, w_004_4334, w_004_4335, w_004_4336, w_004_4338, w_004_4339, w_004_4340, w_004_4342, w_004_4343, w_004_4344, w_004_4345, w_004_4346, w_004_4347, w_004_4348, w_004_4349, w_004_4350, w_004_4351, w_004_4352, w_004_4353, w_004_4354, w_004_4355, w_004_4356, w_004_4357, w_004_4359, w_004_4360, w_004_4361, w_004_4362, w_004_4363, w_004_4364, w_004_4365, w_004_4366, w_004_4367, w_004_4368, w_004_4369, w_004_4370, w_004_4371, w_004_4372, w_004_4373, w_004_4374, w_004_4375, w_004_4376, w_004_4377, w_004_4378, w_004_4380, w_004_4381, w_004_4382, w_004_4383, w_004_4384, w_004_4385, w_004_4386, w_004_4387, w_004_4388, w_004_4390, w_004_4391, w_004_4392, w_004_4393, w_004_4394, w_004_4396, w_004_4397, w_004_4398, w_004_4399, w_004_4400, w_004_4401, w_004_4402, w_004_4403, w_004_4404, w_004_4405, w_004_4406, w_004_4407, w_004_4409, w_004_4410, w_004_4411, w_004_4412, w_004_4413, w_004_4414, w_004_4415, w_004_4416, w_004_4417, w_004_4418, w_004_4420, w_004_4421, w_004_4422, w_004_4423, w_004_4424, w_004_4425, w_004_4427, w_004_4428, w_004_4429, w_004_4430, w_004_4431, w_004_4432, w_004_4433, w_004_4434, w_004_4435, w_004_4436, w_004_4437, w_004_4438, w_004_4439, w_004_4441, w_004_4442, w_004_4443, w_004_4444, w_004_4445, w_004_4446, w_004_4447, w_004_4448, w_004_4449, w_004_4450, w_004_4451, w_004_4452, w_004_4453, w_004_4454, w_004_4457, w_004_4459, w_004_4460, w_004_4461, w_004_4462, w_004_4463, w_004_4464, w_004_4465, w_004_4466, w_004_4467, w_004_4468, w_004_4469, w_004_4471, w_004_4472, w_004_4473, w_004_4474, w_004_4475, w_004_4476, w_004_4478, w_004_4479, w_004_4480, w_004_4481, w_004_4482, w_004_4483, w_004_4484, w_004_4485, w_004_4486, w_004_4487, w_004_4488, w_004_4489, w_004_4490, w_004_4491, w_004_4492, w_004_4494, w_004_4495, w_004_4496, w_004_4497, w_004_4500, w_004_4501, w_004_4502, w_004_4503, w_004_4504, w_004_4505, w_004_4506, w_004_4507, w_004_4508, w_004_4509, w_004_4510, w_004_4511, w_004_4512, w_004_4513, w_004_4514, w_004_4515, w_004_4516, w_004_4517, w_004_4518, w_004_4520, w_004_4521, w_004_4522, w_004_4523, w_004_4524, w_004_4525, w_004_4526, w_004_4527, w_004_4528, w_004_4529, w_004_4530, w_004_4531, w_004_4532, w_004_4533, w_004_4534, w_004_4535, w_004_4537, w_004_4538, w_004_4539, w_004_4540, w_004_4541, w_004_4542, w_004_4543, w_004_4544, w_004_4545, w_004_4546, w_004_4547, w_004_4548, w_004_4549, w_004_4550, w_004_4551, w_004_4552, w_004_4553, w_004_4554, w_004_4555, w_004_4556, w_004_4557, w_004_4558, w_004_4559, w_004_4560, w_004_4561, w_004_4562, w_004_4563, w_004_4564, w_004_4565, w_004_4566, w_004_4568, w_004_4569, w_004_4570, w_004_4571, w_004_4572, w_004_4573, w_004_4574, w_004_4575, w_004_4576, w_004_4577, w_004_4578, w_004_4579, w_004_4581, w_004_4582, w_004_4583, w_004_4586, w_004_4587, w_004_4590, w_004_4591, w_004_4593, w_004_4594, w_004_4595, w_004_4596, w_004_4597, w_004_4598, w_004_4599, w_004_4600, w_004_4601, w_004_4602, w_004_4603, w_004_4604, w_004_4605, w_004_4606, w_004_4607, w_004_4608, w_004_4609, w_004_4610, w_004_4611, w_004_4612, w_004_4613, w_004_4614, w_004_4615, w_004_4616, w_004_4617, w_004_4618, w_004_4619, w_004_4621, w_004_4622, w_004_4623, w_004_4624, w_004_4625, w_004_4626, w_004_4627, w_004_4628, w_004_4629, w_004_4630, w_004_4631, w_004_4632, w_004_4633, w_004_4634, w_004_4635, w_004_4636, w_004_4637, w_004_4638, w_004_4639, w_004_4640, w_004_4641, w_004_4643, w_004_4644, w_004_4645, w_004_4646, w_004_4647, w_004_4648, w_004_4649, w_004_4650, w_004_4651, w_004_4652, w_004_4653, w_004_4655, w_004_4657, w_004_4658, w_004_4659, w_004_4660, w_004_4661, w_004_4662, w_004_4663, w_004_4664, w_004_4665, w_004_4666, w_004_4667, w_004_4668, w_004_4669, w_004_4670, w_004_4671, w_004_4672, w_004_4674, w_004_4675, w_004_4676, w_004_4677, w_004_4678, w_004_4679, w_004_4680, w_004_4681, w_004_4682, w_004_4683, w_004_4684, w_004_4685, w_004_4686, w_004_4687, w_004_4688, w_004_4689, w_004_4690, w_004_4691, w_004_4692, w_004_4693, w_004_4694, w_004_4695, w_004_4696, w_004_4698, w_004_4699, w_004_4701, w_004_4702, w_004_4703, w_004_4704, w_004_4705, w_004_4706, w_004_4708, w_004_4711, w_004_4712, w_004_4713, w_004_4714, w_004_4715, w_004_4716, w_004_4717, w_004_4718, w_004_4719, w_004_4720, w_004_4721, w_004_4722, w_004_4723, w_004_4724, w_004_4725, w_004_4727, w_004_4728, w_004_4729, w_004_4730, w_004_4731, w_004_4732, w_004_4733, w_004_4734, w_004_4735, w_004_4736, w_004_4737, w_004_4738, w_004_4739, w_004_4740, w_004_4741, w_004_4742, w_004_4743, w_004_4744, w_004_4745, w_004_4746, w_004_4748, w_004_4749, w_004_4750, w_004_4752, w_004_4753, w_004_4754, w_004_4756, w_004_4757, w_004_4758, w_004_4759, w_004_4760, w_004_4761, w_004_4762, w_004_4763, w_004_4764, w_004_4765, w_004_4766, w_004_4768, w_004_4769, w_004_4770, w_004_4771, w_004_4772, w_004_4773, w_004_4775, w_004_4776, w_004_4777, w_004_4779;
  wire w_005_000, w_005_001, w_005_002, w_005_003, w_005_004, w_005_005, w_005_006, w_005_007, w_005_008, w_005_009, w_005_010, w_005_011, w_005_012, w_005_013, w_005_014, w_005_015, w_005_016, w_005_017, w_005_018, w_005_019, w_005_020, w_005_021, w_005_022, w_005_023, w_005_024, w_005_025, w_005_026, w_005_027, w_005_028, w_005_029, w_005_030, w_005_031, w_005_032, w_005_033, w_005_034, w_005_035, w_005_036, w_005_037, w_005_038, w_005_039, w_005_040, w_005_041, w_005_042, w_005_043, w_005_044, w_005_045, w_005_046, w_005_047, w_005_048, w_005_049, w_005_050, w_005_051, w_005_052, w_005_053, w_005_054, w_005_055, w_005_056, w_005_057, w_005_058, w_005_059, w_005_060, w_005_061, w_005_062, w_005_063, w_005_064, w_005_065, w_005_066, w_005_067, w_005_068, w_005_069, w_005_070, w_005_071, w_005_072, w_005_073, w_005_074, w_005_075, w_005_076, w_005_077, w_005_078, w_005_079, w_005_080, w_005_081, w_005_082, w_005_083, w_005_084, w_005_085, w_005_086, w_005_087, w_005_088, w_005_089, w_005_090, w_005_091, w_005_092, w_005_093, w_005_094, w_005_095, w_005_096, w_005_097, w_005_098, w_005_099, w_005_100, w_005_101, w_005_102, w_005_103, w_005_104, w_005_105, w_005_106, w_005_107, w_005_108, w_005_109, w_005_110, w_005_111, w_005_112, w_005_113, w_005_114, w_005_115, w_005_116, w_005_117, w_005_118, w_005_119, w_005_120, w_005_121, w_005_122, w_005_123, w_005_124, w_005_125, w_005_126, w_005_127, w_005_128, w_005_129, w_005_130, w_005_131, w_005_132, w_005_133, w_005_134, w_005_135, w_005_136, w_005_137, w_005_138, w_005_139, w_005_140, w_005_141, w_005_142, w_005_143, w_005_144, w_005_145, w_005_146, w_005_147, w_005_148, w_005_149, w_005_150, w_005_151, w_005_152, w_005_153, w_005_154, w_005_155, w_005_156, w_005_157, w_005_158, w_005_159, w_005_160, w_005_161, w_005_162, w_005_163, w_005_164, w_005_165, w_005_166, w_005_167, w_005_168, w_005_169, w_005_170, w_005_171, w_005_172, w_005_173, w_005_174, w_005_175, w_005_176, w_005_177, w_005_178, w_005_179, w_005_180, w_005_181, w_005_182, w_005_183, w_005_184, w_005_185, w_005_186, w_005_187, w_005_188, w_005_189, w_005_190, w_005_191, w_005_192, w_005_193, w_005_194, w_005_195, w_005_196, w_005_197, w_005_198, w_005_199, w_005_200, w_005_201, w_005_202, w_005_203, w_005_204, w_005_205, w_005_206, w_005_207, w_005_208, w_005_209, w_005_210, w_005_211, w_005_212, w_005_213, w_005_214, w_005_215, w_005_216, w_005_217, w_005_218, w_005_219, w_005_220, w_005_221, w_005_222, w_005_223, w_005_224, w_005_225, w_005_226, w_005_227, w_005_228, w_005_229, w_005_230, w_005_231, w_005_232, w_005_233, w_005_234, w_005_235, w_005_236, w_005_237, w_005_238, w_005_239, w_005_240, w_005_241, w_005_242, w_005_243, w_005_244, w_005_245, w_005_246, w_005_247, w_005_248, w_005_249, w_005_250, w_005_251, w_005_252, w_005_253, w_005_254, w_005_255, w_005_256, w_005_257, w_005_258, w_005_259, w_005_260, w_005_261, w_005_262, w_005_263, w_005_264, w_005_265, w_005_266, w_005_267, w_005_268, w_005_269, w_005_270, w_005_271, w_005_272, w_005_273, w_005_274, w_005_275, w_005_276, w_005_277, w_005_278, w_005_279, w_005_280, w_005_281, w_005_282, w_005_283, w_005_284, w_005_285, w_005_286, w_005_287, w_005_288, w_005_289, w_005_290, w_005_291, w_005_292, w_005_293, w_005_294, w_005_295, w_005_296, w_005_297, w_005_298, w_005_299, w_005_300, w_005_301, w_005_302, w_005_303, w_005_304, w_005_305, w_005_306, w_005_307, w_005_308, w_005_309, w_005_310, w_005_311, w_005_312, w_005_313, w_005_314, w_005_315, w_005_316, w_005_317, w_005_318, w_005_319, w_005_320, w_005_321, w_005_322, w_005_323, w_005_324, w_005_325, w_005_326, w_005_327, w_005_328, w_005_329, w_005_330, w_005_331, w_005_332, w_005_333, w_005_334, w_005_335, w_005_336, w_005_337, w_005_338, w_005_339, w_005_340, w_005_341, w_005_342, w_005_343, w_005_344, w_005_345, w_005_346, w_005_347, w_005_348, w_005_349, w_005_350, w_005_351, w_005_352, w_005_353, w_005_354, w_005_355, w_005_356, w_005_357, w_005_358, w_005_359, w_005_360, w_005_361, w_005_362, w_005_363, w_005_364, w_005_365, w_005_366, w_005_367, w_005_368, w_005_369, w_005_370, w_005_371, w_005_372, w_005_373, w_005_374, w_005_375, w_005_376, w_005_377, w_005_378, w_005_379, w_005_380, w_005_381, w_005_382, w_005_383, w_005_384, w_005_385, w_005_386, w_005_387, w_005_388, w_005_389, w_005_390, w_005_391, w_005_392, w_005_393, w_005_394, w_005_395, w_005_396, w_005_397, w_005_398, w_005_399, w_005_400, w_005_401, w_005_402, w_005_403, w_005_404, w_005_405, w_005_406, w_005_407, w_005_408, w_005_409, w_005_410, w_005_411, w_005_412, w_005_413, w_005_414, w_005_415, w_005_416, w_005_417, w_005_418, w_005_419, w_005_420, w_005_421, w_005_422, w_005_423, w_005_424, w_005_425, w_005_426, w_005_427, w_005_428, w_005_429, w_005_430, w_005_431, w_005_432, w_005_433, w_005_434, w_005_435, w_005_436, w_005_437, w_005_438, w_005_439, w_005_440, w_005_441, w_005_442, w_005_443, w_005_444, w_005_445, w_005_446, w_005_447, w_005_448, w_005_449, w_005_450, w_005_451, w_005_452, w_005_453, w_005_454, w_005_455, w_005_456, w_005_457, w_005_458, w_005_459, w_005_460, w_005_461, w_005_462, w_005_463, w_005_464, w_005_465, w_005_466, w_005_467, w_005_468, w_005_469, w_005_470, w_005_471, w_005_472, w_005_473, w_005_474, w_005_475, w_005_476, w_005_477, w_005_478, w_005_479, w_005_480, w_005_481, w_005_482, w_005_483, w_005_484, w_005_485, w_005_486, w_005_487, w_005_488, w_005_489, w_005_490, w_005_491, w_005_492, w_005_493, w_005_494, w_005_495, w_005_496, w_005_497, w_005_498, w_005_499, w_005_500, w_005_501, w_005_502, w_005_503, w_005_504, w_005_505, w_005_506, w_005_507, w_005_508, w_005_509, w_005_510, w_005_511, w_005_512, w_005_513, w_005_514, w_005_515, w_005_516, w_005_517, w_005_518, w_005_519, w_005_520, w_005_521, w_005_522, w_005_523, w_005_524, w_005_525, w_005_526, w_005_527, w_005_528, w_005_529, w_005_530, w_005_531, w_005_532, w_005_533, w_005_534, w_005_535, w_005_536, w_005_537, w_005_538, w_005_539, w_005_540, w_005_541, w_005_542, w_005_543, w_005_544, w_005_545, w_005_546, w_005_547, w_005_548, w_005_549, w_005_550, w_005_551, w_005_552, w_005_553, w_005_554, w_005_555, w_005_556, w_005_557, w_005_558, w_005_559, w_005_560, w_005_561, w_005_562, w_005_563, w_005_564, w_005_565, w_005_566, w_005_567, w_005_568, w_005_569, w_005_570, w_005_571, w_005_572, w_005_573, w_005_574, w_005_575, w_005_576, w_005_577, w_005_578, w_005_579, w_005_580, w_005_581, w_005_582, w_005_583, w_005_584, w_005_585, w_005_586, w_005_587, w_005_588, w_005_589, w_005_590, w_005_591, w_005_592, w_005_593, w_005_594, w_005_595, w_005_596, w_005_597, w_005_598, w_005_599, w_005_600, w_005_601, w_005_602, w_005_603, w_005_604, w_005_606, w_005_607, w_005_608, w_005_609, w_005_610, w_005_611, w_005_612, w_005_613, w_005_614, w_005_615, w_005_616, w_005_617, w_005_618, w_005_619, w_005_620, w_005_621, w_005_622, w_005_623, w_005_624, w_005_625, w_005_626, w_005_627, w_005_628, w_005_629, w_005_630, w_005_631, w_005_632, w_005_633, w_005_634, w_005_635, w_005_636, w_005_637, w_005_638, w_005_639, w_005_640, w_005_641, w_005_642, w_005_643, w_005_644, w_005_645, w_005_646, w_005_647, w_005_648, w_005_649, w_005_650, w_005_651, w_005_652, w_005_653, w_005_654, w_005_655, w_005_656, w_005_657, w_005_658, w_005_659, w_005_660, w_005_661, w_005_662, w_005_663, w_005_664, w_005_665, w_005_666, w_005_667, w_005_668, w_005_669, w_005_670, w_005_671, w_005_672, w_005_673, w_005_674, w_005_675, w_005_676, w_005_677, w_005_678, w_005_679, w_005_680, w_005_681, w_005_682, w_005_683, w_005_684, w_005_685, w_005_686, w_005_687, w_005_688, w_005_689, w_005_690, w_005_691, w_005_692, w_005_693, w_005_694, w_005_695, w_005_696, w_005_697, w_005_698, w_005_699, w_005_700, w_005_701, w_005_702, w_005_703, w_005_704, w_005_705, w_005_706, w_005_707, w_005_708, w_005_709, w_005_710, w_005_711, w_005_712, w_005_713, w_005_714, w_005_715, w_005_716, w_005_717, w_005_718, w_005_719, w_005_720, w_005_721, w_005_722, w_005_723, w_005_724, w_005_725, w_005_726, w_005_727, w_005_728, w_005_729, w_005_730, w_005_731, w_005_732, w_005_733, w_005_734, w_005_735, w_005_736, w_005_737, w_005_738, w_005_739, w_005_740, w_005_741, w_005_742, w_005_743, w_005_744, w_005_745, w_005_746, w_005_747, w_005_748, w_005_749, w_005_750, w_005_751, w_005_752, w_005_753, w_005_754, w_005_755, w_005_756, w_005_757, w_005_758, w_005_759, w_005_760, w_005_761, w_005_762, w_005_763, w_005_764, w_005_765, w_005_766, w_005_767, w_005_768, w_005_769, w_005_770, w_005_771, w_005_772, w_005_773, w_005_774, w_005_775, w_005_776, w_005_777, w_005_778, w_005_779, w_005_780, w_005_781, w_005_782, w_005_783, w_005_784, w_005_785, w_005_786, w_005_787, w_005_788, w_005_789, w_005_790, w_005_791, w_005_792, w_005_793, w_005_794, w_005_795, w_005_796, w_005_797, w_005_798, w_005_799, w_005_800, w_005_801, w_005_802, w_005_803, w_005_804, w_005_805, w_005_806, w_005_807, w_005_808, w_005_809, w_005_810, w_005_811, w_005_812, w_005_813, w_005_814, w_005_815, w_005_816, w_005_817, w_005_818, w_005_819, w_005_820, w_005_821, w_005_822, w_005_823, w_005_824, w_005_825, w_005_826, w_005_827, w_005_828, w_005_829, w_005_830, w_005_831, w_005_832, w_005_833, w_005_834, w_005_835, w_005_836, w_005_837, w_005_838, w_005_839, w_005_840, w_005_841, w_005_842, w_005_843, w_005_844, w_005_845, w_005_846, w_005_847, w_005_848, w_005_849, w_005_850, w_005_851, w_005_852, w_005_853, w_005_854, w_005_855, w_005_856, w_005_857, w_005_858, w_005_859, w_005_860, w_005_861, w_005_862, w_005_863, w_005_864, w_005_865, w_005_866, w_005_867, w_005_868, w_005_869, w_005_870, w_005_871, w_005_872, w_005_873, w_005_874, w_005_875, w_005_876, w_005_877, w_005_878, w_005_879, w_005_880, w_005_881, w_005_882, w_005_883, w_005_884, w_005_885, w_005_886, w_005_887, w_005_888, w_005_889, w_005_890, w_005_891, w_005_892, w_005_893, w_005_894, w_005_895, w_005_896, w_005_897, w_005_898, w_005_899, w_005_900, w_005_901, w_005_902, w_005_903, w_005_904, w_005_905, w_005_906, w_005_907, w_005_908, w_005_909, w_005_910, w_005_911, w_005_912, w_005_913, w_005_914, w_005_915, w_005_916, w_005_917, w_005_918, w_005_919, w_005_920, w_005_921, w_005_922, w_005_923, w_005_924, w_005_925, w_005_926, w_005_927, w_005_928, w_005_929, w_005_930, w_005_931, w_005_932, w_005_933, w_005_934, w_005_935, w_005_936, w_005_937, w_005_938, w_005_939, w_005_940, w_005_941, w_005_942, w_005_943, w_005_944, w_005_945, w_005_946, w_005_947, w_005_948, w_005_949, w_005_950, w_005_951, w_005_952, w_005_953, w_005_954, w_005_955, w_005_956, w_005_957, w_005_958, w_005_959, w_005_960, w_005_961, w_005_962, w_005_963, w_005_964, w_005_965, w_005_966, w_005_967, w_005_968, w_005_969, w_005_970, w_005_971, w_005_972, w_005_973, w_005_974, w_005_975, w_005_976, w_005_977, w_005_978, w_005_979, w_005_980, w_005_981, w_005_982, w_005_983, w_005_984, w_005_985, w_005_986, w_005_987, w_005_988, w_005_989, w_005_990, w_005_991, w_005_992, w_005_993, w_005_994, w_005_995, w_005_996, w_005_997, w_005_998, w_005_999, w_005_1000, w_005_1001, w_005_1002, w_005_1003, w_005_1004, w_005_1005, w_005_1006, w_005_1007, w_005_1008, w_005_1009, w_005_1010, w_005_1011, w_005_1012, w_005_1013, w_005_1014, w_005_1015, w_005_1016, w_005_1017, w_005_1018, w_005_1019, w_005_1020, w_005_1021, w_005_1022, w_005_1023, w_005_1024, w_005_1025, w_005_1026, w_005_1027, w_005_1028, w_005_1029, w_005_1030, w_005_1031, w_005_1032, w_005_1033, w_005_1034, w_005_1035, w_005_1036, w_005_1037, w_005_1038, w_005_1039, w_005_1040, w_005_1041, w_005_1042, w_005_1044, w_005_1045, w_005_1046, w_005_1047, w_005_1048, w_005_1049, w_005_1050, w_005_1051, w_005_1053, w_005_1054, w_005_1055, w_005_1056, w_005_1057, w_005_1058, w_005_1059, w_005_1060, w_005_1061, w_005_1062, w_005_1063, w_005_1064, w_005_1065, w_005_1066, w_005_1067, w_005_1068, w_005_1069, w_005_1070, w_005_1071, w_005_1072, w_005_1073, w_005_1074, w_005_1075, w_005_1076, w_005_1077, w_005_1078, w_005_1079, w_005_1080, w_005_1081, w_005_1082, w_005_1083, w_005_1084, w_005_1085, w_005_1086, w_005_1087, w_005_1088, w_005_1089, w_005_1090, w_005_1091, w_005_1092, w_005_1093, w_005_1094, w_005_1095, w_005_1096, w_005_1097, w_005_1098, w_005_1099, w_005_1100, w_005_1101, w_005_1102, w_005_1103, w_005_1104, w_005_1105, w_005_1106, w_005_1107, w_005_1108, w_005_1109, w_005_1110, w_005_1111, w_005_1112, w_005_1113, w_005_1114, w_005_1115, w_005_1116, w_005_1117, w_005_1118, w_005_1119, w_005_1120, w_005_1121, w_005_1122, w_005_1123, w_005_1124, w_005_1125, w_005_1126, w_005_1127, w_005_1128, w_005_1129, w_005_1130, w_005_1131, w_005_1132, w_005_1133, w_005_1134, w_005_1135, w_005_1136, w_005_1137, w_005_1138, w_005_1139, w_005_1140, w_005_1141, w_005_1142, w_005_1143, w_005_1144, w_005_1145, w_005_1146, w_005_1147, w_005_1148, w_005_1149, w_005_1150, w_005_1151, w_005_1152, w_005_1153, w_005_1154, w_005_1155, w_005_1156, w_005_1157, w_005_1158, w_005_1159, w_005_1160, w_005_1161, w_005_1162, w_005_1163, w_005_1164, w_005_1165, w_005_1166, w_005_1167, w_005_1168, w_005_1169, w_005_1170, w_005_1171, w_005_1172, w_005_1173, w_005_1174, w_005_1175, w_005_1176, w_005_1177, w_005_1178, w_005_1179, w_005_1180, w_005_1181, w_005_1182, w_005_1183, w_005_1184, w_005_1185, w_005_1186, w_005_1187, w_005_1188, w_005_1189, w_005_1190, w_005_1191, w_005_1192, w_005_1193, w_005_1194, w_005_1195, w_005_1196, w_005_1197, w_005_1198, w_005_1199, w_005_1200, w_005_1201, w_005_1202, w_005_1203, w_005_1204, w_005_1205, w_005_1206, w_005_1207, w_005_1208, w_005_1209, w_005_1210, w_005_1211, w_005_1212, w_005_1213, w_005_1214, w_005_1215, w_005_1216, w_005_1217, w_005_1218, w_005_1219, w_005_1220, w_005_1221, w_005_1222, w_005_1223, w_005_1224, w_005_1225, w_005_1226, w_005_1227, w_005_1228, w_005_1229, w_005_1230, w_005_1231, w_005_1232, w_005_1233, w_005_1234, w_005_1235, w_005_1236, w_005_1237, w_005_1238, w_005_1239, w_005_1240, w_005_1241, w_005_1242, w_005_1243, w_005_1244, w_005_1245, w_005_1246, w_005_1247, w_005_1248, w_005_1249, w_005_1250, w_005_1251, w_005_1252, w_005_1253, w_005_1254, w_005_1255, w_005_1256, w_005_1257, w_005_1258, w_005_1259, w_005_1260, w_005_1261, w_005_1262, w_005_1263, w_005_1264, w_005_1265, w_005_1266, w_005_1267, w_005_1268, w_005_1269, w_005_1270, w_005_1271, w_005_1272, w_005_1273, w_005_1274, w_005_1275, w_005_1276, w_005_1277, w_005_1278, w_005_1279, w_005_1280, w_005_1281, w_005_1282, w_005_1283, w_005_1284, w_005_1285, w_005_1286, w_005_1287, w_005_1288, w_005_1289, w_005_1290, w_005_1291, w_005_1292, w_005_1293, w_005_1294, w_005_1295, w_005_1296, w_005_1297, w_005_1298, w_005_1299, w_005_1300, w_005_1301, w_005_1302, w_005_1303, w_005_1304, w_005_1305, w_005_1306, w_005_1307, w_005_1308, w_005_1309, w_005_1310, w_005_1311, w_005_1312, w_005_1313, w_005_1314, w_005_1315, w_005_1316, w_005_1317, w_005_1318, w_005_1319, w_005_1320, w_005_1321, w_005_1322, w_005_1323, w_005_1324, w_005_1325, w_005_1326, w_005_1327, w_005_1328, w_005_1329, w_005_1330, w_005_1331, w_005_1332, w_005_1333, w_005_1334, w_005_1335, w_005_1336, w_005_1337, w_005_1338, w_005_1339, w_005_1340, w_005_1341, w_005_1342, w_005_1343, w_005_1344, w_005_1345, w_005_1346, w_005_1347, w_005_1348, w_005_1349, w_005_1350, w_005_1351, w_005_1352, w_005_1353, w_005_1354, w_005_1355, w_005_1356, w_005_1357, w_005_1358, w_005_1359, w_005_1360, w_005_1361, w_005_1362, w_005_1363, w_005_1364, w_005_1365, w_005_1366, w_005_1367, w_005_1368, w_005_1369, w_005_1370, w_005_1371, w_005_1372, w_005_1373, w_005_1374, w_005_1375, w_005_1376, w_005_1377, w_005_1378, w_005_1379, w_005_1380, w_005_1381, w_005_1382, w_005_1383, w_005_1384, w_005_1385, w_005_1386, w_005_1387, w_005_1388, w_005_1389, w_005_1390, w_005_1391, w_005_1392, w_005_1393, w_005_1394, w_005_1395, w_005_1396, w_005_1397, w_005_1398, w_005_1399, w_005_1400, w_005_1401, w_005_1402, w_005_1403, w_005_1404, w_005_1405, w_005_1406, w_005_1407, w_005_1408, w_005_1409, w_005_1410, w_005_1411, w_005_1412, w_005_1413, w_005_1414, w_005_1415, w_005_1416, w_005_1417, w_005_1418, w_005_1419, w_005_1420, w_005_1421, w_005_1422, w_005_1423, w_005_1424, w_005_1425, w_005_1426, w_005_1427, w_005_1428, w_005_1429, w_005_1430, w_005_1431, w_005_1432, w_005_1433, w_005_1434, w_005_1435, w_005_1436, w_005_1437, w_005_1438, w_005_1439, w_005_1440, w_005_1441, w_005_1442, w_005_1443, w_005_1444, w_005_1445, w_005_1446, w_005_1447, w_005_1448, w_005_1449, w_005_1450, w_005_1451, w_005_1452, w_005_1453, w_005_1454, w_005_1455, w_005_1456, w_005_1457, w_005_1458, w_005_1459, w_005_1460, w_005_1461, w_005_1462, w_005_1463, w_005_1464, w_005_1465, w_005_1466, w_005_1467, w_005_1468, w_005_1469, w_005_1470, w_005_1471, w_005_1472, w_005_1473, w_005_1474, w_005_1475, w_005_1476, w_005_1477, w_005_1478, w_005_1479, w_005_1480, w_005_1481, w_005_1482, w_005_1483, w_005_1484, w_005_1485, w_005_1486, w_005_1487, w_005_1488, w_005_1489, w_005_1490, w_005_1491, w_005_1492, w_005_1493, w_005_1494, w_005_1495, w_005_1496, w_005_1497, w_005_1498, w_005_1499, w_005_1500, w_005_1501, w_005_1502, w_005_1503, w_005_1504, w_005_1505, w_005_1506, w_005_1507, w_005_1508, w_005_1509, w_005_1510, w_005_1511, w_005_1512, w_005_1513, w_005_1514, w_005_1515, w_005_1516, w_005_1517, w_005_1518, w_005_1519, w_005_1520, w_005_1521, w_005_1522, w_005_1523, w_005_1524, w_005_1525, w_005_1526, w_005_1527, w_005_1528, w_005_1529, w_005_1530, w_005_1531, w_005_1532, w_005_1533, w_005_1534, w_005_1535, w_005_1536, w_005_1537, w_005_1538, w_005_1539, w_005_1540, w_005_1541, w_005_1542, w_005_1543, w_005_1544, w_005_1545, w_005_1546, w_005_1547, w_005_1548, w_005_1549, w_005_1550, w_005_1551, w_005_1552, w_005_1553, w_005_1554, w_005_1555, w_005_1556, w_005_1557, w_005_1558, w_005_1559, w_005_1560, w_005_1561, w_005_1562, w_005_1563, w_005_1564, w_005_1565, w_005_1566, w_005_1567, w_005_1568, w_005_1569, w_005_1570, w_005_1571, w_005_1572, w_005_1573, w_005_1574, w_005_1575, w_005_1576, w_005_1577, w_005_1578, w_005_1579, w_005_1580, w_005_1581, w_005_1582, w_005_1583, w_005_1584, w_005_1585, w_005_1586, w_005_1587, w_005_1588, w_005_1589, w_005_1590, w_005_1591, w_005_1592, w_005_1593, w_005_1594, w_005_1595, w_005_1596, w_005_1597, w_005_1598, w_005_1599, w_005_1600, w_005_1601, w_005_1602, w_005_1603, w_005_1604, w_005_1605, w_005_1606, w_005_1607, w_005_1608, w_005_1609, w_005_1611, w_005_1612, w_005_1613, w_005_1614, w_005_1616, w_005_1618, w_005_1619, w_005_1620, w_005_1622;
  wire w_006_000, w_006_001, w_006_002, w_006_003, w_006_004, w_006_005, w_006_006, w_006_007, w_006_008, w_006_009, w_006_010, w_006_011, w_006_013, w_006_014, w_006_015, w_006_016, w_006_017, w_006_018, w_006_019, w_006_020, w_006_021, w_006_022, w_006_023, w_006_024, w_006_025, w_006_026, w_006_027, w_006_028, w_006_029, w_006_030, w_006_031, w_006_032, w_006_033, w_006_034, w_006_035, w_006_036, w_006_037, w_006_038, w_006_039, w_006_040, w_006_041, w_006_042, w_006_043, w_006_044, w_006_045, w_006_046, w_006_047, w_006_048, w_006_049, w_006_050, w_006_051, w_006_052, w_006_053, w_006_054, w_006_055, w_006_056, w_006_057, w_006_058, w_006_059, w_006_060, w_006_061, w_006_062, w_006_064, w_006_065, w_006_066, w_006_067, w_006_068, w_006_069, w_006_070, w_006_071, w_006_072, w_006_073, w_006_074, w_006_077, w_006_078, w_006_079, w_006_080, w_006_081, w_006_082, w_006_083, w_006_084, w_006_085, w_006_086, w_006_087, w_006_088, w_006_089, w_006_090, w_006_091, w_006_092, w_006_093, w_006_094, w_006_095, w_006_096, w_006_097, w_006_098, w_006_099, w_006_100, w_006_101, w_006_102, w_006_103, w_006_104, w_006_105, w_006_106, w_006_107, w_006_108, w_006_109, w_006_110, w_006_111, w_006_112, w_006_113, w_006_114, w_006_115, w_006_116, w_006_117, w_006_118, w_006_119, w_006_120, w_006_121, w_006_122, w_006_123, w_006_124, w_006_125, w_006_126, w_006_127, w_006_128, w_006_129, w_006_130, w_006_131, w_006_132, w_006_133, w_006_134, w_006_135, w_006_136, w_006_137, w_006_138, w_006_139, w_006_140, w_006_141, w_006_142, w_006_144, w_006_145, w_006_146, w_006_147, w_006_148, w_006_149, w_006_150, w_006_151, w_006_152, w_006_153, w_006_154, w_006_155, w_006_156, w_006_157, w_006_158, w_006_159, w_006_161, w_006_162, w_006_163, w_006_164, w_006_165, w_006_166, w_006_167, w_006_168, w_006_169, w_006_170, w_006_171, w_006_172, w_006_173, w_006_174, w_006_175, w_006_176, w_006_177, w_006_178, w_006_179, w_006_180, w_006_181, w_006_182, w_006_183, w_006_184, w_006_185, w_006_186, w_006_187, w_006_188, w_006_189, w_006_190, w_006_191, w_006_192, w_006_193, w_006_194, w_006_195, w_006_196, w_006_197, w_006_198, w_006_199, w_006_200, w_006_201, w_006_202, w_006_203, w_006_204, w_006_205, w_006_206, w_006_207, w_006_208, w_006_209, w_006_210, w_006_211, w_006_212, w_006_213, w_006_214, w_006_215, w_006_216, w_006_217, w_006_218, w_006_219, w_006_220, w_006_221, w_006_222, w_006_223, w_006_224, w_006_225, w_006_226, w_006_227, w_006_228, w_006_229, w_006_230, w_006_231, w_006_232, w_006_233, w_006_234, w_006_235, w_006_236, w_006_237, w_006_238, w_006_239, w_006_240, w_006_241, w_006_242, w_006_243, w_006_244, w_006_245, w_006_246, w_006_247, w_006_248, w_006_249, w_006_250, w_006_251, w_006_252, w_006_253, w_006_254, w_006_255, w_006_257, w_006_258, w_006_259, w_006_260, w_006_261, w_006_262, w_006_263, w_006_264, w_006_265, w_006_266, w_006_267, w_006_268, w_006_269, w_006_270, w_006_271, w_006_272, w_006_273, w_006_274, w_006_275, w_006_276, w_006_277, w_006_278, w_006_279, w_006_280, w_006_281, w_006_282, w_006_283, w_006_284, w_006_285, w_006_286, w_006_288, w_006_289, w_006_290, w_006_291, w_006_292, w_006_293, w_006_294, w_006_295, w_006_296, w_006_297, w_006_298, w_006_299, w_006_300, w_006_301, w_006_302, w_006_303, w_006_304, w_006_305, w_006_306, w_006_307, w_006_308, w_006_309, w_006_310, w_006_311, w_006_312, w_006_313, w_006_314, w_006_315, w_006_316, w_006_317, w_006_318, w_006_319, w_006_320, w_006_321, w_006_322, w_006_323, w_006_324, w_006_325, w_006_326, w_006_327, w_006_328, w_006_329, w_006_330, w_006_331, w_006_332, w_006_333, w_006_334, w_006_335, w_006_336, w_006_337, w_006_338, w_006_339, w_006_340, w_006_341, w_006_342, w_006_343, w_006_344, w_006_345, w_006_346, w_006_347, w_006_348, w_006_349, w_006_350, w_006_351, w_006_352, w_006_353, w_006_354, w_006_355, w_006_356, w_006_357, w_006_358, w_006_359, w_006_360, w_006_361, w_006_362, w_006_363, w_006_364, w_006_365, w_006_366, w_006_367, w_006_368, w_006_369, w_006_370, w_006_371, w_006_372, w_006_373, w_006_374, w_006_375, w_006_376, w_006_377, w_006_378, w_006_379, w_006_380, w_006_381, w_006_382, w_006_384, w_006_385, w_006_386, w_006_387, w_006_388, w_006_389, w_006_390, w_006_391, w_006_392, w_006_393, w_006_394, w_006_395, w_006_396, w_006_397, w_006_398, w_006_399, w_006_400, w_006_401, w_006_402, w_006_403, w_006_404, w_006_405, w_006_406, w_006_407, w_006_408, w_006_409, w_006_410, w_006_411, w_006_412, w_006_413, w_006_414, w_006_415, w_006_416, w_006_417, w_006_418, w_006_419, w_006_420, w_006_421, w_006_422, w_006_424, w_006_425, w_006_426, w_006_427, w_006_428, w_006_429, w_006_430, w_006_431, w_006_432, w_006_433, w_006_434, w_006_435, w_006_436, w_006_437, w_006_438, w_006_439, w_006_440, w_006_441, w_006_442, w_006_443, w_006_444, w_006_445, w_006_446, w_006_447, w_006_448, w_006_449, w_006_450, w_006_451, w_006_452, w_006_453, w_006_454, w_006_455, w_006_456, w_006_457, w_006_458, w_006_459, w_006_460, w_006_461, w_006_462, w_006_463, w_006_464, w_006_465, w_006_466, w_006_467, w_006_468, w_006_469, w_006_470, w_006_471, w_006_472, w_006_473, w_006_474, w_006_475, w_006_476, w_006_477, w_006_478, w_006_480, w_006_481, w_006_482, w_006_483, w_006_484, w_006_485, w_006_486, w_006_487, w_006_488, w_006_489, w_006_490, w_006_491, w_006_492, w_006_493, w_006_494, w_006_495, w_006_496, w_006_498, w_006_499, w_006_500, w_006_501, w_006_502, w_006_503, w_006_504, w_006_505, w_006_506, w_006_508, w_006_509, w_006_511, w_006_512, w_006_513, w_006_514, w_006_515, w_006_516, w_006_517, w_006_518, w_006_519, w_006_520, w_006_521, w_006_522, w_006_523, w_006_524, w_006_525, w_006_526, w_006_527, w_006_528, w_006_529, w_006_531, w_006_532, w_006_533, w_006_534, w_006_535, w_006_536, w_006_537, w_006_538, w_006_539, w_006_540, w_006_541, w_006_542, w_006_543, w_006_544, w_006_545, w_006_546, w_006_547, w_006_548, w_006_549, w_006_550, w_006_551, w_006_552, w_006_553, w_006_554, w_006_555, w_006_556, w_006_557, w_006_558, w_006_559, w_006_560, w_006_561, w_006_562, w_006_563, w_006_564, w_006_565, w_006_566, w_006_567, w_006_568, w_006_569, w_006_570, w_006_571, w_006_572, w_006_573, w_006_574, w_006_575, w_006_576, w_006_577, w_006_578, w_006_579, w_006_580, w_006_581, w_006_582, w_006_584, w_006_585, w_006_586, w_006_587, w_006_588, w_006_589, w_006_590, w_006_591, w_006_592, w_006_593, w_006_594, w_006_595, w_006_596, w_006_597, w_006_598, w_006_599, w_006_600, w_006_601, w_006_602, w_006_603, w_006_604, w_006_605, w_006_606, w_006_607, w_006_608, w_006_609, w_006_610, w_006_611, w_006_612, w_006_613, w_006_614, w_006_615, w_006_616, w_006_617, w_006_618, w_006_619, w_006_620, w_006_621, w_006_622, w_006_623, w_006_624, w_006_625, w_006_626, w_006_627, w_006_628, w_006_629, w_006_630, w_006_631, w_006_632, w_006_633, w_006_634, w_006_635, w_006_636, w_006_637, w_006_638, w_006_639, w_006_640, w_006_641, w_006_642, w_006_643, w_006_644, w_006_645, w_006_646, w_006_647, w_006_648, w_006_649, w_006_650, w_006_651, w_006_652, w_006_653, w_006_654, w_006_655, w_006_656, w_006_657, w_006_658, w_006_659, w_006_660, w_006_661, w_006_662, w_006_663, w_006_664, w_006_665, w_006_666, w_006_667, w_006_668, w_006_669, w_006_670, w_006_671, w_006_672, w_006_673, w_006_674, w_006_675, w_006_676, w_006_677, w_006_678, w_006_679, w_006_680, w_006_681, w_006_682, w_006_683, w_006_684, w_006_685, w_006_686, w_006_687, w_006_689, w_006_690, w_006_691, w_006_692, w_006_693, w_006_694, w_006_695, w_006_696, w_006_697, w_006_698, w_006_699, w_006_700, w_006_701, w_006_702, w_006_703, w_006_704, w_006_705, w_006_706, w_006_707, w_006_708, w_006_709, w_006_710, w_006_711, w_006_712, w_006_713, w_006_714, w_006_715, w_006_716, w_006_717, w_006_718, w_006_719, w_006_720, w_006_721, w_006_722, w_006_723, w_006_724, w_006_725, w_006_726, w_006_727, w_006_728, w_006_729, w_006_730, w_006_731, w_006_732, w_006_733, w_006_734, w_006_735, w_006_736, w_006_737, w_006_738, w_006_739, w_006_741, w_006_742, w_006_743, w_006_744, w_006_745, w_006_746, w_006_747, w_006_748, w_006_750, w_006_751, w_006_752, w_006_753, w_006_754, w_006_755, w_006_756, w_006_757, w_006_758, w_006_759, w_006_760, w_006_761, w_006_762, w_006_763, w_006_764, w_006_765, w_006_766, w_006_767, w_006_768, w_006_769, w_006_770, w_006_771, w_006_772, w_006_773, w_006_774, w_006_775, w_006_776, w_006_777, w_006_778, w_006_779, w_006_780, w_006_781, w_006_782, w_006_783, w_006_784, w_006_785, w_006_786, w_006_787, w_006_788, w_006_789, w_006_790, w_006_791, w_006_792, w_006_793, w_006_794, w_006_795, w_006_796, w_006_797, w_006_798, w_006_799, w_006_800, w_006_801, w_006_802, w_006_803, w_006_804, w_006_805, w_006_806, w_006_807, w_006_808, w_006_809, w_006_810, w_006_811, w_006_812, w_006_813, w_006_814, w_006_815, w_006_816, w_006_817, w_006_818, w_006_819, w_006_820, w_006_821, w_006_822, w_006_823, w_006_824, w_006_825, w_006_826, w_006_827, w_006_828, w_006_829, w_006_830, w_006_831, w_006_832, w_006_833, w_006_834, w_006_835, w_006_836, w_006_837, w_006_838, w_006_839, w_006_840, w_006_841, w_006_842, w_006_843, w_006_844, w_006_845, w_006_846, w_006_847, w_006_848, w_006_849, w_006_850, w_006_851, w_006_853, w_006_854, w_006_855, w_006_856, w_006_857, w_006_858, w_006_859, w_006_860, w_006_861, w_006_862, w_006_863, w_006_864, w_006_865, w_006_866, w_006_867, w_006_868, w_006_869, w_006_870, w_006_871, w_006_872, w_006_873, w_006_874, w_006_875, w_006_876, w_006_877, w_006_878, w_006_879, w_006_880, w_006_881, w_006_882, w_006_883, w_006_884, w_006_885, w_006_886, w_006_887, w_006_888, w_006_889, w_006_890, w_006_891, w_006_892, w_006_893, w_006_894, w_006_895, w_006_896, w_006_897, w_006_898, w_006_899, w_006_900, w_006_901, w_006_902, w_006_903, w_006_904, w_006_905, w_006_906, w_006_907, w_006_908, w_006_909, w_006_910, w_006_911, w_006_912, w_006_913, w_006_914, w_006_915, w_006_916, w_006_917, w_006_918, w_006_919, w_006_920, w_006_921, w_006_922, w_006_923, w_006_924, w_006_925, w_006_926, w_006_927, w_006_928, w_006_929, w_006_930, w_006_931, w_006_932, w_006_933, w_006_934, w_006_935, w_006_936, w_006_937, w_006_938, w_006_939, w_006_940, w_006_941, w_006_942, w_006_943, w_006_945, w_006_946, w_006_947, w_006_948, w_006_949, w_006_950, w_006_951, w_006_952, w_006_953, w_006_954, w_006_955, w_006_956, w_006_957, w_006_958, w_006_959, w_006_960, w_006_961, w_006_962, w_006_963, w_006_964, w_006_965, w_006_966, w_006_967, w_006_968, w_006_969, w_006_970, w_006_971, w_006_972, w_006_973, w_006_974, w_006_975, w_006_976, w_006_977, w_006_978, w_006_979, w_006_980, w_006_981, w_006_982, w_006_983, w_006_984, w_006_985, w_006_986, w_006_987, w_006_988, w_006_989, w_006_990, w_006_991, w_006_992, w_006_993, w_006_994, w_006_995, w_006_996, w_006_997, w_006_998, w_006_999, w_006_1000, w_006_1001, w_006_1002, w_006_1003, w_006_1004, w_006_1005, w_006_1006, w_006_1007, w_006_1009, w_006_1010, w_006_1011, w_006_1012, w_006_1013, w_006_1014, w_006_1015, w_006_1016, w_006_1017, w_006_1018, w_006_1019, w_006_1020, w_006_1021, w_006_1022, w_006_1023, w_006_1024, w_006_1025, w_006_1026, w_006_1027, w_006_1028, w_006_1029, w_006_1030, w_006_1031, w_006_1032, w_006_1033, w_006_1034, w_006_1035, w_006_1036, w_006_1037, w_006_1038, w_006_1039, w_006_1040, w_006_1041, w_006_1042, w_006_1043, w_006_1044, w_006_1045, w_006_1046, w_006_1047, w_006_1048, w_006_1049, w_006_1050, w_006_1051, w_006_1052, w_006_1053, w_006_1054, w_006_1055, w_006_1056, w_006_1057, w_006_1058, w_006_1059, w_006_1060, w_006_1061, w_006_1062, w_006_1063, w_006_1064, w_006_1065, w_006_1066, w_006_1067, w_006_1069, w_006_1070, w_006_1071, w_006_1072, w_006_1073, w_006_1074, w_006_1075, w_006_1076, w_006_1077, w_006_1078, w_006_1079, w_006_1080, w_006_1081, w_006_1082, w_006_1083, w_006_1084, w_006_1085, w_006_1086, w_006_1087, w_006_1088, w_006_1089, w_006_1090, w_006_1091, w_006_1092, w_006_1093, w_006_1094, w_006_1095, w_006_1096, w_006_1097, w_006_1098, w_006_1099, w_006_1100, w_006_1101, w_006_1102, w_006_1103, w_006_1104, w_006_1105, w_006_1106, w_006_1107, w_006_1108, w_006_1109, w_006_1110, w_006_1111, w_006_1112, w_006_1113, w_006_1114, w_006_1115, w_006_1116, w_006_1117, w_006_1118, w_006_1119, w_006_1120, w_006_1121, w_006_1122, w_006_1123, w_006_1124, w_006_1125, w_006_1126, w_006_1127, w_006_1128, w_006_1129, w_006_1130, w_006_1131, w_006_1132, w_006_1133, w_006_1134, w_006_1135, w_006_1136, w_006_1137, w_006_1138, w_006_1139, w_006_1140, w_006_1141, w_006_1142, w_006_1143, w_006_1144, w_006_1145, w_006_1146, w_006_1147, w_006_1148, w_006_1149, w_006_1150, w_006_1151, w_006_1152, w_006_1153, w_006_1154, w_006_1155, w_006_1156, w_006_1157, w_006_1158, w_006_1159, w_006_1160, w_006_1161, w_006_1162, w_006_1163, w_006_1164, w_006_1165, w_006_1166, w_006_1167, w_006_1168, w_006_1169, w_006_1170, w_006_1171, w_006_1172, w_006_1173, w_006_1174, w_006_1175, w_006_1176, w_006_1177, w_006_1178, w_006_1179, w_006_1180, w_006_1181, w_006_1182, w_006_1183, w_006_1184, w_006_1185, w_006_1186, w_006_1187, w_006_1188, w_006_1189, w_006_1190, w_006_1191, w_006_1192, w_006_1193, w_006_1194, w_006_1195, w_006_1196, w_006_1197, w_006_1198, w_006_1199, w_006_1200, w_006_1201, w_006_1202, w_006_1203, w_006_1204, w_006_1205, w_006_1206, w_006_1207, w_006_1208, w_006_1209, w_006_1210, w_006_1211, w_006_1212, w_006_1213, w_006_1214, w_006_1215, w_006_1216, w_006_1217, w_006_1218, w_006_1219, w_006_1220, w_006_1221, w_006_1222, w_006_1223, w_006_1224, w_006_1225, w_006_1226, w_006_1227, w_006_1228, w_006_1229, w_006_1230, w_006_1231, w_006_1232, w_006_1233, w_006_1234, w_006_1235, w_006_1236, w_006_1237, w_006_1238, w_006_1239, w_006_1240, w_006_1241, w_006_1242, w_006_1243, w_006_1244, w_006_1245, w_006_1246, w_006_1247, w_006_1248, w_006_1249, w_006_1250, w_006_1251, w_006_1252, w_006_1253, w_006_1254, w_006_1255, w_006_1256, w_006_1257, w_006_1258, w_006_1259, w_006_1260, w_006_1261, w_006_1262, w_006_1263, w_006_1264, w_006_1265, w_006_1266, w_006_1267, w_006_1268, w_006_1269, w_006_1270, w_006_1271, w_006_1272, w_006_1273, w_006_1274, w_006_1275, w_006_1276, w_006_1277, w_006_1278, w_006_1279, w_006_1280, w_006_1281, w_006_1282, w_006_1283, w_006_1284, w_006_1285, w_006_1286, w_006_1287, w_006_1288, w_006_1289, w_006_1290, w_006_1291, w_006_1292, w_006_1293, w_006_1294, w_006_1295, w_006_1296, w_006_1297, w_006_1298, w_006_1299, w_006_1300, w_006_1301, w_006_1302, w_006_1303, w_006_1304, w_006_1305, w_006_1306, w_006_1307, w_006_1308, w_006_1309, w_006_1310, w_006_1311, w_006_1312, w_006_1313, w_006_1314, w_006_1315, w_006_1316, w_006_1317, w_006_1318, w_006_1319, w_006_1320, w_006_1321, w_006_1322, w_006_1323, w_006_1324, w_006_1326, w_006_1327, w_006_1328, w_006_1329, w_006_1330, w_006_1331, w_006_1332, w_006_1333, w_006_1334, w_006_1335, w_006_1336, w_006_1337, w_006_1338, w_006_1339, w_006_1340, w_006_1341, w_006_1342, w_006_1343, w_006_1344, w_006_1345, w_006_1346, w_006_1347, w_006_1348, w_006_1349, w_006_1350, w_006_1351, w_006_1352, w_006_1353, w_006_1354, w_006_1355, w_006_1356, w_006_1357, w_006_1358, w_006_1359, w_006_1360, w_006_1361, w_006_1362, w_006_1363, w_006_1364, w_006_1365, w_006_1366, w_006_1367, w_006_1368, w_006_1369, w_006_1370, w_006_1371, w_006_1373, w_006_1374, w_006_1375, w_006_1376, w_006_1377, w_006_1378, w_006_1379, w_006_1380, w_006_1381, w_006_1382, w_006_1383, w_006_1384, w_006_1385, w_006_1386, w_006_1387, w_006_1388, w_006_1389, w_006_1390, w_006_1391, w_006_1392, w_006_1393, w_006_1394, w_006_1395, w_006_1396, w_006_1397, w_006_1398, w_006_1399, w_006_1400, w_006_1401, w_006_1402, w_006_1403, w_006_1404, w_006_1405, w_006_1406, w_006_1407, w_006_1408, w_006_1409, w_006_1410, w_006_1411, w_006_1412, w_006_1413, w_006_1414, w_006_1415, w_006_1416, w_006_1417, w_006_1418, w_006_1419, w_006_1420, w_006_1421, w_006_1422, w_006_1423, w_006_1424, w_006_1425, w_006_1426, w_006_1427, w_006_1428, w_006_1429, w_006_1430, w_006_1431, w_006_1432, w_006_1433, w_006_1434, w_006_1435, w_006_1436, w_006_1437, w_006_1438, w_006_1439, w_006_1440, w_006_1441, w_006_1442, w_006_1443, w_006_1444, w_006_1445, w_006_1446, w_006_1447, w_006_1448, w_006_1449, w_006_1450, w_006_1451, w_006_1452, w_006_1453, w_006_1454, w_006_1455, w_006_1456, w_006_1457, w_006_1458, w_006_1459, w_006_1460, w_006_1461, w_006_1462, w_006_1463, w_006_1464, w_006_1465, w_006_1467, w_006_1468, w_006_1469, w_006_1470, w_006_1471, w_006_1472, w_006_1473, w_006_1474, w_006_1475, w_006_1476, w_006_1477, w_006_1478, w_006_1479, w_006_1480, w_006_1481, w_006_1482, w_006_1483, w_006_1484, w_006_1485, w_006_1486, w_006_1487, w_006_1488, w_006_1489, w_006_1490, w_006_1491, w_006_1492, w_006_1493, w_006_1494, w_006_1495, w_006_1496, w_006_1497, w_006_1498, w_006_1499, w_006_1500, w_006_1501, w_006_1502, w_006_1503, w_006_1504, w_006_1505, w_006_1506, w_006_1507, w_006_1508, w_006_1509, w_006_1510, w_006_1511, w_006_1512, w_006_1513, w_006_1514, w_006_1515, w_006_1516, w_006_1517, w_006_1518, w_006_1519, w_006_1520, w_006_1521, w_006_1522, w_006_1523, w_006_1524, w_006_1525, w_006_1526, w_006_1527, w_006_1528, w_006_1529, w_006_1530, w_006_1531, w_006_1532, w_006_1533, w_006_1534, w_006_1535, w_006_1536, w_006_1537, w_006_1538, w_006_1539, w_006_1540, w_006_1541, w_006_1542, w_006_1543, w_006_1544, w_006_1545, w_006_1546, w_006_1547, w_006_1548, w_006_1549, w_006_1550, w_006_1551, w_006_1552, w_006_1553, w_006_1554, w_006_1555, w_006_1556, w_006_1557, w_006_1558, w_006_1559, w_006_1560, w_006_1561, w_006_1562, w_006_1564, w_006_1565, w_006_1566, w_006_1567, w_006_1568, w_006_1569, w_006_1570, w_006_1571, w_006_1572, w_006_1573, w_006_1574, w_006_1575, w_006_1576, w_006_1577, w_006_1578, w_006_1579, w_006_1580, w_006_1581, w_006_1582, w_006_1583, w_006_1584, w_006_1585, w_006_1586, w_006_1587, w_006_1588, w_006_1589, w_006_1590, w_006_1591, w_006_1592, w_006_1593, w_006_1594, w_006_1595, w_006_1596, w_006_1597, w_006_1598, w_006_1599, w_006_1600, w_006_1601, w_006_1602, w_006_1603, w_006_1604, w_006_1605, w_006_1606, w_006_1607, w_006_1608, w_006_1609, w_006_1610, w_006_1611, w_006_1612, w_006_1613, w_006_1614, w_006_1615, w_006_1616, w_006_1617, w_006_1618, w_006_1619, w_006_1620, w_006_1621, w_006_1622, w_006_1623, w_006_1624, w_006_1625, w_006_1626, w_006_1627, w_006_1628, w_006_1629, w_006_1630, w_006_1631, w_006_1632, w_006_1633, w_006_1634, w_006_1635, w_006_1636, w_006_1637, w_006_1638, w_006_1639, w_006_1640, w_006_1641, w_006_1642, w_006_1644, w_006_1645, w_006_1646, w_006_1647, w_006_1648, w_006_1649, w_006_1650, w_006_1651, w_006_1652, w_006_1653, w_006_1654, w_006_1655, w_006_1656, w_006_1657, w_006_1658, w_006_1659, w_006_1660, w_006_1661, w_006_1662, w_006_1663, w_006_1664, w_006_1665, w_006_1666, w_006_1667, w_006_1668, w_006_1669, w_006_1670, w_006_1671, w_006_1672, w_006_1673, w_006_1674, w_006_1675, w_006_1677, w_006_1678, w_006_1679, w_006_1680, w_006_1681, w_006_1682, w_006_1683, w_006_1684, w_006_1685, w_006_1686, w_006_1687, w_006_1688, w_006_1689, w_006_1690, w_006_1691, w_006_1692, w_006_1693, w_006_1694, w_006_1695, w_006_1696, w_006_1697, w_006_1698, w_006_1699, w_006_1700, w_006_1701, w_006_1702, w_006_1703, w_006_1704, w_006_1705, w_006_1706, w_006_1707, w_006_1708, w_006_1709, w_006_1710, w_006_1711, w_006_1712, w_006_1713, w_006_1714, w_006_1715, w_006_1716, w_006_1717, w_006_1718, w_006_1719, w_006_1720, w_006_1721, w_006_1722, w_006_1723, w_006_1724, w_006_1725, w_006_1726, w_006_1727, w_006_1728, w_006_1729, w_006_1730, w_006_1731, w_006_1732, w_006_1733, w_006_1734, w_006_1735, w_006_1736, w_006_1737, w_006_1738, w_006_1739, w_006_1740, w_006_1741, w_006_1742, w_006_1743, w_006_1744, w_006_1745, w_006_1746, w_006_1747, w_006_1748, w_006_1749, w_006_1750, w_006_1751, w_006_1752, w_006_1753, w_006_1754, w_006_1755, w_006_1756, w_006_1757, w_006_1758, w_006_1759, w_006_1760, w_006_1761, w_006_1762, w_006_1763, w_006_1764, w_006_1765, w_006_1766, w_006_1767, w_006_1768, w_006_1769, w_006_1770, w_006_1771, w_006_1772, w_006_1773, w_006_1774, w_006_1775, w_006_1776, w_006_1777, w_006_1778, w_006_1779, w_006_1780, w_006_1781, w_006_1782, w_006_1783, w_006_1784, w_006_1785, w_006_1786, w_006_1787, w_006_1788, w_006_1789, w_006_1790, w_006_1791, w_006_1792, w_006_1793, w_006_1794, w_006_1795, w_006_1796, w_006_1797, w_006_1798, w_006_1799, w_006_1800, w_006_1801, w_006_1802, w_006_1803, w_006_1804, w_006_1805, w_006_1806, w_006_1807, w_006_1808, w_006_1810, w_006_1811, w_006_1812, w_006_1813, w_006_1814, w_006_1815, w_006_1816, w_006_1817, w_006_1818, w_006_1819, w_006_1820, w_006_1821, w_006_1822, w_006_1823, w_006_1824, w_006_1825, w_006_1826, w_006_1827, w_006_1828, w_006_1829, w_006_1830, w_006_1831, w_006_1832, w_006_1833, w_006_1834, w_006_1835, w_006_1836, w_006_1837, w_006_1838, w_006_1839, w_006_1840, w_006_1841, w_006_1842, w_006_1843, w_006_1844, w_006_1845, w_006_1846, w_006_1847, w_006_1848, w_006_1849, w_006_1850, w_006_1851, w_006_1852, w_006_1853, w_006_1854, w_006_1855, w_006_1856, w_006_1857, w_006_1858, w_006_1859, w_006_1860, w_006_1861, w_006_1862, w_006_1863, w_006_1864, w_006_1865, w_006_1866, w_006_1867, w_006_1868, w_006_1869, w_006_1870, w_006_1871, w_006_1872, w_006_1873, w_006_1874, w_006_1875, w_006_1876, w_006_1877, w_006_1878, w_006_1879, w_006_1880, w_006_1881, w_006_1882, w_006_1883, w_006_1884, w_006_1885, w_006_1886, w_006_1887, w_006_1888, w_006_1889, w_006_1890, w_006_1891, w_006_1892, w_006_1893, w_006_1894, w_006_1895, w_006_1896, w_006_1897, w_006_1898, w_006_1899, w_006_1900, w_006_1901, w_006_1902, w_006_1903, w_006_1904, w_006_1905, w_006_1906, w_006_1907, w_006_1908, w_006_1909, w_006_1910, w_006_1911, w_006_1912, w_006_1913, w_006_1914, w_006_1915, w_006_1916, w_006_1917, w_006_1918, w_006_1919, w_006_1920, w_006_1921, w_006_1922, w_006_1923, w_006_1924, w_006_1925, w_006_1926, w_006_1927, w_006_1928, w_006_1929, w_006_1930, w_006_1931, w_006_1932, w_006_1933, w_006_1934, w_006_1935, w_006_1936, w_006_1937, w_006_1938, w_006_1939, w_006_1940, w_006_1941, w_006_1942, w_006_1943, w_006_1944, w_006_1945, w_006_1946, w_006_1947, w_006_1948, w_006_1949, w_006_1950, w_006_1951, w_006_1952, w_006_1953, w_006_1954, w_006_1955, w_006_1956, w_006_1957, w_006_1958, w_006_1959, w_006_1960, w_006_1961, w_006_1962, w_006_1963, w_006_1964, w_006_1965, w_006_1966, w_006_1967, w_006_1968, w_006_1969, w_006_1970, w_006_1971, w_006_1972, w_006_1973, w_006_1974, w_006_1975, w_006_1976, w_006_1977, w_006_1978, w_006_1979, w_006_1980, w_006_1981, w_006_1982, w_006_1983, w_006_1984, w_006_1985, w_006_1986, w_006_1987, w_006_1988, w_006_1989, w_006_1990, w_006_1991, w_006_1992, w_006_1993, w_006_1994, w_006_1995, w_006_1996, w_006_1997, w_006_1998, w_006_1999, w_006_2000, w_006_2001, w_006_2002, w_006_2003, w_006_2004, w_006_2005, w_006_2006, w_006_2007, w_006_2008, w_006_2009, w_006_2010, w_006_2011, w_006_2012, w_006_2013, w_006_2014, w_006_2015, w_006_2016, w_006_2017, w_006_2018, w_006_2019, w_006_2020, w_006_2021, w_006_2022, w_006_2023, w_006_2024, w_006_2025, w_006_2026, w_006_2027, w_006_2028, w_006_2029, w_006_2030, w_006_2031, w_006_2032, w_006_2033, w_006_2034, w_006_2035, w_006_2036, w_006_2037, w_006_2038, w_006_2039, w_006_2040, w_006_2041, w_006_2042, w_006_2043, w_006_2044, w_006_2045, w_006_2046, w_006_2047, w_006_2049, w_006_2050, w_006_2051, w_006_2052, w_006_2053, w_006_2054, w_006_2055, w_006_2056, w_006_2058, w_006_2059, w_006_2060, w_006_2061, w_006_2062, w_006_2063, w_006_2064, w_006_2065, w_006_2066, w_006_2067, w_006_2068, w_006_2069, w_006_2070, w_006_2071, w_006_2072, w_006_2073, w_006_2074, w_006_2075, w_006_2076, w_006_2077, w_006_2078, w_006_2079, w_006_2080, w_006_2081, w_006_2083, w_006_2085, w_006_2086, w_006_2087, w_006_2088, w_006_2089, w_006_2091, w_006_2092, w_006_2093, w_006_2094, w_006_2095, w_006_2096, w_006_2097, w_006_2098, w_006_2100, w_006_2101, w_006_2102, w_006_2103, w_006_2105, w_006_2106, w_006_2107, w_006_2108, w_006_2109, w_006_2111, w_006_2112, w_006_2113, w_006_2114, w_006_2115, w_006_2116, w_006_2117, w_006_2118, w_006_2119, w_006_2121, w_006_2122, w_006_2123, w_006_2124, w_006_2125, w_006_2126, w_006_2127, w_006_2128, w_006_2129, w_006_2130, w_006_2131, w_006_2132, w_006_2133, w_006_2134, w_006_2135, w_006_2138, w_006_2139, w_006_2140, w_006_2141, w_006_2142, w_006_2143, w_006_2144, w_006_2146, w_006_2147, w_006_2148, w_006_2151, w_006_2152, w_006_2153, w_006_2155, w_006_2156, w_006_2157, w_006_2158, w_006_2159, w_006_2160, w_006_2161, w_006_2162, w_006_2163, w_006_2164, w_006_2166, w_006_2167, w_006_2168, w_006_2169, w_006_2170, w_006_2171, w_006_2172, w_006_2173, w_006_2174, w_006_2175, w_006_2176, w_006_2177, w_006_2178, w_006_2179, w_006_2180, w_006_2181, w_006_2182, w_006_2183, w_006_2187, w_006_2188, w_006_2189, w_006_2190, w_006_2191, w_006_2192, w_006_2193, w_006_2194, w_006_2195, w_006_2196, w_006_2197, w_006_2198, w_006_2200, w_006_2203, w_006_2205, w_006_2206, w_006_2207, w_006_2208, w_006_2209, w_006_2210, w_006_2211, w_006_2212, w_006_2213, w_006_2215, w_006_2216, w_006_2217, w_006_2219, w_006_2221, w_006_2222, w_006_2225, w_006_2226, w_006_2227, w_006_2228, w_006_2230, w_006_2231, w_006_2232, w_006_2233, w_006_2234, w_006_2235, w_006_2237, w_006_2238, w_006_2239, w_006_2240, w_006_2241, w_006_2243, w_006_2244, w_006_2245, w_006_2246, w_006_2247, w_006_2248, w_006_2249, w_006_2251, w_006_2252, w_006_2253, w_006_2254, w_006_2256, w_006_2257, w_006_2258, w_006_2260, w_006_2261, w_006_2263, w_006_2264, w_006_2265, w_006_2266, w_006_2267, w_006_2268, w_006_2269, w_006_2270, w_006_2271, w_006_2272, w_006_2273, w_006_2274, w_006_2275, w_006_2276, w_006_2277, w_006_2278, w_006_2279, w_006_2280, w_006_2281, w_006_2282, w_006_2283, w_006_2284, w_006_2285, w_006_2286, w_006_2287, w_006_2289, w_006_2290, w_006_2291, w_006_2292, w_006_2294, w_006_2295, w_006_2296, w_006_2298, w_006_2299, w_006_2300, w_006_2301, w_006_2302, w_006_2303, w_006_2304, w_006_2305, w_006_2306, w_006_2307, w_006_2310, w_006_2311, w_006_2313, w_006_2314, w_006_2315, w_006_2316, w_006_2317, w_006_2318, w_006_2319, w_006_2320, w_006_2321, w_006_2322, w_006_2323, w_006_2324, w_006_2325, w_006_2326, w_006_2328, w_006_2330, w_006_2331, w_006_2332, w_006_2333, w_006_2334, w_006_2336, w_006_2337, w_006_2338, w_006_2339, w_006_2340, w_006_2341, w_006_2342, w_006_2343, w_006_2344, w_006_2345, w_006_2346, w_006_2347, w_006_2348, w_006_2349, w_006_2350, w_006_2351, w_006_2352, w_006_2353, w_006_2354, w_006_2355, w_006_2356, w_006_2357, w_006_2358, w_006_2359, w_006_2360, w_006_2361, w_006_2362, w_006_2363, w_006_2364, w_006_2365, w_006_2366, w_006_2367, w_006_2368, w_006_2369, w_006_2370, w_006_2371, w_006_2372, w_006_2374, w_006_2375, w_006_2376, w_006_2379, w_006_2380, w_006_2381, w_006_2383, w_006_2384, w_006_2385, w_006_2386, w_006_2387, w_006_2388, w_006_2390, w_006_2391, w_006_2392, w_006_2393, w_006_2394, w_006_2396, w_006_2397, w_006_2398, w_006_2399, w_006_2400, w_006_2401, w_006_2404, w_006_2405, w_006_2406, w_006_2407, w_006_2408, w_006_2409, w_006_2410, w_006_2411, w_006_2412, w_006_2413, w_006_2414, w_006_2415, w_006_2416, w_006_2417, w_006_2418, w_006_2419, w_006_2420, w_006_2421, w_006_2423, w_006_2424, w_006_2425, w_006_2426, w_006_2428, w_006_2429, w_006_2430, w_006_2431, w_006_2432, w_006_2433, w_006_2434, w_006_2435, w_006_2436, w_006_2437, w_006_2438, w_006_2439, w_006_2440, w_006_2441, w_006_2442, w_006_2443, w_006_2444, w_006_2445, w_006_2446, w_006_2447, w_006_2448, w_006_2449, w_006_2451, w_006_2453, w_006_2454, w_006_2455, w_006_2456, w_006_2457, w_006_2458, w_006_2460, w_006_2461, w_006_2462, w_006_2463, w_006_2464, w_006_2465, w_006_2466, w_006_2467, w_006_2468, w_006_2469, w_006_2471, w_006_2472, w_006_2473, w_006_2474, w_006_2475, w_006_2476, w_006_2477, w_006_2478, w_006_2479, w_006_2480, w_006_2481, w_006_2482, w_006_2484, w_006_2485, w_006_2486, w_006_2488, w_006_2489, w_006_2490, w_006_2491, w_006_2492, w_006_2493, w_006_2494, w_006_2495, w_006_2496, w_006_2497, w_006_2498, w_006_2499, w_006_2500, w_006_2501, w_006_2502, w_006_2503, w_006_2504, w_006_2505, w_006_2506, w_006_2507, w_006_2509, w_006_2511, w_006_2513, w_006_2514, w_006_2517, w_006_2518, w_006_2519, w_006_2520, w_006_2521, w_006_2525, w_006_2529, w_006_2530, w_006_2531, w_006_2532, w_006_2533, w_006_2535, w_006_2536, w_006_2537, w_006_2538, w_006_2539, w_006_2540, w_006_2541, w_006_2542, w_006_2543, w_006_2544, w_006_2546, w_006_2547, w_006_2548, w_006_2549, w_006_2550, w_006_2551, w_006_2552, w_006_2553, w_006_2554, w_006_2555, w_006_2556, w_006_2557, w_006_2558, w_006_2559, w_006_2561, w_006_2563, w_006_2564, w_006_2565, w_006_2566, w_006_2567, w_006_2568, w_006_2569, w_006_2570, w_006_2571, w_006_2572, w_006_2573, w_006_2574, w_006_2576, w_006_2577, w_006_2578, w_006_2579, w_006_2580, w_006_2582, w_006_2583, w_006_2584, w_006_2585, w_006_2587, w_006_2588, w_006_2589, w_006_2590, w_006_2591, w_006_2592, w_006_2593, w_006_2594, w_006_2595, w_006_2596, w_006_2597, w_006_2598, w_006_2599, w_006_2600, w_006_2601, w_006_2602, w_006_2603, w_006_2604, w_006_2606, w_006_2607, w_006_2608, w_006_2609, w_006_2610, w_006_2611, w_006_2612, w_006_2613, w_006_2614, w_006_2615, w_006_2616, w_006_2618, w_006_2619, w_006_2620, w_006_2621, w_006_2622, w_006_2623, w_006_2624, w_006_2625, w_006_2626, w_006_2627, w_006_2628, w_006_2629, w_006_2630, w_006_2631, w_006_2632, w_006_2633, w_006_2634, w_006_2635, w_006_2636, w_006_2637, w_006_2638, w_006_2640, w_006_2641, w_006_2642, w_006_2643, w_006_2645, w_006_2646, w_006_2647, w_006_2648, w_006_2649, w_006_2650, w_006_2651, w_006_2654, w_006_2656, w_006_2657, w_006_2658, w_006_2659, w_006_2660, w_006_2661, w_006_2662, w_006_2663, w_006_2664, w_006_2665, w_006_2666, w_006_2667, w_006_2669, w_006_2670, w_006_2671, w_006_2672, w_006_2673, w_006_2674, w_006_2675, w_006_2676, w_006_2677, w_006_2678, w_006_2679, w_006_2681, w_006_2682, w_006_2683, w_006_2684, w_006_2685, w_006_2686, w_006_2687, w_006_2688, w_006_2689, w_006_2690, w_006_2691, w_006_2692, w_006_2693, w_006_2695, w_006_2696, w_006_2697, w_006_2698, w_006_2699, w_006_2700, w_006_2701, w_006_2702, w_006_2703, w_006_2704, w_006_2705, w_006_2706, w_006_2707, w_006_2708, w_006_2709, w_006_2710, w_006_2711, w_006_2712, w_006_2713, w_006_2714, w_006_2715, w_006_2717, w_006_2718, w_006_2719, w_006_2720, w_006_2722, w_006_2723, w_006_2724, w_006_2725, w_006_2727, w_006_2728, w_006_2729, w_006_2730, w_006_2731, w_006_2732, w_006_2733, w_006_2735, w_006_2736, w_006_2737, w_006_2738, w_006_2740, w_006_2741, w_006_2743, w_006_2744, w_006_2745, w_006_2746, w_006_2748, w_006_2749, w_006_2750, w_006_2751, w_006_2752, w_006_2753, w_006_2754, w_006_2755, w_006_2756, w_006_2757, w_006_2758, w_006_2760, w_006_2762, w_006_2763, w_006_2764, w_006_2765, w_006_2767, w_006_2768, w_006_2769, w_006_2770, w_006_2771, w_006_2772, w_006_2773, w_006_2775, w_006_2776, w_006_2777, w_006_2778, w_006_2779, w_006_2780, w_006_2783, w_006_2785, w_006_2786, w_006_2788, w_006_2791, w_006_2792, w_006_2793, w_006_2795, w_006_2796, w_006_2797, w_006_2799, w_006_2800, w_006_2801, w_006_2802, w_006_2803, w_006_2804, w_006_2805, w_006_2807, w_006_2808, w_006_2809, w_006_2810, w_006_2812, w_006_2813, w_006_2814, w_006_2816, w_006_2817, w_006_2819, w_006_2821, w_006_2822, w_006_2823, w_006_2824, w_006_2825, w_006_2826, w_006_2827, w_006_2828, w_006_2829, w_006_2830, w_006_2832, w_006_2834, w_006_2835, w_006_2836, w_006_2837, w_006_2838, w_006_2839, w_006_2840, w_006_2841, w_006_2842, w_006_2843, w_006_2844, w_006_2846, w_006_2848, w_006_2849, w_006_2850, w_006_2851, w_006_2852, w_006_2853, w_006_2854, w_006_2855, w_006_2856, w_006_2857, w_006_2858, w_006_2859, w_006_2860, w_006_2861, w_006_2863, w_006_2864, w_006_2865, w_006_2866, w_006_2867, w_006_2868, w_006_2869, w_006_2870, w_006_2872, w_006_2873, w_006_2874, w_006_2875, w_006_2876, w_006_2877, w_006_2878, w_006_2879, w_006_2880, w_006_2882, w_006_2883, w_006_2884, w_006_2886, w_006_2887, w_006_2888, w_006_2889, w_006_2890, w_006_2891, w_006_2892, w_006_2893, w_006_2894, w_006_2896, w_006_2899, w_006_2900, w_006_2901, w_006_2902, w_006_2904, w_006_2905, w_006_2906, w_006_2907, w_006_2908, w_006_2909, w_006_2910, w_006_2911, w_006_2912, w_006_2913, w_006_2914, w_006_2915, w_006_2916, w_006_2917;
  wire w_007_000, w_007_001, w_007_002, w_007_003, w_007_004, w_007_005, w_007_006, w_007_007, w_007_008, w_007_009, w_007_010, w_007_011, w_007_012, w_007_013, w_007_014, w_007_015, w_007_016, w_007_017, w_007_018, w_007_019, w_007_020, w_007_021, w_007_022, w_007_023, w_007_024, w_007_025, w_007_026, w_007_027, w_007_028, w_007_029, w_007_030, w_007_031, w_007_032, w_007_033, w_007_034, w_007_035, w_007_036, w_007_037, w_007_038, w_007_039, w_007_040, w_007_041, w_007_042, w_007_043, w_007_044, w_007_045, w_007_046, w_007_047, w_007_048, w_007_049, w_007_050, w_007_051, w_007_052, w_007_053, w_007_054, w_007_055, w_007_056, w_007_057, w_007_058, w_007_059, w_007_060, w_007_061, w_007_062, w_007_063, w_007_064, w_007_065, w_007_066, w_007_067, w_007_068, w_007_069, w_007_070, w_007_071, w_007_072, w_007_073, w_007_074, w_007_075, w_007_076, w_007_077, w_007_078, w_007_079, w_007_080, w_007_081, w_007_082, w_007_083, w_007_084, w_007_085, w_007_086, w_007_087, w_007_088, w_007_089, w_007_090, w_007_091, w_007_092, w_007_093, w_007_094, w_007_095, w_007_096, w_007_097, w_007_098, w_007_099, w_007_100, w_007_101, w_007_102, w_007_103, w_007_104, w_007_105, w_007_106, w_007_107, w_007_108, w_007_109, w_007_110, w_007_111, w_007_112, w_007_113, w_007_114, w_007_115, w_007_116, w_007_117, w_007_118, w_007_119, w_007_120, w_007_121, w_007_122, w_007_123, w_007_124, w_007_125, w_007_126, w_007_127, w_007_128, w_007_129, w_007_130, w_007_131, w_007_132, w_007_133, w_007_134, w_007_135, w_007_136, w_007_137, w_007_138, w_007_139, w_007_140, w_007_141, w_007_142, w_007_143, w_007_144, w_007_145, w_007_146, w_007_147, w_007_148, w_007_149, w_007_150, w_007_151, w_007_152, w_007_153, w_007_154, w_007_155, w_007_156, w_007_157, w_007_158, w_007_159, w_007_160, w_007_161, w_007_162, w_007_163, w_007_164, w_007_165, w_007_166, w_007_167, w_007_168, w_007_169, w_007_170, w_007_171, w_007_172, w_007_173, w_007_174, w_007_175, w_007_176, w_007_177, w_007_178, w_007_179, w_007_180, w_007_181, w_007_182, w_007_183, w_007_184, w_007_185, w_007_186, w_007_187, w_007_188, w_007_189, w_007_190, w_007_191, w_007_192, w_007_193, w_007_194, w_007_195, w_007_196, w_007_197, w_007_198, w_007_199, w_007_200, w_007_201, w_007_202, w_007_203, w_007_204, w_007_205, w_007_206, w_007_207, w_007_208, w_007_209, w_007_210, w_007_211, w_007_212, w_007_213, w_007_214, w_007_215, w_007_216, w_007_217, w_007_218, w_007_219, w_007_220, w_007_221, w_007_222, w_007_223, w_007_224, w_007_225, w_007_226, w_007_227, w_007_228, w_007_229, w_007_230, w_007_231, w_007_232, w_007_233, w_007_234, w_007_235, w_007_236, w_007_237, w_007_238, w_007_239, w_007_240, w_007_241, w_007_242, w_007_243, w_007_244, w_007_245, w_007_246, w_007_247, w_007_248, w_007_249, w_007_250, w_007_251, w_007_252, w_007_253, w_007_254, w_007_255, w_007_256, w_007_257, w_007_258, w_007_259, w_007_260, w_007_261, w_007_262, w_007_263, w_007_264, w_007_265, w_007_266, w_007_267, w_007_268, w_007_269, w_007_270, w_007_271, w_007_272, w_007_273, w_007_274, w_007_275, w_007_276, w_007_277, w_007_278, w_007_279, w_007_280, w_007_281, w_007_282, w_007_283, w_007_284, w_007_285, w_007_286, w_007_287, w_007_288, w_007_289, w_007_290, w_007_291, w_007_292, w_007_293, w_007_294, w_007_295, w_007_296, w_007_297, w_007_298, w_007_299, w_007_300, w_007_301, w_007_302, w_007_303, w_007_304, w_007_305, w_007_306, w_007_307, w_007_308, w_007_309, w_007_310, w_007_311, w_007_312, w_007_313, w_007_314, w_007_315, w_007_316, w_007_317, w_007_318, w_007_319, w_007_320, w_007_321, w_007_322, w_007_323, w_007_324, w_007_325, w_007_326, w_007_327, w_007_328, w_007_329, w_007_330, w_007_331, w_007_332, w_007_333, w_007_334, w_007_335, w_007_336, w_007_337, w_007_338, w_007_339, w_007_340, w_007_341, w_007_342, w_007_343, w_007_344, w_007_345, w_007_346, w_007_347, w_007_348, w_007_349, w_007_350, w_007_351, w_007_352, w_007_353, w_007_354, w_007_355, w_007_356, w_007_357, w_007_358, w_007_359, w_007_360, w_007_361, w_007_362, w_007_363, w_007_364, w_007_365, w_007_366, w_007_367, w_007_368, w_007_369, w_007_370, w_007_371, w_007_372, w_007_373, w_007_374, w_007_375, w_007_376, w_007_377, w_007_378, w_007_379, w_007_380, w_007_381, w_007_382, w_007_383, w_007_384, w_007_385, w_007_386, w_007_387, w_007_388, w_007_389, w_007_390, w_007_391, w_007_392, w_007_393, w_007_394, w_007_395, w_007_396, w_007_397, w_007_398, w_007_399, w_007_400, w_007_401, w_007_402, w_007_403, w_007_404, w_007_405, w_007_406, w_007_407, w_007_408, w_007_409, w_007_410, w_007_411, w_007_412, w_007_413, w_007_414, w_007_415, w_007_416, w_007_417, w_007_418, w_007_419, w_007_420, w_007_421, w_007_422, w_007_423, w_007_424, w_007_425, w_007_426, w_007_427, w_007_428, w_007_429, w_007_430, w_007_431, w_007_432, w_007_433, w_007_434, w_007_435, w_007_436, w_007_437, w_007_438, w_007_439, w_007_440, w_007_441, w_007_442, w_007_443, w_007_444, w_007_445, w_007_446, w_007_447, w_007_448, w_007_449, w_007_450, w_007_451, w_007_452, w_007_453, w_007_454, w_007_455, w_007_456, w_007_457, w_007_458, w_007_459, w_007_460, w_007_461, w_007_462, w_007_463, w_007_464, w_007_465, w_007_466, w_007_467, w_007_468, w_007_469, w_007_470, w_007_471, w_007_472, w_007_473, w_007_474, w_007_475, w_007_476, w_007_477, w_007_478, w_007_479, w_007_480, w_007_481, w_007_482, w_007_483, w_007_484, w_007_485, w_007_486, w_007_487, w_007_488, w_007_489, w_007_490, w_007_491, w_007_492, w_007_493, w_007_494, w_007_495, w_007_496, w_007_497, w_007_498, w_007_499, w_007_500, w_007_501, w_007_502, w_007_503, w_007_504, w_007_505, w_007_506, w_007_507, w_007_508, w_007_509, w_007_510, w_007_511, w_007_512, w_007_513, w_007_514, w_007_515, w_007_516, w_007_517, w_007_518, w_007_519, w_007_520, w_007_521, w_007_522, w_007_523, w_007_524, w_007_525, w_007_526, w_007_527, w_007_528, w_007_529, w_007_530, w_007_531, w_007_532, w_007_533, w_007_534, w_007_535, w_007_536, w_007_537, w_007_538, w_007_539, w_007_540, w_007_541, w_007_542, w_007_543, w_007_544, w_007_545, w_007_546, w_007_547, w_007_548, w_007_549, w_007_550, w_007_551, w_007_552, w_007_553, w_007_554, w_007_555, w_007_556, w_007_557, w_007_558, w_007_559, w_007_560, w_007_561, w_007_562, w_007_563, w_007_564, w_007_565, w_007_566, w_007_567, w_007_568, w_007_569, w_007_570, w_007_571, w_007_572, w_007_573, w_007_574, w_007_575, w_007_576, w_007_577, w_007_578, w_007_579, w_007_580, w_007_581, w_007_582, w_007_583, w_007_584, w_007_585, w_007_586, w_007_587, w_007_588, w_007_589, w_007_590, w_007_591, w_007_592, w_007_593, w_007_594, w_007_595, w_007_596, w_007_597, w_007_598, w_007_599, w_007_600, w_007_601, w_007_602, w_007_603, w_007_604, w_007_605, w_007_606, w_007_607, w_007_608, w_007_609, w_007_610, w_007_611, w_007_612, w_007_613, w_007_614, w_007_615, w_007_616, w_007_617, w_007_618, w_007_619, w_007_620, w_007_621, w_007_622, w_007_623, w_007_624, w_007_625, w_007_626, w_007_627, w_007_628, w_007_629, w_007_630, w_007_631, w_007_632, w_007_633, w_007_634, w_007_635, w_007_636, w_007_637, w_007_638, w_007_639, w_007_640, w_007_641, w_007_642, w_007_643, w_007_644, w_007_645, w_007_646, w_007_647, w_007_648, w_007_649, w_007_650, w_007_651, w_007_652, w_007_653, w_007_654, w_007_655, w_007_656, w_007_657, w_007_658, w_007_659, w_007_660, w_007_661, w_007_662, w_007_663, w_007_664, w_007_665, w_007_666, w_007_667, w_007_668, w_007_669, w_007_670, w_007_671, w_007_672, w_007_673, w_007_674, w_007_675, w_007_676, w_007_677, w_007_678, w_007_679, w_007_680, w_007_681, w_007_682, w_007_683, w_007_684, w_007_685, w_007_686, w_007_687, w_007_688, w_007_689, w_007_691, w_007_692, w_007_693, w_007_694, w_007_695, w_007_696, w_007_698;
  wire w_008_000, w_008_001, w_008_002, w_008_003, w_008_004, w_008_005, w_008_006, w_008_007, w_008_008, w_008_009, w_008_010, w_008_011, w_008_012, w_008_013, w_008_014, w_008_015, w_008_016, w_008_017, w_008_018, w_008_019, w_008_020, w_008_021, w_008_022, w_008_023, w_008_024, w_008_025, w_008_026, w_008_027, w_008_028, w_008_029, w_008_030, w_008_031, w_008_032, w_008_033, w_008_034, w_008_035, w_008_036, w_008_037, w_008_038, w_008_039, w_008_040, w_008_041, w_008_042, w_008_043, w_008_044, w_008_045, w_008_046, w_008_047, w_008_048, w_008_049, w_008_050, w_008_051, w_008_052, w_008_053, w_008_054, w_008_055, w_008_057, w_008_058, w_008_059, w_008_060, w_008_061, w_008_063, w_008_064, w_008_065, w_008_066, w_008_067, w_008_068, w_008_069, w_008_070, w_008_071, w_008_072, w_008_073, w_008_074, w_008_075, w_008_076, w_008_077, w_008_078, w_008_080, w_008_081, w_008_082, w_008_083, w_008_084, w_008_085, w_008_086, w_008_087, w_008_088, w_008_089, w_008_090, w_008_091, w_008_092, w_008_093, w_008_094, w_008_095, w_008_096, w_008_097, w_008_098, w_008_099, w_008_100, w_008_101, w_008_102, w_008_103, w_008_104, w_008_105, w_008_106, w_008_107, w_008_108, w_008_109, w_008_110, w_008_111, w_008_112, w_008_113, w_008_114, w_008_115, w_008_116, w_008_117, w_008_118, w_008_119, w_008_120, w_008_121, w_008_122, w_008_123, w_008_124, w_008_125, w_008_126, w_008_129, w_008_130, w_008_131, w_008_132, w_008_133, w_008_134, w_008_135, w_008_136, w_008_137, w_008_138, w_008_139, w_008_140, w_008_141, w_008_142, w_008_143, w_008_144, w_008_145, w_008_146, w_008_147, w_008_148, w_008_149, w_008_150, w_008_151, w_008_152, w_008_153, w_008_154, w_008_155, w_008_156, w_008_157, w_008_158, w_008_159, w_008_160, w_008_161, w_008_162, w_008_163, w_008_164, w_008_165, w_008_166, w_008_167, w_008_168, w_008_169, w_008_170, w_008_171, w_008_172, w_008_173, w_008_174, w_008_175, w_008_176, w_008_178, w_008_179, w_008_180, w_008_181, w_008_182, w_008_183, w_008_184, w_008_185, w_008_186, w_008_187, w_008_188, w_008_189, w_008_190, w_008_191, w_008_192, w_008_193, w_008_194, w_008_195, w_008_196, w_008_197, w_008_198, w_008_199, w_008_200, w_008_201, w_008_202, w_008_203, w_008_204, w_008_205, w_008_206, w_008_207, w_008_208, w_008_209, w_008_210, w_008_211, w_008_212, w_008_213, w_008_214, w_008_215, w_008_216, w_008_217, w_008_218, w_008_219, w_008_220, w_008_221, w_008_222, w_008_223, w_008_224, w_008_225, w_008_226, w_008_227, w_008_228, w_008_229, w_008_230, w_008_231, w_008_232, w_008_233, w_008_234, w_008_235, w_008_236, w_008_237, w_008_238, w_008_239, w_008_240, w_008_241, w_008_242, w_008_243, w_008_244, w_008_245, w_008_246, w_008_247, w_008_248, w_008_250, w_008_251, w_008_252, w_008_253, w_008_254, w_008_255, w_008_256, w_008_257, w_008_258, w_008_259, w_008_260, w_008_261, w_008_262, w_008_263, w_008_264, w_008_265, w_008_266, w_008_267, w_008_268, w_008_269, w_008_270, w_008_271, w_008_272, w_008_273, w_008_274, w_008_275, w_008_276, w_008_277, w_008_278, w_008_279, w_008_280, w_008_281, w_008_282, w_008_283, w_008_284, w_008_285, w_008_286, w_008_287, w_008_288, w_008_289, w_008_290, w_008_291, w_008_292, w_008_293, w_008_294, w_008_295, w_008_296, w_008_297, w_008_298, w_008_299, w_008_300, w_008_301, w_008_302, w_008_303, w_008_304, w_008_305, w_008_307, w_008_308, w_008_309, w_008_310, w_008_311, w_008_312, w_008_313, w_008_315, w_008_316, w_008_317, w_008_318, w_008_319, w_008_320, w_008_321, w_008_322, w_008_323, w_008_324, w_008_325, w_008_326, w_008_327, w_008_328, w_008_329, w_008_330, w_008_331, w_008_332, w_008_333, w_008_334, w_008_335, w_008_336, w_008_337, w_008_338, w_008_339, w_008_340, w_008_341, w_008_342, w_008_343, w_008_344, w_008_345, w_008_346, w_008_347, w_008_348, w_008_349, w_008_350, w_008_351, w_008_352, w_008_353, w_008_355, w_008_356, w_008_357, w_008_358, w_008_359, w_008_360, w_008_361, w_008_362, w_008_363, w_008_364, w_008_365, w_008_366, w_008_367, w_008_368, w_008_369, w_008_370, w_008_371, w_008_372, w_008_373, w_008_374, w_008_375, w_008_376, w_008_377, w_008_378, w_008_379, w_008_380, w_008_381, w_008_382, w_008_383, w_008_384, w_008_385, w_008_386, w_008_387, w_008_388, w_008_389, w_008_391, w_008_392, w_008_393, w_008_394, w_008_395, w_008_396, w_008_397, w_008_398, w_008_399, w_008_400, w_008_401, w_008_402, w_008_403, w_008_404, w_008_405, w_008_406, w_008_407, w_008_408, w_008_409, w_008_410, w_008_411, w_008_412, w_008_413, w_008_414, w_008_415, w_008_416, w_008_417, w_008_418, w_008_419, w_008_420, w_008_421, w_008_422, w_008_423, w_008_424, w_008_425, w_008_426, w_008_427, w_008_428, w_008_430, w_008_431, w_008_432, w_008_433, w_008_434, w_008_435, w_008_436, w_008_437, w_008_438, w_008_439, w_008_440, w_008_441, w_008_442, w_008_443, w_008_444, w_008_445, w_008_446, w_008_447, w_008_448, w_008_449, w_008_450, w_008_451, w_008_452, w_008_453, w_008_454, w_008_455, w_008_456, w_008_457, w_008_458, w_008_459, w_008_460, w_008_461, w_008_462, w_008_463, w_008_464, w_008_465, w_008_466, w_008_467, w_008_468, w_008_469, w_008_470, w_008_471, w_008_472, w_008_473, w_008_474, w_008_475, w_008_476, w_008_477, w_008_478, w_008_479, w_008_480, w_008_481, w_008_482, w_008_483, w_008_484, w_008_485, w_008_486, w_008_487, w_008_488, w_008_489, w_008_490, w_008_491, w_008_492, w_008_493, w_008_494, w_008_495, w_008_496, w_008_497, w_008_498, w_008_499, w_008_500, w_008_501, w_008_502, w_008_503, w_008_505, w_008_506, w_008_507, w_008_508, w_008_509, w_008_510, w_008_511, w_008_512, w_008_514, w_008_515, w_008_516, w_008_517, w_008_518, w_008_519, w_008_520, w_008_521, w_008_522, w_008_523, w_008_524, w_008_525, w_008_527, w_008_528, w_008_529, w_008_530, w_008_531, w_008_532, w_008_533, w_008_534, w_008_535, w_008_536, w_008_537, w_008_538, w_008_539, w_008_540, w_008_541, w_008_542, w_008_543, w_008_544, w_008_545, w_008_546, w_008_547, w_008_548, w_008_549, w_008_550, w_008_551, w_008_552, w_008_553, w_008_554, w_008_555, w_008_556, w_008_557, w_008_558, w_008_559, w_008_560, w_008_561, w_008_562, w_008_563, w_008_564, w_008_565, w_008_566, w_008_567, w_008_568, w_008_569, w_008_570, w_008_571, w_008_572, w_008_573, w_008_574, w_008_575, w_008_576, w_008_577, w_008_578, w_008_580, w_008_581, w_008_582, w_008_583, w_008_584, w_008_585, w_008_586, w_008_587, w_008_588, w_008_589, w_008_590, w_008_591, w_008_592, w_008_593, w_008_594, w_008_595, w_008_596, w_008_597, w_008_598, w_008_599, w_008_600, w_008_601, w_008_602, w_008_603, w_008_604, w_008_605, w_008_606, w_008_607, w_008_608, w_008_609, w_008_610, w_008_611, w_008_612, w_008_613, w_008_614, w_008_615, w_008_616, w_008_617, w_008_618, w_008_619, w_008_620, w_008_621, w_008_622, w_008_623, w_008_624, w_008_625, w_008_626, w_008_627, w_008_628, w_008_629, w_008_630, w_008_631, w_008_632, w_008_633, w_008_634, w_008_635, w_008_636, w_008_637, w_008_638, w_008_639, w_008_640, w_008_641, w_008_642, w_008_643, w_008_644, w_008_645, w_008_646, w_008_647, w_008_648, w_008_649, w_008_650, w_008_651, w_008_652, w_008_653, w_008_654, w_008_655, w_008_657, w_008_658, w_008_659, w_008_660, w_008_661, w_008_662, w_008_663, w_008_664, w_008_665, w_008_666, w_008_667, w_008_668, w_008_669, w_008_670, w_008_671, w_008_672, w_008_673, w_008_675, w_008_676, w_008_677, w_008_678, w_008_679, w_008_680, w_008_681, w_008_682, w_008_683, w_008_684, w_008_685, w_008_686, w_008_687, w_008_688, w_008_689, w_008_690, w_008_691, w_008_692, w_008_693, w_008_694, w_008_695, w_008_696, w_008_697, w_008_698, w_008_699, w_008_700, w_008_701, w_008_702, w_008_703, w_008_704, w_008_705, w_008_706, w_008_707, w_008_708, w_008_709, w_008_710, w_008_711, w_008_712, w_008_713, w_008_714, w_008_715, w_008_716, w_008_717, w_008_718, w_008_719, w_008_720, w_008_721, w_008_722, w_008_723, w_008_724, w_008_725, w_008_726, w_008_727, w_008_728, w_008_729, w_008_730, w_008_731, w_008_732, w_008_733, w_008_734, w_008_735, w_008_736, w_008_737, w_008_738, w_008_739, w_008_740, w_008_741, w_008_742, w_008_743, w_008_744, w_008_745, w_008_746, w_008_747, w_008_748, w_008_749, w_008_750, w_008_751, w_008_752, w_008_753, w_008_754, w_008_755, w_008_756, w_008_757, w_008_758, w_008_759, w_008_760, w_008_761, w_008_762, w_008_763, w_008_764, w_008_765, w_008_766, w_008_767, w_008_768, w_008_769, w_008_770, w_008_771, w_008_772, w_008_773, w_008_774, w_008_775, w_008_776, w_008_777, w_008_778, w_008_779, w_008_780, w_008_781, w_008_782, w_008_783, w_008_784, w_008_785, w_008_786, w_008_788, w_008_789, w_008_790, w_008_791, w_008_792, w_008_793, w_008_795, w_008_796, w_008_797, w_008_798, w_008_799, w_008_800, w_008_801, w_008_802, w_008_803, w_008_804, w_008_805, w_008_806, w_008_807, w_008_808, w_008_809, w_008_810, w_008_811, w_008_812, w_008_813, w_008_814, w_008_815, w_008_816, w_008_818, w_008_819, w_008_820, w_008_821, w_008_822, w_008_823, w_008_824, w_008_825, w_008_826, w_008_827, w_008_828, w_008_829, w_008_830, w_008_831, w_008_832, w_008_833, w_008_834, w_008_835, w_008_836, w_008_837, w_008_838, w_008_839, w_008_840, w_008_841, w_008_842, w_008_843, w_008_844, w_008_845, w_008_846, w_008_847, w_008_848, w_008_849, w_008_850, w_008_851, w_008_852, w_008_853, w_008_854, w_008_855, w_008_856, w_008_857, w_008_858, w_008_859, w_008_860, w_008_861, w_008_862, w_008_863, w_008_864, w_008_865, w_008_866, w_008_867, w_008_868, w_008_869, w_008_870, w_008_871, w_008_872, w_008_873, w_008_874, w_008_875, w_008_876, w_008_878, w_008_879, w_008_880, w_008_881, w_008_882, w_008_883, w_008_884, w_008_885, w_008_886, w_008_887, w_008_888, w_008_889, w_008_890, w_008_891, w_008_892, w_008_893, w_008_894, w_008_895, w_008_896, w_008_897, w_008_898, w_008_899, w_008_900, w_008_901, w_008_902, w_008_903, w_008_904, w_008_905, w_008_906, w_008_907, w_008_908, w_008_909, w_008_910, w_008_911, w_008_912, w_008_913, w_008_914, w_008_915, w_008_916, w_008_917, w_008_918, w_008_919, w_008_920, w_008_921, w_008_922, w_008_923, w_008_924, w_008_925, w_008_926, w_008_927, w_008_928, w_008_930, w_008_931, w_008_932, w_008_933, w_008_934, w_008_935, w_008_936, w_008_938, w_008_939, w_008_940, w_008_941, w_008_942, w_008_943, w_008_944, w_008_945, w_008_946, w_008_947, w_008_948, w_008_949, w_008_951, w_008_952, w_008_953, w_008_954, w_008_955, w_008_956, w_008_957, w_008_958, w_008_960, w_008_961, w_008_962, w_008_963, w_008_964, w_008_965, w_008_966, w_008_967, w_008_968, w_008_969, w_008_970, w_008_971, w_008_972, w_008_973, w_008_974, w_008_975, w_008_976, w_008_977, w_008_978, w_008_979, w_008_980, w_008_981, w_008_982, w_008_983, w_008_984, w_008_985, w_008_986, w_008_987, w_008_988, w_008_989, w_008_990, w_008_991, w_008_992, w_008_993, w_008_994, w_008_995, w_008_996, w_008_997, w_008_998, w_008_999, w_008_1000, w_008_1001, w_008_1002, w_008_1003, w_008_1004, w_008_1005, w_008_1006, w_008_1007, w_008_1008, w_008_1009, w_008_1010, w_008_1011, w_008_1012, w_008_1013, w_008_1014, w_008_1015, w_008_1016, w_008_1017, w_008_1018, w_008_1019, w_008_1020, w_008_1021, w_008_1022, w_008_1023, w_008_1024, w_008_1025, w_008_1026, w_008_1027, w_008_1028, w_008_1029, w_008_1030, w_008_1031, w_008_1032, w_008_1033, w_008_1034, w_008_1035, w_008_1036, w_008_1037, w_008_1038, w_008_1039, w_008_1040, w_008_1041, w_008_1042, w_008_1043, w_008_1044, w_008_1045, w_008_1046, w_008_1047, w_008_1048, w_008_1049, w_008_1050, w_008_1051, w_008_1052, w_008_1053, w_008_1054, w_008_1055, w_008_1056, w_008_1057, w_008_1058, w_008_1059, w_008_1060, w_008_1061, w_008_1062, w_008_1063, w_008_1064, w_008_1065, w_008_1066, w_008_1067, w_008_1068, w_008_1069, w_008_1070, w_008_1071, w_008_1072, w_008_1073, w_008_1074, w_008_1075, w_008_1076, w_008_1077, w_008_1078, w_008_1079, w_008_1080, w_008_1081, w_008_1082, w_008_1083, w_008_1084, w_008_1085, w_008_1086, w_008_1087, w_008_1088, w_008_1089, w_008_1090, w_008_1091, w_008_1092, w_008_1093, w_008_1094, w_008_1095, w_008_1096, w_008_1097, w_008_1099, w_008_1100, w_008_1101, w_008_1102, w_008_1103, w_008_1104, w_008_1105, w_008_1106, w_008_1107, w_008_1108, w_008_1109, w_008_1110, w_008_1111, w_008_1112, w_008_1113, w_008_1114, w_008_1115, w_008_1116, w_008_1117, w_008_1118, w_008_1119, w_008_1120, w_008_1121, w_008_1122, w_008_1123, w_008_1124, w_008_1125, w_008_1126, w_008_1127, w_008_1128, w_008_1129, w_008_1130, w_008_1131, w_008_1132, w_008_1133, w_008_1134, w_008_1135, w_008_1136, w_008_1137, w_008_1138, w_008_1139, w_008_1140, w_008_1141, w_008_1142, w_008_1143, w_008_1144, w_008_1145, w_008_1146, w_008_1147, w_008_1148, w_008_1149, w_008_1150, w_008_1151, w_008_1152, w_008_1153, w_008_1154, w_008_1155, w_008_1156, w_008_1157, w_008_1158, w_008_1159, w_008_1160, w_008_1161, w_008_1162, w_008_1163, w_008_1164, w_008_1165, w_008_1166, w_008_1167, w_008_1168, w_008_1169, w_008_1170, w_008_1171, w_008_1172, w_008_1173, w_008_1174, w_008_1175, w_008_1176, w_008_1177, w_008_1178, w_008_1179, w_008_1180, w_008_1181, w_008_1182, w_008_1183, w_008_1184, w_008_1185, w_008_1186, w_008_1187, w_008_1188, w_008_1189, w_008_1190, w_008_1191, w_008_1192, w_008_1193, w_008_1194, w_008_1195, w_008_1196, w_008_1197, w_008_1198, w_008_1199, w_008_1200, w_008_1201, w_008_1202, w_008_1203, w_008_1204, w_008_1205, w_008_1206, w_008_1207, w_008_1209, w_008_1210, w_008_1211, w_008_1212, w_008_1213, w_008_1214, w_008_1215, w_008_1216, w_008_1217, w_008_1218, w_008_1220, w_008_1221, w_008_1222, w_008_1223, w_008_1224, w_008_1225, w_008_1226, w_008_1227, w_008_1228, w_008_1229, w_008_1230, w_008_1231, w_008_1232, w_008_1233, w_008_1234, w_008_1235, w_008_1236, w_008_1237, w_008_1238, w_008_1240, w_008_1241, w_008_1242, w_008_1243, w_008_1244, w_008_1245, w_008_1246, w_008_1247, w_008_1248, w_008_1249, w_008_1250, w_008_1251, w_008_1252, w_008_1253, w_008_1254, w_008_1255, w_008_1256, w_008_1257, w_008_1258, w_008_1259, w_008_1260, w_008_1261, w_008_1262, w_008_1263, w_008_1264, w_008_1265, w_008_1266, w_008_1267, w_008_1268, w_008_1269, w_008_1270, w_008_1271, w_008_1272, w_008_1273, w_008_1274, w_008_1275, w_008_1276, w_008_1277, w_008_1278, w_008_1279, w_008_1280, w_008_1281, w_008_1282, w_008_1283, w_008_1285, w_008_1286, w_008_1287, w_008_1288, w_008_1289, w_008_1290, w_008_1291, w_008_1292, w_008_1293, w_008_1294, w_008_1295, w_008_1296, w_008_1297, w_008_1298, w_008_1299, w_008_1300, w_008_1301, w_008_1302, w_008_1303, w_008_1304, w_008_1305, w_008_1306, w_008_1307, w_008_1308, w_008_1309, w_008_1310, w_008_1311, w_008_1312, w_008_1313, w_008_1314, w_008_1315, w_008_1316, w_008_1317, w_008_1318, w_008_1319, w_008_1320, w_008_1321, w_008_1322, w_008_1323, w_008_1324, w_008_1325, w_008_1326, w_008_1327, w_008_1328, w_008_1329, w_008_1330, w_008_1331, w_008_1332, w_008_1333, w_008_1334, w_008_1335, w_008_1336, w_008_1337, w_008_1338, w_008_1339, w_008_1340, w_008_1341, w_008_1342, w_008_1343, w_008_1344, w_008_1345, w_008_1346, w_008_1347, w_008_1348, w_008_1349, w_008_1350, w_008_1351, w_008_1352, w_008_1353, w_008_1354, w_008_1355, w_008_1356, w_008_1357, w_008_1358, w_008_1359, w_008_1360, w_008_1361, w_008_1362, w_008_1363, w_008_1364, w_008_1365, w_008_1366, w_008_1367, w_008_1368, w_008_1369, w_008_1370, w_008_1371, w_008_1372, w_008_1373, w_008_1374, w_008_1375, w_008_1376, w_008_1377, w_008_1378, w_008_1379, w_008_1380, w_008_1381, w_008_1382, w_008_1383, w_008_1384, w_008_1385, w_008_1386, w_008_1387, w_008_1388, w_008_1389, w_008_1390, w_008_1391, w_008_1392, w_008_1394, w_008_1395, w_008_1396, w_008_1397, w_008_1398, w_008_1399, w_008_1400, w_008_1401, w_008_1402, w_008_1403, w_008_1404, w_008_1405, w_008_1406, w_008_1407, w_008_1408, w_008_1409, w_008_1410, w_008_1411, w_008_1412, w_008_1413, w_008_1414, w_008_1415, w_008_1416, w_008_1417, w_008_1418, w_008_1419, w_008_1420, w_008_1421, w_008_1422, w_008_1423, w_008_1424, w_008_1425, w_008_1426, w_008_1427, w_008_1428, w_008_1429, w_008_1430, w_008_1431, w_008_1432, w_008_1433, w_008_1434, w_008_1435, w_008_1436, w_008_1437, w_008_1438, w_008_1439, w_008_1440, w_008_1441, w_008_1442, w_008_1443, w_008_1444, w_008_1445, w_008_1446, w_008_1447, w_008_1448, w_008_1449, w_008_1450, w_008_1451, w_008_1452, w_008_1453, w_008_1454, w_008_1455, w_008_1456, w_008_1457, w_008_1458, w_008_1459, w_008_1460, w_008_1461, w_008_1462, w_008_1463, w_008_1464, w_008_1465, w_008_1467, w_008_1468, w_008_1469, w_008_1470, w_008_1471, w_008_1472, w_008_1473, w_008_1474, w_008_1475, w_008_1476, w_008_1477, w_008_1478, w_008_1479, w_008_1480, w_008_1481, w_008_1482, w_008_1483, w_008_1484, w_008_1485, w_008_1486, w_008_1487, w_008_1488, w_008_1489, w_008_1490, w_008_1491, w_008_1492, w_008_1493, w_008_1494, w_008_1495, w_008_1496, w_008_1497, w_008_1498, w_008_1499, w_008_1500, w_008_1501, w_008_1502, w_008_1503, w_008_1504, w_008_1505, w_008_1506, w_008_1507, w_008_1508, w_008_1509, w_008_1510, w_008_1511, w_008_1512, w_008_1513, w_008_1514, w_008_1515, w_008_1516, w_008_1517, w_008_1518, w_008_1519, w_008_1520, w_008_1521, w_008_1522, w_008_1523, w_008_1524, w_008_1525, w_008_1526, w_008_1527, w_008_1528, w_008_1529, w_008_1530, w_008_1531, w_008_1532, w_008_1533, w_008_1534, w_008_1535, w_008_1536, w_008_1537, w_008_1538, w_008_1539, w_008_1540, w_008_1541, w_008_1542, w_008_1543, w_008_1544, w_008_1545, w_008_1546, w_008_1547, w_008_1548, w_008_1549, w_008_1550, w_008_1551, w_008_1552, w_008_1553, w_008_1554, w_008_1555, w_008_1556, w_008_1557, w_008_1558, w_008_1559, w_008_1560, w_008_1561, w_008_1562, w_008_1563, w_008_1564, w_008_1565, w_008_1566, w_008_1567, w_008_1568, w_008_1569, w_008_1570, w_008_1571, w_008_1572, w_008_1573, w_008_1574, w_008_1575, w_008_1576, w_008_1577, w_008_1578, w_008_1579, w_008_1580, w_008_1581, w_008_1582, w_008_1584, w_008_1585, w_008_1586, w_008_1587, w_008_1588, w_008_1589, w_008_1590, w_008_1591, w_008_1592, w_008_1593, w_008_1594, w_008_1595, w_008_1596, w_008_1597, w_008_1598, w_008_1599, w_008_1600, w_008_1601, w_008_1602, w_008_1603, w_008_1604, w_008_1605, w_008_1606, w_008_1607, w_008_1608, w_008_1609, w_008_1610, w_008_1611, w_008_1612, w_008_1613, w_008_1614, w_008_1615, w_008_1616, w_008_1617, w_008_1618, w_008_1619, w_008_1620, w_008_1621, w_008_1622, w_008_1623, w_008_1624, w_008_1627, w_008_1628, w_008_1629, w_008_1630, w_008_1631, w_008_1632, w_008_1633, w_008_1634, w_008_1635, w_008_1636, w_008_1637, w_008_1638, w_008_1639, w_008_1640, w_008_1642, w_008_1643, w_008_1644, w_008_1645, w_008_1646, w_008_1647, w_008_1648, w_008_1650, w_008_1651, w_008_1652, w_008_1653, w_008_1654, w_008_1655, w_008_1656, w_008_1657, w_008_1658, w_008_1659, w_008_1660, w_008_1661, w_008_1662, w_008_1663, w_008_1664, w_008_1665, w_008_1666, w_008_1667, w_008_1669, w_008_1670, w_008_1671, w_008_1672, w_008_1673, w_008_1674, w_008_1675, w_008_1676, w_008_1677, w_008_1678, w_008_1679, w_008_1680, w_008_1681, w_008_1682, w_008_1683, w_008_1684, w_008_1685, w_008_1686, w_008_1687, w_008_1688, w_008_1689, w_008_1690, w_008_1691, w_008_1692, w_008_1693, w_008_1694, w_008_1695, w_008_1696, w_008_1697, w_008_1698, w_008_1699, w_008_1700, w_008_1701, w_008_1702, w_008_1703, w_008_1704, w_008_1705, w_008_1706, w_008_1707, w_008_1708, w_008_1709, w_008_1710, w_008_1711, w_008_1712, w_008_1713, w_008_1714, w_008_1715, w_008_1716, w_008_1717, w_008_1718, w_008_1719, w_008_1720, w_008_1721, w_008_1722, w_008_1723, w_008_1724, w_008_1725, w_008_1726, w_008_1727, w_008_1728, w_008_1729, w_008_1731, w_008_1732, w_008_1733, w_008_1734, w_008_1735, w_008_1736, w_008_1737, w_008_1738, w_008_1739, w_008_1740, w_008_1741, w_008_1742, w_008_1743, w_008_1744, w_008_1745, w_008_1746, w_008_1747, w_008_1748, w_008_1750, w_008_1751, w_008_1752, w_008_1753, w_008_1754, w_008_1755, w_008_1756, w_008_1757, w_008_1758, w_008_1759, w_008_1760, w_008_1761, w_008_1762, w_008_1763, w_008_1764, w_008_1765, w_008_1766, w_008_1767, w_008_1768, w_008_1769, w_008_1770, w_008_1771, w_008_1772, w_008_1773, w_008_1774, w_008_1775, w_008_1776, w_008_1777, w_008_1778, w_008_1779, w_008_1780, w_008_1781, w_008_1783, w_008_1784, w_008_1785, w_008_1786, w_008_1787, w_008_1788, w_008_1789, w_008_1790, w_008_1791, w_008_1792, w_008_1793, w_008_1794, w_008_1795, w_008_1796, w_008_1797, w_008_1798, w_008_1799, w_008_1800, w_008_1801, w_008_1802, w_008_1803, w_008_1804, w_008_1805, w_008_1806, w_008_1807, w_008_1808, w_008_1809, w_008_1811, w_008_1812, w_008_1813, w_008_1814, w_008_1815, w_008_1816, w_008_1817, w_008_1818, w_008_1820, w_008_1821, w_008_1822, w_008_1823, w_008_1824, w_008_1825, w_008_1826, w_008_1827, w_008_1828, w_008_1829, w_008_1830, w_008_1831, w_008_1832, w_008_1833, w_008_1834, w_008_1835, w_008_1836, w_008_1837, w_008_1838, w_008_1839, w_008_1840, w_008_1841, w_008_1842, w_008_1843, w_008_1844, w_008_1845, w_008_1846, w_008_1847, w_008_1848, w_008_1849, w_008_1850, w_008_1851, w_008_1852, w_008_1853, w_008_1854, w_008_1855, w_008_1856, w_008_1857, w_008_1858, w_008_1859, w_008_1860, w_008_1861, w_008_1862, w_008_1863, w_008_1864, w_008_1865, w_008_1866, w_008_1868, w_008_1869, w_008_1870, w_008_1871, w_008_1872, w_008_1873, w_008_1874, w_008_1875, w_008_1876, w_008_1877, w_008_1878, w_008_1879, w_008_1880, w_008_1881, w_008_1882, w_008_1883, w_008_1886, w_008_1887, w_008_1888, w_008_1889, w_008_1890, w_008_1891, w_008_1892, w_008_1893, w_008_1894, w_008_1895, w_008_1896, w_008_1897, w_008_1898, w_008_1899, w_008_1900, w_008_1901, w_008_1902, w_008_1903, w_008_1904, w_008_1905, w_008_1906, w_008_1907, w_008_1908, w_008_1909, w_008_1910, w_008_1911, w_008_1912, w_008_1913, w_008_1914, w_008_1915, w_008_1916, w_008_1917, w_008_1918, w_008_1919, w_008_1921, w_008_1922, w_008_1923, w_008_1924, w_008_1925, w_008_1926, w_008_1927, w_008_1928, w_008_1930, w_008_1931, w_008_1932, w_008_1933, w_008_1934, w_008_1935, w_008_1936, w_008_1937, w_008_1938, w_008_1939, w_008_1940, w_008_1941, w_008_1942, w_008_1943, w_008_1944, w_008_1945, w_008_1946, w_008_1947, w_008_1948, w_008_1949, w_008_1950, w_008_1951, w_008_1952, w_008_1953, w_008_1954, w_008_1955, w_008_1956, w_008_1957, w_008_1958, w_008_1959, w_008_1960, w_008_1961, w_008_1962, w_008_1963, w_008_1964, w_008_1965, w_008_1966, w_008_1967, w_008_1968, w_008_1969, w_008_1970, w_008_1971, w_008_1972, w_008_1973, w_008_1974, w_008_1975, w_008_1976, w_008_1977, w_008_1978, w_008_1979, w_008_1980, w_008_1981, w_008_1982, w_008_1983, w_008_1984, w_008_1985, w_008_1986, w_008_1987, w_008_1988, w_008_1989, w_008_1990, w_008_1991, w_008_1992, w_008_1993, w_008_1994, w_008_1995, w_008_1996, w_008_1997, w_008_1998, w_008_1999, w_008_2000, w_008_2001, w_008_2002, w_008_2003, w_008_2004, w_008_2006, w_008_2007, w_008_2008, w_008_2009, w_008_2010, w_008_2011, w_008_2012, w_008_2013, w_008_2014, w_008_2015, w_008_2016, w_008_2017, w_008_2018, w_008_2019, w_008_2020, w_008_2021, w_008_2022, w_008_2023, w_008_2024, w_008_2025, w_008_2026, w_008_2027, w_008_2028, w_008_2029, w_008_2030, w_008_2031, w_008_2032, w_008_2033, w_008_2034, w_008_2035, w_008_2036, w_008_2037, w_008_2038, w_008_2039, w_008_2040, w_008_2041, w_008_2042, w_008_2043, w_008_2044, w_008_2045, w_008_2046, w_008_2047, w_008_2048, w_008_2049, w_008_2050, w_008_2051, w_008_2052, w_008_2053, w_008_2054, w_008_2055, w_008_2056, w_008_2057, w_008_2058, w_008_2059, w_008_2060, w_008_2061, w_008_2062, w_008_2063, w_008_2064, w_008_2065, w_008_2066, w_008_2067, w_008_2068, w_008_2069, w_008_2070, w_008_2071, w_008_2072, w_008_2073, w_008_2074, w_008_2075, w_008_2076, w_008_2077, w_008_2078, w_008_2079, w_008_2080, w_008_2081, w_008_2082, w_008_2083, w_008_2084, w_008_2085, w_008_2086, w_008_2087, w_008_2088, w_008_2089, w_008_2090, w_008_2091, w_008_2092, w_008_2093, w_008_2095, w_008_2096, w_008_2097, w_008_2098, w_008_2099, w_008_2100, w_008_2101, w_008_2102, w_008_2103, w_008_2104, w_008_2105, w_008_2106, w_008_2107, w_008_2108, w_008_2109, w_008_2110, w_008_2111, w_008_2112, w_008_2113, w_008_2114, w_008_2115, w_008_2116, w_008_2117, w_008_2118, w_008_2119, w_008_2120, w_008_2121, w_008_2122, w_008_2123, w_008_2124, w_008_2125, w_008_2126, w_008_2127, w_008_2128, w_008_2129, w_008_2130, w_008_2131, w_008_2132, w_008_2133, w_008_2134, w_008_2135, w_008_2136, w_008_2137, w_008_2138, w_008_2139, w_008_2140, w_008_2141, w_008_2142, w_008_2143, w_008_2144, w_008_2145, w_008_2146, w_008_2147, w_008_2148, w_008_2149, w_008_2150, w_008_2151, w_008_2152, w_008_2153, w_008_2154, w_008_2155, w_008_2156, w_008_2157, w_008_2158, w_008_2159, w_008_2160, w_008_2161, w_008_2162, w_008_2163, w_008_2164, w_008_2165, w_008_2166, w_008_2167, w_008_2168, w_008_2169, w_008_2170, w_008_2171, w_008_2172, w_008_2173, w_008_2174, w_008_2175, w_008_2176, w_008_2177, w_008_2178, w_008_2179, w_008_2180, w_008_2181, w_008_2182, w_008_2183, w_008_2184, w_008_2185, w_008_2187, w_008_2188, w_008_2189, w_008_2190, w_008_2191, w_008_2192, w_008_2193, w_008_2194, w_008_2195, w_008_2196, w_008_2197, w_008_2198, w_008_2199, w_008_2200, w_008_2201, w_008_2202, w_008_2203, w_008_2204, w_008_2205, w_008_2206, w_008_2207, w_008_2208, w_008_2209, w_008_2210, w_008_2211, w_008_2212, w_008_2213, w_008_2214, w_008_2215, w_008_2216, w_008_2217, w_008_2218, w_008_2220, w_008_2221, w_008_2222, w_008_2223, w_008_2224, w_008_2225, w_008_2226, w_008_2227, w_008_2228, w_008_2229, w_008_2230, w_008_2232, w_008_2233, w_008_2234, w_008_2235, w_008_2236, w_008_2237, w_008_2238, w_008_2239, w_008_2240, w_008_2241, w_008_2242, w_008_2243, w_008_2244, w_008_2245, w_008_2246, w_008_2247, w_008_2248, w_008_2251, w_008_2252, w_008_2253, w_008_2254, w_008_2255, w_008_2256, w_008_2257, w_008_2258, w_008_2259, w_008_2260, w_008_2261, w_008_2262, w_008_2263, w_008_2264, w_008_2265, w_008_2266, w_008_2267, w_008_2269, w_008_2270, w_008_2271, w_008_2272, w_008_2273, w_008_2274, w_008_2275, w_008_2276, w_008_2277, w_008_2278, w_008_2279, w_008_2280, w_008_2282, w_008_2283, w_008_2284, w_008_2285, w_008_2286, w_008_2287, w_008_2288, w_008_2289, w_008_2290, w_008_2291, w_008_2292, w_008_2293, w_008_2294, w_008_2295, w_008_2296, w_008_2297, w_008_2298, w_008_2299, w_008_2300, w_008_2301, w_008_2302, w_008_2303, w_008_2304, w_008_2305, w_008_2306, w_008_2307, w_008_2308, w_008_2309, w_008_2310, w_008_2311, w_008_2312, w_008_2313, w_008_2314, w_008_2315, w_008_2316, w_008_2317, w_008_2319, w_008_2320, w_008_2321, w_008_2322, w_008_2323, w_008_2324, w_008_2325, w_008_2326, w_008_2328, w_008_2329, w_008_2330, w_008_2331, w_008_2332, w_008_2333, w_008_2334, w_008_2335, w_008_2336, w_008_2337, w_008_2338, w_008_2339, w_008_2340, w_008_2341, w_008_2342, w_008_2343, w_008_2344, w_008_2345, w_008_2346, w_008_2347, w_008_2349, w_008_2350, w_008_2351, w_008_2352, w_008_2353, w_008_2354, w_008_2355, w_008_2356, w_008_2357, w_008_2358, w_008_2359, w_008_2360, w_008_2361, w_008_2362, w_008_2363, w_008_2364, w_008_2365, w_008_2366, w_008_2367, w_008_2368, w_008_2369, w_008_2370, w_008_2371, w_008_2373, w_008_2374, w_008_2375, w_008_2376, w_008_2377, w_008_2378, w_008_2379, w_008_2380, w_008_2381, w_008_2382, w_008_2383, w_008_2384, w_008_2385, w_008_2386, w_008_2387, w_008_2388, w_008_2389, w_008_2390, w_008_2391, w_008_2392, w_008_2393, w_008_2394, w_008_2395, w_008_2396, w_008_2397, w_008_2398, w_008_2399, w_008_2400, w_008_2401, w_008_2402, w_008_2404, w_008_2405, w_008_2406, w_008_2407, w_008_2408, w_008_2409, w_008_2410, w_008_2411, w_008_2412, w_008_2413, w_008_2414, w_008_2415, w_008_2416, w_008_2417, w_008_2418, w_008_2419, w_008_2420, w_008_2421, w_008_2422, w_008_2423, w_008_2424, w_008_2425, w_008_2426, w_008_2427, w_008_2428, w_008_2429, w_008_2430, w_008_2431, w_008_2432, w_008_2433, w_008_2434, w_008_2435, w_008_2436, w_008_2437, w_008_2438, w_008_2439, w_008_2440, w_008_2441, w_008_2442, w_008_2443, w_008_2444, w_008_2445, w_008_2446, w_008_2447, w_008_2448, w_008_2449, w_008_2450, w_008_2451, w_008_2452, w_008_2453, w_008_2454, w_008_2455, w_008_2456, w_008_2457, w_008_2458, w_008_2459, w_008_2461, w_008_2462, w_008_2463, w_008_2464, w_008_2465, w_008_2466, w_008_2467, w_008_2468, w_008_2470, w_008_2471, w_008_2472, w_008_2473, w_008_2474, w_008_2475, w_008_2476, w_008_2477, w_008_2478, w_008_2479, w_008_2480, w_008_2481, w_008_2482, w_008_2483, w_008_2484, w_008_2485, w_008_2486, w_008_2488, w_008_2489, w_008_2490, w_008_2491, w_008_2493, w_008_2494, w_008_2496, w_008_2497, w_008_2499, w_008_2500, w_008_2501, w_008_2502, w_008_2503, w_008_2504, w_008_2505, w_008_2506, w_008_2507, w_008_2510, w_008_2511, w_008_2513, w_008_2515, w_008_2516, w_008_2517, w_008_2518, w_008_2519, w_008_2520, w_008_2521, w_008_2522, w_008_2523, w_008_2525, w_008_2527, w_008_2528, w_008_2529, w_008_2530, w_008_2531, w_008_2532, w_008_2533, w_008_2534, w_008_2535, w_008_2536, w_008_2537, w_008_2538, w_008_2540, w_008_2542, w_008_2543, w_008_2544, w_008_2545, w_008_2547, w_008_2548, w_008_2549, w_008_2552, w_008_2554, w_008_2556, w_008_2557, w_008_2558, w_008_2559, w_008_2560, w_008_2561, w_008_2562, w_008_2563, w_008_2564, w_008_2565, w_008_2566, w_008_2567, w_008_2568, w_008_2570, w_008_2571;
  wire w_009_000, w_009_001, w_009_002, w_009_003, w_009_005, w_009_006, w_009_007, w_009_008, w_009_009, w_009_010, w_009_011, w_009_012, w_009_013, w_009_014, w_009_015, w_009_017, w_009_018, w_009_019, w_009_020, w_009_021, w_009_022, w_009_023, w_009_024, w_009_025, w_009_026, w_009_027, w_009_028, w_009_029, w_009_030, w_009_031, w_009_032, w_009_033, w_009_034, w_009_035, w_009_036, w_009_037, w_009_038, w_009_039, w_009_040, w_009_041, w_009_042, w_009_043, w_009_044, w_009_045, w_009_046, w_009_047, w_009_048, w_009_049, w_009_050, w_009_051, w_009_052, w_009_053, w_009_054, w_009_055, w_009_056, w_009_057, w_009_058, w_009_059, w_009_060, w_009_062, w_009_063, w_009_064, w_009_065, w_009_066, w_009_067, w_009_068, w_009_069, w_009_070, w_009_071, w_009_072, w_009_074, w_009_075, w_009_076, w_009_077, w_009_078, w_009_079, w_009_080, w_009_081, w_009_082, w_009_083, w_009_084, w_009_085, w_009_086, w_009_087, w_009_088, w_009_089, w_009_090, w_009_091, w_009_092, w_009_093, w_009_094, w_009_095, w_009_096, w_009_097, w_009_098, w_009_099, w_009_100, w_009_101, w_009_102, w_009_103, w_009_104, w_009_105, w_009_106, w_009_107, w_009_108, w_009_109, w_009_110, w_009_111, w_009_112, w_009_113, w_009_114, w_009_115, w_009_116, w_009_117, w_009_118, w_009_119, w_009_120, w_009_121, w_009_122, w_009_123, w_009_124, w_009_125, w_009_126, w_009_127, w_009_128, w_009_130, w_009_131, w_009_132, w_009_133, w_009_134, w_009_135, w_009_136, w_009_137, w_009_139, w_009_140, w_009_141, w_009_142, w_009_143, w_009_144, w_009_145, w_009_146, w_009_147, w_009_148, w_009_149, w_009_150, w_009_151, w_009_152, w_009_153, w_009_154, w_009_155, w_009_156, w_009_157, w_009_158, w_009_159, w_009_160, w_009_161, w_009_162, w_009_163, w_009_164, w_009_165, w_009_166, w_009_167, w_009_168, w_009_169, w_009_170, w_009_171, w_009_172, w_009_173, w_009_174, w_009_175, w_009_176, w_009_177, w_009_178, w_009_179, w_009_180, w_009_181, w_009_182, w_009_183, w_009_184, w_009_185, w_009_186, w_009_187, w_009_188, w_009_189, w_009_190, w_009_191, w_009_192, w_009_193, w_009_194, w_009_195, w_009_196, w_009_197, w_009_198, w_009_199, w_009_200, w_009_201, w_009_202, w_009_203, w_009_204, w_009_205, w_009_206, w_009_207, w_009_208, w_009_209, w_009_210, w_009_211, w_009_212, w_009_213, w_009_214, w_009_215, w_009_216, w_009_217, w_009_218, w_009_219, w_009_220, w_009_221, w_009_222, w_009_223, w_009_224, w_009_225, w_009_226, w_009_227, w_009_228, w_009_229, w_009_230, w_009_231, w_009_232, w_009_233, w_009_234, w_009_235, w_009_236, w_009_237, w_009_238, w_009_239, w_009_240, w_009_241, w_009_242, w_009_243, w_009_244, w_009_245, w_009_246, w_009_247, w_009_248, w_009_249, w_009_250, w_009_251, w_009_252, w_009_253, w_009_254, w_009_255, w_009_256, w_009_257, w_009_258, w_009_259, w_009_260, w_009_261, w_009_262, w_009_263, w_009_264, w_009_265, w_009_266, w_009_267, w_009_268, w_009_269, w_009_270, w_009_271, w_009_272, w_009_273, w_009_274, w_009_275, w_009_276, w_009_277, w_009_278, w_009_279, w_009_280, w_009_282, w_009_283, w_009_284, w_009_285, w_009_286, w_009_287, w_009_288, w_009_289, w_009_290, w_009_291, w_009_292, w_009_293, w_009_294, w_009_295, w_009_296, w_009_297, w_009_298, w_009_299, w_009_300, w_009_301, w_009_303, w_009_304, w_009_305, w_009_306, w_009_307, w_009_308, w_009_309, w_009_310, w_009_311, w_009_312, w_009_313, w_009_314, w_009_315, w_009_316, w_009_317, w_009_318, w_009_319, w_009_320, w_009_321, w_009_322, w_009_323, w_009_324, w_009_325, w_009_326, w_009_327, w_009_328, w_009_330, w_009_331, w_009_332, w_009_333, w_009_334, w_009_335, w_009_336, w_009_337, w_009_338, w_009_339, w_009_340, w_009_341, w_009_343, w_009_344, w_009_345, w_009_346, w_009_347, w_009_348, w_009_349, w_009_350, w_009_351, w_009_352, w_009_353, w_009_354, w_009_356, w_009_357, w_009_358, w_009_359, w_009_360, w_009_361, w_009_362, w_009_363, w_009_364, w_009_365, w_009_366, w_009_367, w_009_368, w_009_369, w_009_370, w_009_371, w_009_372, w_009_373, w_009_374, w_009_375, w_009_376, w_009_377, w_009_378, w_009_379, w_009_381, w_009_382, w_009_383, w_009_384, w_009_385, w_009_386, w_009_387, w_009_388, w_009_389, w_009_390, w_009_391, w_009_392, w_009_393, w_009_395, w_009_396, w_009_397, w_009_398, w_009_399, w_009_400, w_009_401, w_009_402, w_009_403, w_009_404, w_009_405, w_009_406, w_009_407, w_009_408, w_009_409, w_009_410, w_009_411, w_009_412, w_009_413, w_009_414, w_009_415, w_009_416, w_009_417, w_009_418, w_009_419, w_009_420, w_009_421, w_009_422, w_009_423, w_009_424, w_009_425, w_009_426, w_009_427, w_009_428, w_009_429, w_009_430, w_009_431, w_009_432, w_009_433, w_009_434, w_009_435, w_009_436, w_009_437, w_009_438, w_009_439, w_009_440, w_009_441, w_009_442, w_009_443, w_009_444, w_009_445, w_009_446, w_009_447, w_009_448, w_009_449, w_009_450, w_009_451, w_009_452, w_009_453, w_009_454, w_009_455, w_009_456, w_009_457, w_009_458, w_009_459, w_009_460, w_009_461, w_009_462, w_009_463, w_009_464, w_009_465, w_009_466, w_009_467, w_009_468, w_009_469, w_009_470, w_009_471, w_009_472, w_009_473, w_009_474, w_009_475, w_009_476, w_009_477, w_009_478, w_009_479, w_009_480, w_009_481, w_009_482, w_009_483, w_009_484, w_009_485, w_009_486, w_009_487, w_009_488, w_009_489, w_009_490, w_009_491, w_009_492, w_009_493, w_009_494, w_009_495, w_009_496, w_009_497, w_009_498, w_009_499, w_009_500, w_009_501, w_009_502, w_009_503, w_009_504, w_009_505, w_009_506, w_009_507, w_009_508, w_009_509, w_009_510, w_009_511, w_009_512, w_009_513, w_009_514, w_009_515, w_009_516, w_009_517, w_009_518, w_009_519, w_009_520, w_009_521, w_009_522, w_009_523, w_009_524, w_009_525, w_009_526, w_009_527, w_009_528, w_009_529, w_009_530, w_009_531, w_009_532, w_009_533, w_009_534, w_009_535, w_009_536, w_009_537, w_009_538, w_009_539, w_009_541, w_009_543, w_009_544, w_009_545, w_009_546, w_009_547, w_009_549, w_009_550, w_009_551, w_009_552, w_009_553, w_009_554, w_009_555, w_009_556, w_009_557, w_009_558, w_009_559, w_009_560, w_009_561, w_009_562, w_009_563, w_009_564, w_009_565, w_009_566, w_009_567, w_009_568, w_009_569, w_009_570, w_009_571, w_009_572, w_009_573, w_009_574, w_009_575, w_009_576, w_009_577, w_009_578, w_009_579, w_009_580, w_009_581, w_009_582, w_009_583, w_009_584, w_009_585, w_009_586, w_009_587, w_009_588, w_009_589, w_009_590, w_009_591, w_009_592, w_009_593, w_009_594, w_009_595, w_009_596, w_009_597, w_009_598, w_009_599, w_009_600, w_009_601, w_009_602, w_009_603, w_009_604, w_009_605, w_009_606, w_009_607, w_009_608, w_009_609, w_009_610, w_009_611, w_009_612, w_009_613, w_009_614, w_009_615, w_009_616, w_009_617, w_009_618, w_009_619, w_009_620, w_009_621, w_009_622, w_009_623, w_009_624, w_009_625, w_009_626, w_009_627, w_009_628, w_009_629, w_009_630, w_009_631, w_009_632, w_009_633, w_009_634, w_009_635, w_009_636, w_009_637, w_009_638, w_009_639, w_009_640, w_009_641, w_009_642, w_009_643, w_009_644, w_009_645, w_009_646, w_009_647, w_009_648, w_009_649, w_009_650, w_009_651, w_009_652, w_009_653, w_009_654, w_009_655, w_009_656, w_009_657, w_009_658, w_009_659, w_009_660, w_009_661, w_009_662, w_009_663, w_009_664, w_009_665, w_009_666, w_009_667, w_009_668, w_009_669, w_009_670, w_009_671, w_009_672, w_009_673, w_009_674, w_009_675, w_009_676, w_009_677, w_009_678, w_009_679, w_009_680, w_009_681, w_009_682, w_009_683, w_009_684, w_009_685, w_009_686, w_009_687, w_009_688, w_009_690, w_009_691, w_009_692, w_009_693, w_009_694, w_009_695, w_009_696, w_009_697, w_009_698, w_009_699, w_009_700, w_009_701, w_009_702, w_009_703, w_009_704, w_009_705, w_009_706, w_009_707, w_009_708, w_009_709, w_009_710, w_009_711, w_009_712, w_009_713, w_009_714, w_009_715, w_009_716, w_009_717, w_009_718, w_009_719, w_009_720, w_009_721, w_009_722, w_009_723, w_009_724, w_009_725, w_009_726, w_009_727, w_009_728, w_009_729, w_009_730, w_009_731, w_009_732, w_009_733, w_009_734, w_009_735, w_009_736, w_009_737, w_009_738, w_009_739, w_009_740, w_009_741, w_009_742, w_009_743, w_009_744, w_009_745, w_009_746, w_009_747, w_009_748, w_009_749, w_009_750, w_009_751, w_009_752, w_009_753, w_009_754, w_009_755, w_009_756, w_009_757, w_009_758, w_009_759, w_009_760, w_009_761, w_009_762, w_009_763, w_009_764, w_009_765, w_009_766, w_009_767, w_009_768, w_009_769, w_009_770, w_009_771, w_009_772, w_009_773, w_009_774, w_009_775, w_009_776, w_009_777, w_009_778, w_009_779, w_009_780, w_009_781, w_009_782, w_009_783, w_009_784, w_009_785, w_009_786, w_009_787, w_009_788, w_009_789, w_009_790, w_009_791, w_009_792, w_009_793, w_009_794, w_009_795, w_009_796, w_009_797, w_009_798, w_009_799, w_009_800, w_009_801, w_009_802, w_009_803, w_009_804, w_009_805, w_009_806, w_009_807, w_009_808, w_009_810, w_009_811, w_009_812, w_009_813, w_009_814, w_009_815, w_009_816, w_009_817, w_009_818, w_009_819, w_009_820, w_009_822, w_009_823, w_009_824, w_009_825, w_009_826, w_009_827, w_009_829, w_009_830, w_009_831, w_009_832, w_009_833, w_009_834, w_009_835, w_009_836, w_009_837, w_009_838, w_009_839, w_009_840, w_009_841, w_009_842, w_009_843, w_009_844, w_009_845, w_009_846, w_009_847, w_009_848, w_009_849, w_009_850, w_009_851, w_009_852, w_009_853, w_009_854, w_009_855, w_009_856, w_009_857, w_009_858, w_009_859, w_009_860, w_009_861, w_009_862, w_009_863, w_009_864, w_009_865, w_009_866, w_009_867, w_009_868, w_009_869, w_009_870, w_009_871, w_009_872, w_009_873, w_009_874, w_009_875, w_009_876, w_009_877, w_009_878, w_009_879, w_009_880, w_009_881, w_009_882, w_009_884, w_009_885, w_009_887, w_009_888, w_009_889, w_009_890, w_009_891, w_009_892, w_009_893, w_009_894, w_009_895, w_009_896, w_009_897, w_009_898, w_009_899, w_009_900, w_009_901, w_009_902, w_009_903, w_009_905, w_009_906, w_009_908, w_009_909, w_009_910, w_009_911, w_009_912, w_009_913, w_009_914, w_009_915, w_009_916, w_009_918, w_009_919, w_009_920, w_009_921, w_009_922, w_009_923, w_009_924, w_009_925, w_009_926, w_009_927, w_009_928, w_009_929, w_009_930, w_009_931, w_009_932, w_009_933, w_009_934, w_009_935, w_009_936, w_009_937, w_009_938, w_009_939, w_009_940, w_009_941, w_009_942, w_009_943, w_009_944, w_009_945, w_009_946, w_009_947, w_009_948, w_009_949, w_009_950, w_009_951, w_009_952, w_009_953, w_009_954, w_009_955, w_009_956, w_009_957, w_009_958, w_009_960, w_009_961, w_009_962, w_009_963, w_009_964, w_009_965, w_009_966, w_009_967, w_009_968, w_009_969, w_009_970, w_009_971, w_009_972, w_009_973, w_009_974, w_009_975, w_009_977, w_009_978, w_009_979, w_009_980, w_009_981, w_009_982, w_009_983, w_009_984, w_009_985, w_009_986, w_009_987, w_009_988, w_009_989, w_009_990, w_009_991, w_009_992, w_009_993, w_009_994, w_009_995, w_009_997, w_009_998, w_009_999, w_009_1000, w_009_1001, w_009_1002, w_009_1003, w_009_1004, w_009_1005, w_009_1006, w_009_1007, w_009_1008, w_009_1009, w_009_1010, w_009_1011, w_009_1012, w_009_1013, w_009_1014, w_009_1015, w_009_1016, w_009_1017, w_009_1018, w_009_1019, w_009_1020, w_009_1021, w_009_1022, w_009_1023, w_009_1024, w_009_1025, w_009_1026, w_009_1027, w_009_1028, w_009_1029, w_009_1030, w_009_1031, w_009_1033, w_009_1034, w_009_1035, w_009_1036, w_009_1037, w_009_1038, w_009_1039, w_009_1040, w_009_1041, w_009_1042, w_009_1043, w_009_1044, w_009_1045, w_009_1046, w_009_1047, w_009_1048, w_009_1049, w_009_1050, w_009_1051, w_009_1052, w_009_1053, w_009_1054, w_009_1055, w_009_1056, w_009_1057, w_009_1058, w_009_1059, w_009_1060, w_009_1061, w_009_1062, w_009_1063, w_009_1064, w_009_1065, w_009_1066, w_009_1067, w_009_1069, w_009_1071, w_009_1072, w_009_1073, w_009_1074, w_009_1075, w_009_1076, w_009_1077, w_009_1078, w_009_1079, w_009_1080, w_009_1081, w_009_1082, w_009_1083, w_009_1084, w_009_1085, w_009_1086, w_009_1087, w_009_1088, w_009_1089, w_009_1090, w_009_1091, w_009_1092, w_009_1093, w_009_1094, w_009_1095, w_009_1096, w_009_1097, w_009_1098, w_009_1099, w_009_1100, w_009_1101, w_009_1102, w_009_1103, w_009_1104, w_009_1105, w_009_1106, w_009_1107, w_009_1108, w_009_1109, w_009_1110, w_009_1111, w_009_1112, w_009_1113, w_009_1114, w_009_1115, w_009_1116, w_009_1117, w_009_1118, w_009_1119, w_009_1120, w_009_1121, w_009_1122, w_009_1123, w_009_1124, w_009_1126, w_009_1127, w_009_1128, w_009_1129, w_009_1130, w_009_1131, w_009_1132, w_009_1133, w_009_1134, w_009_1135, w_009_1136, w_009_1137, w_009_1138, w_009_1139, w_009_1140, w_009_1141, w_009_1142, w_009_1143, w_009_1144, w_009_1145, w_009_1146, w_009_1147, w_009_1148, w_009_1149, w_009_1150, w_009_1151, w_009_1152, w_009_1153, w_009_1154, w_009_1155, w_009_1156, w_009_1157, w_009_1158, w_009_1159, w_009_1160, w_009_1161, w_009_1162, w_009_1163, w_009_1164, w_009_1166, w_009_1167, w_009_1168, w_009_1169, w_009_1170, w_009_1171, w_009_1173, w_009_1174, w_009_1175, w_009_1176, w_009_1177, w_009_1178, w_009_1179, w_009_1180, w_009_1181, w_009_1182, w_009_1183, w_009_1184, w_009_1185, w_009_1186, w_009_1187, w_009_1188, w_009_1189, w_009_1190, w_009_1191, w_009_1192, w_009_1193, w_009_1194, w_009_1195, w_009_1196, w_009_1197, w_009_1199, w_009_1200, w_009_1201, w_009_1202, w_009_1203, w_009_1204, w_009_1205, w_009_1206, w_009_1207, w_009_1208, w_009_1209, w_009_1210, w_009_1211, w_009_1212, w_009_1213, w_009_1214, w_009_1215, w_009_1216, w_009_1217, w_009_1218, w_009_1219, w_009_1220, w_009_1221, w_009_1222, w_009_1223, w_009_1224, w_009_1225, w_009_1226, w_009_1227, w_009_1228, w_009_1229, w_009_1230, w_009_1231, w_009_1232, w_009_1233, w_009_1234, w_009_1235, w_009_1236, w_009_1237, w_009_1238, w_009_1239, w_009_1240, w_009_1241, w_009_1242, w_009_1243, w_009_1244, w_009_1245, w_009_1246, w_009_1248, w_009_1249, w_009_1250, w_009_1251, w_009_1252, w_009_1253, w_009_1254, w_009_1255, w_009_1256, w_009_1257, w_009_1258, w_009_1259, w_009_1260, w_009_1261, w_009_1262, w_009_1263, w_009_1264, w_009_1265, w_009_1266, w_009_1267, w_009_1268, w_009_1269, w_009_1270, w_009_1271, w_009_1272, w_009_1273, w_009_1274, w_009_1275, w_009_1276, w_009_1277, w_009_1278, w_009_1279, w_009_1280, w_009_1281, w_009_1282, w_009_1283, w_009_1284, w_009_1285, w_009_1286, w_009_1287, w_009_1288, w_009_1289, w_009_1291, w_009_1292, w_009_1293, w_009_1294, w_009_1295, w_009_1296, w_009_1297, w_009_1298, w_009_1299, w_009_1300, w_009_1301, w_009_1302, w_009_1303, w_009_1304, w_009_1305, w_009_1306, w_009_1307, w_009_1308, w_009_1309, w_009_1310, w_009_1311, w_009_1312, w_009_1313, w_009_1314, w_009_1315, w_009_1316, w_009_1317, w_009_1318, w_009_1319, w_009_1320, w_009_1321, w_009_1322, w_009_1323, w_009_1324, w_009_1325, w_009_1326, w_009_1327, w_009_1328, w_009_1329, w_009_1330, w_009_1331, w_009_1332, w_009_1333, w_009_1334, w_009_1335, w_009_1336, w_009_1337, w_009_1338, w_009_1339, w_009_1340, w_009_1341, w_009_1342, w_009_1343, w_009_1344, w_009_1345, w_009_1346, w_009_1347, w_009_1348, w_009_1349, w_009_1350, w_009_1351, w_009_1352, w_009_1353, w_009_1354, w_009_1355, w_009_1356, w_009_1357, w_009_1358, w_009_1359, w_009_1360, w_009_1361, w_009_1362, w_009_1363, w_009_1364, w_009_1365, w_009_1366, w_009_1367, w_009_1368, w_009_1369, w_009_1370, w_009_1371, w_009_1372, w_009_1373, w_009_1374, w_009_1375, w_009_1376, w_009_1377, w_009_1378, w_009_1379, w_009_1380, w_009_1381, w_009_1382, w_009_1383, w_009_1384, w_009_1385, w_009_1386, w_009_1387, w_009_1388, w_009_1389, w_009_1390, w_009_1391, w_009_1392, w_009_1393, w_009_1394, w_009_1395, w_009_1396, w_009_1397, w_009_1398, w_009_1399, w_009_1400, w_009_1401, w_009_1403, w_009_1404, w_009_1405, w_009_1406, w_009_1407, w_009_1408, w_009_1409, w_009_1410, w_009_1411, w_009_1412, w_009_1413, w_009_1414, w_009_1415, w_009_1416, w_009_1417, w_009_1418, w_009_1419, w_009_1420, w_009_1421, w_009_1422, w_009_1423, w_009_1424, w_009_1425, w_009_1426, w_009_1427, w_009_1428, w_009_1429, w_009_1430, w_009_1431, w_009_1432, w_009_1433, w_009_1434, w_009_1435, w_009_1436, w_009_1437, w_009_1438, w_009_1439, w_009_1440, w_009_1441, w_009_1442, w_009_1443, w_009_1444, w_009_1445, w_009_1447, w_009_1448, w_009_1449, w_009_1450, w_009_1451, w_009_1452, w_009_1453, w_009_1454, w_009_1455, w_009_1456, w_009_1457, w_009_1458, w_009_1459, w_009_1460, w_009_1461, w_009_1462, w_009_1463, w_009_1464, w_009_1465, w_009_1466, w_009_1467, w_009_1468, w_009_1470, w_009_1472, w_009_1473, w_009_1474, w_009_1475, w_009_1476, w_009_1477, w_009_1478, w_009_1479, w_009_1480, w_009_1481, w_009_1483, w_009_1484, w_009_1485, w_009_1486, w_009_1487, w_009_1488, w_009_1489, w_009_1490, w_009_1491, w_009_1492, w_009_1493, w_009_1494, w_009_1495, w_009_1496, w_009_1497, w_009_1498, w_009_1499, w_009_1500, w_009_1501, w_009_1502, w_009_1503, w_009_1504, w_009_1505, w_009_1506, w_009_1507, w_009_1508, w_009_1509, w_009_1510, w_009_1511, w_009_1513, w_009_1514, w_009_1515, w_009_1516, w_009_1517, w_009_1518, w_009_1519, w_009_1520, w_009_1521, w_009_1522, w_009_1523, w_009_1524, w_009_1525, w_009_1526, w_009_1527, w_009_1528, w_009_1529, w_009_1530, w_009_1531, w_009_1532, w_009_1533, w_009_1534, w_009_1535, w_009_1536, w_009_1537, w_009_1538, w_009_1540, w_009_1541, w_009_1542, w_009_1543, w_009_1544, w_009_1545, w_009_1546, w_009_1547, w_009_1548, w_009_1549, w_009_1550, w_009_1551, w_009_1552, w_009_1553, w_009_1554, w_009_1555, w_009_1556, w_009_1557, w_009_1558, w_009_1559, w_009_1560, w_009_1561, w_009_1562, w_009_1563, w_009_1564, w_009_1565, w_009_1566, w_009_1567, w_009_1568, w_009_1569, w_009_1570, w_009_1572, w_009_1573, w_009_1574, w_009_1575, w_009_1576, w_009_1577, w_009_1578, w_009_1579, w_009_1580, w_009_1581, w_009_1582, w_009_1583, w_009_1584, w_009_1585, w_009_1586, w_009_1587, w_009_1588, w_009_1589, w_009_1590, w_009_1591, w_009_1592, w_009_1593, w_009_1595, w_009_1596, w_009_1597, w_009_1598, w_009_1599, w_009_1600, w_009_1601, w_009_1602, w_009_1603, w_009_1604, w_009_1605, w_009_1606, w_009_1607, w_009_1608, w_009_1609, w_009_1610, w_009_1612, w_009_1613, w_009_1614, w_009_1615, w_009_1616, w_009_1617, w_009_1619, w_009_1620, w_009_1621, w_009_1622, w_009_1623, w_009_1624, w_009_1625, w_009_1626, w_009_1627, w_009_1628, w_009_1629, w_009_1630, w_009_1631, w_009_1632, w_009_1633, w_009_1634, w_009_1635, w_009_1636, w_009_1637, w_009_1638, w_009_1642, w_009_1643, w_009_1644, w_009_1645, w_009_1646, w_009_1647, w_009_1648, w_009_1649, w_009_1650, w_009_1651, w_009_1652, w_009_1653, w_009_1654, w_009_1655, w_009_1656, w_009_1657, w_009_1658, w_009_1659, w_009_1660, w_009_1661, w_009_1662, w_009_1663, w_009_1664, w_009_1665, w_009_1666, w_009_1667, w_009_1668, w_009_1669, w_009_1670, w_009_1671, w_009_1672, w_009_1673, w_009_1674, w_009_1675, w_009_1676, w_009_1677, w_009_1678, w_009_1679, w_009_1680, w_009_1681, w_009_1682, w_009_1683, w_009_1684, w_009_1685, w_009_1686, w_009_1687, w_009_1688, w_009_1689, w_009_1690, w_009_1691, w_009_1692, w_009_1693, w_009_1694, w_009_1695, w_009_1696, w_009_1697, w_009_1698, w_009_1699, w_009_1700, w_009_1701, w_009_1702, w_009_1703, w_009_1704, w_009_1705, w_009_1706, w_009_1707, w_009_1708, w_009_1709, w_009_1710, w_009_1711, w_009_1712, w_009_1713, w_009_1714, w_009_1715, w_009_1716, w_009_1717, w_009_1718, w_009_1719, w_009_1720, w_009_1721, w_009_1722, w_009_1723, w_009_1724, w_009_1725, w_009_1726, w_009_1727, w_009_1728, w_009_1729, w_009_1730, w_009_1731, w_009_1732, w_009_1733, w_009_1734, w_009_1735, w_009_1736, w_009_1737, w_009_1738, w_009_1739, w_009_1740, w_009_1741, w_009_1742, w_009_1743, w_009_1744, w_009_1746, w_009_1747, w_009_1748, w_009_1749, w_009_1750, w_009_1751, w_009_1752, w_009_1753, w_009_1754, w_009_1755, w_009_1756, w_009_1757, w_009_1758, w_009_1759, w_009_1760, w_009_1761, w_009_1762, w_009_1763, w_009_1764, w_009_1765, w_009_1766, w_009_1767, w_009_1768, w_009_1769, w_009_1770, w_009_1771, w_009_1772, w_009_1773, w_009_1774, w_009_1775, w_009_1776, w_009_1777, w_009_1778, w_009_1779, w_009_1780, w_009_1781, w_009_1782, w_009_1783, w_009_1785, w_009_1786, w_009_1787, w_009_1788, w_009_1789, w_009_1790, w_009_1791, w_009_1792, w_009_1793, w_009_1794, w_009_1795, w_009_1796, w_009_1797, w_009_1798, w_009_1799, w_009_1800, w_009_1801, w_009_1802, w_009_1803, w_009_1804, w_009_1805, w_009_1806, w_009_1807, w_009_1808, w_009_1809, w_009_1810, w_009_1811, w_009_1812, w_009_1813, w_009_1814, w_009_1815, w_009_1816, w_009_1817, w_009_1818, w_009_1819, w_009_1820, w_009_1822, w_009_1823, w_009_1824, w_009_1825, w_009_1826, w_009_1827, w_009_1828, w_009_1830, w_009_1831, w_009_1833, w_009_1834, w_009_1835, w_009_1836, w_009_1837, w_009_1838, w_009_1839, w_009_1840, w_009_1841, w_009_1842, w_009_1843, w_009_1844, w_009_1845, w_009_1846, w_009_1847, w_009_1848, w_009_1849, w_009_1850, w_009_1851, w_009_1852, w_009_1853, w_009_1854, w_009_1855, w_009_1856, w_009_1857, w_009_1858, w_009_1859, w_009_1860, w_009_1861, w_009_1862, w_009_1863, w_009_1864, w_009_1865, w_009_1866, w_009_1867, w_009_1868, w_009_1869, w_009_1870, w_009_1871, w_009_1872, w_009_1873, w_009_1874, w_009_1875, w_009_1876, w_009_1878, w_009_1879, w_009_1880, w_009_1881, w_009_1882, w_009_1883, w_009_1884, w_009_1885, w_009_1886, w_009_1887, w_009_1888, w_009_1889, w_009_1890, w_009_1891, w_009_1893, w_009_1894, w_009_1895, w_009_1896, w_009_1897, w_009_1898, w_009_1899, w_009_1900, w_009_1901, w_009_1902, w_009_1903, w_009_1904, w_009_1905, w_009_1906, w_009_1907, w_009_1908, w_009_1909, w_009_1910, w_009_1911, w_009_1912, w_009_1913, w_009_1914, w_009_1915, w_009_1916, w_009_1917, w_009_1918, w_009_1919, w_009_1920, w_009_1921, w_009_1922, w_009_1923, w_009_1924, w_009_1925, w_009_1926, w_009_1927, w_009_1928, w_009_1929, w_009_1930, w_009_1931, w_009_1932, w_009_1933, w_009_1934, w_009_1935, w_009_1936, w_009_1937, w_009_1938, w_009_1939, w_009_1940, w_009_1941, w_009_1942, w_009_1943, w_009_1944, w_009_1945, w_009_1946, w_009_1947, w_009_1948, w_009_1949, w_009_1951, w_009_1952, w_009_1953, w_009_1954, w_009_1955, w_009_1956, w_009_1957, w_009_1958, w_009_1959, w_009_1960, w_009_1961, w_009_1962, w_009_1963, w_009_1964, w_009_1965, w_009_1966, w_009_1967, w_009_1968, w_009_1969, w_009_1970, w_009_1971, w_009_1972, w_009_1973, w_009_1974, w_009_1975, w_009_1976, w_009_1977, w_009_1978, w_009_1979, w_009_1980, w_009_1981, w_009_1982, w_009_1983, w_009_1984, w_009_1985, w_009_1986, w_009_1988, w_009_1989, w_009_1990, w_009_1991, w_009_1992, w_009_1993, w_009_1994, w_009_1995, w_009_1996, w_009_1997, w_009_1998, w_009_1999, w_009_2000, w_009_2001, w_009_2002, w_009_2003, w_009_2004, w_009_2005, w_009_2006, w_009_2007, w_009_2009, w_009_2010, w_009_2011, w_009_2012, w_009_2013, w_009_2014, w_009_2015, w_009_2016, w_009_2017, w_009_2018, w_009_2019, w_009_2020, w_009_2021, w_009_2022, w_009_2023, w_009_2024, w_009_2025, w_009_2026, w_009_2027, w_009_2028, w_009_2029, w_009_2030, w_009_2031, w_009_2032, w_009_2033, w_009_2034, w_009_2035, w_009_2036, w_009_2037, w_009_2038, w_009_2039, w_009_2040, w_009_2041, w_009_2042, w_009_2043, w_009_2045, w_009_2046, w_009_2047, w_009_2048, w_009_2049, w_009_2050, w_009_2051, w_009_2052, w_009_2053, w_009_2054, w_009_2055, w_009_2056, w_009_2057, w_009_2058, w_009_2059, w_009_2060, w_009_2061, w_009_2062, w_009_2063, w_009_2064, w_009_2065, w_009_2066, w_009_2067, w_009_2068, w_009_2069, w_009_2070, w_009_2071, w_009_2072, w_009_2073, w_009_2074, w_009_2075, w_009_2076, w_009_2077, w_009_2078, w_009_2079, w_009_2080, w_009_2081, w_009_2082, w_009_2083, w_009_2084, w_009_2085, w_009_2086, w_009_2087, w_009_2088, w_009_2089, w_009_2090, w_009_2091, w_009_2092, w_009_2093, w_009_2094, w_009_2095, w_009_2096, w_009_2097, w_009_2098, w_009_2099, w_009_2100, w_009_2103, w_009_2104, w_009_2105, w_009_2106, w_009_2107, w_009_2108, w_009_2109, w_009_2110, w_009_2111, w_009_2112, w_009_2113, w_009_2114, w_009_2115, w_009_2116, w_009_2117, w_009_2118, w_009_2119, w_009_2121, w_009_2122, w_009_2123, w_009_2124, w_009_2125, w_009_2127, w_009_2128, w_009_2130, w_009_2131, w_009_2132, w_009_2133, w_009_2134, w_009_2135, w_009_2136, w_009_2137, w_009_2138, w_009_2139, w_009_2140, w_009_2141, w_009_2142, w_009_2143, w_009_2144, w_009_2145, w_009_2146, w_009_2147, w_009_2148, w_009_2149, w_009_2150, w_009_2151, w_009_2152, w_009_2153, w_009_2154, w_009_2155, w_009_2156, w_009_2158, w_009_2159, w_009_2160, w_009_2161, w_009_2162, w_009_2163, w_009_2164, w_009_2165, w_009_2166, w_009_2167, w_009_2168, w_009_2169, w_009_2170, w_009_2171, w_009_2172, w_009_2173, w_009_2174, w_009_2175, w_009_2176, w_009_2177, w_009_2178, w_009_2179, w_009_2180, w_009_2181, w_009_2182, w_009_2183, w_009_2184, w_009_2186, w_009_2187, w_009_2188, w_009_2189, w_009_2190, w_009_2191, w_009_2192, w_009_2193, w_009_2194, w_009_2195, w_009_2196, w_009_2197, w_009_2198, w_009_2199, w_009_2200, w_009_2201, w_009_2202, w_009_2203, w_009_2204, w_009_2205, w_009_2206, w_009_2207, w_009_2208, w_009_2209, w_009_2210, w_009_2211, w_009_2212, w_009_2213, w_009_2214, w_009_2215, w_009_2216, w_009_2217, w_009_2218, w_009_2219, w_009_2220, w_009_2221, w_009_2222, w_009_2223, w_009_2224, w_009_2225, w_009_2226, w_009_2227, w_009_2228, w_009_2229, w_009_2230, w_009_2231, w_009_2232, w_009_2233, w_009_2234, w_009_2235, w_009_2236, w_009_2237, w_009_2238, w_009_2239, w_009_2240, w_009_2241, w_009_2243, w_009_2244, w_009_2245, w_009_2246, w_009_2247, w_009_2248, w_009_2249, w_009_2250, w_009_2252, w_009_2253, w_009_2254, w_009_2255, w_009_2256, w_009_2257, w_009_2258, w_009_2259, w_009_2260, w_009_2261, w_009_2262, w_009_2263, w_009_2264, w_009_2265, w_009_2266, w_009_2267, w_009_2268, w_009_2269, w_009_2270, w_009_2271, w_009_2272, w_009_2273, w_009_2274, w_009_2275, w_009_2276, w_009_2277, w_009_2278, w_009_2279, w_009_2280, w_009_2281, w_009_2282, w_009_2283, w_009_2284, w_009_2285, w_009_2286, w_009_2287, w_009_2288, w_009_2289, w_009_2290, w_009_2291, w_009_2292, w_009_2293, w_009_2294, w_009_2295, w_009_2296, w_009_2297, w_009_2298, w_009_2299, w_009_2300, w_009_2301, w_009_2302, w_009_2303, w_009_2304, w_009_2305, w_009_2306, w_009_2307, w_009_2308, w_009_2309, w_009_2310, w_009_2311, w_009_2312, w_009_2313, w_009_2314, w_009_2315, w_009_2316, w_009_2317, w_009_2318, w_009_2319, w_009_2320, w_009_2321, w_009_2322, w_009_2324, w_009_2325, w_009_2326, w_009_2327, w_009_2328, w_009_2329, w_009_2330, w_009_2331, w_009_2332, w_009_2333, w_009_2334, w_009_2335, w_009_2336, w_009_2337, w_009_2338, w_009_2339, w_009_2340, w_009_2341, w_009_2342, w_009_2344, w_009_2345, w_009_2346, w_009_2347, w_009_2348, w_009_2349, w_009_2350, w_009_2351, w_009_2352, w_009_2353, w_009_2354, w_009_2355, w_009_2356, w_009_2357, w_009_2358, w_009_2359, w_009_2360, w_009_2361, w_009_2362, w_009_2363, w_009_2364, w_009_2365, w_009_2366, w_009_2367, w_009_2369, w_009_2370, w_009_2371, w_009_2372, w_009_2373, w_009_2374, w_009_2375, w_009_2376, w_009_2377, w_009_2378, w_009_2379, w_009_2380, w_009_2381, w_009_2382, w_009_2383, w_009_2384, w_009_2385, w_009_2386, w_009_2387, w_009_2388, w_009_2389, w_009_2390, w_009_2391, w_009_2392, w_009_2393, w_009_2394, w_009_2395, w_009_2396, w_009_2397, w_009_2398, w_009_2399, w_009_2400, w_009_2401, w_009_2402, w_009_2403, w_009_2404, w_009_2405, w_009_2406, w_009_2407, w_009_2408, w_009_2409, w_009_2410, w_009_2411, w_009_2412, w_009_2413, w_009_2414, w_009_2415, w_009_2416, w_009_2417, w_009_2418, w_009_2419, w_009_2421, w_009_2424, w_009_2425, w_009_2426, w_009_2427, w_009_2428, w_009_2429, w_009_2431, w_009_2432, w_009_2436, w_009_2437, w_009_2438, w_009_2439, w_009_2440, w_009_2441, w_009_2443, w_009_2444, w_009_2445, w_009_2446, w_009_2449, w_009_2450, w_009_2451, w_009_2452, w_009_2453, w_009_2454, w_009_2455, w_009_2456, w_009_2457, w_009_2458, w_009_2459, w_009_2460, w_009_2461, w_009_2462, w_009_2463, w_009_2464, w_009_2465, w_009_2466, w_009_2468, w_009_2471, w_009_2472, w_009_2473, w_009_2474, w_009_2475, w_009_2477, w_009_2478, w_009_2479, w_009_2480, w_009_2481, w_009_2482, w_009_2483, w_009_2484, w_009_2486, w_009_2488, w_009_2489, w_009_2490, w_009_2491, w_009_2492, w_009_2493, w_009_2495, w_009_2496, w_009_2497, w_009_2499, w_009_2500, w_009_2501, w_009_2503, w_009_2504, w_009_2505, w_009_2506, w_009_2507, w_009_2508, w_009_2510, w_009_2511, w_009_2512, w_009_2513, w_009_2514, w_009_2515, w_009_2516, w_009_2517, w_009_2518, w_009_2519, w_009_2522, w_009_2523, w_009_2524, w_009_2526, w_009_2527, w_009_2528, w_009_2530, w_009_2531, w_009_2532, w_009_2533, w_009_2534, w_009_2535, w_009_2536, w_009_2537, w_009_2538, w_009_2539, w_009_2540, w_009_2541, w_009_2543, w_009_2545, w_009_2546, w_009_2547, w_009_2548, w_009_2549, w_009_2550, w_009_2552, w_009_2553, w_009_2554, w_009_2555, w_009_2556, w_009_2557, w_009_2558, w_009_2559, w_009_2560, w_009_2561, w_009_2562, w_009_2563, w_009_2564, w_009_2566, w_009_2567, w_009_2568, w_009_2569, w_009_2570, w_009_2572, w_009_2574, w_009_2575, w_009_2576, w_009_2577, w_009_2578, w_009_2579, w_009_2581, w_009_2582, w_009_2583, w_009_2584, w_009_2585, w_009_2586, w_009_2587, w_009_2588, w_009_2590;
  wire w_010_000, w_010_001, w_010_002, w_010_003, w_010_004, w_010_005, w_010_006, w_010_007, w_010_008, w_010_009, w_010_010, w_010_011, w_010_012, w_010_013, w_010_014, w_010_015, w_010_016, w_010_017, w_010_018, w_010_019, w_010_020, w_010_021, w_010_022, w_010_023, w_010_024, w_010_025, w_010_026, w_010_027, w_010_028, w_010_029, w_010_030, w_010_031, w_010_032, w_010_033, w_010_034, w_010_035, w_010_036, w_010_037, w_010_038, w_010_039, w_010_040, w_010_041, w_010_042, w_010_043, w_010_044, w_010_045, w_010_046, w_010_047, w_010_048, w_010_049, w_010_050, w_010_051, w_010_052, w_010_053, w_010_054, w_010_055, w_010_056, w_010_057, w_010_058, w_010_059, w_010_060, w_010_061, w_010_062, w_010_063, w_010_064, w_010_065, w_010_066, w_010_067, w_010_068, w_010_069, w_010_070, w_010_071, w_010_072, w_010_073, w_010_074, w_010_075, w_010_076, w_010_077, w_010_078, w_010_079, w_010_080, w_010_081, w_010_082, w_010_083, w_010_084, w_010_085, w_010_086, w_010_087, w_010_088, w_010_089, w_010_090, w_010_091, w_010_092, w_010_093, w_010_094, w_010_095, w_010_096, w_010_097, w_010_098, w_010_099, w_010_100, w_010_101, w_010_102, w_010_103, w_010_104, w_010_105, w_010_106, w_010_107, w_010_108, w_010_109, w_010_110, w_010_111, w_010_112, w_010_113, w_010_114, w_010_115, w_010_116, w_010_117, w_010_118, w_010_119, w_010_120, w_010_121, w_010_122, w_010_123, w_010_124, w_010_125, w_010_126, w_010_127, w_010_128, w_010_129, w_010_130, w_010_131, w_010_132, w_010_133, w_010_134, w_010_135, w_010_136, w_010_137, w_010_138, w_010_139, w_010_140, w_010_141, w_010_142, w_010_143, w_010_144, w_010_145, w_010_146, w_010_147, w_010_148, w_010_149, w_010_150, w_010_151, w_010_152, w_010_153, w_010_154, w_010_155, w_010_156, w_010_157, w_010_158, w_010_159, w_010_160, w_010_161, w_010_162, w_010_163, w_010_164, w_010_165, w_010_166, w_010_167, w_010_168, w_010_169, w_010_170, w_010_171, w_010_172, w_010_173, w_010_174, w_010_175, w_010_176, w_010_177, w_010_178, w_010_179, w_010_180, w_010_181, w_010_182, w_010_183, w_010_184, w_010_185, w_010_186, w_010_187, w_010_188, w_010_189, w_010_190, w_010_191, w_010_192, w_010_193, w_010_194, w_010_195, w_010_196, w_010_197, w_010_198, w_010_199, w_010_200, w_010_201, w_010_202, w_010_203, w_010_204, w_010_205, w_010_206, w_010_207, w_010_208, w_010_209, w_010_210, w_010_211, w_010_212, w_010_213, w_010_214, w_010_215, w_010_216, w_010_217, w_010_218, w_010_219, w_010_220, w_010_221, w_010_222, w_010_223, w_010_224, w_010_225, w_010_226, w_010_227, w_010_228, w_010_229, w_010_230, w_010_231, w_010_232, w_010_233, w_010_234, w_010_235, w_010_236, w_010_237, w_010_238, w_010_239, w_010_240, w_010_241, w_010_242, w_010_243, w_010_244, w_010_245, w_010_246, w_010_247, w_010_248, w_010_249, w_010_250, w_010_251, w_010_252, w_010_253, w_010_254, w_010_255, w_010_256, w_010_257, w_010_258, w_010_259, w_010_260, w_010_261, w_010_262, w_010_263, w_010_264, w_010_265, w_010_266, w_010_267, w_010_268, w_010_269, w_010_270, w_010_271, w_010_272, w_010_273, w_010_274, w_010_275, w_010_276, w_010_277, w_010_278, w_010_279, w_010_280, w_010_281, w_010_282, w_010_283, w_010_284, w_010_285, w_010_286, w_010_287, w_010_288, w_010_289, w_010_290, w_010_291, w_010_292, w_010_293, w_010_294, w_010_295, w_010_296, w_010_297, w_010_298, w_010_299, w_010_300, w_010_301, w_010_302, w_010_303, w_010_304, w_010_305, w_010_306, w_010_307, w_010_308, w_010_309, w_010_310, w_010_311, w_010_312, w_010_313, w_010_314, w_010_315, w_010_316, w_010_317, w_010_318, w_010_319, w_010_320, w_010_321, w_010_322, w_010_323, w_010_324, w_010_325, w_010_326, w_010_327, w_010_328, w_010_329, w_010_330, w_010_331, w_010_332, w_010_333, w_010_334, w_010_335, w_010_336, w_010_337, w_010_338, w_010_339, w_010_340, w_010_341, w_010_342, w_010_343, w_010_344, w_010_345, w_010_346, w_010_347, w_010_348, w_010_349, w_010_350, w_010_351, w_010_352, w_010_353, w_010_354, w_010_355, w_010_356, w_010_357, w_010_358, w_010_359, w_010_360, w_010_361, w_010_362, w_010_363, w_010_364, w_010_365, w_010_366, w_010_367, w_010_368, w_010_369, w_010_370, w_010_371, w_010_372, w_010_373, w_010_374, w_010_375, w_010_376, w_010_377, w_010_378, w_010_379, w_010_380, w_010_381, w_010_382, w_010_383, w_010_384, w_010_385, w_010_386, w_010_387, w_010_388, w_010_389, w_010_390, w_010_391, w_010_392, w_010_393, w_010_394, w_010_395, w_010_396, w_010_397, w_010_398, w_010_399, w_010_400, w_010_401, w_010_402, w_010_403, w_010_404, w_010_405, w_010_406, w_010_407, w_010_408, w_010_409, w_010_410, w_010_411, w_010_412, w_010_413, w_010_414, w_010_415, w_010_416, w_010_417, w_010_418, w_010_419, w_010_420, w_010_421, w_010_422, w_010_423, w_010_424, w_010_425, w_010_426, w_010_427, w_010_428, w_010_429, w_010_430, w_010_431, w_010_432, w_010_433, w_010_434, w_010_435, w_010_436, w_010_437, w_010_438, w_010_439, w_010_440, w_010_441, w_010_442, w_010_443, w_010_444, w_010_445, w_010_446, w_010_447, w_010_448, w_010_449, w_010_450, w_010_451, w_010_452, w_010_453, w_010_454, w_010_455, w_010_456, w_010_457, w_010_458, w_010_459, w_010_460, w_010_461, w_010_462, w_010_463, w_010_464, w_010_465, w_010_466, w_010_467, w_010_468, w_010_469, w_010_470, w_010_471, w_010_472, w_010_473, w_010_474, w_010_475, w_010_476, w_010_477, w_010_478, w_010_479, w_010_480, w_010_481, w_010_482, w_010_483, w_010_484, w_010_485, w_010_486, w_010_487, w_010_488, w_010_489, w_010_490, w_010_491, w_010_492, w_010_493, w_010_494, w_010_495, w_010_496, w_010_497, w_010_498, w_010_499, w_010_500, w_010_501, w_010_502, w_010_503, w_010_504, w_010_505, w_010_506, w_010_507, w_010_508, w_010_509, w_010_510, w_010_511, w_010_512, w_010_513, w_010_514, w_010_515, w_010_516, w_010_517, w_010_518, w_010_519, w_010_520, w_010_521, w_010_522, w_010_523, w_010_524, w_010_525, w_010_526, w_010_527, w_010_528, w_010_529, w_010_530, w_010_531, w_010_532, w_010_533, w_010_534, w_010_535, w_010_536, w_010_537, w_010_538, w_010_539, w_010_540, w_010_541, w_010_542, w_010_543, w_010_544, w_010_545, w_010_546, w_010_547, w_010_548, w_010_549, w_010_550, w_010_551, w_010_552, w_010_553, w_010_554, w_010_555, w_010_556, w_010_557, w_010_558, w_010_559, w_010_560, w_010_561, w_010_562, w_010_563, w_010_564, w_010_565, w_010_566, w_010_567, w_010_568, w_010_569, w_010_570, w_010_571, w_010_572, w_010_573, w_010_574, w_010_575, w_010_576, w_010_577, w_010_578, w_010_579, w_010_580, w_010_581, w_010_582, w_010_583, w_010_584, w_010_585, w_010_586, w_010_587, w_010_588, w_010_589, w_010_590, w_010_591, w_010_592, w_010_593, w_010_594, w_010_595, w_010_596, w_010_597, w_010_598, w_010_599, w_010_600, w_010_601, w_010_602, w_010_603, w_010_604, w_010_605, w_010_606, w_010_607, w_010_608, w_010_609, w_010_610, w_010_611, w_010_612, w_010_613, w_010_614, w_010_615, w_010_616, w_010_617, w_010_618, w_010_619, w_010_620, w_010_621, w_010_622, w_010_623, w_010_624, w_010_625, w_010_626, w_010_627, w_010_628, w_010_629, w_010_630, w_010_631, w_010_632, w_010_633, w_010_634, w_010_635, w_010_636, w_010_637, w_010_638, w_010_639, w_010_640, w_010_641, w_010_642, w_010_643, w_010_644, w_010_645, w_010_646, w_010_647, w_010_648, w_010_649, w_010_650, w_010_651, w_010_652, w_010_653, w_010_654, w_010_655, w_010_656, w_010_657;
  wire w_011_000, w_011_001, w_011_002, w_011_003, w_011_004, w_011_005, w_011_006, w_011_007, w_011_008, w_011_009, w_011_010, w_011_011, w_011_012, w_011_013, w_011_014, w_011_015, w_011_016, w_011_017, w_011_018, w_011_019, w_011_020, w_011_021, w_011_022, w_011_023, w_011_024, w_011_025, w_011_026, w_011_027, w_011_028, w_011_029, w_011_030, w_011_031, w_011_032, w_011_033, w_011_034, w_011_035, w_011_036, w_011_037, w_011_038, w_011_039, w_011_040, w_011_041, w_011_042, w_011_043, w_011_044, w_011_045, w_011_046, w_011_047, w_011_048, w_011_049, w_011_050, w_011_051, w_011_052, w_011_053, w_011_054, w_011_055, w_011_056, w_011_057, w_011_059, w_011_060, w_011_061, w_011_062, w_011_063, w_011_064, w_011_065, w_011_066, w_011_067, w_011_069, w_011_070, w_011_071, w_011_072, w_011_073, w_011_074, w_011_075, w_011_076, w_011_077, w_011_078, w_011_079, w_011_080, w_011_081, w_011_082, w_011_083, w_011_084, w_011_085, w_011_086, w_011_087, w_011_088, w_011_089, w_011_090, w_011_091, w_011_092, w_011_093, w_011_094, w_011_095, w_011_096, w_011_097, w_011_098, w_011_099, w_011_100, w_011_101, w_011_102, w_011_103, w_011_104, w_011_105, w_011_106, w_011_107, w_011_108, w_011_109, w_011_110, w_011_111, w_011_112, w_011_113, w_011_114, w_011_115, w_011_117, w_011_118, w_011_119, w_011_120, w_011_121, w_011_122, w_011_123, w_011_124, w_011_125, w_011_126, w_011_127, w_011_128, w_011_129, w_011_130, w_011_131, w_011_132, w_011_133, w_011_134, w_011_136, w_011_137, w_011_138, w_011_139, w_011_140, w_011_141, w_011_142, w_011_143, w_011_144, w_011_145, w_011_146, w_011_147, w_011_148, w_011_149, w_011_150, w_011_151, w_011_152, w_011_153, w_011_154, w_011_155, w_011_156, w_011_157, w_011_158, w_011_159, w_011_160, w_011_161, w_011_162, w_011_163, w_011_164, w_011_165, w_011_166, w_011_167, w_011_168, w_011_169, w_011_170, w_011_171, w_011_172, w_011_173, w_011_174, w_011_175, w_011_176, w_011_177, w_011_178, w_011_179, w_011_180, w_011_181, w_011_182, w_011_183, w_011_184, w_011_185, w_011_186, w_011_187, w_011_188, w_011_189, w_011_190, w_011_191, w_011_192, w_011_193, w_011_194, w_011_195, w_011_196, w_011_197, w_011_198, w_011_199, w_011_200, w_011_201, w_011_202, w_011_203, w_011_204, w_011_205, w_011_206, w_011_207, w_011_208, w_011_209, w_011_210, w_011_211, w_011_212, w_011_213, w_011_214, w_011_215, w_011_216, w_011_217, w_011_218, w_011_219, w_011_220, w_011_221, w_011_222, w_011_223, w_011_224, w_011_225, w_011_226, w_011_227, w_011_228, w_011_229, w_011_230, w_011_231, w_011_232, w_011_233, w_011_234, w_011_235, w_011_236, w_011_237, w_011_238, w_011_239, w_011_240, w_011_241, w_011_242, w_011_243, w_011_244, w_011_245, w_011_246, w_011_247, w_011_248, w_011_249, w_011_250, w_011_251, w_011_252, w_011_253, w_011_255, w_011_256, w_011_257, w_011_258, w_011_259, w_011_260, w_011_261, w_011_262, w_011_263, w_011_264, w_011_265, w_011_266, w_011_267, w_011_268, w_011_269, w_011_270, w_011_271, w_011_272, w_011_273, w_011_274, w_011_275, w_011_276, w_011_277, w_011_278, w_011_279, w_011_280, w_011_281, w_011_282, w_011_283, w_011_284, w_011_285, w_011_286, w_011_287, w_011_288, w_011_289, w_011_290, w_011_291, w_011_292, w_011_293, w_011_294, w_011_295, w_011_296, w_011_297, w_011_298, w_011_299, w_011_300, w_011_301, w_011_302, w_011_303, w_011_304, w_011_305, w_011_306, w_011_307, w_011_308, w_011_309, w_011_310, w_011_311, w_011_312, w_011_313, w_011_314, w_011_315, w_011_316, w_011_317, w_011_318, w_011_319, w_011_320, w_011_321, w_011_322, w_011_323, w_011_324, w_011_325, w_011_326, w_011_327, w_011_328, w_011_329, w_011_330, w_011_331, w_011_332, w_011_333, w_011_334, w_011_335, w_011_336, w_011_337, w_011_338, w_011_339, w_011_340, w_011_341, w_011_342, w_011_343, w_011_344, w_011_345, w_011_346, w_011_347, w_011_348, w_011_349, w_011_350, w_011_351, w_011_352, w_011_353, w_011_354, w_011_355, w_011_356, w_011_357, w_011_358, w_011_359, w_011_360, w_011_361, w_011_362, w_011_363, w_011_364, w_011_365, w_011_366, w_011_367, w_011_368, w_011_369, w_011_370, w_011_371, w_011_372, w_011_374, w_011_375, w_011_376, w_011_377, w_011_378, w_011_379, w_011_380, w_011_381, w_011_382, w_011_383, w_011_384, w_011_385, w_011_386, w_011_387, w_011_388, w_011_389, w_011_391, w_011_392, w_011_393, w_011_394, w_011_395, w_011_397, w_011_398, w_011_399, w_011_400, w_011_401, w_011_402, w_011_403, w_011_404, w_011_405, w_011_406, w_011_407, w_011_408, w_011_409, w_011_410, w_011_411, w_011_412, w_011_413, w_011_414, w_011_415, w_011_416, w_011_417, w_011_418, w_011_419, w_011_420, w_011_421, w_011_422, w_011_423, w_011_424, w_011_425, w_011_426, w_011_427, w_011_428, w_011_429, w_011_430, w_011_431, w_011_432, w_011_433, w_011_434, w_011_435, w_011_436, w_011_437, w_011_438, w_011_439, w_011_440, w_011_441, w_011_442, w_011_443, w_011_444, w_011_445, w_011_446, w_011_447, w_011_448, w_011_449, w_011_450, w_011_451, w_011_452, w_011_453, w_011_454, w_011_455, w_011_456, w_011_457, w_011_458, w_011_459, w_011_460, w_011_461, w_011_462, w_011_463, w_011_464, w_011_465, w_011_466, w_011_467, w_011_468, w_011_469, w_011_471, w_011_472, w_011_473, w_011_474, w_011_475, w_011_476, w_011_477, w_011_478, w_011_479, w_011_480, w_011_481, w_011_482, w_011_483, w_011_484, w_011_485, w_011_486, w_011_487, w_011_488, w_011_489, w_011_490, w_011_491, w_011_492, w_011_493, w_011_495, w_011_496, w_011_497, w_011_498, w_011_499, w_011_500, w_011_501, w_011_502, w_011_503, w_011_504, w_011_505, w_011_506, w_011_507, w_011_508, w_011_509, w_011_510, w_011_511, w_011_512, w_011_514, w_011_515, w_011_516, w_011_517, w_011_518, w_011_519, w_011_520, w_011_521, w_011_522, w_011_523, w_011_524, w_011_525, w_011_526, w_011_527, w_011_528, w_011_529, w_011_530, w_011_531, w_011_532, w_011_533, w_011_534, w_011_535, w_011_536, w_011_537, w_011_538, w_011_539, w_011_540, w_011_541, w_011_543, w_011_544, w_011_545, w_011_546, w_011_547, w_011_548, w_011_549, w_011_550, w_011_551, w_011_552, w_011_553, w_011_555, w_011_556, w_011_557, w_011_558, w_011_559, w_011_560, w_011_561, w_011_562, w_011_563, w_011_564, w_011_565, w_011_566, w_011_567, w_011_568, w_011_569, w_011_570, w_011_571, w_011_572, w_011_573, w_011_574, w_011_575, w_011_576, w_011_577, w_011_578, w_011_579, w_011_580, w_011_581, w_011_582, w_011_583, w_011_584, w_011_585, w_011_586, w_011_587, w_011_588, w_011_589, w_011_590, w_011_591, w_011_592, w_011_593, w_011_594, w_011_595, w_011_596, w_011_597, w_011_598, w_011_599, w_011_600, w_011_601, w_011_602, w_011_603, w_011_604, w_011_605, w_011_606, w_011_608, w_011_609, w_011_610, w_011_611, w_011_612, w_011_613, w_011_614, w_011_615, w_011_616, w_011_617, w_011_618, w_011_619, w_011_620, w_011_621, w_011_622, w_011_623, w_011_624, w_011_625, w_011_626, w_011_627, w_011_628, w_011_630, w_011_632, w_011_633, w_011_634, w_011_635, w_011_636, w_011_637, w_011_638, w_011_639, w_011_640, w_011_641, w_011_642, w_011_643, w_011_644, w_011_645, w_011_646, w_011_647, w_011_648, w_011_649, w_011_650, w_011_651, w_011_652, w_011_653, w_011_654, w_011_655, w_011_656, w_011_657, w_011_658, w_011_659, w_011_660, w_011_661, w_011_662, w_011_663, w_011_664, w_011_665, w_011_666, w_011_667, w_011_668, w_011_669, w_011_670, w_011_671, w_011_672, w_011_673, w_011_674, w_011_675, w_011_676, w_011_677, w_011_678, w_011_679, w_011_680, w_011_681, w_011_682, w_011_683, w_011_684, w_011_685, w_011_686, w_011_687, w_011_688, w_011_689, w_011_690, w_011_691, w_011_692, w_011_693, w_011_694, w_011_695, w_011_696, w_011_697, w_011_698, w_011_699, w_011_700, w_011_701, w_011_702, w_011_703, w_011_704, w_011_705, w_011_706, w_011_707, w_011_709, w_011_710, w_011_711, w_011_712, w_011_713, w_011_714, w_011_715, w_011_716, w_011_717, w_011_718, w_011_719, w_011_720, w_011_721, w_011_722, w_011_723, w_011_724, w_011_725, w_011_726, w_011_727, w_011_728, w_011_729, w_011_730, w_011_731, w_011_732, w_011_733, w_011_734, w_011_735, w_011_736, w_011_737, w_011_738, w_011_739, w_011_740, w_011_741, w_011_742, w_011_743, w_011_744, w_011_745, w_011_746, w_011_747, w_011_748, w_011_749, w_011_750, w_011_751, w_011_752, w_011_753, w_011_754, w_011_755, w_011_756, w_011_757, w_011_758, w_011_759, w_011_760, w_011_762, w_011_763, w_011_764, w_011_765, w_011_766, w_011_767, w_011_768, w_011_769, w_011_770, w_011_771, w_011_772, w_011_773, w_011_774, w_011_775, w_011_776, w_011_777, w_011_778, w_011_779, w_011_780, w_011_781, w_011_782, w_011_783, w_011_784, w_011_785, w_011_786, w_011_787, w_011_788, w_011_789, w_011_790, w_011_791, w_011_792, w_011_793, w_011_795, w_011_796, w_011_797, w_011_798, w_011_799, w_011_800, w_011_801, w_011_802, w_011_803, w_011_804, w_011_805, w_011_806, w_011_807, w_011_808, w_011_809, w_011_810, w_011_812, w_011_813, w_011_814, w_011_815, w_011_816, w_011_817, w_011_818, w_011_819, w_011_820, w_011_821, w_011_822, w_011_823, w_011_824, w_011_825, w_011_826, w_011_827, w_011_828, w_011_829, w_011_831, w_011_832, w_011_833, w_011_834, w_011_835, w_011_836, w_011_837, w_011_838, w_011_839, w_011_840, w_011_841, w_011_842, w_011_843, w_011_844, w_011_845, w_011_846, w_011_847, w_011_848, w_011_849, w_011_850, w_011_851, w_011_852, w_011_853, w_011_854, w_011_855, w_011_856, w_011_857, w_011_858, w_011_859, w_011_860, w_011_861, w_011_862, w_011_863, w_011_864, w_011_865, w_011_866, w_011_867, w_011_869, w_011_870, w_011_871, w_011_872, w_011_873, w_011_874, w_011_875, w_011_876, w_011_877, w_011_879, w_011_880, w_011_882, w_011_883, w_011_884, w_011_885, w_011_886, w_011_887, w_011_888, w_011_889, w_011_890, w_011_891, w_011_892, w_011_893, w_011_894, w_011_896, w_011_899, w_011_900, w_011_901, w_011_902, w_011_903, w_011_904, w_011_905, w_011_906, w_011_907, w_011_908, w_011_910, w_011_911, w_011_912, w_011_913, w_011_914, w_011_915, w_011_916, w_011_917, w_011_918, w_011_919, w_011_920, w_011_921, w_011_922, w_011_923, w_011_924, w_011_925, w_011_926, w_011_927, w_011_928, w_011_929, w_011_930, w_011_931, w_011_932, w_011_933, w_011_934, w_011_935, w_011_936, w_011_937, w_011_938, w_011_939, w_011_940, w_011_941, w_011_942, w_011_943, w_011_944, w_011_945, w_011_946, w_011_947, w_011_948, w_011_949, w_011_950, w_011_951, w_011_952, w_011_953, w_011_954, w_011_955, w_011_956, w_011_957, w_011_958, w_011_959, w_011_960, w_011_961, w_011_962, w_011_963, w_011_964, w_011_965, w_011_967, w_011_968, w_011_969, w_011_970, w_011_971, w_011_972, w_011_973, w_011_974, w_011_975, w_011_976, w_011_977, w_011_978, w_011_979, w_011_980, w_011_981, w_011_982, w_011_983, w_011_984, w_011_985, w_011_986, w_011_987, w_011_988, w_011_989, w_011_990, w_011_991, w_011_992, w_011_993, w_011_994, w_011_995, w_011_996, w_011_997, w_011_998, w_011_999, w_011_1000, w_011_1001, w_011_1002, w_011_1003, w_011_1004, w_011_1005, w_011_1006, w_011_1007, w_011_1008, w_011_1010, w_011_1011, w_011_1012, w_011_1013, w_011_1014, w_011_1015, w_011_1016, w_011_1017, w_011_1018, w_011_1019, w_011_1020, w_011_1021, w_011_1022, w_011_1023, w_011_1024, w_011_1025, w_011_1026, w_011_1027, w_011_1028, w_011_1029, w_011_1030, w_011_1031, w_011_1033, w_011_1034, w_011_1035, w_011_1036, w_011_1037, w_011_1038, w_011_1039, w_011_1040, w_011_1041, w_011_1042, w_011_1043, w_011_1044, w_011_1045, w_011_1046, w_011_1047, w_011_1048, w_011_1049, w_011_1051, w_011_1053, w_011_1054, w_011_1055, w_011_1056, w_011_1057, w_011_1058, w_011_1059, w_011_1060, w_011_1061, w_011_1062, w_011_1063, w_011_1064, w_011_1065, w_011_1066, w_011_1067, w_011_1068, w_011_1069, w_011_1070, w_011_1072, w_011_1073, w_011_1074, w_011_1075, w_011_1076, w_011_1077, w_011_1078, w_011_1079, w_011_1080, w_011_1081, w_011_1082, w_011_1083, w_011_1084, w_011_1085, w_011_1086, w_011_1087, w_011_1088, w_011_1089, w_011_1090, w_011_1091, w_011_1092, w_011_1093, w_011_1094, w_011_1095, w_011_1096, w_011_1097, w_011_1098, w_011_1099, w_011_1100, w_011_1101, w_011_1103, w_011_1105, w_011_1106, w_011_1107, w_011_1108, w_011_1109, w_011_1110, w_011_1111, w_011_1112, w_011_1113, w_011_1114, w_011_1115, w_011_1117, w_011_1118, w_011_1119, w_011_1120, w_011_1121, w_011_1122, w_011_1123, w_011_1124, w_011_1126, w_011_1127, w_011_1128, w_011_1130, w_011_1131, w_011_1132, w_011_1133, w_011_1134, w_011_1135, w_011_1136, w_011_1137, w_011_1138, w_011_1139, w_011_1140, w_011_1141, w_011_1142, w_011_1143, w_011_1144, w_011_1145, w_011_1146, w_011_1147, w_011_1149, w_011_1150, w_011_1151, w_011_1152, w_011_1153, w_011_1154, w_011_1155, w_011_1156, w_011_1157, w_011_1158, w_011_1159, w_011_1160, w_011_1161, w_011_1162, w_011_1163, w_011_1164, w_011_1165, w_011_1166, w_011_1167, w_011_1168, w_011_1170, w_011_1171, w_011_1172, w_011_1173, w_011_1174, w_011_1175, w_011_1177, w_011_1178, w_011_1179, w_011_1180, w_011_1181, w_011_1182, w_011_1183, w_011_1184, w_011_1185, w_011_1186, w_011_1187, w_011_1188, w_011_1189, w_011_1190, w_011_1191, w_011_1192, w_011_1193, w_011_1194, w_011_1195, w_011_1196, w_011_1197, w_011_1198, w_011_1199, w_011_1200, w_011_1202, w_011_1203, w_011_1204, w_011_1205, w_011_1206, w_011_1207, w_011_1208, w_011_1209, w_011_1210, w_011_1211, w_011_1212, w_011_1213, w_011_1214, w_011_1215, w_011_1216, w_011_1217, w_011_1218, w_011_1219, w_011_1220, w_011_1221, w_011_1223, w_011_1224, w_011_1225, w_011_1226, w_011_1227, w_011_1228, w_011_1229, w_011_1230, w_011_1231, w_011_1232, w_011_1233, w_011_1234, w_011_1235, w_011_1236, w_011_1237, w_011_1238, w_011_1239, w_011_1240, w_011_1241, w_011_1242, w_011_1243, w_011_1244, w_011_1245, w_011_1246, w_011_1247, w_011_1248, w_011_1249, w_011_1250, w_011_1251, w_011_1252, w_011_1253, w_011_1254, w_011_1255, w_011_1256, w_011_1257, w_011_1258, w_011_1259, w_011_1260, w_011_1261, w_011_1262, w_011_1263, w_011_1264, w_011_1265, w_011_1266, w_011_1267, w_011_1268, w_011_1269, w_011_1270, w_011_1271, w_011_1272, w_011_1273, w_011_1274, w_011_1275, w_011_1276, w_011_1277, w_011_1278, w_011_1279, w_011_1280, w_011_1281, w_011_1282, w_011_1283, w_011_1284, w_011_1285, w_011_1286, w_011_1287, w_011_1288, w_011_1289, w_011_1291, w_011_1292, w_011_1293, w_011_1294, w_011_1295, w_011_1296, w_011_1297, w_011_1298, w_011_1299, w_011_1300, w_011_1301, w_011_1303, w_011_1304, w_011_1305, w_011_1306, w_011_1307, w_011_1308, w_011_1309, w_011_1310, w_011_1311, w_011_1312, w_011_1313, w_011_1314, w_011_1315, w_011_1316, w_011_1317, w_011_1318, w_011_1319, w_011_1320, w_011_1321, w_011_1322, w_011_1323, w_011_1324, w_011_1325, w_011_1326, w_011_1327, w_011_1328, w_011_1329, w_011_1330, w_011_1331, w_011_1332, w_011_1333, w_011_1334, w_011_1335, w_011_1336, w_011_1337, w_011_1338, w_011_1339, w_011_1340, w_011_1341, w_011_1342, w_011_1343, w_011_1344, w_011_1345, w_011_1346, w_011_1347, w_011_1348, w_011_1349, w_011_1350, w_011_1351, w_011_1352, w_011_1353, w_011_1354, w_011_1355, w_011_1356, w_011_1357, w_011_1358, w_011_1359, w_011_1360, w_011_1361, w_011_1362, w_011_1363, w_011_1364, w_011_1365, w_011_1366, w_011_1367, w_011_1368, w_011_1369, w_011_1370, w_011_1371, w_011_1372, w_011_1373, w_011_1374, w_011_1375, w_011_1376, w_011_1377, w_011_1378, w_011_1379, w_011_1380, w_011_1381, w_011_1382, w_011_1383, w_011_1384, w_011_1385, w_011_1386, w_011_1387, w_011_1388, w_011_1389, w_011_1390, w_011_1392, w_011_1393, w_011_1394, w_011_1395, w_011_1396, w_011_1397, w_011_1398, w_011_1399, w_011_1400, w_011_1401, w_011_1402, w_011_1403, w_011_1404, w_011_1405, w_011_1406, w_011_1408, w_011_1409, w_011_1410, w_011_1411, w_011_1412, w_011_1413, w_011_1414, w_011_1415, w_011_1416, w_011_1417, w_011_1418, w_011_1419, w_011_1420, w_011_1421, w_011_1422, w_011_1423, w_011_1424, w_011_1425, w_011_1426, w_011_1427, w_011_1428, w_011_1429, w_011_1430, w_011_1431, w_011_1432, w_011_1433, w_011_1434, w_011_1435, w_011_1436, w_011_1437, w_011_1438, w_011_1439, w_011_1440, w_011_1441, w_011_1442, w_011_1443, w_011_1444, w_011_1445, w_011_1446, w_011_1447, w_011_1448, w_011_1449, w_011_1450, w_011_1451, w_011_1452, w_011_1453, w_011_1454, w_011_1455, w_011_1456, w_011_1457, w_011_1458, w_011_1459, w_011_1460, w_011_1461, w_011_1462, w_011_1463, w_011_1464, w_011_1465, w_011_1466, w_011_1467, w_011_1468, w_011_1469, w_011_1470, w_011_1471, w_011_1472, w_011_1473, w_011_1474, w_011_1475, w_011_1476, w_011_1477, w_011_1478, w_011_1479, w_011_1480, w_011_1481, w_011_1482, w_011_1483, w_011_1484, w_011_1485, w_011_1486, w_011_1487, w_011_1488, w_011_1489, w_011_1490, w_011_1491, w_011_1492, w_011_1493, w_011_1494, w_011_1495, w_011_1496, w_011_1497, w_011_1498, w_011_1499, w_011_1500, w_011_1501, w_011_1502, w_011_1503, w_011_1504, w_011_1505, w_011_1506, w_011_1508, w_011_1509, w_011_1510, w_011_1511, w_011_1512, w_011_1513, w_011_1514, w_011_1515, w_011_1516, w_011_1517, w_011_1518, w_011_1519, w_011_1520, w_011_1521, w_011_1522, w_011_1523, w_011_1524, w_011_1525, w_011_1526, w_011_1527, w_011_1528, w_011_1529, w_011_1530, w_011_1531, w_011_1532, w_011_1533, w_011_1534, w_011_1535, w_011_1536, w_011_1537, w_011_1538, w_011_1539, w_011_1541, w_011_1542, w_011_1543, w_011_1544, w_011_1545, w_011_1546, w_011_1547, w_011_1548, w_011_1549, w_011_1550, w_011_1551, w_011_1552, w_011_1553, w_011_1554, w_011_1555, w_011_1556, w_011_1557, w_011_1558, w_011_1559, w_011_1562, w_011_1563, w_011_1564, w_011_1565, w_011_1566, w_011_1567, w_011_1569, w_011_1570, w_011_1571, w_011_1572, w_011_1573, w_011_1574, w_011_1575, w_011_1576, w_011_1577, w_011_1578, w_011_1579, w_011_1580, w_011_1581, w_011_1582, w_011_1583, w_011_1584, w_011_1585, w_011_1586, w_011_1587, w_011_1588, w_011_1589, w_011_1590, w_011_1591, w_011_1592, w_011_1593, w_011_1594, w_011_1595, w_011_1596, w_011_1597, w_011_1598, w_011_1599, w_011_1600, w_011_1601, w_011_1602, w_011_1603, w_011_1604, w_011_1605, w_011_1606, w_011_1607, w_011_1608, w_011_1609, w_011_1611, w_011_1612, w_011_1613, w_011_1614, w_011_1616, w_011_1617, w_011_1618, w_011_1619, w_011_1620, w_011_1621, w_011_1622, w_011_1623, w_011_1624, w_011_1625, w_011_1626, w_011_1627, w_011_1628, w_011_1629, w_011_1630, w_011_1631, w_011_1632, w_011_1634, w_011_1635, w_011_1636, w_011_1637, w_011_1638, w_011_1639, w_011_1640, w_011_1641, w_011_1642, w_011_1643, w_011_1644, w_011_1645, w_011_1646, w_011_1647, w_011_1648, w_011_1649, w_011_1650, w_011_1651, w_011_1652, w_011_1653, w_011_1654, w_011_1655, w_011_1656, w_011_1657, w_011_1659, w_011_1660, w_011_1661, w_011_1662, w_011_1663, w_011_1664, w_011_1665, w_011_1666, w_011_1667, w_011_1668, w_011_1669, w_011_1670, w_011_1671, w_011_1672, w_011_1673, w_011_1674, w_011_1675, w_011_1676, w_011_1677, w_011_1678, w_011_1679, w_011_1681, w_011_1682, w_011_1683, w_011_1685, w_011_1686, w_011_1687, w_011_1688, w_011_1689, w_011_1691, w_011_1692, w_011_1693, w_011_1694, w_011_1695, w_011_1696, w_011_1697, w_011_1698, w_011_1699, w_011_1700, w_011_1701, w_011_1702, w_011_1703, w_011_1704, w_011_1705, w_011_1707, w_011_1708, w_011_1709, w_011_1710, w_011_1711, w_011_1712, w_011_1713, w_011_1714, w_011_1715, w_011_1716, w_011_1717, w_011_1718, w_011_1719, w_011_1720, w_011_1721, w_011_1722, w_011_1723, w_011_1724, w_011_1725, w_011_1726, w_011_1727, w_011_1728, w_011_1729, w_011_1730, w_011_1731, w_011_1732, w_011_1733, w_011_1734, w_011_1735, w_011_1737, w_011_1738, w_011_1739, w_011_1740, w_011_1741, w_011_1742, w_011_1743, w_011_1744, w_011_1745, w_011_1747, w_011_1748, w_011_1749, w_011_1750, w_011_1751, w_011_1752, w_011_1753, w_011_1754, w_011_1755, w_011_1756, w_011_1757, w_011_1758, w_011_1759, w_011_1760, w_011_1761, w_011_1762, w_011_1763, w_011_1764, w_011_1765, w_011_1766, w_011_1767, w_011_1768, w_011_1769, w_011_1770, w_011_1771, w_011_1772, w_011_1773, w_011_1774, w_011_1775, w_011_1776, w_011_1777, w_011_1779, w_011_1780, w_011_1781, w_011_1782, w_011_1783, w_011_1784, w_011_1785, w_011_1786, w_011_1787, w_011_1788, w_011_1789, w_011_1790, w_011_1791, w_011_1792, w_011_1793, w_011_1795, w_011_1796, w_011_1797, w_011_1798, w_011_1799, w_011_1800, w_011_1801, w_011_1802, w_011_1803, w_011_1804, w_011_1805, w_011_1806, w_011_1807, w_011_1808, w_011_1809, w_011_1810, w_011_1811, w_011_1812, w_011_1813, w_011_1814, w_011_1815, w_011_1816, w_011_1817, w_011_1818, w_011_1819, w_011_1820, w_011_1821, w_011_1822, w_011_1823, w_011_1824, w_011_1825, w_011_1826, w_011_1827, w_011_1828, w_011_1829, w_011_1830, w_011_1831, w_011_1832, w_011_1833, w_011_1834, w_011_1836, w_011_1837, w_011_1838, w_011_1839, w_011_1840, w_011_1841, w_011_1842, w_011_1843, w_011_1844, w_011_1845, w_011_1846, w_011_1847, w_011_1848, w_011_1849, w_011_1850, w_011_1851, w_011_1852, w_011_1853, w_011_1854, w_011_1855, w_011_1856, w_011_1858, w_011_1859, w_011_1860, w_011_1861, w_011_1862, w_011_1863, w_011_1864, w_011_1865, w_011_1866, w_011_1867, w_011_1869, w_011_1870, w_011_1871, w_011_1872, w_011_1873, w_011_1874, w_011_1875, w_011_1876, w_011_1877, w_011_1878, w_011_1879, w_011_1880, w_011_1881, w_011_1882, w_011_1883, w_011_1884, w_011_1885, w_011_1886, w_011_1887, w_011_1888, w_011_1891, w_011_1892, w_011_1893, w_011_1894, w_011_1895, w_011_1896, w_011_1897, w_011_1898, w_011_1899, w_011_1900, w_011_1901, w_011_1902, w_011_1903, w_011_1904, w_011_1905, w_011_1906, w_011_1907, w_011_1908, w_011_1909, w_011_1910, w_011_1911, w_011_1912, w_011_1913, w_011_1914, w_011_1915, w_011_1916, w_011_1917, w_011_1918, w_011_1920, w_011_1921, w_011_1922, w_011_1924, w_011_1925, w_011_1926, w_011_1927, w_011_1928, w_011_1929, w_011_1930, w_011_1931, w_011_1932, w_011_1933, w_011_1934, w_011_1935, w_011_1936, w_011_1937, w_011_1938, w_011_1939, w_011_1940, w_011_1941, w_011_1942, w_011_1943, w_011_1944, w_011_1945, w_011_1946, w_011_1947, w_011_1948, w_011_1951, w_011_1952, w_011_1953, w_011_1954, w_011_1955, w_011_1956, w_011_1957, w_011_1959, w_011_1960, w_011_1961, w_011_1962, w_011_1963, w_011_1964, w_011_1966, w_011_1967, w_011_1968, w_011_1969, w_011_1970, w_011_1971, w_011_1972, w_011_1973, w_011_1975, w_011_1976, w_011_1977, w_011_1978, w_011_1979, w_011_1980, w_011_1981, w_011_1982, w_011_1983, w_011_1984, w_011_1985, w_011_1986, w_011_1987, w_011_1988, w_011_1990, w_011_1991, w_011_1992, w_011_1993, w_011_1994, w_011_1995, w_011_1996, w_011_1997, w_011_1998, w_011_1999, w_011_2000, w_011_2001, w_011_2002, w_011_2003, w_011_2004, w_011_2005, w_011_2006, w_011_2007, w_011_2008, w_011_2009, w_011_2010, w_011_2011, w_011_2013, w_011_2014, w_011_2015, w_011_2016, w_011_2017, w_011_2018, w_011_2019, w_011_2020, w_011_2021, w_011_2022, w_011_2023, w_011_2024, w_011_2025, w_011_2026, w_011_2027, w_011_2028, w_011_2029, w_011_2030, w_011_2031, w_011_2032, w_011_2033, w_011_2034, w_011_2035, w_011_2036, w_011_2037, w_011_2038, w_011_2039, w_011_2040, w_011_2041, w_011_2042, w_011_2043, w_011_2044, w_011_2046, w_011_2047, w_011_2048, w_011_2049, w_011_2050, w_011_2051, w_011_2052, w_011_2053, w_011_2054, w_011_2055, w_011_2056, w_011_2057, w_011_2058, w_011_2060, w_011_2061, w_011_2062, w_011_2063, w_011_2064, w_011_2065, w_011_2066, w_011_2067, w_011_2068, w_011_2069, w_011_2070, w_011_2071, w_011_2072, w_011_2073, w_011_2074, w_011_2075, w_011_2076, w_011_2077, w_011_2078, w_011_2079, w_011_2080, w_011_2081, w_011_2082, w_011_2083, w_011_2084, w_011_2085, w_011_2086, w_011_2087, w_011_2088, w_011_2089, w_011_2090, w_011_2091, w_011_2092, w_011_2093, w_011_2094, w_011_2095, w_011_2096, w_011_2097, w_011_2098, w_011_2099, w_011_2100, w_011_2101, w_011_2102, w_011_2103, w_011_2104, w_011_2105, w_011_2106, w_011_2107, w_011_2108, w_011_2109, w_011_2110, w_011_2111, w_011_2112, w_011_2113, w_011_2114, w_011_2115, w_011_2116, w_011_2117, w_011_2118, w_011_2119, w_011_2120, w_011_2122, w_011_2123, w_011_2124, w_011_2125, w_011_2126, w_011_2128, w_011_2129, w_011_2130, w_011_2131, w_011_2132, w_011_2133, w_011_2134, w_011_2135, w_011_2136, w_011_2138, w_011_2139, w_011_2140, w_011_2141, w_011_2142, w_011_2143, w_011_2144, w_011_2146, w_011_2147, w_011_2148, w_011_2149, w_011_2150, w_011_2151, w_011_2152, w_011_2153, w_011_2154, w_011_2155, w_011_2156, w_011_2157, w_011_2158, w_011_2159, w_011_2161, w_011_2162, w_011_2163, w_011_2164, w_011_2165, w_011_2166, w_011_2167, w_011_2168, w_011_2169, w_011_2170, w_011_2171, w_011_2172, w_011_2173, w_011_2174, w_011_2175, w_011_2176, w_011_2177, w_011_2178, w_011_2179, w_011_2180, w_011_2181, w_011_2182, w_011_2183, w_011_2184, w_011_2187, w_011_2188, w_011_2189, w_011_2190, w_011_2191, w_011_2192, w_011_2193, w_011_2194, w_011_2195, w_011_2196, w_011_2197, w_011_2198, w_011_2199, w_011_2200, w_011_2201, w_011_2202, w_011_2203, w_011_2204, w_011_2205, w_011_2206, w_011_2207, w_011_2209, w_011_2210, w_011_2211, w_011_2212, w_011_2213, w_011_2215, w_011_2216, w_011_2217, w_011_2218, w_011_2219, w_011_2220, w_011_2221, w_011_2222, w_011_2223, w_011_2224, w_011_2225, w_011_2226, w_011_2227, w_011_2228, w_011_2229, w_011_2230, w_011_2231, w_011_2232, w_011_2233, w_011_2234, w_011_2236, w_011_2237, w_011_2238, w_011_2239, w_011_2240, w_011_2241, w_011_2242, w_011_2243, w_011_2244, w_011_2245, w_011_2246, w_011_2247, w_011_2248, w_011_2249, w_011_2250, w_011_2251, w_011_2252, w_011_2253, w_011_2254, w_011_2255, w_011_2256, w_011_2257, w_011_2258, w_011_2259, w_011_2260, w_011_2261, w_011_2262, w_011_2263, w_011_2264, w_011_2265, w_011_2266, w_011_2267, w_011_2269, w_011_2270, w_011_2271, w_011_2272, w_011_2273, w_011_2274, w_011_2275, w_011_2276, w_011_2277, w_011_2278, w_011_2279, w_011_2280, w_011_2281, w_011_2282, w_011_2283, w_011_2284, w_011_2285, w_011_2286, w_011_2287, w_011_2288, w_011_2289, w_011_2290, w_011_2291, w_011_2292, w_011_2293, w_011_2294, w_011_2295, w_011_2296, w_011_2297, w_011_2299, w_011_2300, w_011_2301, w_011_2302, w_011_2303, w_011_2304, w_011_2305, w_011_2306, w_011_2307, w_011_2308, w_011_2309, w_011_2310, w_011_2311, w_011_2312, w_011_2313, w_011_2314, w_011_2315, w_011_2316, w_011_2317, w_011_2318, w_011_2319, w_011_2320, w_011_2321, w_011_2322, w_011_2323, w_011_2324, w_011_2325, w_011_2326, w_011_2327, w_011_2328;
  wire w_012_000, w_012_001, w_012_002, w_012_003, w_012_004, w_012_005, w_012_006, w_012_007, w_012_008, w_012_009, w_012_010, w_012_011, w_012_012, w_012_013, w_012_014, w_012_015, w_012_016, w_012_017, w_012_018, w_012_019, w_012_020, w_012_021, w_012_022, w_012_023, w_012_024, w_012_025, w_012_026, w_012_027, w_012_028, w_012_029, w_012_030, w_012_031, w_012_032, w_012_033, w_012_034, w_012_035, w_012_036, w_012_037, w_012_038, w_012_039, w_012_040, w_012_041, w_012_042, w_012_043, w_012_044, w_012_045, w_012_046, w_012_047, w_012_048, w_012_049, w_012_050, w_012_051, w_012_052, w_012_053, w_012_054, w_012_055, w_012_056, w_012_057, w_012_058, w_012_059, w_012_060, w_012_061, w_012_062, w_012_063, w_012_064, w_012_065, w_012_066, w_012_067, w_012_068, w_012_069, w_012_070, w_012_071, w_012_072, w_012_073, w_012_074, w_012_075, w_012_076, w_012_077, w_012_078, w_012_079, w_012_080, w_012_081, w_012_082, w_012_083, w_012_084, w_012_085, w_012_086, w_012_087, w_012_088, w_012_089, w_012_090, w_012_091, w_012_092, w_012_093, w_012_094, w_012_095, w_012_096, w_012_097, w_012_098, w_012_099, w_012_100, w_012_101, w_012_102, w_012_103, w_012_104, w_012_105, w_012_106, w_012_107, w_012_108, w_012_109, w_012_110, w_012_111, w_012_112, w_012_113, w_012_114, w_012_115, w_012_116, w_012_117, w_012_118, w_012_119, w_012_120, w_012_121, w_012_122, w_012_123, w_012_124, w_012_125, w_012_126, w_012_127, w_012_128, w_012_129, w_012_130, w_012_131, w_012_132, w_012_133, w_012_134, w_012_135, w_012_136, w_012_137, w_012_138, w_012_139, w_012_140, w_012_141, w_012_142, w_012_143, w_012_144, w_012_145, w_012_146, w_012_147, w_012_148, w_012_149, w_012_150, w_012_151, w_012_152, w_012_153, w_012_154, w_012_155, w_012_156, w_012_157, w_012_158, w_012_159, w_012_160, w_012_161, w_012_162, w_012_163, w_012_164, w_012_165, w_012_166, w_012_167, w_012_168, w_012_169, w_012_170, w_012_171, w_012_172, w_012_173, w_012_174, w_012_175, w_012_176, w_012_177, w_012_178, w_012_179, w_012_180, w_012_181, w_012_182, w_012_183, w_012_184, w_012_185, w_012_186, w_012_187, w_012_188, w_012_189, w_012_190, w_012_191, w_012_192, w_012_193, w_012_194, w_012_195, w_012_196, w_012_197, w_012_198, w_012_199, w_012_200, w_012_201, w_012_202, w_012_203, w_012_204, w_012_205, w_012_206, w_012_207, w_012_208, w_012_209, w_012_210, w_012_211, w_012_212, w_012_213, w_012_214, w_012_215, w_012_216, w_012_217, w_012_218, w_012_219, w_012_220, w_012_221, w_012_222, w_012_223, w_012_224, w_012_225, w_012_226, w_012_227, w_012_228, w_012_229, w_012_230, w_012_231, w_012_232, w_012_233, w_012_234, w_012_235, w_012_236, w_012_237, w_012_238, w_012_239, w_012_240, w_012_241, w_012_242, w_012_243, w_012_244, w_012_245, w_012_246, w_012_247, w_012_248, w_012_249, w_012_250, w_012_251, w_012_252, w_012_253, w_012_254, w_012_255, w_012_256, w_012_257, w_012_258, w_012_259, w_012_260, w_012_261, w_012_262, w_012_263, w_012_264, w_012_265, w_012_266, w_012_267, w_012_268, w_012_269, w_012_270, w_012_271, w_012_272, w_012_273, w_012_274, w_012_275, w_012_276, w_012_277, w_012_278, w_012_279, w_012_280, w_012_281, w_012_282, w_012_283, w_012_284, w_012_285, w_012_286, w_012_287, w_012_288, w_012_289, w_012_290, w_012_291, w_012_292, w_012_293, w_012_294, w_012_295, w_012_296, w_012_297, w_012_298, w_012_299, w_012_300, w_012_301, w_012_302, w_012_303, w_012_304, w_012_305, w_012_306, w_012_307, w_012_308, w_012_309, w_012_310, w_012_311, w_012_312, w_012_313, w_012_314, w_012_315, w_012_316, w_012_317, w_012_318, w_012_319, w_012_320, w_012_321, w_012_322, w_012_323, w_012_324, w_012_325, w_012_326, w_012_327, w_012_328, w_012_329, w_012_330, w_012_331, w_012_332, w_012_333, w_012_334, w_012_335, w_012_336, w_012_337, w_012_338, w_012_339, w_012_340, w_012_341, w_012_342, w_012_343, w_012_344, w_012_345, w_012_346, w_012_347, w_012_348, w_012_349, w_012_350, w_012_351, w_012_352, w_012_353, w_012_354, w_012_355, w_012_356, w_012_357, w_012_358, w_012_359, w_012_360, w_012_361, w_012_362, w_012_363, w_012_364, w_012_365, w_012_366, w_012_367, w_012_368, w_012_369, w_012_370, w_012_371, w_012_372, w_012_373, w_012_374, w_012_375, w_012_376, w_012_377, w_012_378, w_012_379, w_012_380, w_012_381, w_012_382, w_012_383, w_012_384, w_012_385, w_012_386, w_012_387, w_012_388, w_012_389, w_012_390, w_012_391, w_012_392, w_012_393, w_012_394, w_012_395, w_012_396, w_012_397, w_012_398, w_012_399, w_012_400, w_012_401, w_012_402, w_012_403, w_012_404, w_012_405, w_012_406, w_012_407, w_012_408, w_012_409, w_012_410, w_012_411, w_012_412, w_012_413, w_012_414, w_012_415, w_012_416, w_012_417, w_012_418, w_012_419, w_012_420, w_012_421, w_012_422, w_012_423, w_012_424, w_012_425, w_012_426, w_012_427, w_012_428, w_012_429, w_012_430, w_012_431, w_012_432, w_012_433, w_012_434, w_012_435, w_012_436, w_012_437, w_012_438, w_012_439, w_012_440, w_012_441, w_012_442, w_012_443, w_012_444, w_012_445, w_012_446, w_012_447, w_012_448, w_012_449, w_012_450, w_012_451, w_012_452, w_012_453, w_012_454, w_012_455, w_012_456, w_012_457, w_012_458, w_012_459, w_012_460, w_012_461, w_012_462, w_012_463, w_012_464, w_012_465, w_012_466, w_012_467, w_012_468, w_012_469, w_012_470, w_012_471, w_012_472, w_012_473, w_012_474, w_012_475, w_012_476, w_012_477, w_012_478, w_012_479, w_012_480, w_012_481, w_012_482, w_012_483, w_012_484, w_012_485, w_012_486, w_012_487, w_012_488, w_012_489, w_012_490, w_012_491, w_012_492, w_012_493, w_012_494, w_012_495, w_012_496, w_012_497, w_012_498, w_012_499, w_012_500, w_012_501, w_012_502, w_012_503, w_012_504, w_012_505, w_012_506, w_012_507, w_012_508, w_012_509, w_012_510, w_012_511, w_012_512, w_012_513, w_012_514, w_012_515, w_012_516, w_012_517, w_012_518, w_012_519, w_012_520, w_012_521, w_012_522, w_012_523, w_012_524, w_012_525, w_012_526, w_012_527, w_012_528, w_012_529, w_012_530, w_012_531, w_012_532, w_012_533, w_012_534, w_012_535, w_012_536, w_012_537, w_012_538, w_012_539, w_012_540, w_012_541, w_012_542, w_012_543, w_012_544, w_012_545, w_012_546, w_012_547, w_012_548, w_012_549, w_012_550, w_012_551, w_012_552, w_012_553, w_012_554, w_012_555, w_012_556, w_012_557, w_012_558, w_012_559, w_012_560, w_012_561, w_012_562, w_012_563, w_012_564, w_012_565, w_012_566, w_012_567, w_012_568, w_012_569, w_012_570, w_012_571, w_012_572, w_012_573, w_012_574, w_012_575, w_012_576, w_012_577, w_012_578, w_012_579, w_012_580, w_012_581, w_012_582, w_012_583, w_012_584, w_012_585, w_012_586, w_012_587, w_012_588, w_012_589, w_012_590, w_012_591, w_012_592, w_012_593, w_012_594, w_012_595, w_012_596, w_012_597, w_012_598, w_012_599, w_012_600, w_012_601, w_012_602, w_012_603, w_012_604, w_012_605, w_012_606, w_012_607, w_012_608, w_012_609, w_012_610, w_012_611, w_012_612, w_012_613, w_012_614, w_012_615, w_012_616, w_012_617, w_012_618, w_012_619, w_012_620, w_012_621, w_012_622, w_012_623, w_012_624, w_012_625, w_012_626, w_012_627, w_012_628, w_012_629, w_012_630, w_012_631, w_012_632, w_012_633, w_012_634, w_012_635, w_012_636, w_012_637, w_012_638, w_012_639, w_012_640, w_012_641, w_012_642, w_012_643, w_012_644, w_012_645, w_012_646, w_012_647, w_012_648, w_012_649, w_012_650, w_012_651, w_012_652, w_012_653, w_012_654, w_012_655, w_012_656, w_012_657, w_012_658, w_012_659, w_012_660, w_012_661, w_012_662, w_012_663, w_012_664, w_012_665, w_012_666, w_012_667, w_012_668, w_012_669, w_012_670, w_012_671, w_012_672, w_012_673, w_012_674, w_012_675, w_012_676, w_012_677, w_012_678, w_012_679, w_012_680, w_012_681, w_012_682, w_012_683, w_012_684, w_012_685, w_012_686, w_012_687, w_012_688, w_012_689, w_012_690, w_012_691, w_012_692, w_012_693, w_012_694, w_012_695, w_012_696, w_012_697, w_012_698, w_012_699, w_012_700, w_012_701, w_012_702, w_012_703, w_012_704, w_012_705, w_012_706, w_012_707, w_012_708, w_012_709, w_012_710, w_012_711, w_012_712, w_012_713, w_012_714, w_012_715, w_012_716, w_012_717, w_012_718, w_012_719, w_012_720, w_012_721, w_012_722, w_012_723, w_012_724, w_012_725, w_012_726, w_012_727, w_012_728, w_012_729, w_012_730, w_012_731, w_012_732, w_012_733, w_012_734, w_012_735, w_012_736, w_012_737, w_012_738, w_012_739, w_012_740, w_012_741, w_012_742, w_012_743, w_012_744, w_012_745, w_012_746, w_012_747, w_012_748, w_012_749, w_012_750, w_012_751, w_012_752, w_012_753, w_012_754, w_012_755, w_012_756, w_012_757, w_012_758, w_012_759, w_012_760, w_012_761, w_012_762, w_012_763, w_012_764, w_012_765, w_012_766, w_012_767, w_012_768, w_012_769, w_012_770, w_012_771, w_012_772, w_012_773, w_012_774, w_012_775, w_012_776, w_012_777, w_012_778, w_012_779, w_012_780, w_012_781, w_012_782, w_012_783, w_012_784, w_012_785, w_012_786, w_012_787, w_012_788, w_012_789, w_012_790, w_012_791, w_012_792, w_012_793, w_012_794, w_012_795, w_012_796, w_012_797, w_012_798, w_012_799, w_012_800, w_012_801, w_012_802, w_012_803, w_012_804, w_012_805, w_012_806, w_012_807, w_012_808, w_012_809, w_012_810, w_012_811, w_012_812, w_012_813, w_012_814, w_012_815, w_012_816, w_012_817, w_012_818, w_012_819, w_012_820, w_012_821, w_012_822, w_012_823, w_012_824, w_012_825, w_012_826, w_012_827, w_012_828, w_012_829, w_012_830, w_012_831, w_012_832, w_012_833, w_012_834, w_012_835, w_012_836, w_012_837, w_012_838, w_012_839, w_012_840, w_012_841, w_012_842, w_012_843, w_012_844, w_012_845, w_012_846, w_012_847, w_012_848, w_012_849, w_012_850, w_012_851, w_012_852, w_012_853, w_012_854, w_012_855, w_012_856, w_012_857, w_012_858, w_012_859, w_012_860, w_012_861, w_012_862, w_012_863, w_012_864, w_012_865, w_012_866, w_012_867, w_012_868, w_012_869, w_012_870, w_012_871, w_012_872, w_012_873, w_012_874, w_012_875, w_012_876, w_012_877, w_012_878, w_012_879, w_012_880, w_012_881, w_012_882, w_012_883, w_012_884, w_012_885, w_012_886, w_012_887, w_012_888, w_012_889, w_012_890, w_012_891, w_012_892, w_012_893, w_012_894, w_012_895, w_012_896, w_012_897, w_012_898, w_012_899, w_012_900, w_012_901, w_012_902, w_012_903, w_012_904, w_012_905, w_012_906, w_012_907, w_012_908, w_012_909, w_012_910, w_012_911, w_012_912, w_012_913, w_012_914, w_012_915, w_012_916, w_012_917, w_012_918, w_012_919, w_012_920, w_012_921, w_012_922, w_012_923, w_012_924, w_012_925;
  wire w_013_000, w_013_001, w_013_002, w_013_003, w_013_004, w_013_005, w_013_006, w_013_007, w_013_008, w_013_009, w_013_010, w_013_011, w_013_012, w_013_013, w_013_014, w_013_015, w_013_016, w_013_017, w_013_018, w_013_019, w_013_021, w_013_022, w_013_023, w_013_024, w_013_025, w_013_026, w_013_027, w_013_028, w_013_029, w_013_031, w_013_032, w_013_033, w_013_034, w_013_035, w_013_036, w_013_037, w_013_039, w_013_040, w_013_041, w_013_042, w_013_043, w_013_044, w_013_045, w_013_046, w_013_047, w_013_048, w_013_049, w_013_052, w_013_053, w_013_054, w_013_055, w_013_056, w_013_057, w_013_058, w_013_059, w_013_060, w_013_061, w_013_062, w_013_063, w_013_064, w_013_065, w_013_066, w_013_067, w_013_068, w_013_069, w_013_070, w_013_071, w_013_072, w_013_074, w_013_075, w_013_076, w_013_077, w_013_078, w_013_079, w_013_080, w_013_081, w_013_082, w_013_083, w_013_084, w_013_085, w_013_086, w_013_087, w_013_088, w_013_089, w_013_090, w_013_091, w_013_092, w_013_093, w_013_094, w_013_095, w_013_096, w_013_097, w_013_098, w_013_099, w_013_101, w_013_102, w_013_103, w_013_104, w_013_105, w_013_106, w_013_107, w_013_108, w_013_109, w_013_110, w_013_111, w_013_112, w_013_113, w_013_114, w_013_115, w_013_116, w_013_117, w_013_118, w_013_119, w_013_120, w_013_121, w_013_123, w_013_124, w_013_125, w_013_127, w_013_128, w_013_129, w_013_130, w_013_131, w_013_132, w_013_133, w_013_134, w_013_135, w_013_136, w_013_138, w_013_141, w_013_142, w_013_143, w_013_144, w_013_145, w_013_146, w_013_147, w_013_148, w_013_149, w_013_150, w_013_151, w_013_152, w_013_153, w_013_154, w_013_155, w_013_156, w_013_157, w_013_158, w_013_159, w_013_160, w_013_161, w_013_162, w_013_163, w_013_164, w_013_165, w_013_166, w_013_167, w_013_168, w_013_172, w_013_173, w_013_174, w_013_175, w_013_176, w_013_177, w_013_178, w_013_179, w_013_181, w_013_182, w_013_183, w_013_184, w_013_186, w_013_187, w_013_188, w_013_189, w_013_190, w_013_191, w_013_192, w_013_193, w_013_194, w_013_195, w_013_196, w_013_197, w_013_198, w_013_199, w_013_201, w_013_202, w_013_203, w_013_204, w_013_205, w_013_206, w_013_209, w_013_210, w_013_211, w_013_212, w_013_213, w_013_214, w_013_215, w_013_217, w_013_218, w_013_219, w_013_220, w_013_221, w_013_222, w_013_223, w_013_224, w_013_225, w_013_226, w_013_227, w_013_228, w_013_229, w_013_230, w_013_231, w_013_232, w_013_233, w_013_234, w_013_235, w_013_236, w_013_237, w_013_238, w_013_239, w_013_240, w_013_241, w_013_242, w_013_243, w_013_244, w_013_245, w_013_246, w_013_247, w_013_248, w_013_249, w_013_251, w_013_252, w_013_253, w_013_254, w_013_255, w_013_256, w_013_257, w_013_258, w_013_259, w_013_260, w_013_261, w_013_262, w_013_263, w_013_264, w_013_265, w_013_266, w_013_267, w_013_268, w_013_269, w_013_270, w_013_271, w_013_272, w_013_273, w_013_274, w_013_275, w_013_276, w_013_277, w_013_278, w_013_279, w_013_280, w_013_281, w_013_282, w_013_283, w_013_284, w_013_285, w_013_286, w_013_287, w_013_288, w_013_289, w_013_290, w_013_291, w_013_292, w_013_293, w_013_294, w_013_295, w_013_296, w_013_297, w_013_299, w_013_300, w_013_301, w_013_302, w_013_303, w_013_304, w_013_305, w_013_306, w_013_308, w_013_309, w_013_310, w_013_311, w_013_312, w_013_313, w_013_314, w_013_315, w_013_316, w_013_317, w_013_318, w_013_319, w_013_320, w_013_321, w_013_322, w_013_323, w_013_324, w_013_325, w_013_326, w_013_328, w_013_329, w_013_330, w_013_331, w_013_332, w_013_333, w_013_334, w_013_335, w_013_336, w_013_337, w_013_338, w_013_339, w_013_340, w_013_341, w_013_342, w_013_343, w_013_344, w_013_345, w_013_346, w_013_347, w_013_348, w_013_349, w_013_350, w_013_351, w_013_352, w_013_353, w_013_354, w_013_355, w_013_356, w_013_357, w_013_358, w_013_359, w_013_360, w_013_361, w_013_362, w_013_363, w_013_364, w_013_365, w_013_366, w_013_367, w_013_369, w_013_370, w_013_371, w_013_372, w_013_373, w_013_374, w_013_375, w_013_376, w_013_377, w_013_378, w_013_379, w_013_380, w_013_381, w_013_382, w_013_383, w_013_384, w_013_385, w_013_386, w_013_387, w_013_388, w_013_389, w_013_390, w_013_391, w_013_392, w_013_393, w_013_394, w_013_395, w_013_396, w_013_397, w_013_399, w_013_400, w_013_401, w_013_402, w_013_403, w_013_404, w_013_406, w_013_407, w_013_408, w_013_409, w_013_410, w_013_411, w_013_412, w_013_413, w_013_414, w_013_415, w_013_416, w_013_417, w_013_418, w_013_419, w_013_420, w_013_421, w_013_422, w_013_423, w_013_424, w_013_425, w_013_426, w_013_428, w_013_429, w_013_430, w_013_431, w_013_432, w_013_433, w_013_434, w_013_435, w_013_437, w_013_438, w_013_439, w_013_440, w_013_441, w_013_442, w_013_443, w_013_444, w_013_445, w_013_446, w_013_447, w_013_448, w_013_449, w_013_450, w_013_451, w_013_452, w_013_453, w_013_454, w_013_455, w_013_456, w_013_457, w_013_458, w_013_459, w_013_460, w_013_461, w_013_462, w_013_463, w_013_464, w_013_465, w_013_466, w_013_467, w_013_468, w_013_469, w_013_470, w_013_471, w_013_472, w_013_473, w_013_474, w_013_475, w_013_476, w_013_477, w_013_478, w_013_479, w_013_480, w_013_481, w_013_482, w_013_483, w_013_484, w_013_485, w_013_486, w_013_487, w_013_488, w_013_489, w_013_490, w_013_491, w_013_492, w_013_493, w_013_494, w_013_495, w_013_496, w_013_497, w_013_498, w_013_500, w_013_501, w_013_502, w_013_503, w_013_504, w_013_505, w_013_506, w_013_507, w_013_508, w_013_509, w_013_510, w_013_511, w_013_512, w_013_513, w_013_514, w_013_515, w_013_516, w_013_518, w_013_519, w_013_520, w_013_521, w_013_522, w_013_523, w_013_524, w_013_525, w_013_526, w_013_527, w_013_528, w_013_529, w_013_530, w_013_531, w_013_532, w_013_533, w_013_534, w_013_535, w_013_536, w_013_537, w_013_538, w_013_539, w_013_540, w_013_541, w_013_542, w_013_543, w_013_544, w_013_545, w_013_546, w_013_547, w_013_548, w_013_549, w_013_550, w_013_551, w_013_552, w_013_553, w_013_554, w_013_555, w_013_556, w_013_557, w_013_558, w_013_559, w_013_560, w_013_561, w_013_562, w_013_564, w_013_565, w_013_566, w_013_567, w_013_568, w_013_569, w_013_570, w_013_571, w_013_573, w_013_574, w_013_575, w_013_576, w_013_577, w_013_578, w_013_579, w_013_580, w_013_581, w_013_583, w_013_584, w_013_585, w_013_586, w_013_587, w_013_588, w_013_589, w_013_590, w_013_591, w_013_592, w_013_593, w_013_595, w_013_596, w_013_597, w_013_598, w_013_599, w_013_600, w_013_601, w_013_602, w_013_603, w_013_604, w_013_605, w_013_606, w_013_607, w_013_608, w_013_609, w_013_610, w_013_611, w_013_612, w_013_613, w_013_615, w_013_616, w_013_617, w_013_618, w_013_619, w_013_620, w_013_621, w_013_622, w_013_623, w_013_624, w_013_625, w_013_626, w_013_627, w_013_628, w_013_629, w_013_630, w_013_631, w_013_632, w_013_633, w_013_634, w_013_635, w_013_637, w_013_638, w_013_639, w_013_640, w_013_641, w_013_642, w_013_643, w_013_644, w_013_645, w_013_646, w_013_647, w_013_649, w_013_650, w_013_651, w_013_652, w_013_653, w_013_654, w_013_655, w_013_656, w_013_657, w_013_658, w_013_659, w_013_660, w_013_661, w_013_662, w_013_663, w_013_664, w_013_665, w_013_666, w_013_667, w_013_668, w_013_669, w_013_670, w_013_671, w_013_673, w_013_674, w_013_676, w_013_677, w_013_678, w_013_679, w_013_680, w_013_681, w_013_682, w_013_683, w_013_684, w_013_685, w_013_686, w_013_687, w_013_688, w_013_689, w_013_690, w_013_691, w_013_692, w_013_693, w_013_694, w_013_695, w_013_696, w_013_697, w_013_698, w_013_699, w_013_700, w_013_701, w_013_702, w_013_703, w_013_704, w_013_705, w_013_706, w_013_707, w_013_708, w_013_709, w_013_710, w_013_711, w_013_712, w_013_713, w_013_714, w_013_715, w_013_716, w_013_717, w_013_718, w_013_719, w_013_720, w_013_721, w_013_722, w_013_723, w_013_724, w_013_725, w_013_726, w_013_727, w_013_728, w_013_729, w_013_730, w_013_731, w_013_733, w_013_734, w_013_735, w_013_736, w_013_737, w_013_738, w_013_739, w_013_740, w_013_741, w_013_743, w_013_744, w_013_745, w_013_746, w_013_747, w_013_748, w_013_749, w_013_750, w_013_751, w_013_752, w_013_753, w_013_754, w_013_755, w_013_756, w_013_757, w_013_758, w_013_759, w_013_760, w_013_761, w_013_762, w_013_763, w_013_764, w_013_765, w_013_766, w_013_767, w_013_768, w_013_769, w_013_770, w_013_771, w_013_772, w_013_773, w_013_774, w_013_775, w_013_776, w_013_777, w_013_778, w_013_779, w_013_780, w_013_781, w_013_782, w_013_783, w_013_784, w_013_785, w_013_786, w_013_787, w_013_788, w_013_789, w_013_790, w_013_791, w_013_792, w_013_793, w_013_794, w_013_795, w_013_796, w_013_797, w_013_798, w_013_799, w_013_800, w_013_801, w_013_802, w_013_803, w_013_804, w_013_805, w_013_806, w_013_807, w_013_808, w_013_809, w_013_810, w_013_811, w_013_812, w_013_813, w_013_814, w_013_815, w_013_816, w_013_817, w_013_818, w_013_819, w_013_820, w_013_821, w_013_822, w_013_823, w_013_824, w_013_825, w_013_826, w_013_828, w_013_829, w_013_830, w_013_831, w_013_832, w_013_833, w_013_834, w_013_835, w_013_836, w_013_838, w_013_839, w_013_840, w_013_841, w_013_842, w_013_844, w_013_845, w_013_846, w_013_847, w_013_848, w_013_849, w_013_850, w_013_851, w_013_852, w_013_853, w_013_855, w_013_856, w_013_857, w_013_858, w_013_859, w_013_860, w_013_861, w_013_862, w_013_863, w_013_864, w_013_865, w_013_866, w_013_867, w_013_868, w_013_869, w_013_870, w_013_871, w_013_872, w_013_873, w_013_874, w_013_875, w_013_876, w_013_877, w_013_878, w_013_879, w_013_880, w_013_881, w_013_882, w_013_883, w_013_884, w_013_885, w_013_886, w_013_887, w_013_888, w_013_889, w_013_890, w_013_891, w_013_892, w_013_893, w_013_894, w_013_895, w_013_896, w_013_897, w_013_898, w_013_899, w_013_900, w_013_901, w_013_902, w_013_903, w_013_904, w_013_905, w_013_906, w_013_907, w_013_908, w_013_909, w_013_911, w_013_912, w_013_913, w_013_914, w_013_915, w_013_916, w_013_917, w_013_918, w_013_919, w_013_920, w_013_921, w_013_922, w_013_923, w_013_924, w_013_925, w_013_926, w_013_927, w_013_928, w_013_929, w_013_930, w_013_931, w_013_932, w_013_933, w_013_934, w_013_935, w_013_936, w_013_937, w_013_938, w_013_939, w_013_940, w_013_941, w_013_942, w_013_943, w_013_944, w_013_945, w_013_946, w_013_947, w_013_948, w_013_949, w_013_950, w_013_952, w_013_953, w_013_954, w_013_956, w_013_957, w_013_958, w_013_959, w_013_960, w_013_961, w_013_962, w_013_963, w_013_964, w_013_965, w_013_966, w_013_967, w_013_968, w_013_969, w_013_970, w_013_971, w_013_972, w_013_973, w_013_974, w_013_975, w_013_976, w_013_977, w_013_978, w_013_979, w_013_980, w_013_981, w_013_982, w_013_984, w_013_985, w_013_986, w_013_987, w_013_988, w_013_989, w_013_990, w_013_991, w_013_992, w_013_993, w_013_994, w_013_996, w_013_997, w_013_998, w_013_999, w_013_1000, w_013_1001, w_013_1002, w_013_1003, w_013_1005, w_013_1006, w_013_1007, w_013_1008, w_013_1009, w_013_1010, w_013_1011, w_013_1012, w_013_1013, w_013_1014, w_013_1015, w_013_1016, w_013_1017, w_013_1018, w_013_1019, w_013_1020, w_013_1021, w_013_1022, w_013_1023, w_013_1024, w_013_1025, w_013_1026, w_013_1027, w_013_1028, w_013_1029, w_013_1030, w_013_1031, w_013_1032, w_013_1033, w_013_1034, w_013_1035, w_013_1036, w_013_1037, w_013_1038, w_013_1039, w_013_1040, w_013_1041, w_013_1042, w_013_1043, w_013_1044, w_013_1045, w_013_1046, w_013_1047, w_013_1048, w_013_1049, w_013_1051, w_013_1053, w_013_1054, w_013_1055, w_013_1056, w_013_1057, w_013_1058, w_013_1059, w_013_1060, w_013_1061, w_013_1062, w_013_1063, w_013_1064, w_013_1065, w_013_1067, w_013_1068, w_013_1069, w_013_1070, w_013_1071, w_013_1072, w_013_1073, w_013_1074, w_013_1075, w_013_1076, w_013_1077, w_013_1078, w_013_1079, w_013_1080, w_013_1081, w_013_1082, w_013_1083, w_013_1084, w_013_1085, w_013_1086, w_013_1087, w_013_1088, w_013_1089, w_013_1090, w_013_1091, w_013_1092, w_013_1093, w_013_1094, w_013_1095, w_013_1096, w_013_1097, w_013_1098, w_013_1099, w_013_1100, w_013_1101, w_013_1102, w_013_1103, w_013_1104, w_013_1105, w_013_1106, w_013_1107, w_013_1108, w_013_1109, w_013_1110, w_013_1111, w_013_1112, w_013_1113, w_013_1114, w_013_1115, w_013_1116, w_013_1117, w_013_1118, w_013_1119, w_013_1120, w_013_1121, w_013_1122, w_013_1123, w_013_1124, w_013_1125, w_013_1126, w_013_1127, w_013_1128, w_013_1129, w_013_1130, w_013_1131, w_013_1132, w_013_1133, w_013_1134, w_013_1135, w_013_1136, w_013_1137, w_013_1138, w_013_1139, w_013_1140, w_013_1141, w_013_1142, w_013_1143, w_013_1144, w_013_1145, w_013_1146, w_013_1147, w_013_1148, w_013_1149, w_013_1150, w_013_1151, w_013_1152, w_013_1153, w_013_1154, w_013_1155, w_013_1156, w_013_1157, w_013_1158, w_013_1159, w_013_1160, w_013_1161, w_013_1162, w_013_1163, w_013_1164, w_013_1165, w_013_1166, w_013_1167, w_013_1168, w_013_1169, w_013_1170, w_013_1171, w_013_1172, w_013_1173, w_013_1174, w_013_1175, w_013_1176, w_013_1177, w_013_1178, w_013_1179, w_013_1180, w_013_1181, w_013_1182, w_013_1183, w_013_1185, w_013_1186, w_013_1187, w_013_1188, w_013_1189, w_013_1191, w_013_1192, w_013_1193, w_013_1194, w_013_1195, w_013_1196, w_013_1197, w_013_1198, w_013_1199, w_013_1200, w_013_1201, w_013_1202, w_013_1203, w_013_1204, w_013_1205, w_013_1206, w_013_1207, w_013_1208, w_013_1209, w_013_1210, w_013_1211, w_013_1212, w_013_1213, w_013_1214, w_013_1215, w_013_1216, w_013_1217, w_013_1218, w_013_1219, w_013_1220, w_013_1221, w_013_1222, w_013_1223, w_013_1224, w_013_1225, w_013_1226, w_013_1227, w_013_1228, w_013_1229, w_013_1230, w_013_1231, w_013_1232, w_013_1233, w_013_1234, w_013_1235, w_013_1236, w_013_1237, w_013_1238, w_013_1239, w_013_1240, w_013_1241, w_013_1242, w_013_1243, w_013_1244, w_013_1245, w_013_1246, w_013_1247, w_013_1248, w_013_1249, w_013_1250, w_013_1251, w_013_1252, w_013_1253, w_013_1254, w_013_1255, w_013_1256, w_013_1257, w_013_1258, w_013_1259, w_013_1260, w_013_1261, w_013_1262, w_013_1263, w_013_1264, w_013_1265, w_013_1266, w_013_1267, w_013_1268, w_013_1269, w_013_1270, w_013_1271, w_013_1272, w_013_1273, w_013_1274, w_013_1275, w_013_1276, w_013_1277, w_013_1278, w_013_1279, w_013_1280, w_013_1281, w_013_1282, w_013_1283, w_013_1284, w_013_1285, w_013_1286, w_013_1287, w_013_1288, w_013_1289, w_013_1290, w_013_1291, w_013_1292, w_013_1293, w_013_1294, w_013_1295, w_013_1296, w_013_1297, w_013_1298, w_013_1299, w_013_1300, w_013_1301, w_013_1302, w_013_1303, w_013_1304, w_013_1305, w_013_1306, w_013_1307, w_013_1308, w_013_1309, w_013_1310, w_013_1311, w_013_1312, w_013_1313, w_013_1314, w_013_1315, w_013_1316, w_013_1317, w_013_1318, w_013_1319, w_013_1320, w_013_1321, w_013_1322, w_013_1323, w_013_1324, w_013_1325, w_013_1326, w_013_1327, w_013_1329, w_013_1330, w_013_1331, w_013_1332, w_013_1333, w_013_1334, w_013_1335, w_013_1336, w_013_1337, w_013_1338, w_013_1339, w_013_1340, w_013_1341, w_013_1342, w_013_1343, w_013_1344, w_013_1345, w_013_1347, w_013_1348, w_013_1349, w_013_1350, w_013_1351, w_013_1353, w_013_1354, w_013_1355, w_013_1356, w_013_1357, w_013_1358, w_013_1359, w_013_1361, w_013_1362, w_013_1363, w_013_1364, w_013_1365, w_013_1366, w_013_1367, w_013_1368, w_013_1370, w_013_1372, w_013_1373, w_013_1374, w_013_1375, w_013_1376, w_013_1377, w_013_1378, w_013_1379, w_013_1380, w_013_1381, w_013_1383, w_013_1385, w_013_1386, w_013_1387, w_013_1390, w_013_1391, w_013_1392, w_013_1393, w_013_1394, w_013_1395, w_013_1396, w_013_1397, w_013_1399, w_013_1400, w_013_1401, w_013_1402, w_013_1403, w_013_1404, w_013_1405, w_013_1406, w_013_1408, w_013_1409, w_013_1410, w_013_1411, w_013_1412, w_013_1414, w_013_1415, w_013_1416, w_013_1417, w_013_1418, w_013_1419, w_013_1421, w_013_1422, w_013_1423, w_013_1425, w_013_1426, w_013_1427, w_013_1428, w_013_1429, w_013_1431, w_013_1432, w_013_1436, w_013_1437, w_013_1439, w_013_1440, w_013_1442, w_013_1443, w_013_1444, w_013_1446, w_013_1447, w_013_1448, w_013_1449, w_013_1452, w_013_1453, w_013_1454, w_013_1456, w_013_1457, w_013_1458, w_013_1459, w_013_1460, w_013_1461, w_013_1462, w_013_1463, w_013_1464, w_013_1465, w_013_1467, w_013_1469, w_013_1470, w_013_1472, w_013_1473, w_013_1474, w_013_1475, w_013_1476, w_013_1477, w_013_1479, w_013_1480, w_013_1482, w_013_1483, w_013_1484, w_013_1485, w_013_1486, w_013_1487, w_013_1488, w_013_1491, w_013_1492, w_013_1493, w_013_1497, w_013_1499, w_013_1500, w_013_1501, w_013_1502, w_013_1503, w_013_1504, w_013_1505, w_013_1507, w_013_1508, w_013_1509, w_013_1510, w_013_1511, w_013_1512, w_013_1514, w_013_1515, w_013_1516, w_013_1517, w_013_1518, w_013_1519, w_013_1520, w_013_1521, w_013_1522, w_013_1523, w_013_1524, w_013_1525, w_013_1526, w_013_1527, w_013_1529, w_013_1531, w_013_1532, w_013_1533, w_013_1534, w_013_1537, w_013_1538, w_013_1539, w_013_1540, w_013_1541, w_013_1542, w_013_1543, w_013_1544, w_013_1545, w_013_1546, w_013_1547, w_013_1550, w_013_1552, w_013_1554, w_013_1555, w_013_1556, w_013_1557, w_013_1558, w_013_1559, w_013_1560, w_013_1561, w_013_1562, w_013_1563, w_013_1564, w_013_1565, w_013_1566, w_013_1568, w_013_1569, w_013_1571, w_013_1573, w_013_1574, w_013_1575, w_013_1578, w_013_1579, w_013_1580, w_013_1581, w_013_1582, w_013_1583, w_013_1584, w_013_1585, w_013_1586, w_013_1587, w_013_1589, w_013_1590, w_013_1592, w_013_1593, w_013_1594, w_013_1596, w_013_1597, w_013_1598, w_013_1599, w_013_1600, w_013_1601, w_013_1602, w_013_1603, w_013_1604, w_013_1605, w_013_1606, w_013_1608, w_013_1609, w_013_1610, w_013_1612, w_013_1613, w_013_1614, w_013_1615, w_013_1616, w_013_1617, w_013_1618, w_013_1619, w_013_1621, w_013_1623, w_013_1625, w_013_1626, w_013_1627, w_013_1628, w_013_1629, w_013_1631, w_013_1632, w_013_1634, w_013_1635, w_013_1636, w_013_1637, w_013_1638, w_013_1639, w_013_1640, w_013_1641, w_013_1644, w_013_1645, w_013_1648, w_013_1649, w_013_1650, w_013_1652, w_013_1653, w_013_1654, w_013_1655, w_013_1656, w_013_1657, w_013_1658, w_013_1659, w_013_1660, w_013_1661, w_013_1662, w_013_1663, w_013_1664, w_013_1665, w_013_1666, w_013_1667, w_013_1668, w_013_1669, w_013_1671, w_013_1672, w_013_1673, w_013_1675, w_013_1676, w_013_1677, w_013_1678, w_013_1679, w_013_1680, w_013_1681, w_013_1682, w_013_1683, w_013_1684, w_013_1685, w_013_1686, w_013_1687, w_013_1688, w_013_1689, w_013_1690, w_013_1691, w_013_1692, w_013_1693, w_013_1694, w_013_1695, w_013_1696, w_013_1697, w_013_1698, w_013_1699, w_013_1700, w_013_1701, w_013_1702, w_013_1703, w_013_1704, w_013_1705, w_013_1706, w_013_1707, w_013_1708, w_013_1709, w_013_1712, w_013_1713, w_013_1715, w_013_1717, w_013_1718, w_013_1719, w_013_1720, w_013_1721, w_013_1722, w_013_1724, w_013_1725, w_013_1726, w_013_1727, w_013_1728, w_013_1729, w_013_1730, w_013_1731, w_013_1732, w_013_1733, w_013_1734, w_013_1735, w_013_1737, w_013_1738, w_013_1739, w_013_1740, w_013_1741, w_013_1743, w_013_1744, w_013_1745, w_013_1746, w_013_1747, w_013_1748, w_013_1749, w_013_1750, w_013_1751, w_013_1752, w_013_1753, w_013_1755, w_013_1756, w_013_1757, w_013_1758, w_013_1759, w_013_1760, w_013_1761, w_013_1762, w_013_1763, w_013_1764, w_013_1766, w_013_1767, w_013_1768, w_013_1770, w_013_1771, w_013_1772, w_013_1773, w_013_1774, w_013_1775, w_013_1776, w_013_1777, w_013_1779, w_013_1780, w_013_1784, w_013_1785, w_013_1787, w_013_1788, w_013_1791, w_013_1792, w_013_1793, w_013_1795, w_013_1796, w_013_1798, w_013_1799, w_013_1800, w_013_1801, w_013_1802, w_013_1803, w_013_1804, w_013_1805, w_013_1806, w_013_1807, w_013_1808, w_013_1809, w_013_1813, w_013_1814, w_013_1815, w_013_1817, w_013_1818, w_013_1819, w_013_1820, w_013_1821, w_013_1822, w_013_1823, w_013_1825, w_013_1826, w_013_1827, w_013_1828, w_013_1829, w_013_1830, w_013_1831, w_013_1833, w_013_1834, w_013_1835, w_013_1836, w_013_1837, w_013_1838, w_013_1839, w_013_1840, w_013_1841, w_013_1843, w_013_1845, w_013_1846, w_013_1847, w_013_1848, w_013_1849, w_013_1853, w_013_1854, w_013_1855, w_013_1856, w_013_1857, w_013_1858, w_013_1859, w_013_1860, w_013_1861, w_013_1862, w_013_1863, w_013_1864, w_013_1865, w_013_1866, w_013_1867, w_013_1868, w_013_1870, w_013_1871, w_013_1873, w_013_1874, w_013_1875, w_013_1876, w_013_1878, w_013_1879, w_013_1880, w_013_1881, w_013_1882, w_013_1883, w_013_1884, w_013_1887, w_013_1888, w_013_1889, w_013_1890, w_013_1891, w_013_1892, w_013_1893, w_013_1894, w_013_1895, w_013_1896, w_013_1897, w_013_1898, w_013_1901, w_013_1902, w_013_1903, w_013_1905, w_013_1906, w_013_1907, w_013_1909, w_013_1910, w_013_1914, w_013_1915, w_013_1917, w_013_1918, w_013_1919, w_013_1920, w_013_1921, w_013_1922, w_013_1923, w_013_1924, w_013_1925, w_013_1926, w_013_1930, w_013_1931, w_013_1932, w_013_1933, w_013_1934, w_013_1935, w_013_1936, w_013_1937, w_013_1938, w_013_1939, w_013_1940, w_013_1942, w_013_1944, w_013_1945, w_013_1946, w_013_1947, w_013_1949, w_013_1950, w_013_1951, w_013_1952, w_013_1953, w_013_1954, w_013_1955, w_013_1956, w_013_1958, w_013_1959, w_013_1960, w_013_1961, w_013_1962, w_013_1963, w_013_1964, w_013_1965, w_013_1966, w_013_1967, w_013_1968, w_013_1969, w_013_1971, w_013_1973, w_013_1975, w_013_1976, w_013_1977, w_013_1978, w_013_1979, w_013_1980, w_013_1982, w_013_1983, w_013_1984, w_013_1986, w_013_1987, w_013_1989, w_013_1990, w_013_1991, w_013_1992, w_013_1993, w_013_1995, w_013_1996, w_013_1997, w_013_1998, w_013_1999, w_013_2000, w_013_2001, w_013_2002, w_013_2003, w_013_2005, w_013_2006, w_013_2007, w_013_2009, w_013_2010, w_013_2011, w_013_2012, w_013_2014, w_013_2015, w_013_2016, w_013_2018, w_013_2020, w_013_2022, w_013_2023, w_013_2025, w_013_2026, w_013_2027, w_013_2028, w_013_2030, w_013_2031, w_013_2032, w_013_2033, w_013_2034, w_013_2035, w_013_2038, w_013_2039, w_013_2043, w_013_2044, w_013_2045, w_013_2046, w_013_2047, w_013_2048, w_013_2049, w_013_2050, w_013_2051, w_013_2053, w_013_2054, w_013_2056, w_013_2058, w_013_2059, w_013_2060, w_013_2062, w_013_2064, w_013_2065, w_013_2066, w_013_2067, w_013_2068, w_013_2069, w_013_2070, w_013_2071, w_013_2072, w_013_2073, w_013_2074, w_013_2075, w_013_2076, w_013_2077, w_013_2078, w_013_2079, w_013_2080, w_013_2081, w_013_2082, w_013_2084, w_013_2085, w_013_2086, w_013_2087, w_013_2089, w_013_2090, w_013_2091, w_013_2092, w_013_2093, w_013_2094, w_013_2095, w_013_2096, w_013_2099, w_013_2100, w_013_2101, w_013_2103, w_013_2104, w_013_2105, w_013_2106, w_013_2107, w_013_2109, w_013_2110, w_013_2111, w_013_2112, w_013_2113, w_013_2115, w_013_2117, w_013_2118, w_013_2120, w_013_2121, w_013_2122, w_013_2124, w_013_2125, w_013_2126, w_013_2127, w_013_2128, w_013_2130, w_013_2132, w_013_2133, w_013_2134, w_013_2135, w_013_2136, w_013_2137, w_013_2138, w_013_2139, w_013_2140, w_013_2141, w_013_2142, w_013_2143, w_013_2144, w_013_2145, w_013_2147, w_013_2148, w_013_2149, w_013_2150, w_013_2151, w_013_2152, w_013_2153, w_013_2155, w_013_2157, w_013_2159, w_013_2161, w_013_2162, w_013_2163, w_013_2165, w_013_2166, w_013_2167, w_013_2169, w_013_2170, w_013_2171, w_013_2172, w_013_2173, w_013_2174, w_013_2175, w_013_2176, w_013_2178, w_013_2179, w_013_2180, w_013_2181, w_013_2182, w_013_2183, w_013_2184, w_013_2187, w_013_2189, w_013_2190, w_013_2191, w_013_2192, w_013_2193, w_013_2194, w_013_2195, w_013_2196, w_013_2197, w_013_2198, w_013_2199, w_013_2200, w_013_2201, w_013_2202, w_013_2203, w_013_2204, w_013_2205, w_013_2206, w_013_2208, w_013_2209, w_013_2210, w_013_2211, w_013_2213, w_013_2214, w_013_2215, w_013_2216, w_013_2217, w_013_2219, w_013_2221, w_013_2222, w_013_2223, w_013_2224, w_013_2225, w_013_2226, w_013_2227, w_013_2228, w_013_2229, w_013_2230, w_013_2231, w_013_2232, w_013_2233, w_013_2234, w_013_2235, w_013_2236, w_013_2237, w_013_2238, w_013_2239, w_013_2241, w_013_2242, w_013_2243, w_013_2244, w_013_2245, w_013_2246, w_013_2247, w_013_2249, w_013_2250, w_013_2251, w_013_2253, w_013_2254, w_013_2255, w_013_2256, w_013_2258, w_013_2259, w_013_2260, w_013_2261, w_013_2262, w_013_2263, w_013_2264, w_013_2265, w_013_2268, w_013_2269, w_013_2270, w_013_2271, w_013_2272, w_013_2276, w_013_2277, w_013_2278, w_013_2279, w_013_2281, w_013_2282, w_013_2283, w_013_2284, w_013_2285, w_013_2286, w_013_2287, w_013_2288, w_013_2289, w_013_2290, w_013_2291, w_013_2292, w_013_2293, w_013_2294, w_013_2296, w_013_2297, w_013_2298, w_013_2299, w_013_2300, w_013_2301, w_013_2302, w_013_2303, w_013_2304, w_013_2305, w_013_2306, w_013_2308, w_013_2309, w_013_2311, w_013_2312, w_013_2313, w_013_2314, w_013_2315, w_013_2316, w_013_2317, w_013_2319, w_013_2320, w_013_2321, w_013_2323, w_013_2325, w_013_2326, w_013_2327, w_013_2328, w_013_2330, w_013_2332, w_013_2333, w_013_2334, w_013_2335, w_013_2336, w_013_2337, w_013_2338, w_013_2339, w_013_2340, w_013_2341, w_013_2342, w_013_2343, w_013_2344, w_013_2345, w_013_2346, w_013_2348, w_013_2349, w_013_2350, w_013_2351, w_013_2352, w_013_2353, w_013_2354, w_013_2355, w_013_2356, w_013_2357, w_013_2358, w_013_2359, w_013_2360, w_013_2361, w_013_2362, w_013_2363, w_013_2365, w_013_2367, w_013_2369, w_013_2370, w_013_2372, w_013_2373, w_013_2374, w_013_2375, w_013_2376, w_013_2378, w_013_2379, w_013_2381, w_013_2382, w_013_2383, w_013_2384, w_013_2385, w_013_2386, w_013_2388, w_013_2391, w_013_2392, w_013_2393, w_013_2394, w_013_2395, w_013_2396, w_013_2397, w_013_2398, w_013_2399, w_013_2401, w_013_2402, w_013_2403, w_013_2404, w_013_2405, w_013_2407, w_013_2408, w_013_2411, w_013_2413, w_013_2415, w_013_2417, w_013_2419, w_013_2420, w_013_2421, w_013_2423, w_013_2424, w_013_2425, w_013_2426, w_013_2428, w_013_2429, w_013_2430, w_013_2431, w_013_2432, w_013_2433, w_013_2434, w_013_2435, w_013_2436, w_013_2437, w_013_2438, w_013_2439, w_013_2440, w_013_2441, w_013_2442, w_013_2443, w_013_2445, w_013_2446, w_013_2447, w_013_2448, w_013_2449, w_013_2451, w_013_2452, w_013_2453, w_013_2454, w_013_2455, w_013_2456, w_013_2457, w_013_2458, w_013_2459, w_013_2461, w_013_2462, w_013_2463, w_013_2464, w_013_2465, w_013_2466, w_013_2467, w_013_2468, w_013_2469, w_013_2470, w_013_2474, w_013_2476, w_013_2477, w_013_2478, w_013_2479, w_013_2480, w_013_2481, w_013_2482, w_013_2483, w_013_2484, w_013_2485, w_013_2486, w_013_2487, w_013_2490, w_013_2492, w_013_2493, w_013_2494, w_013_2496, w_013_2497, w_013_2498, w_013_2499, w_013_2500, w_013_2501, w_013_2502, w_013_2504, w_013_2506, w_013_2507, w_013_2508, w_013_2509, w_013_2510, w_013_2512, w_013_2513, w_013_2514, w_013_2516, w_013_2517, w_013_2518, w_013_2519, w_013_2522, w_013_2523, w_013_2524, w_013_2526, w_013_2527, w_013_2529, w_013_2530, w_013_2531, w_013_2532, w_013_2533, w_013_2534, w_013_2535, w_013_2536, w_013_2537, w_013_2538, w_013_2539, w_013_2540, w_013_2541, w_013_2542, w_013_2543, w_013_2545, w_013_2547, w_013_2548, w_013_2549, w_013_2550, w_013_2551, w_013_2552, w_013_2553, w_013_2555, w_013_2556, w_013_2557, w_013_2559, w_013_2560, w_013_2563, w_013_2564, w_013_2565, w_013_2566, w_013_2567, w_013_2569, w_013_2570, w_013_2571, w_013_2572, w_013_2573, w_013_2574, w_013_2575, w_013_2576, w_013_2578, w_013_2579, w_013_2581, w_013_2582, w_013_2584, w_013_2585, w_013_2587, w_013_2590, w_013_2592, w_013_2593, w_013_2594, w_013_2595, w_013_2597, w_013_2598, w_013_2599, w_013_2600, w_013_2601, w_013_2602, w_013_2604, w_013_2605, w_013_2606, w_013_2607, w_013_2609, w_013_2611, w_013_2612, w_013_2613, w_013_2614, w_013_2615, w_013_2618, w_013_2619, w_013_2620, w_013_2621, w_013_2622, w_013_2624, w_013_2626, w_013_2627, w_013_2628, w_013_2630, w_013_2631, w_013_2632, w_013_2633, w_013_2636, w_013_2640, w_013_2642, w_013_2643, w_013_2644, w_013_2645, w_013_2646, w_013_2647, w_013_2649, w_013_2650, w_013_2651, w_013_2653, w_013_2654, w_013_2656, w_013_2657, w_013_2659, w_013_2660, w_013_2661, w_013_2662, w_013_2663, w_013_2664, w_013_2665, w_013_2666, w_013_2667, w_013_2668, w_013_2669, w_013_2670, w_013_2671, w_013_2673, w_013_2674, w_013_2675, w_013_2676, w_013_2677, w_013_2678, w_013_2680, w_013_2682, w_013_2683, w_013_2684, w_013_2685, w_013_2686, w_013_2687, w_013_2688, w_013_2690, w_013_2691, w_013_2692, w_013_2693, w_013_2694, w_013_2695, w_013_2697, w_013_2698, w_013_2699, w_013_2700, w_013_2701, w_013_2703, w_013_2704, w_013_2705, w_013_2706, w_013_2707, w_013_2708, w_013_2711, w_013_2712, w_013_2713, w_013_2714, w_013_2715, w_013_2716, w_013_2717, w_013_2718, w_013_2719, w_013_2720, w_013_2721, w_013_2722, w_013_2723, w_013_2724, w_013_2725, w_013_2726, w_013_2728, w_013_2730, w_013_2731, w_013_2732, w_013_2734, w_013_2736, w_013_2738, w_013_2739, w_013_2740, w_013_2741, w_013_2742, w_013_2743, w_013_2744, w_013_2745, w_013_2746, w_013_2748, w_013_2749, w_013_2750, w_013_2752, w_013_2753, w_013_2754, w_013_2755, w_013_2756, w_013_2757, w_013_2758, w_013_2759, w_013_2760, w_013_2761, w_013_2762, w_013_2763, w_013_2764, w_013_2765, w_013_2766, w_013_2767, w_013_2769, w_013_2770, w_013_2773, w_013_2774, w_013_2775, w_013_2776, w_013_2778, w_013_2779, w_013_2780, w_013_2781, w_013_2783, w_013_2784, w_013_2785, w_013_2787, w_013_2789, w_013_2790, w_013_2791, w_013_2792, w_013_2793, w_013_2795, w_013_2796, w_013_2797, w_013_2798, w_013_2799, w_013_2800, w_013_2801, w_013_2802, w_013_2803, w_013_2805, w_013_2806, w_013_2808, w_013_2809, w_013_2810, w_013_2811, w_013_2812, w_013_2813, w_013_2814, w_013_2815, w_013_2816, w_013_2818, w_013_2819, w_013_2820, w_013_2821, w_013_2822, w_013_2824, w_013_2825, w_013_2829, w_013_2831, w_013_2833, w_013_2835, w_013_2836, w_013_2837, w_013_2838, w_013_2839, w_013_2840, w_013_2842, w_013_2843, w_013_2844, w_013_2845, w_013_2846, w_013_2847, w_013_2848, w_013_2851, w_013_2852, w_013_2853, w_013_2854, w_013_2855, w_013_2856, w_013_2859, w_013_2861, w_013_2862, w_013_2863, w_013_2864, w_013_2865, w_013_2866, w_013_2867, w_013_2868, w_013_2869, w_013_2870, w_013_2872, w_013_2874, w_013_2878, w_013_2881, w_013_2882, w_013_2883, w_013_2884, w_013_2885, w_013_2888, w_013_2890, w_013_2891, w_013_2892, w_013_2893, w_013_2894, w_013_2895, w_013_2896, w_013_2897, w_013_2898, w_013_2900, w_013_2902, w_013_2903, w_013_2904, w_013_2907, w_013_2908, w_013_2909, w_013_2910, w_013_2912, w_013_2913, w_013_2915, w_013_2916, w_013_2917, w_013_2918, w_013_2919, w_013_2920, w_013_2921, w_013_2922, w_013_2925, w_013_2926, w_013_2927, w_013_2928, w_013_2930, w_013_2931, w_013_2932, w_013_2933, w_013_2934, w_013_2936, w_013_2937, w_013_2938, w_013_2941, w_013_2943, w_013_2944, w_013_2945, w_013_2946, w_013_2947, w_013_2948, w_013_2949, w_013_2950, w_013_2952, w_013_2953, w_013_2956, w_013_2957, w_013_2958, w_013_2959, w_013_2960, w_013_2961, w_013_2962, w_013_2963, w_013_2964, w_013_2965, w_013_2966, w_013_2967, w_013_2968, w_013_2969, w_013_2970, w_013_2971, w_013_2974, w_013_2975, w_013_2976, w_013_2977, w_013_2978, w_013_2979, w_013_2980, w_013_2982, w_013_2983, w_013_2984, w_013_2985, w_013_2986, w_013_2987, w_013_2991, w_013_2993, w_013_2994, w_013_2995, w_013_2996, w_013_2997, w_013_2999, w_013_3001, w_013_3002, w_013_3003, w_013_3006, w_013_3007, w_013_3008, w_013_3009, w_013_3010, w_013_3011, w_013_3012, w_013_3013, w_013_3014, w_013_3015, w_013_3016, w_013_3018, w_013_3019, w_013_3020, w_013_3021, w_013_3022, w_013_3023, w_013_3025, w_013_3026, w_013_3027, w_013_3028, w_013_3029, w_013_3030, w_013_3032, w_013_3034, w_013_3035, w_013_3036, w_013_3037, w_013_3038, w_013_3039, w_013_3041, w_013_3042, w_013_3043, w_013_3044, w_013_3045, w_013_3046, w_013_3047, w_013_3048, w_013_3049, w_013_3050, w_013_3051, w_013_3052, w_013_3053, w_013_3055, w_013_3056, w_013_3058, w_013_3059, w_013_3060, w_013_3061, w_013_3062, w_013_3063, w_013_3065, w_013_3067, w_013_3068, w_013_3069, w_013_3070, w_013_3071, w_013_3072, w_013_3074, w_013_3075, w_013_3076, w_013_3077, w_013_3079, w_013_3080, w_013_3084, w_013_3085, w_013_3087, w_013_3088, w_013_3091, w_013_3093, w_013_3094, w_013_3095, w_013_3096, w_013_3098, w_013_3100, w_013_3101, w_013_3102, w_013_3103, w_013_3105, w_013_3106, w_013_3107, w_013_3108, w_013_3109, w_013_3110, w_013_3111, w_013_3112, w_013_3113, w_013_3114, w_013_3115, w_013_3116, w_013_3117, w_013_3118, w_013_3119, w_013_3120, w_013_3121, w_013_3122, w_013_3123, w_013_3124, w_013_3127, w_013_3128, w_013_3129, w_013_3130, w_013_3132, w_013_3134, w_013_3137, w_013_3138, w_013_3139, w_013_3142, w_013_3143, w_013_3146, w_013_3147, w_013_3149, w_013_3150, w_013_3151, w_013_3152, w_013_3153, w_013_3154, w_013_3155, w_013_3156, w_013_3157, w_013_3158, w_013_3159, w_013_3160, w_013_3162, w_013_3163, w_013_3164, w_013_3165, w_013_3166, w_013_3168, w_013_3169, w_013_3170, w_013_3171, w_013_3176, w_013_3177, w_013_3178, w_013_3179, w_013_3181, w_013_3183, w_013_3186, w_013_3187, w_013_3190, w_013_3191, w_013_3192, w_013_3193, w_013_3195, w_013_3196, w_013_3198, w_013_3203, w_013_3204, w_013_3205, w_013_3206, w_013_3207, w_013_3210, w_013_3211, w_013_3212, w_013_3213, w_013_3214, w_013_3216, w_013_3217, w_013_3218, w_013_3219, w_013_3222, w_013_3226, w_013_3227, w_013_3228, w_013_3229, w_013_3230, w_013_3233, w_013_3234, w_013_3235, w_013_3236, w_013_3237, w_013_3238, w_013_3239, w_013_3240, w_013_3241, w_013_3242, w_013_3244, w_013_3245, w_013_3248, w_013_3249, w_013_3250, w_013_3251, w_013_3254, w_013_3255, w_013_3256, w_013_3257, w_013_3258, w_013_3259, w_013_3260, w_013_3261, w_013_3262, w_013_3263, w_013_3264, w_013_3265, w_013_3266, w_013_3267, w_013_3268, w_013_3270, w_013_3271, w_013_3272, w_013_3274, w_013_3275, w_013_3276, w_013_3277, w_013_3278, w_013_3279, w_013_3280, w_013_3281, w_013_3282, w_013_3284, w_013_3285, w_013_3286, w_013_3287, w_013_3288, w_013_3289, w_013_3290, w_013_3291, w_013_3292, w_013_3293, w_013_3294, w_013_3295, w_013_3296, w_013_3297, w_013_3298, w_013_3299, w_013_3300, w_013_3302, w_013_3303, w_013_3304, w_013_3305, w_013_3306, w_013_3308, w_013_3309, w_013_3310, w_013_3311, w_013_3312, w_013_3314, w_013_3315, w_013_3317, w_013_3319, w_013_3320, w_013_3321, w_013_3322, w_013_3323, w_013_3324, w_013_3326, w_013_3327, w_013_3330, w_013_3333, w_013_3334, w_013_3336, w_013_3337, w_013_3338, w_013_3339, w_013_3340, w_013_3341, w_013_3342, w_013_3347, w_013_3348, w_013_3350, w_013_3351, w_013_3352, w_013_3353, w_013_3355, w_013_3356, w_013_3358, w_013_3359, w_013_3361, w_013_3362, w_013_3363, w_013_3364, w_013_3365, w_013_3366, w_013_3367, w_013_3368, w_013_3369, w_013_3370, w_013_3371, w_013_3373, w_013_3374, w_013_3376, w_013_3377, w_013_3378, w_013_3379, w_013_3381, w_013_3384, w_013_3385, w_013_3386, w_013_3387, w_013_3388, w_013_3389, w_013_3390, w_013_3391, w_013_3393, w_013_3394, w_013_3395, w_013_3396, w_013_3397, w_013_3398, w_013_3399, w_013_3401, w_013_3403, w_013_3404, w_013_3405, w_013_3406, w_013_3407, w_013_3408, w_013_3409, w_013_3410, w_013_3412, w_013_3413, w_013_3415, w_013_3416, w_013_3417, w_013_3418, w_013_3419, w_013_3420, w_013_3422, w_013_3423, w_013_3424, w_013_3426, w_013_3427, w_013_3428, w_013_3429, w_013_3430, w_013_3431, w_013_3432, w_013_3433, w_013_3436, w_013_3437, w_013_3438, w_013_3439, w_013_3440, w_013_3441, w_013_3442, w_013_3443, w_013_3444, w_013_3445, w_013_3447, w_013_3448, w_013_3449, w_013_3450, w_013_3451, w_013_3452, w_013_3453, w_013_3454, w_013_3455, w_013_3456, w_013_3457, w_013_3458, w_013_3459, w_013_3460, w_013_3461, w_013_3462, w_013_3463, w_013_3464, w_013_3466, w_013_3468, w_013_3469, w_013_3470, w_013_3471, w_013_3472, w_013_3473, w_013_3474, w_013_3475, w_013_3476, w_013_3477, w_013_3479, w_013_3480, w_013_3481, w_013_3482, w_013_3483, w_013_3484, w_013_3485, w_013_3486, w_013_3487, w_013_3488, w_013_3490, w_013_3491, w_013_3492, w_013_3493, w_013_3494, w_013_3495, w_013_3497, w_013_3499, w_013_3500, w_013_3501, w_013_3502, w_013_3503, w_013_3505, w_013_3506, w_013_3508, w_013_3509, w_013_3510, w_013_3511, w_013_3512, w_013_3513, w_013_3514, w_013_3517, w_013_3518, w_013_3520, w_013_3521, w_013_3522, w_013_3523, w_013_3524, w_013_3525, w_013_3526, w_013_3527, w_013_3528, w_013_3529, w_013_3530, w_013_3531, w_013_3532, w_013_3533, w_013_3534, w_013_3537, w_013_3538, w_013_3539, w_013_3540, w_013_3541, w_013_3542, w_013_3543, w_013_3545, w_013_3546, w_013_3547, w_013_3548, w_013_3549, w_013_3551, w_013_3552, w_013_3553, w_013_3554, w_013_3555, w_013_3558, w_013_3559, w_013_3560, w_013_3561, w_013_3562, w_013_3563, w_013_3564, w_013_3565, w_013_3566, w_013_3567, w_013_3568, w_013_3569, w_013_3570, w_013_3571, w_013_3573, w_013_3574, w_013_3575, w_013_3576, w_013_3577, w_013_3578, w_013_3579, w_013_3580, w_013_3581, w_013_3583, w_013_3584, w_013_3586, w_013_3588, w_013_3590, w_013_3591, w_013_3592, w_013_3593, w_013_3594, w_013_3596, w_013_3597, w_013_3598, w_013_3599, w_013_3601, w_013_3602, w_013_3603, w_013_3604, w_013_3605, w_013_3606, w_013_3607, w_013_3608, w_013_3609, w_013_3610, w_013_3611, w_013_3612, w_013_3613, w_013_3614, w_013_3615, w_013_3617, w_013_3618, w_013_3619, w_013_3620, w_013_3622, w_013_3623, w_013_3625, w_013_3626, w_013_3627, w_013_3628, w_013_3629, w_013_3630, w_013_3632, w_013_3633, w_013_3634, w_013_3635, w_013_3636, w_013_3637, w_013_3638, w_013_3639, w_013_3640, w_013_3641, w_013_3642, w_013_3644, w_013_3647, w_013_3648, w_013_3649, w_013_3650, w_013_3651, w_013_3652, w_013_3653, w_013_3654;
  wire w_014_000, w_014_001, w_014_002, w_014_003, w_014_004, w_014_005, w_014_006, w_014_007, w_014_009, w_014_010, w_014_012, w_014_013, w_014_015, w_014_016, w_014_017, w_014_018, w_014_019, w_014_020, w_014_022, w_014_023, w_014_024, w_014_025, w_014_026, w_014_027, w_014_028, w_014_029, w_014_030, w_014_031, w_014_032, w_014_033, w_014_034, w_014_035, w_014_037, w_014_038, w_014_039, w_014_040, w_014_041, w_014_042, w_014_043, w_014_044, w_014_045, w_014_046, w_014_047, w_014_048, w_014_049, w_014_050, w_014_051, w_014_052, w_014_054, w_014_055, w_014_056, w_014_057, w_014_058, w_014_059, w_014_060, w_014_061, w_014_062, w_014_063, w_014_064, w_014_065, w_014_066, w_014_067, w_014_068, w_014_069, w_014_070, w_014_071, w_014_072, w_014_073, w_014_074, w_014_075, w_014_076, w_014_078, w_014_079, w_014_080, w_014_081, w_014_082, w_014_083, w_014_085, w_014_086, w_014_087, w_014_088, w_014_089, w_014_090, w_014_091, w_014_092, w_014_093, w_014_094, w_014_095, w_014_096, w_014_097, w_014_098, w_014_100, w_014_101, w_014_102, w_014_103, w_014_105, w_014_106, w_014_107, w_014_108, w_014_109, w_014_110, w_014_111, w_014_112, w_014_113, w_014_114, w_014_115, w_014_116, w_014_117, w_014_118, w_014_119, w_014_120, w_014_121, w_014_122, w_014_123, w_014_124, w_014_126, w_014_127, w_014_128, w_014_129, w_014_130, w_014_131, w_014_132, w_014_133, w_014_134, w_014_135, w_014_136, w_014_137, w_014_138, w_014_139, w_014_140, w_014_141, w_014_143, w_014_144, w_014_145, w_014_146, w_014_147, w_014_148, w_014_149, w_014_150, w_014_151, w_014_152, w_014_153, w_014_154, w_014_155, w_014_156, w_014_157, w_014_158, w_014_159, w_014_160, w_014_161, w_014_162, w_014_163, w_014_164, w_014_165, w_014_166, w_014_167, w_014_168, w_014_169, w_014_170, w_014_171, w_014_172, w_014_173, w_014_174, w_014_175, w_014_177, w_014_178, w_014_179, w_014_180, w_014_181, w_014_182, w_014_183, w_014_184, w_014_185, w_014_186, w_014_187, w_014_188, w_014_189, w_014_190, w_014_191, w_014_192, w_014_193, w_014_194, w_014_195, w_014_196, w_014_197, w_014_198, w_014_199, w_014_201, w_014_202, w_014_203, w_014_204, w_014_205, w_014_206, w_014_207, w_014_208, w_014_209, w_014_210, w_014_211, w_014_212, w_014_213, w_014_214, w_014_215, w_014_216, w_014_217, w_014_218, w_014_219, w_014_220, w_014_221, w_014_222, w_014_224, w_014_225, w_014_226, w_014_227, w_014_228, w_014_229, w_014_230, w_014_231, w_014_232, w_014_233, w_014_234, w_014_235, w_014_236, w_014_237, w_014_238, w_014_239, w_014_240, w_014_241, w_014_242, w_014_243, w_014_244, w_014_245, w_014_246, w_014_247, w_014_248, w_014_249, w_014_250, w_014_251, w_014_252, w_014_253, w_014_254, w_014_255, w_014_256, w_014_257, w_014_258, w_014_259, w_014_260, w_014_261, w_014_262, w_014_263, w_014_264, w_014_265, w_014_266, w_014_267, w_014_268, w_014_269, w_014_270, w_014_271, w_014_272, w_014_273, w_014_274, w_014_275, w_014_276, w_014_277, w_014_278, w_014_279, w_014_280, w_014_281, w_014_282, w_014_283, w_014_284, w_014_285, w_014_286, w_014_287, w_014_288, w_014_289, w_014_290, w_014_291, w_014_292, w_014_293, w_014_294, w_014_295, w_014_296, w_014_297, w_014_298, w_014_299, w_014_300, w_014_301, w_014_302, w_014_303, w_014_304, w_014_305, w_014_306, w_014_307, w_014_308, w_014_309, w_014_310, w_014_311, w_014_312, w_014_313, w_014_314, w_014_315, w_014_316, w_014_317, w_014_318, w_014_319, w_014_320, w_014_321, w_014_322, w_014_323, w_014_324, w_014_325, w_014_326, w_014_327, w_014_328, w_014_329, w_014_330, w_014_331, w_014_332, w_014_333, w_014_335, w_014_336, w_014_337, w_014_338, w_014_339, w_014_340, w_014_341, w_014_342, w_014_343, w_014_344, w_014_345, w_014_346, w_014_347, w_014_348, w_014_349, w_014_350, w_014_351, w_014_352, w_014_353, w_014_354, w_014_355, w_014_356, w_014_357, w_014_358, w_014_359, w_014_361, w_014_362, w_014_363, w_014_364, w_014_365, w_014_366, w_014_367, w_014_368, w_014_369, w_014_370, w_014_371, w_014_372, w_014_373, w_014_375, w_014_376, w_014_377, w_014_379, w_014_380, w_014_381, w_014_382, w_014_383, w_014_384, w_014_385, w_014_386, w_014_388, w_014_389, w_014_390, w_014_391, w_014_392, w_014_393, w_014_394, w_014_395, w_014_396, w_014_397, w_014_398, w_014_399, w_014_400, w_014_401, w_014_402, w_014_403, w_014_404, w_014_405, w_014_406, w_014_407, w_014_408, w_014_409, w_014_410, w_014_411, w_014_412, w_014_413, w_014_414, w_014_415, w_014_416, w_014_417, w_014_418, w_014_419, w_014_420, w_014_421, w_014_422, w_014_423, w_014_424, w_014_425, w_014_426, w_014_427, w_014_428, w_014_429, w_014_430, w_014_431, w_014_432, w_014_433, w_014_434, w_014_435, w_014_436, w_014_437, w_014_438, w_014_439, w_014_440, w_014_441, w_014_442, w_014_443, w_014_444, w_014_445, w_014_446, w_014_447, w_014_448, w_014_449, w_014_450, w_014_451, w_014_452, w_014_453, w_014_454, w_014_455, w_014_456, w_014_457, w_014_458, w_014_459, w_014_460, w_014_461, w_014_462, w_014_463, w_014_464, w_014_465, w_014_466, w_014_467, w_014_468, w_014_469, w_014_470, w_014_471, w_014_472, w_014_473, w_014_474, w_014_475, w_014_476, w_014_477, w_014_478, w_014_479, w_014_480, w_014_482, w_014_483, w_014_484, w_014_485, w_014_486, w_014_487, w_014_488, w_014_489, w_014_490, w_014_491, w_014_492, w_014_493, w_014_494, w_014_495, w_014_496, w_014_497, w_014_498, w_014_499, w_014_500, w_014_501, w_014_502, w_014_503, w_014_504, w_014_505, w_014_506, w_014_507, w_014_508, w_014_510, w_014_511, w_014_512, w_014_513, w_014_514, w_014_515, w_014_516, w_014_518, w_014_519, w_014_520, w_014_521, w_014_522, w_014_523, w_014_524, w_014_525, w_014_526, w_014_527, w_014_528, w_014_529, w_014_530, w_014_531, w_014_532, w_014_533, w_014_535, w_014_536, w_014_537, w_014_538, w_014_539, w_014_540, w_014_541, w_014_542, w_014_543, w_014_544, w_014_546, w_014_547, w_014_549, w_014_550, w_014_551, w_014_552, w_014_553, w_014_554, w_014_555, w_014_556, w_014_557, w_014_558, w_014_559, w_014_560, w_014_561, w_014_562, w_014_563, w_014_564, w_014_565, w_014_566, w_014_567, w_014_568, w_014_569, w_014_570, w_014_571, w_014_572, w_014_573, w_014_574, w_014_575, w_014_576, w_014_577, w_014_578, w_014_579, w_014_580, w_014_581, w_014_582, w_014_583, w_014_584, w_014_585, w_014_586, w_014_587, w_014_588, w_014_589, w_014_590, w_014_592, w_014_593, w_014_594, w_014_595, w_014_596, w_014_598, w_014_599, w_014_600, w_014_601, w_014_602, w_014_603, w_014_604, w_014_605, w_014_606, w_014_607, w_014_608, w_014_609, w_014_610, w_014_611, w_014_612, w_014_613, w_014_614, w_014_615, w_014_616, w_014_617, w_014_618, w_014_619, w_014_620, w_014_621, w_014_622, w_014_623, w_014_624, w_014_625, w_014_626, w_014_627, w_014_628, w_014_629, w_014_630, w_014_631, w_014_632, w_014_633, w_014_634, w_014_635, w_014_636, w_014_637, w_014_639, w_014_640, w_014_641, w_014_642, w_014_643, w_014_644, w_014_646, w_014_647, w_014_648, w_014_649, w_014_650, w_014_651, w_014_652, w_014_653, w_014_654, w_014_655, w_014_656, w_014_657, w_014_658, w_014_659, w_014_660, w_014_661, w_014_662, w_014_663, w_014_664, w_014_665, w_014_666, w_014_667, w_014_669, w_014_670, w_014_671, w_014_672, w_014_673, w_014_674, w_014_675, w_014_676, w_014_677, w_014_678, w_014_679, w_014_680, w_014_681, w_014_682, w_014_683, w_014_684, w_014_685, w_014_686, w_014_687, w_014_688, w_014_689, w_014_690, w_014_691, w_014_693, w_014_694, w_014_695, w_014_696, w_014_697, w_014_698, w_014_699, w_014_700, w_014_701, w_014_702, w_014_703, w_014_704, w_014_705, w_014_706, w_014_707, w_014_708, w_014_709, w_014_710, w_014_711, w_014_712, w_014_713, w_014_714, w_014_715, w_014_716, w_014_717, w_014_718, w_014_719, w_014_720, w_014_721, w_014_722, w_014_723, w_014_724, w_014_725, w_014_726, w_014_727, w_014_728, w_014_729, w_014_730, w_014_732, w_014_733, w_014_734, w_014_735, w_014_736, w_014_737, w_014_739, w_014_740, w_014_741, w_014_742, w_014_743, w_014_744, w_014_745, w_014_746, w_014_747, w_014_748, w_014_749, w_014_750, w_014_751, w_014_752, w_014_753, w_014_754, w_014_755, w_014_756, w_014_757, w_014_759, w_014_760, w_014_761, w_014_762, w_014_763, w_014_764, w_014_765, w_014_766, w_014_767, w_014_768, w_014_769, w_014_770, w_014_771, w_014_772, w_014_773, w_014_774, w_014_775, w_014_776, w_014_777, w_014_778, w_014_779, w_014_780, w_014_781, w_014_782, w_014_783, w_014_784, w_014_785, w_014_786, w_014_787, w_014_788, w_014_789, w_014_791, w_014_792, w_014_794, w_014_795, w_014_796, w_014_797, w_014_798, w_014_799, w_014_800, w_014_801, w_014_802, w_014_803, w_014_804, w_014_805, w_014_806, w_014_807, w_014_808, w_014_809, w_014_810, w_014_811, w_014_812, w_014_813, w_014_814, w_014_815, w_014_816, w_014_817, w_014_818, w_014_819, w_014_820, w_014_821, w_014_823, w_014_824, w_014_825, w_014_826, w_014_827, w_014_828, w_014_829, w_014_830, w_014_831, w_014_832, w_014_833, w_014_834, w_014_835, w_014_836, w_014_837, w_014_838, w_014_839, w_014_840, w_014_841, w_014_842, w_014_843, w_014_844, w_014_845, w_014_846, w_014_847, w_014_848, w_014_849, w_014_850, w_014_851, w_014_852, w_014_853, w_014_854, w_014_855, w_014_856, w_014_857, w_014_858, w_014_859, w_014_860, w_014_861, w_014_862, w_014_863, w_014_864, w_014_865, w_014_866, w_014_867, w_014_868, w_014_869, w_014_870, w_014_871, w_014_872, w_014_873, w_014_874, w_014_875, w_014_876, w_014_877, w_014_878, w_014_879, w_014_880, w_014_881, w_014_882, w_014_883, w_014_884, w_014_885, w_014_886, w_014_887, w_014_888, w_014_889, w_014_890, w_014_891, w_014_892, w_014_893, w_014_894, w_014_895, w_014_897, w_014_898, w_014_899, w_014_900, w_014_901, w_014_902, w_014_904, w_014_905, w_014_906, w_014_907, w_014_908, w_014_909, w_014_910, w_014_911, w_014_912, w_014_913, w_014_914, w_014_915, w_014_916, w_014_917, w_014_918, w_014_920, w_014_921, w_014_922, w_014_923, w_014_924, w_014_925, w_014_926, w_014_927, w_014_928, w_014_929, w_014_930, w_014_931, w_014_932, w_014_933, w_014_934, w_014_935, w_014_936, w_014_937, w_014_938, w_014_939, w_014_940, w_014_941, w_014_942, w_014_943, w_014_944, w_014_945, w_014_946, w_014_947, w_014_948, w_014_949, w_014_951, w_014_952, w_014_953, w_014_954, w_014_955, w_014_956, w_014_957, w_014_958, w_014_959, w_014_961, w_014_963, w_014_964, w_014_966, w_014_967, w_014_968, w_014_969, w_014_970, w_014_971, w_014_972, w_014_973, w_014_974, w_014_975, w_014_976, w_014_977, w_014_978, w_014_979, w_014_980, w_014_981, w_014_982, w_014_983, w_014_984, w_014_985, w_014_986, w_014_987, w_014_988, w_014_989, w_014_990, w_014_991, w_014_992, w_014_993, w_014_994, w_014_995, w_014_996, w_014_997, w_014_998, w_014_999, w_014_1000, w_014_1001, w_014_1002, w_014_1003, w_014_1004, w_014_1005, w_014_1006, w_014_1007, w_014_1008, w_014_1009, w_014_1010, w_014_1011, w_014_1012, w_014_1013, w_014_1014, w_014_1015, w_014_1016, w_014_1017, w_014_1018, w_014_1019, w_014_1020, w_014_1021, w_014_1022, w_014_1023, w_014_1024, w_014_1026, w_014_1027, w_014_1028, w_014_1029, w_014_1030, w_014_1031, w_014_1032, w_014_1033, w_014_1034, w_014_1035, w_014_1036, w_014_1037, w_014_1038, w_014_1039, w_014_1040, w_014_1041, w_014_1042, w_014_1043, w_014_1044, w_014_1045, w_014_1046, w_014_1047, w_014_1048, w_014_1049, w_014_1050, w_014_1052, w_014_1053, w_014_1054, w_014_1055, w_014_1056, w_014_1057, w_014_1058, w_014_1059, w_014_1060, w_014_1061, w_014_1062, w_014_1063, w_014_1064, w_014_1065, w_014_1066, w_014_1067, w_014_1068, w_014_1070, w_014_1071, w_014_1072, w_014_1073, w_014_1074, w_014_1075, w_014_1076, w_014_1077, w_014_1078, w_014_1079, w_014_1081, w_014_1082, w_014_1083, w_014_1084, w_014_1085, w_014_1086, w_014_1087, w_014_1088, w_014_1089, w_014_1090, w_014_1091, w_014_1092, w_014_1093, w_014_1094, w_014_1095, w_014_1096, w_014_1098, w_014_1100, w_014_1101, w_014_1102, w_014_1103, w_014_1104, w_014_1105, w_014_1106, w_014_1107, w_014_1108, w_014_1109, w_014_1110, w_014_1111, w_014_1112, w_014_1113, w_014_1114, w_014_1115, w_014_1116, w_014_1117, w_014_1119, w_014_1120, w_014_1121, w_014_1122, w_014_1123, w_014_1124, w_014_1126, w_014_1127, w_014_1128, w_014_1129, w_014_1130, w_014_1131, w_014_1132, w_014_1133, w_014_1135, w_014_1136, w_014_1138, w_014_1139, w_014_1140, w_014_1141, w_014_1143, w_014_1144, w_014_1145, w_014_1146, w_014_1147, w_014_1148, w_014_1149, w_014_1150, w_014_1151, w_014_1152, w_014_1153, w_014_1154, w_014_1156, w_014_1157, w_014_1158, w_014_1159, w_014_1160, w_014_1161, w_014_1162, w_014_1163, w_014_1164, w_014_1165, w_014_1166, w_014_1167, w_014_1168, w_014_1169, w_014_1170, w_014_1171, w_014_1172, w_014_1173, w_014_1174, w_014_1175, w_014_1176, w_014_1177, w_014_1178, w_014_1179, w_014_1180, w_014_1181, w_014_1182, w_014_1183, w_014_1184, w_014_1185, w_014_1186, w_014_1187, w_014_1188, w_014_1189, w_014_1190, w_014_1191, w_014_1192, w_014_1193, w_014_1194, w_014_1195, w_014_1196, w_014_1197, w_014_1198, w_014_1199, w_014_1200, w_014_1201, w_014_1202, w_014_1203, w_014_1204, w_014_1205, w_014_1206, w_014_1207, w_014_1208, w_014_1209, w_014_1210, w_014_1211, w_014_1212, w_014_1213, w_014_1214, w_014_1215, w_014_1216, w_014_1217, w_014_1218, w_014_1219, w_014_1220, w_014_1221, w_014_1222, w_014_1223, w_014_1225, w_014_1226, w_014_1227, w_014_1228, w_014_1229, w_014_1230, w_014_1232, w_014_1233, w_014_1234, w_014_1235, w_014_1236, w_014_1237, w_014_1238, w_014_1239, w_014_1240, w_014_1241, w_014_1242, w_014_1243, w_014_1244, w_014_1245, w_014_1246, w_014_1247, w_014_1248, w_014_1249, w_014_1250, w_014_1251, w_014_1252, w_014_1253, w_014_1254, w_014_1255, w_014_1256, w_014_1257, w_014_1258, w_014_1259, w_014_1260, w_014_1261, w_014_1262, w_014_1263, w_014_1264, w_014_1265, w_014_1266, w_014_1267, w_014_1268, w_014_1269, w_014_1270, w_014_1272, w_014_1273, w_014_1274, w_014_1275, w_014_1276, w_014_1277, w_014_1278, w_014_1279, w_014_1280, w_014_1281, w_014_1282, w_014_1283, w_014_1284, w_014_1285, w_014_1286, w_014_1288, w_014_1289, w_014_1290, w_014_1291, w_014_1292, w_014_1294, w_014_1295, w_014_1297, w_014_1298, w_014_1299, w_014_1300, w_014_1301, w_014_1302, w_014_1303, w_014_1305, w_014_1306, w_014_1307, w_014_1308, w_014_1309, w_014_1310, w_014_1311, w_014_1312, w_014_1313, w_014_1314, w_014_1315, w_014_1316, w_014_1317, w_014_1318, w_014_1319, w_014_1320, w_014_1321, w_014_1322, w_014_1323, w_014_1324, w_014_1325, w_014_1326, w_014_1327, w_014_1328, w_014_1329, w_014_1330, w_014_1331, w_014_1332, w_014_1334, w_014_1335, w_014_1336, w_014_1337, w_014_1338, w_014_1340, w_014_1341, w_014_1342, w_014_1343, w_014_1345, w_014_1347, w_014_1348, w_014_1349, w_014_1350, w_014_1351, w_014_1352, w_014_1353, w_014_1354, w_014_1355, w_014_1356, w_014_1357, w_014_1358, w_014_1359, w_014_1360, w_014_1361, w_014_1362, w_014_1363, w_014_1364, w_014_1365, w_014_1366, w_014_1368, w_014_1369, w_014_1370, w_014_1371, w_014_1372, w_014_1373, w_014_1374, w_014_1375, w_014_1376, w_014_1377, w_014_1378, w_014_1379, w_014_1381, w_014_1383, w_014_1384, w_014_1385, w_014_1386, w_014_1387, w_014_1388, w_014_1389, w_014_1390, w_014_1391, w_014_1392, w_014_1393, w_014_1394, w_014_1395, w_014_1396, w_014_1397, w_014_1398, w_014_1399, w_014_1400, w_014_1401, w_014_1402, w_014_1403, w_014_1404, w_014_1405, w_014_1406, w_014_1407, w_014_1408, w_014_1409, w_014_1410, w_014_1411, w_014_1412, w_014_1413, w_014_1414, w_014_1415, w_014_1416, w_014_1417, w_014_1418, w_014_1419, w_014_1420, w_014_1421, w_014_1422, w_014_1423, w_014_1424, w_014_1426, w_014_1427, w_014_1428, w_014_1429, w_014_1430, w_014_1431, w_014_1432, w_014_1433, w_014_1434, w_014_1435, w_014_1436, w_014_1437, w_014_1438, w_014_1439, w_014_1440, w_014_1441, w_014_1442, w_014_1443, w_014_1444, w_014_1445, w_014_1446, w_014_1447, w_014_1448, w_014_1449, w_014_1450, w_014_1451, w_014_1452, w_014_1453, w_014_1454, w_014_1455, w_014_1456, w_014_1457, w_014_1458, w_014_1459, w_014_1460, w_014_1461, w_014_1462, w_014_1463, w_014_1465, w_014_1466, w_014_1467, w_014_1468, w_014_1469, w_014_1470, w_014_1471, w_014_1472, w_014_1473, w_014_1474, w_014_1475, w_014_1476, w_014_1477, w_014_1478, w_014_1479, w_014_1480, w_014_1481, w_014_1482, w_014_1483, w_014_1484, w_014_1485, w_014_1486, w_014_1487, w_014_1488, w_014_1489, w_014_1490, w_014_1491, w_014_1492, w_014_1493, w_014_1494, w_014_1495, w_014_1496, w_014_1497, w_014_1498, w_014_1499, w_014_1500, w_014_1501, w_014_1502, w_014_1503, w_014_1504, w_014_1505, w_014_1506, w_014_1507, w_014_1508, w_014_1509, w_014_1510, w_014_1511, w_014_1512, w_014_1513, w_014_1514, w_014_1515, w_014_1516, w_014_1517, w_014_1518, w_014_1519, w_014_1520, w_014_1521, w_014_1522, w_014_1523, w_014_1524, w_014_1525, w_014_1526, w_014_1527, w_014_1529, w_014_1530, w_014_1531, w_014_1532, w_014_1533, w_014_1534, w_014_1535, w_014_1536, w_014_1537, w_014_1538, w_014_1539, w_014_1540, w_014_1541, w_014_1542, w_014_1543, w_014_1544, w_014_1545, w_014_1546, w_014_1547, w_014_1548, w_014_1549, w_014_1550, w_014_1551, w_014_1552, w_014_1553, w_014_1554, w_014_1555, w_014_1556, w_014_1557, w_014_1558, w_014_1559, w_014_1560, w_014_1561, w_014_1562, w_014_1564, w_014_1565, w_014_1567, w_014_1568, w_014_1569, w_014_1570, w_014_1571, w_014_1572, w_014_1573, w_014_1574, w_014_1575, w_014_1576, w_014_1577, w_014_1578, w_014_1579, w_014_1580, w_014_1581, w_014_1582, w_014_1584, w_014_1585, w_014_1586, w_014_1587, w_014_1588, w_014_1589, w_014_1590, w_014_1591, w_014_1592, w_014_1593, w_014_1594, w_014_1595, w_014_1596, w_014_1597, w_014_1598, w_014_1599, w_014_1600, w_014_1601, w_014_1602, w_014_1603, w_014_1604, w_014_1605, w_014_1606, w_014_1607, w_014_1608, w_014_1609, w_014_1610, w_014_1611, w_014_1612, w_014_1613, w_014_1614, w_014_1615, w_014_1616, w_014_1617, w_014_1618, w_014_1619, w_014_1621, w_014_1622, w_014_1623, w_014_1624, w_014_1625, w_014_1626, w_014_1627, w_014_1628, w_014_1629, w_014_1630, w_014_1631, w_014_1632, w_014_1633, w_014_1634, w_014_1635, w_014_1636, w_014_1637, w_014_1638, w_014_1639, w_014_1640, w_014_1641, w_014_1642, w_014_1643, w_014_1644, w_014_1645, w_014_1646, w_014_1647, w_014_1648, w_014_1649, w_014_1650, w_014_1651, w_014_1652, w_014_1653, w_014_1654, w_014_1655, w_014_1656, w_014_1657, w_014_1658, w_014_1659, w_014_1660, w_014_1661, w_014_1662, w_014_1663, w_014_1664, w_014_1665, w_014_1666, w_014_1667, w_014_1668, w_014_1669, w_014_1670, w_014_1671, w_014_1672, w_014_1673, w_014_1674, w_014_1675, w_014_1676, w_014_1677, w_014_1678, w_014_1679, w_014_1680, w_014_1681, w_014_1682, w_014_1683, w_014_1684, w_014_1685, w_014_1686, w_014_1687, w_014_1688, w_014_1690, w_014_1691, w_014_1692, w_014_1694, w_014_1695, w_014_1696, w_014_1697, w_014_1698, w_014_1699, w_014_1700, w_014_1701, w_014_1703, w_014_1704, w_014_1705, w_014_1706, w_014_1707, w_014_1708, w_014_1709, w_014_1710, w_014_1711, w_014_1712, w_014_1713, w_014_1714, w_014_1715, w_014_1716, w_014_1717, w_014_1718, w_014_1719, w_014_1720, w_014_1721, w_014_1722, w_014_1723, w_014_1724, w_014_1725, w_014_1727, w_014_1728, w_014_1729, w_014_1730, w_014_1731, w_014_1732, w_014_1733, w_014_1734, w_014_1735, w_014_1736, w_014_1737, w_014_1738, w_014_1739, w_014_1740, w_014_1741, w_014_1742, w_014_1743, w_014_1744, w_014_1745, w_014_1746, w_014_1747, w_014_1748, w_014_1749, w_014_1750, w_014_1751, w_014_1752, w_014_1753, w_014_1754, w_014_1755, w_014_1756, w_014_1759, w_014_1760, w_014_1761, w_014_1762, w_014_1763, w_014_1764, w_014_1765, w_014_1766, w_014_1767, w_014_1768, w_014_1769, w_014_1770, w_014_1771, w_014_1772, w_014_1773, w_014_1774, w_014_1775, w_014_1776, w_014_1777, w_014_1778, w_014_1779, w_014_1780, w_014_1781, w_014_1782, w_014_1783, w_014_1784, w_014_1785, w_014_1786, w_014_1788, w_014_1789, w_014_1790, w_014_1791, w_014_1792, w_014_1793, w_014_1794, w_014_1796, w_014_1797, w_014_1798, w_014_1801, w_014_1802, w_014_1803, w_014_1804, w_014_1805, w_014_1806, w_014_1807, w_014_1808, w_014_1809, w_014_1811, w_014_1813, w_014_1815, w_014_1816, w_014_1817, w_014_1818, w_014_1819, w_014_1820, w_014_1821, w_014_1822, w_014_1823, w_014_1824, w_014_1825, w_014_1826, w_014_1828, w_014_1829, w_014_1830, w_014_1832, w_014_1833, w_014_1834, w_014_1836, w_014_1837, w_014_1839, w_014_1840, w_014_1841, w_014_1843, w_014_1844, w_014_1845, w_014_1846, w_014_1848, w_014_1849, w_014_1850, w_014_1852, w_014_1853, w_014_1855, w_014_1858, w_014_1859, w_014_1860, w_014_1863, w_014_1864, w_014_1866, w_014_1867, w_014_1868, w_014_1869, w_014_1870, w_014_1872, w_014_1874, w_014_1875, w_014_1876, w_014_1877, w_014_1878, w_014_1879, w_014_1880, w_014_1881, w_014_1882, w_014_1883, w_014_1884, w_014_1885, w_014_1886, w_014_1887, w_014_1889, w_014_1890, w_014_1891, w_014_1892, w_014_1893, w_014_1894, w_014_1895, w_014_1896, w_014_1897, w_014_1898, w_014_1899, w_014_1900, w_014_1901, w_014_1904, w_014_1905, w_014_1907, w_014_1908, w_014_1909, w_014_1910, w_014_1912, w_014_1914, w_014_1915, w_014_1916, w_014_1919, w_014_1920, w_014_1921, w_014_1922, w_014_1923, w_014_1924, w_014_1925, w_014_1926, w_014_1928, w_014_1929, w_014_1930, w_014_1931, w_014_1932, w_014_1933, w_014_1934, w_014_1935, w_014_1936, w_014_1937, w_014_1939, w_014_1940, w_014_1941, w_014_1942, w_014_1944, w_014_1945, w_014_1946, w_014_1948, w_014_1950, w_014_1951, w_014_1952, w_014_1953, w_014_1954, w_014_1955, w_014_1956, w_014_1957, w_014_1958, w_014_1959, w_014_1960, w_014_1961, w_014_1962, w_014_1963, w_014_1964, w_014_1966, w_014_1967, w_014_1968, w_014_1970, w_014_1971, w_014_1972, w_014_1975, w_014_1976, w_014_1977, w_014_1978, w_014_1979, w_014_1980, w_014_1981, w_014_1982, w_014_1983, w_014_1984, w_014_1985, w_014_1987, w_014_1988, w_014_1990, w_014_1991, w_014_1992, w_014_1993, w_014_1994, w_014_1995, w_014_1996, w_014_1997, w_014_2000, w_014_2001, w_014_2002, w_014_2003, w_014_2004, w_014_2005, w_014_2006, w_014_2007, w_014_2008, w_014_2009, w_014_2010, w_014_2011, w_014_2012, w_014_2013, w_014_2015, w_014_2016, w_014_2017, w_014_2018, w_014_2019, w_014_2020, w_014_2021, w_014_2023, w_014_2024, w_014_2025, w_014_2026, w_014_2028, w_014_2030, w_014_2031, w_014_2032, w_014_2033, w_014_2034, w_014_2035, w_014_2036, w_014_2037, w_014_2038, w_014_2039, w_014_2040, w_014_2042, w_014_2043, w_014_2045, w_014_2046, w_014_2047, w_014_2048, w_014_2049, w_014_2051, w_014_2052, w_014_2053, w_014_2055, w_014_2056, w_014_2057, w_014_2058, w_014_2059, w_014_2060, w_014_2061, w_014_2065, w_014_2066, w_014_2068, w_014_2069, w_014_2070, w_014_2072, w_014_2074, w_014_2075, w_014_2076, w_014_2077, w_014_2078, w_014_2080, w_014_2081, w_014_2082, w_014_2083, w_014_2084, w_014_2086, w_014_2087, w_014_2088, w_014_2090, w_014_2091, w_014_2092, w_014_2093, w_014_2094, w_014_2095, w_014_2096, w_014_2097, w_014_2098, w_014_2099, w_014_2100, w_014_2101, w_014_2102, w_014_2103, w_014_2105, w_014_2106, w_014_2107, w_014_2109, w_014_2110, w_014_2111, w_014_2113, w_014_2114, w_014_2116, w_014_2117, w_014_2118, w_014_2119, w_014_2122, w_014_2123, w_014_2125, w_014_2126, w_014_2127, w_014_2128, w_014_2131, w_014_2132, w_014_2133, w_014_2134, w_014_2137, w_014_2138, w_014_2139, w_014_2140, w_014_2141, w_014_2143, w_014_2144, w_014_2145, w_014_2146, w_014_2147, w_014_2148, w_014_2149, w_014_2150, w_014_2151, w_014_2153, w_014_2154, w_014_2155, w_014_2156, w_014_2157, w_014_2158, w_014_2159, w_014_2160, w_014_2161, w_014_2162, w_014_2163, w_014_2165, w_014_2168, w_014_2169, w_014_2170, w_014_2171, w_014_2173, w_014_2174, w_014_2176, w_014_2177, w_014_2179, w_014_2180, w_014_2181, w_014_2183, w_014_2185, w_014_2186, w_014_2187, w_014_2189, w_014_2190, w_014_2191, w_014_2192, w_014_2193, w_014_2195, w_014_2196, w_014_2200, w_014_2201, w_014_2202, w_014_2203, w_014_2204, w_014_2206, w_014_2207, w_014_2209, w_014_2210, w_014_2211, w_014_2212, w_014_2213, w_014_2214, w_014_2217, w_014_2220, w_014_2221, w_014_2222, w_014_2223, w_014_2224, w_014_2225, w_014_2226, w_014_2227, w_014_2228, w_014_2229, w_014_2231, w_014_2232, w_014_2233, w_014_2235, w_014_2236, w_014_2239, w_014_2240, w_014_2241, w_014_2242, w_014_2243, w_014_2244, w_014_2245, w_014_2246, w_014_2247, w_014_2250, w_014_2251, w_014_2252, w_014_2253, w_014_2254, w_014_2256, w_014_2257, w_014_2258, w_014_2260, w_014_2261, w_014_2263, w_014_2264, w_014_2265, w_014_2267, w_014_2270, w_014_2271, w_014_2274, w_014_2275, w_014_2276, w_014_2277, w_014_2278, w_014_2279, w_014_2282, w_014_2283, w_014_2284, w_014_2286, w_014_2287, w_014_2288, w_014_2290, w_014_2292, w_014_2293, w_014_2296, w_014_2298, w_014_2299, w_014_2301, w_014_2302, w_014_2303, w_014_2306, w_014_2307, w_014_2308, w_014_2311, w_014_2312, w_014_2314, w_014_2315, w_014_2316, w_014_2317, w_014_2318, w_014_2319, w_014_2320, w_014_2321, w_014_2322, w_014_2325, w_014_2326, w_014_2327, w_014_2328, w_014_2330, w_014_2331, w_014_2332, w_014_2334, w_014_2335, w_014_2336, w_014_2337, w_014_2338, w_014_2339, w_014_2341, w_014_2342, w_014_2343, w_014_2344, w_014_2345, w_014_2347, w_014_2348, w_014_2349, w_014_2350, w_014_2351, w_014_2352, w_014_2354, w_014_2355, w_014_2357, w_014_2358, w_014_2359, w_014_2360, w_014_2361, w_014_2362, w_014_2363, w_014_2364, w_014_2366, w_014_2368, w_014_2369, w_014_2370, w_014_2371, w_014_2374, w_014_2375, w_014_2376, w_014_2377, w_014_2379, w_014_2380, w_014_2382, w_014_2383, w_014_2384, w_014_2387, w_014_2388, w_014_2389, w_014_2390, w_014_2391, w_014_2392, w_014_2394, w_014_2396, w_014_2397, w_014_2398, w_014_2399, w_014_2402, w_014_2403, w_014_2404, w_014_2405, w_014_2406, w_014_2407, w_014_2409, w_014_2412, w_014_2413, w_014_2414, w_014_2415, w_014_2416, w_014_2417, w_014_2418, w_014_2419, w_014_2420, w_014_2421, w_014_2422, w_014_2423, w_014_2425, w_014_2427, w_014_2429, w_014_2430, w_014_2431, w_014_2432, w_014_2435, w_014_2437, w_014_2438, w_014_2440, w_014_2441, w_014_2442, w_014_2443, w_014_2444, w_014_2445, w_014_2448, w_014_2449, w_014_2451, w_014_2454, w_014_2455, w_014_2456, w_014_2457, w_014_2458, w_014_2459, w_014_2460, w_014_2461, w_014_2462, w_014_2464, w_014_2465, w_014_2466, w_014_2467, w_014_2468, w_014_2469, w_014_2471, w_014_2473, w_014_2474, w_014_2475, w_014_2476, w_014_2477, w_014_2478, w_014_2479, w_014_2480, w_014_2481, w_014_2483, w_014_2484, w_014_2485, w_014_2486, w_014_2487, w_014_2488, w_014_2489, w_014_2490, w_014_2491, w_014_2492, w_014_2495, w_014_2497, w_014_2498, w_014_2499, w_014_2500, w_014_2501, w_014_2502, w_014_2503, w_014_2505, w_014_2506, w_014_2507, w_014_2508, w_014_2509, w_014_2512, w_014_2513, w_014_2514, w_014_2515, w_014_2516, w_014_2517, w_014_2518, w_014_2519, w_014_2520, w_014_2521, w_014_2524, w_014_2525, w_014_2526, w_014_2527, w_014_2528, w_014_2530, w_014_2531, w_014_2532, w_014_2533, w_014_2534, w_014_2536, w_014_2537, w_014_2538, w_014_2539, w_014_2540, w_014_2541, w_014_2543, w_014_2545, w_014_2546, w_014_2547, w_014_2549, w_014_2550, w_014_2551, w_014_2553, w_014_2556, w_014_2557, w_014_2559, w_014_2560, w_014_2561, w_014_2562, w_014_2565, w_014_2566, w_014_2567, w_014_2571, w_014_2572, w_014_2573, w_014_2574, w_014_2575, w_014_2577, w_014_2578, w_014_2580, w_014_2581, w_014_2583, w_014_2585, w_014_2587, w_014_2589, w_014_2590, w_014_2591, w_014_2592, w_014_2593, w_014_2596, w_014_2597, w_014_2601, w_014_2602, w_014_2604, w_014_2607, w_014_2608, w_014_2609, w_014_2610, w_014_2611, w_014_2612, w_014_2613, w_014_2614, w_014_2615, w_014_2616, w_014_2617, w_014_2619, w_014_2620, w_014_2621, w_014_2622, w_014_2623, w_014_2624, w_014_2625, w_014_2626, w_014_2627, w_014_2628, w_014_2629, w_014_2631, w_014_2632, w_014_2633, w_014_2634, w_014_2636, w_014_2637, w_014_2638, w_014_2639, w_014_2640, w_014_2641, w_014_2642, w_014_2643, w_014_2644, w_014_2645, w_014_2646, w_014_2647, w_014_2648, w_014_2649, w_014_2650, w_014_2651, w_014_2652, w_014_2653, w_014_2654, w_014_2655, w_014_2657, w_014_2658, w_014_2659, w_014_2661, w_014_2662, w_014_2663, w_014_2664, w_014_2665, w_014_2666, w_014_2667, w_014_2668, w_014_2669, w_014_2671, w_014_2674, w_014_2675, w_014_2676, w_014_2677, w_014_2678, w_014_2679, w_014_2680, w_014_2681, w_014_2683, w_014_2684, w_014_2685, w_014_2686, w_014_2687, w_014_2689, w_014_2690, w_014_2691, w_014_2692, w_014_2693, w_014_2694, w_014_2695, w_014_2696, w_014_2697, w_014_2698, w_014_2699, w_014_2700, w_014_2701, w_014_2702, w_014_2705, w_014_2706, w_014_2707, w_014_2708, w_014_2711, w_014_2712, w_014_2713, w_014_2714, w_014_2715, w_014_2716, w_014_2717, w_014_2718, w_014_2719, w_014_2720, w_014_2721, w_014_2722, w_014_2723, w_014_2724, w_014_2725, w_014_2726, w_014_2727, w_014_2728, w_014_2729, w_014_2730, w_014_2731, w_014_2733, w_014_2734, w_014_2735, w_014_2737, w_014_2738, w_014_2740, w_014_2743, w_014_2745, w_014_2746, w_014_2747, w_014_2752, w_014_2754, w_014_2755, w_014_2756, w_014_2758, w_014_2759, w_014_2760, w_014_2762, w_014_2763, w_014_2765, w_014_2767, w_014_2768, w_014_2770, w_014_2771, w_014_2772, w_014_2773, w_014_2774, w_014_2775, w_014_2776, w_014_2778, w_014_2779, w_014_2780, w_014_2782, w_014_2783, w_014_2784, w_014_2785, w_014_2786, w_014_2788, w_014_2789, w_014_2790, w_014_2792, w_014_2794, w_014_2796, w_014_2798, w_014_2799, w_014_2800, w_014_2801, w_014_2804, w_014_2805, w_014_2806, w_014_2807, w_014_2810, w_014_2811, w_014_2812, w_014_2813, w_014_2814, w_014_2815, w_014_2816, w_014_2817, w_014_2820, w_014_2821, w_014_2822, w_014_2823, w_014_2824, w_014_2825, w_014_2826, w_014_2827, w_014_2828, w_014_2829, w_014_2830, w_014_2831, w_014_2832, w_014_2833, w_014_2834, w_014_2836, w_014_2837, w_014_2838, w_014_2839, w_014_2840, w_014_2841, w_014_2843, w_014_2844, w_014_2845, w_014_2846, w_014_2847, w_014_2848, w_014_2849, w_014_2850, w_014_2851, w_014_2852, w_014_2854, w_014_2856, w_014_2857, w_014_2858, w_014_2859, w_014_2861, w_014_2862, w_014_2863, w_014_2864, w_014_2865, w_014_2866, w_014_2867, w_014_2870, w_014_2872, w_014_2873, w_014_2874, w_014_2875, w_014_2876, w_014_2878, w_014_2879, w_014_2880, w_014_2881, w_014_2882, w_014_2883, w_014_2884, w_014_2885, w_014_2886, w_014_2887, w_014_2888, w_014_2889, w_014_2891, w_014_2892, w_014_2894, w_014_2895, w_014_2896, w_014_2897, w_014_2898, w_014_2899, w_014_2900, w_014_2901, w_014_2902, w_014_2904, w_014_2905, w_014_2906, w_014_2907, w_014_2908, w_014_2909, w_014_2910, w_014_2911, w_014_2912, w_014_2913, w_014_2914, w_014_2915, w_014_2916, w_014_2918, w_014_2919, w_014_2920, w_014_2921, w_014_2922, w_014_2925, w_014_2926, w_014_2927, w_014_2928, w_014_2930, w_014_2932, w_014_2933, w_014_2934, w_014_2935, w_014_2936, w_014_2937, w_014_2938, w_014_2939, w_014_2940, w_014_2941, w_014_2942, w_014_2943, w_014_2944, w_014_2945, w_014_2946, w_014_2947, w_014_2948, w_014_2949, w_014_2950, w_014_2951, w_014_2952, w_014_2953, w_014_2954, w_014_2955, w_014_2957, w_014_2958, w_014_2959, w_014_2960, w_014_2961, w_014_2962, w_014_2963, w_014_2964, w_014_2966, w_014_2969, w_014_2970, w_014_2971, w_014_2972, w_014_2974, w_014_2975, w_014_2976, w_014_2977, w_014_2978, w_014_2981, w_014_2982, w_014_2983, w_014_2984, w_014_2986, w_014_2987, w_014_2988, w_014_2989, w_014_2990, w_014_2991, w_014_2992, w_014_2994, w_014_2995, w_014_2997, w_014_2999, w_014_3001, w_014_3002, w_014_3003, w_014_3004, w_014_3006, w_014_3007, w_014_3008, w_014_3009, w_014_3010, w_014_3012, w_014_3014, w_014_3015, w_014_3017, w_014_3018, w_014_3020, w_014_3021, w_014_3022, w_014_3023, w_014_3024, w_014_3025, w_014_3026, w_014_3027, w_014_3028, w_014_3029, w_014_3030, w_014_3031, w_014_3032, w_014_3033, w_014_3035, w_014_3037, w_014_3039, w_014_3040, w_014_3041, w_014_3042, w_014_3044, w_014_3046, w_014_3047, w_014_3048, w_014_3049, w_014_3050, w_014_3051, w_014_3052, w_014_3053, w_014_3054, w_014_3055, w_014_3056, w_014_3057, w_014_3058, w_014_3059, w_014_3061, w_014_3062, w_014_3063, w_014_3064, w_014_3065, w_014_3066, w_014_3068, w_014_3069, w_014_3070, w_014_3071, w_014_3072, w_014_3073, w_014_3074, w_014_3075, w_014_3076, w_014_3077, w_014_3078, w_014_3079, w_014_3081, w_014_3083, w_014_3085, w_014_3086, w_014_3087, w_014_3088, w_014_3089, w_014_3090, w_014_3091, w_014_3093, w_014_3094, w_014_3095, w_014_3096, w_014_3097, w_014_3098, w_014_3099, w_014_3101, w_014_3103, w_014_3104, w_014_3105, w_014_3106, w_014_3107, w_014_3109, w_014_3110, w_014_3112, w_014_3113, w_014_3114, w_014_3115, w_014_3117, w_014_3118, w_014_3119, w_014_3120, w_014_3121, w_014_3122, w_014_3123, w_014_3124, w_014_3126, w_014_3127, w_014_3128, w_014_3129, w_014_3130, w_014_3131, w_014_3132, w_014_3133, w_014_3134, w_014_3135, w_014_3136, w_014_3137, w_014_3138, w_014_3139, w_014_3140, w_014_3141, w_014_3143, w_014_3144, w_014_3145, w_014_3148, w_014_3149, w_014_3151, w_014_3154, w_014_3155, w_014_3156, w_014_3157, w_014_3160, w_014_3162, w_014_3165, w_014_3167, w_014_3168, w_014_3169, w_014_3170, w_014_3171, w_014_3172, w_014_3173, w_014_3174, w_014_3175, w_014_3177, w_014_3178, w_014_3179, w_014_3180, w_014_3182, w_014_3184, w_014_3185, w_014_3186, w_014_3187, w_014_3188, w_014_3189, w_014_3190, w_014_3192, w_014_3193, w_014_3194, w_014_3195, w_014_3196, w_014_3197, w_014_3198, w_014_3199, w_014_3201;
  wire w_015_000, w_015_001, w_015_002, w_015_003, w_015_004, w_015_005, w_015_006, w_015_007, w_015_008, w_015_009, w_015_011, w_015_012, w_015_013, w_015_014, w_015_015, w_015_016, w_015_017, w_015_018, w_015_019, w_015_020, w_015_021, w_015_022, w_015_023, w_015_024, w_015_025, w_015_026, w_015_027, w_015_028, w_015_029, w_015_030, w_015_031, w_015_032, w_015_033, w_015_034, w_015_035, w_015_036, w_015_037, w_015_039, w_015_040, w_015_041, w_015_042, w_015_044, w_015_045, w_015_046, w_015_047, w_015_048, w_015_049, w_015_050, w_015_051, w_015_052, w_015_053, w_015_054, w_015_056, w_015_058, w_015_059, w_015_061, w_015_062, w_015_063, w_015_064, w_015_065, w_015_069, w_015_070, w_015_072, w_015_073, w_015_074, w_015_075, w_015_076, w_015_077, w_015_079, w_015_080, w_015_081, w_015_082, w_015_084, w_015_087, w_015_088, w_015_089, w_015_091, w_015_092, w_015_094, w_015_095, w_015_096, w_015_097, w_015_098, w_015_099, w_015_101, w_015_102, w_015_103, w_015_104, w_015_105, w_015_107, w_015_108, w_015_109, w_015_110, w_015_111, w_015_112, w_015_113, w_015_114, w_015_115, w_015_116, w_015_117, w_015_118, w_015_119, w_015_120, w_015_122, w_015_123, w_015_124, w_015_125, w_015_126, w_015_127, w_015_128, w_015_130, w_015_132, w_015_133, w_015_135, w_015_136, w_015_137, w_015_138, w_015_140, w_015_141, w_015_143, w_015_144, w_015_145, w_015_146, w_015_147, w_015_148, w_015_149, w_015_150, w_015_151, w_015_152, w_015_153, w_015_154, w_015_155, w_015_157, w_015_158, w_015_159, w_015_160, w_015_161, w_015_162, w_015_164, w_015_165, w_015_166, w_015_168, w_015_170, w_015_171, w_015_172, w_015_173, w_015_174, w_015_175, w_015_176, w_015_178, w_015_180, w_015_182, w_015_183, w_015_184, w_015_185, w_015_186, w_015_187, w_015_189, w_015_191, w_015_192, w_015_193, w_015_194, w_015_195, w_015_196, w_015_197, w_015_198, w_015_199, w_015_200, w_015_201, w_015_202, w_015_203, w_015_204, w_015_205, w_015_206, w_015_207, w_015_208, w_015_209, w_015_210, w_015_211, w_015_212, w_015_213, w_015_217, w_015_218, w_015_219, w_015_220, w_015_221, w_015_222, w_015_223, w_015_224, w_015_225, w_015_227, w_015_228, w_015_229, w_015_230, w_015_231, w_015_232, w_015_234, w_015_235, w_015_236, w_015_238, w_015_239, w_015_240, w_015_241, w_015_242, w_015_243, w_015_244, w_015_245, w_015_246, w_015_247, w_015_248, w_015_249, w_015_250, w_015_251, w_015_252, w_015_253, w_015_254, w_015_255, w_015_257, w_015_258, w_015_259, w_015_262, w_015_263, w_015_264, w_015_266, w_015_267, w_015_268, w_015_269, w_015_270, w_015_271, w_015_272, w_015_273, w_015_274, w_015_275, w_015_276, w_015_277, w_015_280, w_015_281, w_015_282, w_015_283, w_015_284, w_015_285, w_015_286, w_015_288, w_015_289, w_015_290, w_015_291, w_015_292, w_015_294, w_015_295, w_015_296, w_015_297, w_015_298, w_015_299, w_015_300, w_015_302, w_015_303, w_015_305, w_015_308, w_015_309, w_015_310, w_015_312, w_015_313, w_015_316, w_015_317, w_015_319, w_015_321, w_015_322, w_015_324, w_015_325, w_015_327, w_015_329, w_015_330, w_015_332, w_015_334, w_015_335, w_015_337, w_015_341, w_015_342, w_015_343, w_015_344, w_015_345, w_015_346, w_015_349, w_015_350, w_015_351, w_015_353, w_015_354, w_015_355, w_015_357, w_015_358, w_015_359, w_015_361, w_015_362, w_015_363, w_015_364, w_015_365, w_015_366, w_015_367, w_015_368, w_015_369, w_015_372, w_015_373, w_015_374, w_015_375, w_015_376, w_015_377, w_015_378, w_015_380, w_015_381, w_015_382, w_015_383, w_015_384, w_015_386, w_015_387, w_015_388, w_015_389, w_015_390, w_015_391, w_015_392, w_015_395, w_015_396, w_015_397, w_015_398, w_015_399, w_015_400, w_015_402, w_015_403, w_015_404, w_015_407, w_015_408, w_015_409, w_015_410, w_015_411, w_015_412, w_015_413, w_015_414, w_015_415, w_015_416, w_015_417, w_015_418, w_015_420, w_015_422, w_015_424, w_015_425, w_015_426, w_015_427, w_015_429, w_015_431, w_015_433, w_015_434, w_015_435, w_015_436, w_015_443, w_015_444, w_015_445, w_015_446, w_015_448, w_015_449, w_015_450, w_015_451, w_015_452, w_015_453, w_015_454, w_015_456, w_015_459, w_015_460, w_015_462, w_015_463, w_015_464, w_015_466, w_015_467, w_015_468, w_015_469, w_015_471, w_015_472, w_015_473, w_015_474, w_015_475, w_015_476, w_015_477, w_015_478, w_015_479, w_015_481, w_015_482, w_015_483, w_015_485, w_015_486, w_015_487, w_015_488, w_015_489, w_015_491, w_015_492, w_015_494, w_015_496, w_015_497, w_015_499, w_015_500, w_015_501, w_015_503, w_015_504, w_015_505, w_015_507, w_015_508, w_015_509, w_015_510, w_015_511, w_015_512, w_015_513, w_015_514, w_015_515, w_015_517, w_015_518, w_015_519, w_015_520, w_015_521, w_015_523, w_015_524, w_015_525, w_015_527, w_015_528, w_015_531, w_015_533, w_015_534, w_015_536, w_015_537, w_015_538, w_015_540, w_015_541, w_015_542, w_015_544, w_015_545, w_015_546, w_015_547, w_015_548, w_015_549, w_015_550, w_015_551, w_015_552, w_015_553, w_015_554, w_015_555, w_015_556, w_015_558, w_015_559, w_015_561, w_015_566, w_015_567, w_015_568, w_015_569, w_015_571, w_015_572, w_015_573, w_015_575, w_015_576, w_015_577, w_015_579, w_015_580, w_015_581, w_015_582, w_015_583, w_015_584, w_015_585, w_015_586, w_015_589, w_015_591, w_015_592, w_015_593, w_015_594, w_015_595, w_015_598, w_015_599, w_015_600, w_015_601, w_015_602, w_015_603, w_015_605, w_015_606, w_015_608, w_015_609, w_015_610, w_015_611, w_015_612, w_015_613, w_015_614, w_015_615, w_015_616, w_015_617, w_015_618, w_015_621, w_015_622, w_015_626, w_015_627, w_015_629, w_015_630, w_015_631, w_015_632, w_015_634, w_015_635, w_015_636, w_015_637, w_015_638, w_015_639, w_015_640, w_015_641, w_015_643, w_015_644, w_015_646, w_015_649, w_015_651, w_015_652, w_015_653, w_015_655, w_015_656, w_015_657, w_015_658, w_015_659, w_015_660, w_015_661, w_015_663, w_015_665, w_015_666, w_015_667, w_015_668, w_015_671, w_015_672, w_015_673, w_015_674, w_015_675, w_015_677, w_015_679, w_015_680, w_015_682, w_015_683, w_015_684, w_015_685, w_015_686, w_015_687, w_015_688, w_015_689, w_015_690, w_015_691, w_015_692, w_015_693, w_015_695, w_015_696, w_015_697, w_015_698, w_015_699, w_015_700, w_015_701, w_015_702, w_015_703, w_015_704, w_015_705, w_015_706, w_015_707, w_015_709, w_015_710, w_015_711, w_015_712, w_015_715, w_015_716, w_015_717, w_015_718, w_015_721, w_015_722, w_015_723, w_015_724, w_015_726, w_015_727, w_015_728, w_015_730, w_015_731, w_015_732, w_015_734, w_015_735, w_015_736, w_015_737, w_015_738, w_015_741, w_015_743, w_015_744, w_015_745, w_015_747, w_015_748, w_015_749, w_015_750, w_015_751, w_015_752, w_015_754, w_015_755, w_015_757, w_015_758, w_015_762, w_015_763, w_015_764, w_015_765, w_015_766, w_015_767, w_015_768, w_015_769, w_015_770, w_015_771, w_015_777, w_015_778, w_015_779, w_015_781, w_015_782, w_015_783, w_015_784, w_015_786, w_015_787, w_015_791, w_015_792, w_015_793, w_015_794, w_015_795, w_015_796, w_015_798, w_015_800, w_015_801, w_015_802, w_015_803, w_015_804, w_015_807, w_015_808, w_015_809, w_015_810, w_015_814, w_015_815, w_015_816, w_015_817, w_015_818, w_015_819, w_015_821, w_015_823, w_015_824, w_015_825, w_015_826, w_015_827, w_015_828, w_015_829, w_015_830, w_015_831, w_015_832, w_015_833, w_015_834, w_015_835, w_015_836, w_015_838, w_015_839, w_015_840, w_015_842, w_015_843, w_015_844, w_015_846, w_015_847, w_015_848, w_015_849, w_015_850, w_015_852, w_015_853, w_015_854, w_015_855, w_015_856, w_015_857, w_015_858, w_015_859, w_015_863, w_015_864, w_015_866, w_015_868, w_015_869, w_015_870, w_015_872, w_015_874, w_015_875, w_015_876, w_015_877, w_015_878, w_015_879, w_015_880, w_015_882, w_015_883, w_015_884, w_015_885, w_015_886, w_015_888, w_015_889, w_015_890, w_015_891, w_015_892, w_015_893, w_015_894, w_015_895, w_015_896, w_015_897, w_015_898, w_015_899, w_015_900, w_015_901, w_015_902, w_015_904, w_015_906, w_015_907, w_015_909, w_015_910, w_015_911, w_015_912, w_015_913, w_015_918, w_015_920, w_015_923, w_015_924, w_015_925, w_015_928, w_015_932, w_015_933, w_015_934, w_015_936, w_015_937, w_015_941, w_015_942, w_015_943, w_015_948, w_015_949, w_015_950, w_015_954, w_015_955, w_015_956, w_015_957, w_015_959, w_015_960, w_015_961, w_015_962, w_015_963, w_015_964, w_015_965, w_015_966, w_015_967, w_015_968, w_015_969, w_015_971, w_015_972, w_015_973, w_015_974, w_015_975, w_015_977, w_015_978, w_015_979, w_015_981, w_015_983, w_015_985, w_015_986, w_015_987, w_015_989, w_015_990, w_015_991, w_015_992, w_015_994, w_015_995, w_015_996, w_015_997, w_015_998, w_015_999, w_015_1000, w_015_1001, w_015_1002, w_015_1004, w_015_1005, w_015_1006, w_015_1007, w_015_1009, w_015_1012, w_015_1013, w_015_1014, w_015_1015, w_015_1018, w_015_1019, w_015_1020, w_015_1021, w_015_1023, w_015_1024, w_015_1025, w_015_1026, w_015_1027, w_015_1028, w_015_1029, w_015_1030, w_015_1031, w_015_1033, w_015_1034, w_015_1035, w_015_1036, w_015_1037, w_015_1038, w_015_1039, w_015_1040, w_015_1046, w_015_1047, w_015_1048, w_015_1049, w_015_1050, w_015_1051, w_015_1052, w_015_1053, w_015_1054, w_015_1055, w_015_1056, w_015_1058, w_015_1059, w_015_1060, w_015_1061, w_015_1063, w_015_1064, w_015_1065, w_015_1066, w_015_1068, w_015_1069, w_015_1070, w_015_1072, w_015_1073, w_015_1076, w_015_1077, w_015_1078, w_015_1079, w_015_1081, w_015_1082, w_015_1083, w_015_1084, w_015_1085, w_015_1086, w_015_1087, w_015_1088, w_015_1089, w_015_1091, w_015_1092, w_015_1093, w_015_1094, w_015_1095, w_015_1096, w_015_1097, w_015_1098, w_015_1099, w_015_1102, w_015_1103, w_015_1104, w_015_1105, w_015_1106, w_015_1107, w_015_1109, w_015_1110, w_015_1111, w_015_1112, w_015_1113, w_015_1114, w_015_1116, w_015_1118, w_015_1119, w_015_1120, w_015_1121, w_015_1122, w_015_1123, w_015_1125, w_015_1126, w_015_1129, w_015_1130, w_015_1131, w_015_1132, w_015_1133, w_015_1134, w_015_1135, w_015_1136, w_015_1138, w_015_1139, w_015_1140, w_015_1141, w_015_1142, w_015_1144, w_015_1145, w_015_1146, w_015_1147, w_015_1148, w_015_1149, w_015_1150, w_015_1151, w_015_1152, w_015_1154, w_015_1155, w_015_1156, w_015_1157, w_015_1158, w_015_1159, w_015_1160, w_015_1161, w_015_1163, w_015_1164, w_015_1165, w_015_1166, w_015_1167, w_015_1168, w_015_1169, w_015_1170, w_015_1173, w_015_1174, w_015_1176, w_015_1177, w_015_1178, w_015_1179, w_015_1181, w_015_1182, w_015_1183, w_015_1184, w_015_1186, w_015_1187, w_015_1189, w_015_1191, w_015_1193, w_015_1194, w_015_1196, w_015_1197, w_015_1198, w_015_1199, w_015_1200, w_015_1201, w_015_1202, w_015_1203, w_015_1204, w_015_1205, w_015_1209, w_015_1210, w_015_1211, w_015_1212, w_015_1213, w_015_1214, w_015_1215, w_015_1216, w_015_1217, w_015_1218, w_015_1219, w_015_1221, w_015_1222, w_015_1223, w_015_1224, w_015_1225, w_015_1226, w_015_1227, w_015_1228, w_015_1229, w_015_1230, w_015_1231, w_015_1232, w_015_1233, w_015_1234, w_015_1235, w_015_1236, w_015_1237, w_015_1238, w_015_1239, w_015_1240, w_015_1242, w_015_1243, w_015_1244, w_015_1246, w_015_1247, w_015_1248, w_015_1249, w_015_1251, w_015_1252, w_015_1253, w_015_1254, w_015_1255, w_015_1256, w_015_1257, w_015_1258, w_015_1260, w_015_1261, w_015_1262, w_015_1263, w_015_1264, w_015_1265, w_015_1269, w_015_1270, w_015_1271, w_015_1272, w_015_1274, w_015_1275, w_015_1277, w_015_1279, w_015_1280, w_015_1281, w_015_1282, w_015_1287, w_015_1288, w_015_1289, w_015_1292, w_015_1293, w_015_1294, w_015_1295, w_015_1296, w_015_1297, w_015_1298, w_015_1299, w_015_1300, w_015_1302, w_015_1303, w_015_1305, w_015_1306, w_015_1308, w_015_1309, w_015_1310, w_015_1311, w_015_1312, w_015_1313, w_015_1315, w_015_1318, w_015_1319, w_015_1320, w_015_1321, w_015_1323, w_015_1324, w_015_1326, w_015_1327, w_015_1329, w_015_1330, w_015_1332, w_015_1333, w_015_1334, w_015_1336, w_015_1338, w_015_1339, w_015_1340, w_015_1342, w_015_1343, w_015_1344, w_015_1345, w_015_1346, w_015_1347, w_015_1348, w_015_1349, w_015_1350, w_015_1351, w_015_1352, w_015_1354, w_015_1356, w_015_1358, w_015_1359, w_015_1360, w_015_1361, w_015_1362, w_015_1363, w_015_1364, w_015_1365, w_015_1366, w_015_1367, w_015_1369, w_015_1371, w_015_1372, w_015_1373, w_015_1374, w_015_1377, w_015_1378, w_015_1379, w_015_1380, w_015_1381, w_015_1383, w_015_1384, w_015_1385, w_015_1387, w_015_1388, w_015_1390, w_015_1391, w_015_1392, w_015_1393, w_015_1394, w_015_1395, w_015_1396, w_015_1397, w_015_1398, w_015_1399, w_015_1400, w_015_1402, w_015_1404, w_015_1405, w_015_1406, w_015_1407, w_015_1408, w_015_1409, w_015_1411, w_015_1413, w_015_1414, w_015_1415, w_015_1417, w_015_1418, w_015_1419, w_015_1420, w_015_1421, w_015_1422, w_015_1423, w_015_1424, w_015_1425, w_015_1427, w_015_1429, w_015_1430, w_015_1431, w_015_1433, w_015_1437, w_015_1440, w_015_1441, w_015_1442, w_015_1444, w_015_1445, w_015_1446, w_015_1449, w_015_1450, w_015_1451, w_015_1452, w_015_1453, w_015_1454, w_015_1455, w_015_1457, w_015_1458, w_015_1459, w_015_1460, w_015_1461, w_015_1462, w_015_1463, w_015_1467, w_015_1468, w_015_1469, w_015_1472, w_015_1473, w_015_1474, w_015_1476, w_015_1477, w_015_1478, w_015_1479, w_015_1480, w_015_1482, w_015_1485, w_015_1487, w_015_1488, w_015_1489, w_015_1490, w_015_1491, w_015_1492, w_015_1493, w_015_1494, w_015_1495, w_015_1496, w_015_1497, w_015_1499, w_015_1500, w_015_1501, w_015_1502, w_015_1503, w_015_1504, w_015_1508, w_015_1510, w_015_1512, w_015_1513, w_015_1514, w_015_1515, w_015_1516, w_015_1517, w_015_1518, w_015_1519, w_015_1520, w_015_1521, w_015_1522, w_015_1523, w_015_1524, w_015_1525, w_015_1526, w_015_1528, w_015_1529, w_015_1530, w_015_1531, w_015_1532, w_015_1533, w_015_1534, w_015_1535, w_015_1537, w_015_1538, w_015_1539, w_015_1544, w_015_1545, w_015_1546, w_015_1549, w_015_1552, w_015_1555, w_015_1556, w_015_1557, w_015_1558, w_015_1559, w_015_1561, w_015_1562, w_015_1563, w_015_1564, w_015_1565, w_015_1566, w_015_1568, w_015_1569, w_015_1573, w_015_1574, w_015_1575, w_015_1576, w_015_1577, w_015_1578, w_015_1579, w_015_1580, w_015_1581, w_015_1582, w_015_1584, w_015_1585, w_015_1586, w_015_1587, w_015_1588, w_015_1589, w_015_1591, w_015_1592, w_015_1594, w_015_1597, w_015_1598, w_015_1599, w_015_1600, w_015_1601, w_015_1602, w_015_1603, w_015_1604, w_015_1605, w_015_1608, w_015_1609, w_015_1612, w_015_1613, w_015_1615, w_015_1616, w_015_1617, w_015_1618, w_015_1619, w_015_1621, w_015_1626, w_015_1627, w_015_1628, w_015_1629, w_015_1630, w_015_1631, w_015_1632, w_015_1633, w_015_1634, w_015_1637, w_015_1638, w_015_1639, w_015_1641, w_015_1642, w_015_1643, w_015_1644, w_015_1646, w_015_1648, w_015_1650, w_015_1651, w_015_1652, w_015_1653, w_015_1654, w_015_1655, w_015_1656, w_015_1657, w_015_1658, w_015_1659, w_015_1661, w_015_1665, w_015_1671, w_015_1672, w_015_1673, w_015_1674, w_015_1675, w_015_1676, w_015_1677, w_015_1678, w_015_1679, w_015_1680, w_015_1681, w_015_1683, w_015_1684, w_015_1685, w_015_1686, w_015_1688, w_015_1689, w_015_1692, w_015_1693, w_015_1694, w_015_1696, w_015_1697, w_015_1698, w_015_1699, w_015_1700, w_015_1702, w_015_1703, w_015_1704, w_015_1705, w_015_1708, w_015_1709, w_015_1710, w_015_1711, w_015_1712, w_015_1713, w_015_1715, w_015_1716, w_015_1717, w_015_1718, w_015_1720, w_015_1721, w_015_1723, w_015_1724, w_015_1725, w_015_1726, w_015_1727, w_015_1728, w_015_1729, w_015_1730, w_015_1733, w_015_1735, w_015_1736, w_015_1737, w_015_1738, w_015_1739, w_015_1741, w_015_1742, w_015_1744, w_015_1745, w_015_1746, w_015_1747, w_015_1749, w_015_1750, w_015_1751, w_015_1752, w_015_1755, w_015_1756, w_015_1757, w_015_1759, w_015_1760, w_015_1761, w_015_1762, w_015_1764, w_015_1765, w_015_1766, w_015_1767, w_015_1769, w_015_1770, w_015_1771, w_015_1772, w_015_1773, w_015_1774, w_015_1775, w_015_1776, w_015_1777, w_015_1778, w_015_1779, w_015_1780, w_015_1781, w_015_1782, w_015_1783, w_015_1784, w_015_1786, w_015_1787, w_015_1788, w_015_1789, w_015_1790, w_015_1791, w_015_1792, w_015_1793, w_015_1794, w_015_1795, w_015_1797, w_015_1798, w_015_1799, w_015_1801, w_015_1802, w_015_1803, w_015_1804, w_015_1805, w_015_1806, w_015_1807, w_015_1808, w_015_1809, w_015_1810, w_015_1811, w_015_1813, w_015_1814, w_015_1815, w_015_1816, w_015_1817, w_015_1818, w_015_1819, w_015_1820, w_015_1821, w_015_1822, w_015_1824, w_015_1825, w_015_1827, w_015_1828, w_015_1829, w_015_1831, w_015_1832, w_015_1833, w_015_1834, w_015_1835, w_015_1836, w_015_1838, w_015_1840, w_015_1841, w_015_1845, w_015_1846, w_015_1848, w_015_1850, w_015_1853, w_015_1854, w_015_1855, w_015_1856, w_015_1857, w_015_1858, w_015_1861, w_015_1862, w_015_1863, w_015_1864, w_015_1865, w_015_1866, w_015_1867, w_015_1868, w_015_1869, w_015_1870, w_015_1871, w_015_1872, w_015_1873, w_015_1875, w_015_1877, w_015_1879, w_015_1881, w_015_1882, w_015_1883, w_015_1885, w_015_1886, w_015_1888, w_015_1891, w_015_1892, w_015_1895, w_015_1896, w_015_1897, w_015_1899, w_015_1900, w_015_1902, w_015_1903, w_015_1904, w_015_1905, w_015_1906, w_015_1907, w_015_1908, w_015_1909, w_015_1910, w_015_1912, w_015_1913, w_015_1914, w_015_1915, w_015_1917, w_015_1920, w_015_1921, w_015_1922, w_015_1924, w_015_1925, w_015_1926, w_015_1927, w_015_1929, w_015_1930, w_015_1932, w_015_1933, w_015_1935, w_015_1936, w_015_1938, w_015_1939, w_015_1940, w_015_1941, w_015_1942, w_015_1943, w_015_1946, w_015_1947, w_015_1948, w_015_1949, w_015_1950, w_015_1951, w_015_1952, w_015_1953, w_015_1955, w_015_1956, w_015_1957, w_015_1959, w_015_1960, w_015_1962, w_015_1963, w_015_1964, w_015_1965, w_015_1966, w_015_1969, w_015_1970, w_015_1971, w_015_1972, w_015_1973, w_015_1974, w_015_1975, w_015_1976, w_015_1977, w_015_1978, w_015_1980, w_015_1981, w_015_1982, w_015_1983, w_015_1984, w_015_1985, w_015_1986, w_015_1987, w_015_1988, w_015_1989, w_015_1991, w_015_1992, w_015_1995, w_015_1996, w_015_1997, w_015_1999, w_015_2000, w_015_2002, w_015_2003, w_015_2004, w_015_2005, w_015_2006, w_015_2010, w_015_2011, w_015_2012, w_015_2013, w_015_2015, w_015_2016, w_015_2017, w_015_2018, w_015_2019, w_015_2020, w_015_2021, w_015_2023, w_015_2025, w_015_2026, w_015_2027, w_015_2028, w_015_2029, w_015_2030, w_015_2033, w_015_2034, w_015_2036, w_015_2037, w_015_2038, w_015_2040, w_015_2044, w_015_2045, w_015_2047, w_015_2048, w_015_2049, w_015_2052, w_015_2054, w_015_2055, w_015_2056, w_015_2057, w_015_2058, w_015_2061, w_015_2062, w_015_2063, w_015_2064, w_015_2065, w_015_2066, w_015_2068, w_015_2069, w_015_2070, w_015_2071, w_015_2072, w_015_2073, w_015_2074, w_015_2075, w_015_2076, w_015_2077, w_015_2078, w_015_2080, w_015_2081, w_015_2082, w_015_2085, w_015_2086, w_015_2087, w_015_2088, w_015_2089, w_015_2090, w_015_2091, w_015_2092, w_015_2093, w_015_2094, w_015_2096, w_015_2097, w_015_2098, w_015_2099, w_015_2101, w_015_2102, w_015_2103, w_015_2104, w_015_2105, w_015_2107, w_015_2108, w_015_2109, w_015_2110, w_015_2112, w_015_2113, w_015_2114, w_015_2115, w_015_2116, w_015_2118, w_015_2120, w_015_2121, w_015_2122, w_015_2124, w_015_2125, w_015_2126, w_015_2127, w_015_2128, w_015_2130, w_015_2131, w_015_2132, w_015_2133, w_015_2134, w_015_2135, w_015_2136, w_015_2137, w_015_2139, w_015_2141, w_015_2142, w_015_2143, w_015_2144, w_015_2146, w_015_2148, w_015_2149, w_015_2150, w_015_2151, w_015_2152, w_015_2153, w_015_2154, w_015_2155, w_015_2159, w_015_2160, w_015_2162, w_015_2163, w_015_2165, w_015_2167, w_015_2169, w_015_2170, w_015_2171, w_015_2174, w_015_2175, w_015_2176, w_015_2179, w_015_2181, w_015_2182, w_015_2183, w_015_2184, w_015_2185, w_015_2186, w_015_2187, w_015_2188, w_015_2190, w_015_2192, w_015_2193, w_015_2194, w_015_2195, w_015_2197, w_015_2199, w_015_2200, w_015_2203, w_015_2204, w_015_2205, w_015_2206, w_015_2207, w_015_2209, w_015_2210, w_015_2212, w_015_2213, w_015_2214, w_015_2215, w_015_2216, w_015_2219, w_015_2220, w_015_2221, w_015_2222, w_015_2224, w_015_2225, w_015_2226, w_015_2227, w_015_2229, w_015_2230, w_015_2231, w_015_2232, w_015_2233, w_015_2234, w_015_2235, w_015_2236, w_015_2237, w_015_2238, w_015_2240, w_015_2242, w_015_2244, w_015_2245, w_015_2246, w_015_2247, w_015_2248, w_015_2249, w_015_2250, w_015_2251, w_015_2252, w_015_2254, w_015_2256, w_015_2257, w_015_2259, w_015_2262, w_015_2263, w_015_2264, w_015_2265, w_015_2266, w_015_2267, w_015_2268, w_015_2269, w_015_2270, w_015_2271, w_015_2272, w_015_2275, w_015_2276, w_015_2277, w_015_2278, w_015_2279, w_015_2280, w_015_2281, w_015_2282, w_015_2284, w_015_2285, w_015_2286, w_015_2287, w_015_2288, w_015_2289, w_015_2290, w_015_2293, w_015_2294, w_015_2296, w_015_2298, w_015_2299, w_015_2302, w_015_2303, w_015_2304, w_015_2305, w_015_2306, w_015_2307, w_015_2308, w_015_2309, w_015_2310, w_015_2311, w_015_2312, w_015_2313, w_015_2314, w_015_2315, w_015_2318, w_015_2319, w_015_2321, w_015_2324, w_015_2325, w_015_2327, w_015_2328, w_015_2329, w_015_2330, w_015_2331, w_015_2332, w_015_2333, w_015_2335, w_015_2336, w_015_2337, w_015_2338, w_015_2339, w_015_2340, w_015_2341, w_015_2342, w_015_2343, w_015_2344, w_015_2346, w_015_2347, w_015_2349, w_015_2351, w_015_2352, w_015_2353, w_015_2354, w_015_2355, w_015_2357, w_015_2358, w_015_2361, w_015_2362, w_015_2363, w_015_2364, w_015_2366, w_015_2367, w_015_2368, w_015_2369, w_015_2371, w_015_2373, w_015_2374, w_015_2376, w_015_2378, w_015_2379, w_015_2380, w_015_2381, w_015_2382, w_015_2383, w_015_2384, w_015_2385, w_015_2389, w_015_2390, w_015_2391, w_015_2392, w_015_2394, w_015_2395, w_015_2396, w_015_2397, w_015_2398, w_015_2399, w_015_2400, w_015_2401, w_015_2403, w_015_2404, w_015_2406, w_015_2407, w_015_2408, w_015_2409, w_015_2412, w_015_2413, w_015_2415, w_015_2417, w_015_2418, w_015_2419, w_015_2421, w_015_2422, w_015_2423, w_015_2424, w_015_2427, w_015_2428, w_015_2430, w_015_2432, w_015_2434, w_015_2435, w_015_2436, w_015_2437, w_015_2438, w_015_2439, w_015_2440, w_015_2441, w_015_2444, w_015_2445, w_015_2447, w_015_2448, w_015_2449, w_015_2451, w_015_2452, w_015_2453, w_015_2456, w_015_2458, w_015_2459, w_015_2462, w_015_2463, w_015_2465, w_015_2467, w_015_2468, w_015_2469, w_015_2470, w_015_2471, w_015_2472, w_015_2473, w_015_2476, w_015_2477, w_015_2478, w_015_2480, w_015_2481, w_015_2482, w_015_2483, w_015_2484, w_015_2485, w_015_2488, w_015_2489, w_015_2490, w_015_2492, w_015_2493, w_015_2494, w_015_2495, w_015_2498, w_015_2499, w_015_2500, w_015_2501, w_015_2502, w_015_2503, w_015_2506, w_015_2507, w_015_2512, w_015_2514, w_015_2515, w_015_2516, w_015_2518, w_015_2519, w_015_2520, w_015_2521, w_015_2522, w_015_2523, w_015_2524, w_015_2526, w_015_2528, w_015_2529, w_015_2530, w_015_2531, w_015_2532, w_015_2533, w_015_2534, w_015_2536, w_015_2537, w_015_2540, w_015_2542, w_015_2543, w_015_2544, w_015_2545, w_015_2546, w_015_2547, w_015_2548, w_015_2549, w_015_2550, w_015_2551, w_015_2552, w_015_2553, w_015_2554, w_015_2555, w_015_2556, w_015_2557, w_015_2558, w_015_2559, w_015_2560, w_015_2561, w_015_2562, w_015_2563, w_015_2564, w_015_2565, w_015_2566, w_015_2567, w_015_2568, w_015_2573, w_015_2575, w_015_2576, w_015_2577, w_015_2578, w_015_2579, w_015_2580, w_015_2582, w_015_2583, w_015_2584, w_015_2586, w_015_2589, w_015_2590, w_015_2591, w_015_2592, w_015_2593, w_015_2594, w_015_2595, w_015_2596, w_015_2597, w_015_2598, w_015_2600, w_015_2601, w_015_2602, w_015_2603, w_015_2604, w_015_2605, w_015_2607, w_015_2608, w_015_2609, w_015_2610, w_015_2611, w_015_2612, w_015_2614, w_015_2615, w_015_2616, w_015_2617, w_015_2619, w_015_2620, w_015_2621, w_015_2624, w_015_2625, w_015_2626, w_015_2627, w_015_2629, w_015_2631, w_015_2632, w_015_2633, w_015_2634, w_015_2636, w_015_2637, w_015_2638, w_015_2641, w_015_2642, w_015_2643, w_015_2644, w_015_2645, w_015_2646, w_015_2648, w_015_2650, w_015_2653, w_015_2654, w_015_2655, w_015_2656, w_015_2657, w_015_2658, w_015_2660, w_015_2661, w_015_2662, w_015_2663, w_015_2666, w_015_2667, w_015_2669, w_015_2670, w_015_2672, w_015_2673, w_015_2674, w_015_2675, w_015_2676, w_015_2677, w_015_2680, w_015_2681, w_015_2683, w_015_2686, w_015_2688, w_015_2690, w_015_2691, w_015_2695, w_015_2696, w_015_2697, w_015_2699, w_015_2700, w_015_2701, w_015_2703, w_015_2704, w_015_2706, w_015_2707, w_015_2708, w_015_2709, w_015_2710, w_015_2711, w_015_2712, w_015_2713, w_015_2714, w_015_2716, w_015_2717, w_015_2719, w_015_2720, w_015_2721, w_015_2722, w_015_2723, w_015_2724, w_015_2727, w_015_2728, w_015_2729, w_015_2730, w_015_2731, w_015_2733, w_015_2734, w_015_2737, w_015_2738, w_015_2739, w_015_2741, w_015_2742, w_015_2743, w_015_2745, w_015_2746, w_015_2747, w_015_2748, w_015_2749, w_015_2750, w_015_2751, w_015_2752, w_015_2753, w_015_2756, w_015_2757, w_015_2758, w_015_2759, w_015_2760, w_015_2761, w_015_2762, w_015_2763, w_015_2764, w_015_2765, w_015_2766, w_015_2768, w_015_2769, w_015_2772, w_015_2773, w_015_2774, w_015_2775, w_015_2776, w_015_2777, w_015_2778, w_015_2779, w_015_2780, w_015_2781, w_015_2782, w_015_2786, w_015_2788, w_015_2789, w_015_2790, w_015_2792, w_015_2793, w_015_2794, w_015_2795, w_015_2796, w_015_2797, w_015_2801, w_015_2802, w_015_2803, w_015_2804, w_015_2805, w_015_2806, w_015_2807, w_015_2809, w_015_2813, w_015_2814, w_015_2815, w_015_2818, w_015_2820, w_015_2823, w_015_2824, w_015_2825, w_015_2826, w_015_2827, w_015_2828, w_015_2829, w_015_2830, w_015_2831, w_015_2832, w_015_2833, w_015_2835, w_015_2836, w_015_2837, w_015_2838, w_015_2840, w_015_2841, w_015_2843, w_015_2844, w_015_2845, w_015_2846, w_015_2848, w_015_2849, w_015_2850, w_015_2853, w_015_2854, w_015_2855, w_015_2856, w_015_2858, w_015_2860, w_015_2861, w_015_2863, w_015_2864, w_015_2865, w_015_2866, w_015_2867, w_015_2868, w_015_2869, w_015_2870, w_015_2871, w_015_2872, w_015_2873, w_015_2874, w_015_2877, w_015_2879, w_015_2880, w_015_2884, w_015_2885, w_015_2886, w_015_2887, w_015_2889, w_015_2890, w_015_2891, w_015_2892, w_015_2893, w_015_2894, w_015_2895, w_015_2896, w_015_2897, w_015_2898, w_015_2900, w_015_2902, w_015_2906, w_015_2907, w_015_2911, w_015_2912, w_015_2914, w_015_2915, w_015_2916, w_015_2917, w_015_2918, w_015_2919, w_015_2920, w_015_2922, w_015_2923, w_015_2924, w_015_2925, w_015_2927, w_015_2930, w_015_2931, w_015_2932, w_015_2933, w_015_2935, w_015_2936, w_015_2937, w_015_2938, w_015_2939, w_015_2940, w_015_2941, w_015_2942, w_015_2943, w_015_2945, w_015_2948, w_015_2949, w_015_2950, w_015_2953, w_015_2954, w_015_2955, w_015_2956, w_015_2960, w_015_2962, w_015_2963, w_015_2964, w_015_2967, w_015_2968, w_015_2969, w_015_2970, w_015_2971, w_015_2972, w_015_2973, w_015_2974, w_015_2975, w_015_2976, w_015_2978, w_015_2979, w_015_2981, w_015_2982, w_015_2983, w_015_2985, w_015_2986, w_015_2987, w_015_2988, w_015_2989, w_015_2990, w_015_2991, w_015_2992, w_015_2993, w_015_2996, w_015_2997, w_015_2998, w_015_2999, w_015_3000, w_015_3001, w_015_3002, w_015_3007, w_015_3008, w_015_3011, w_015_3012, w_015_3013, w_015_3014, w_015_3015, w_015_3016, w_015_3017, w_015_3018, w_015_3019, w_015_3020, w_015_3021, w_015_3022, w_015_3023, w_015_3026, w_015_3028, w_015_3029, w_015_3030, w_015_3031, w_015_3032, w_015_3033, w_015_3034, w_015_3035, w_015_3036, w_015_3037, w_015_3038, w_015_3039, w_015_3041, w_015_3042, w_015_3045, w_015_3046, w_015_3047, w_015_3048, w_015_3049, w_015_3051, w_015_3052, w_015_3053, w_015_3054, w_015_3056, w_015_3057, w_015_3058, w_015_3062, w_015_3063, w_015_3064, w_015_3065, w_015_3066, w_015_3067, w_015_3068, w_015_3069, w_015_3071, w_015_3072, w_015_3073, w_015_3074, w_015_3075, w_015_3076, w_015_3078, w_015_3079, w_015_3080, w_015_3082, w_015_3083, w_015_3084, w_015_3085, w_015_3086, w_015_3087, w_015_3088, w_015_3090, w_015_3092, w_015_3096, w_015_3097, w_015_3098, w_015_3099, w_015_3100, w_015_3101, w_015_3102, w_015_3103, w_015_3104, w_015_3105, w_015_3106, w_015_3107, w_015_3108, w_015_3109, w_015_3110, w_015_3111, w_015_3112, w_015_3114, w_015_3115, w_015_3116, w_015_3117, w_015_3118, w_015_3119, w_015_3120, w_015_3121, w_015_3122, w_015_3125, w_015_3126, w_015_3128, w_015_3131, w_015_3134, w_015_3135, w_015_3137, w_015_3138, w_015_3139, w_015_3141, w_015_3142, w_015_3143, w_015_3144, w_015_3146, w_015_3147, w_015_3148, w_015_3149, w_015_3150, w_015_3151, w_015_3152, w_015_3153, w_015_3154, w_015_3155, w_015_3156, w_015_3157, w_015_3158, w_015_3159, w_015_3160, w_015_3161, w_015_3163, w_015_3164, w_015_3165, w_015_3166, w_015_3167, w_015_3169, w_015_3171, w_015_3172, w_015_3173, w_015_3174, w_015_3175, w_015_3177, w_015_3178, w_015_3179, w_015_3180, w_015_3182, w_015_3183, w_015_3184, w_015_3185, w_015_3186, w_015_3187, w_015_3188, w_015_3189, w_015_3190, w_015_3191, w_015_3192, w_015_3194, w_015_3197, w_015_3198, w_015_3199, w_015_3200, w_015_3201, w_015_3204, w_015_3205, w_015_3207, w_015_3208, w_015_3210, w_015_3211, w_015_3212, w_015_3213, w_015_3214, w_015_3215, w_015_3216, w_015_3218, w_015_3219, w_015_3220, w_015_3221, w_015_3222, w_015_3223, w_015_3224, w_015_3225, w_015_3226, w_015_3229, w_015_3230, w_015_3233, w_015_3234, w_015_3236, w_015_3237, w_015_3238, w_015_3239, w_015_3242, w_015_3243, w_015_3244, w_015_3245, w_015_3246, w_015_3247, w_015_3248, w_015_3250, w_015_3252, w_015_3254, w_015_3256, w_015_3257, w_015_3260, w_015_3261, w_015_3262, w_015_3263, w_015_3264, w_015_3265, w_015_3266, w_015_3267, w_015_3269, w_015_3270, w_015_3271, w_015_3272, w_015_3273, w_015_3277, w_015_3279, w_015_3280, w_015_3281, w_015_3282, w_015_3283, w_015_3285, w_015_3288, w_015_3289, w_015_3290, w_015_3291, w_015_3292, w_015_3293, w_015_3294, w_015_3295, w_015_3296, w_015_3297, w_015_3298, w_015_3301, w_015_3304, w_015_3305, w_015_3306, w_015_3307, w_015_3308, w_015_3311, w_015_3312, w_015_3313, w_015_3314, w_015_3315, w_015_3317, w_015_3321, w_015_3323, w_015_3324, w_015_3325, w_015_3326, w_015_3327, w_015_3330, w_015_3331, w_015_3334, w_015_3336, w_015_3337, w_015_3338, w_015_3340, w_015_3344, w_015_3345, w_015_3346, w_015_3348, w_015_3350, w_015_3351, w_015_3352, w_015_3353, w_015_3354, w_015_3355, w_015_3356, w_015_3357, w_015_3358, w_015_3360, w_015_3361, w_015_3362, w_015_3364, w_015_3365, w_015_3370, w_015_3371, w_015_3374, w_015_3375, w_015_3379, w_015_3381, w_015_3383, w_015_3384, w_015_3386, w_015_3387, w_015_3388, w_015_3392, w_015_3393, w_015_3395, w_015_3397, w_015_3398, w_015_3399, w_015_3400, w_015_3401, w_015_3402, w_015_3405, w_015_3406, w_015_3407, w_015_3408, w_015_3409, w_015_3410, w_015_3411, w_015_3412, w_015_3413, w_015_3414, w_015_3415, w_015_3417, w_015_3418, w_015_3419, w_015_3420, w_015_3421, w_015_3422, w_015_3423, w_015_3424, w_015_3427, w_015_3428, w_015_3429, w_015_3430, w_015_3431, w_015_3432, w_015_3436, w_015_3437, w_015_3439, w_015_3440, w_015_3441, w_015_3442, w_015_3444, w_015_3445, w_015_3447, w_015_3448, w_015_3449, w_015_3450, w_015_3451, w_015_3453, w_015_3454, w_015_3455, w_015_3456, w_015_3457, w_015_3458, w_015_3459, w_015_3460, w_015_3461, w_015_3462, w_015_3467, w_015_3469, w_015_3470, w_015_3471, w_015_3472, w_015_3473, w_015_3474, w_015_3475, w_015_3476, w_015_3477, w_015_3478, w_015_3480, w_015_3481, w_015_3483, w_015_3485, w_015_3486, w_015_3488, w_015_3491, w_015_3492, w_015_3493, w_015_3494, w_015_3495, w_015_3497, w_015_3498, w_015_3499, w_015_3500, w_015_3501, w_015_3504, w_015_3505, w_015_3506, w_015_3507, w_015_3509, w_015_3511, w_015_3512, w_015_3513, w_015_3514, w_015_3515, w_015_3516, w_015_3517, w_015_3518, w_015_3519, w_015_3520, w_015_3522, w_015_3523, w_015_3524, w_015_3526, w_015_3527, w_015_3528, w_015_3529, w_015_3532, w_015_3534, w_015_3536, w_015_3537, w_015_3538, w_015_3539, w_015_3540, w_015_3541, w_015_3542, w_015_3543, w_015_3544, w_015_3545, w_015_3546, w_015_3547, w_015_3549, w_015_3551, w_015_3552, w_015_3553, w_015_3554, w_015_3555, w_015_3557, w_015_3558, w_015_3559, w_015_3560, w_015_3561, w_015_3562, w_015_3564, w_015_3565, w_015_3566, w_015_3567, w_015_3568, w_015_3569, w_015_3572, w_015_3573, w_015_3574, w_015_3575, w_015_3576, w_015_3577, w_015_3579, w_015_3580, w_015_3583, w_015_3584, w_015_3585, w_015_3586, w_015_3587, w_015_3588, w_015_3589, w_015_3591, w_015_3592, w_015_3594, w_015_3596, w_015_3597, w_015_3601, w_015_3602, w_015_3603, w_015_3605, w_015_3606, w_015_3607, w_015_3608, w_015_3609, w_015_3611, w_015_3612, w_015_3613, w_015_3614, w_015_3615, w_015_3616, w_015_3617, w_015_3620, w_015_3623, w_015_3624, w_015_3625, w_015_3626, w_015_3627, w_015_3628, w_015_3629, w_015_3630, w_015_3631, w_015_3632, w_015_3633, w_015_3634, w_015_3635, w_015_3637, w_015_3638, w_015_3639, w_015_3640, w_015_3641, w_015_3642, w_015_3643, w_015_3644, w_015_3646, w_015_3647, w_015_3648, w_015_3649, w_015_3650, w_015_3651, w_015_3652, w_015_3656, w_015_3657, w_015_3658, w_015_3662, w_015_3663, w_015_3664, w_015_3665, w_015_3666, w_015_3667, w_015_3671, w_015_3672, w_015_3674, w_015_3675, w_015_3676, w_015_3677, w_015_3680, w_015_3681, w_015_3682, w_015_3683, w_015_3684, w_015_3686, w_015_3687, w_015_3688, w_015_3689, w_015_3691, w_015_3692, w_015_3693, w_015_3694, w_015_3695, w_015_3697, w_015_3698, w_015_3699, w_015_3700, w_015_3701, w_015_3702, w_015_3704, w_015_3705, w_015_3706, w_015_3709, w_015_3711, w_015_3713, w_015_3714, w_015_3716, w_015_3717, w_015_3718, w_015_3719, w_015_3722, w_015_3725, w_015_3726, w_015_3727, w_015_3728, w_015_3730, w_015_3731, w_015_3732, w_015_3733, w_015_3737, w_015_3738, w_015_3739, w_015_3740, w_015_3743, w_015_3744, w_015_3745, w_015_3746, w_015_3747, w_015_3748, w_015_3750, w_015_3751, w_015_3752, w_015_3753, w_015_3755, w_015_3756, w_015_3758, w_015_3759, w_015_3761, w_015_3765, w_015_3767, w_015_3768, w_015_3769, w_015_3770, w_015_3771, w_015_3772, w_015_3773, w_015_3774, w_015_3775, w_015_3777, w_015_3779, w_015_3780, w_015_3781, w_015_3782, w_015_3783, w_015_3787, w_015_3788, w_015_3789, w_015_3790, w_015_3791, w_015_3793, w_015_3794, w_015_3795, w_015_3797, w_015_3798, w_015_3799, w_015_3800, w_015_3801, w_015_3802, w_015_3803, w_015_3804, w_015_3805, w_015_3807, w_015_3808, w_015_3809, w_015_3811, w_015_3812, w_015_3813, w_015_3814, w_015_3815, w_015_3816, w_015_3817, w_015_3818, w_015_3819, w_015_3820, w_015_3821, w_015_3822, w_015_3823, w_015_3825, w_015_3826, w_015_3828, w_015_3829, w_015_3830, w_015_3831, w_015_3833, w_015_3834, w_015_3835, w_015_3836, w_015_3837, w_015_3839, w_015_3841, w_015_3842, w_015_3843, w_015_3844, w_015_3845, w_015_3846, w_015_3847, w_015_3848, w_015_3849, w_015_3850, w_015_3851, w_015_3852, w_015_3853, w_015_3854, w_015_3856, w_015_3857, w_015_3859, w_015_3861, w_015_3862, w_015_3865, w_015_3866, w_015_3867, w_015_3868, w_015_3869, w_015_3871, w_015_3872, w_015_3873, w_015_3874, w_015_3875, w_015_3876, w_015_3877, w_015_3878, w_015_3879, w_015_3880, w_015_3881, w_015_3882, w_015_3883, w_015_3884, w_015_3885, w_015_3886, w_015_3887, w_015_3889, w_015_3890, w_015_3891, w_015_3892, w_015_3893, w_015_3894, w_015_3895, w_015_3896, w_015_3897, w_015_3899, w_015_3902, w_015_3904, w_015_3905, w_015_3906, w_015_3908, w_015_3909, w_015_3910, w_015_3911, w_015_3912, w_015_3913, w_015_3914, w_015_3915, w_015_3916, w_015_3918, w_015_3919, w_015_3920, w_015_3921, w_015_3922, w_015_3923, w_015_3924, w_015_3925, w_015_3927, w_015_3928, w_015_3930, w_015_3933, w_015_3934, w_015_3936, w_015_3937, w_015_3938, w_015_3939, w_015_3941, w_015_3943, w_015_3944, w_015_3945, w_015_3947, w_015_3948, w_015_3950, w_015_3951, w_015_3953, w_015_3954, w_015_3955, w_015_3956, w_015_3957, w_015_3959, w_015_3961, w_015_3962, w_015_3963, w_015_3964, w_015_3965, w_015_3966, w_015_3967, w_015_3968, w_015_3969, w_015_3970, w_015_3971, w_015_3973, w_015_3975, w_015_3976, w_015_3977, w_015_3979, w_015_3980, w_015_3981, w_015_3982, w_015_3983, w_015_3984, w_015_3985, w_015_3986, w_015_3987, w_015_3988, w_015_3989, w_015_3991, w_015_3992, w_015_3995, w_015_3996, w_015_3997, w_015_3998, w_015_3999, w_015_4000, w_015_4002, w_015_4003, w_015_4004, w_015_4005, w_015_4007, w_015_4008, w_015_4010, w_015_4011, w_015_4012, w_015_4013, w_015_4014, w_015_4015, w_015_4016, w_015_4018, w_015_4019, w_015_4020, w_015_4021, w_015_4022, w_015_4024, w_015_4025, w_015_4026, w_015_4027, w_015_4031, w_015_4033, w_015_4034, w_015_4035, w_015_4036, w_015_4040, w_015_4041, w_015_4043, w_015_4044, w_015_4045, w_015_4046, w_015_4047, w_015_4048, w_015_4049, w_015_4051, w_015_4052, w_015_4053, w_015_4055, w_015_4057, w_015_4059, w_015_4061, w_015_4063, w_015_4064, w_015_4065, w_015_4066, w_015_4067, w_015_4068, w_015_4069, w_015_4070, w_015_4072, w_015_4073, w_015_4074, w_015_4075, w_015_4076, w_015_4077, w_015_4078, w_015_4079, w_015_4080, w_015_4081, w_015_4082, w_015_4083, w_015_4085, w_015_4087, w_015_4088, w_015_4090, w_015_4091, w_015_4092, w_015_4094, w_015_4095, w_015_4097, w_015_4098, w_015_4100, w_015_4102, w_015_4103, w_015_4104, w_015_4105, w_015_4106, w_015_4107, w_015_4108, w_015_4109, w_015_4110, w_015_4111, w_015_4112, w_015_4114, w_015_4116, w_015_4117, w_015_4118, w_015_4119, w_015_4120, w_015_4121, w_015_4122, w_015_4123, w_015_4125, w_015_4126, w_015_4127, w_015_4128, w_015_4129, w_015_4130, w_015_4131, w_015_4132, w_015_4133, w_015_4134, w_015_4135, w_015_4136, w_015_4137, w_015_4142, w_015_4144, w_015_4145, w_015_4146, w_015_4147, w_015_4149, w_015_4150, w_015_4151, w_015_4152, w_015_4154, w_015_4155, w_015_4157, w_015_4159, w_015_4160, w_015_4161, w_015_4163, w_015_4166, w_015_4168, w_015_4169, w_015_4170, w_015_4171, w_015_4172, w_015_4173, w_015_4174, w_015_4175, w_015_4176, w_015_4177, w_015_4178, w_015_4179, w_015_4180, w_015_4181, w_015_4182, w_015_4183, w_015_4186, w_015_4188, w_015_4189, w_015_4190, w_015_4191, w_015_4195, w_015_4196, w_015_4197, w_015_4198, w_015_4199, w_015_4200, w_015_4203, w_015_4204, w_015_4205, w_015_4206, w_015_4207, w_015_4208, w_015_4209, w_015_4210, w_015_4212, w_015_4213, w_015_4214, w_015_4215, w_015_4216, w_015_4217, w_015_4218, w_015_4220, w_015_4223, w_015_4224, w_015_4225, w_015_4226, w_015_4227, w_015_4229, w_015_4230, w_015_4231, w_015_4232, w_015_4234, w_015_4235, w_015_4236, w_015_4237, w_015_4242, w_015_4244, w_015_4246, w_015_4247, w_015_4248, w_015_4249, w_015_4251, w_015_4252, w_015_4253, w_015_4254, w_015_4255, w_015_4256, w_015_4257, w_015_4258, w_015_4259, w_015_4260, w_015_4261, w_015_4263, w_015_4266, w_015_4267, w_015_4268, w_015_4269, w_015_4270, w_015_4271, w_015_4272, w_015_4273, w_015_4274, w_015_4275, w_015_4276, w_015_4279, w_015_4280, w_015_4282, w_015_4283, w_015_4284, w_015_4285, w_015_4286, w_015_4287, w_015_4288, w_015_4292, w_015_4293, w_015_4294, w_015_4295, w_015_4296, w_015_4297, w_015_4298, w_015_4299, w_015_4300, w_015_4301, w_015_4304, w_015_4305, w_015_4306, w_015_4307, w_015_4309, w_015_4310, w_015_4311, w_015_4312, w_015_4315, w_015_4316, w_015_4317, w_015_4318, w_015_4320, w_015_4321, w_015_4323, w_015_4324, w_015_4325, w_015_4327, w_015_4328, w_015_4329, w_015_4330, w_015_4331, w_015_4332, w_015_4333, w_015_4334, w_015_4336, w_015_4337, w_015_4338, w_015_4339, w_015_4340, w_015_4341, w_015_4342, w_015_4344, w_015_4345, w_015_4346, w_015_4347, w_015_4348, w_015_4349, w_015_4350, w_015_4351, w_015_4353, w_015_4354, w_015_4355, w_015_4356, w_015_4358, w_015_4359, w_015_4360, w_015_4361, w_015_4362, w_015_4363, w_015_4364, w_015_4365, w_015_4366, w_015_4368, w_015_4369, w_015_4371, w_015_4372, w_015_4373, w_015_4374, w_015_4375, w_015_4376, w_015_4378, w_015_4379, w_015_4380, w_015_4381, w_015_4383, w_015_4384, w_015_4385, w_015_4386, w_015_4390, w_015_4391, w_015_4392, w_015_4393, w_015_4394, w_015_4396, w_015_4397, w_015_4398, w_015_4399, w_015_4400, w_015_4401, w_015_4402, w_015_4403, w_015_4404, w_015_4406, w_015_4408, w_015_4409, w_015_4410, w_015_4411, w_015_4415, w_015_4416, w_015_4417, w_015_4418, w_015_4419, w_015_4421, w_015_4422, w_015_4423, w_015_4424, w_015_4426, w_015_4427, w_015_4429, w_015_4430, w_015_4431, w_015_4434, w_015_4435, w_015_4437, w_015_4439, w_015_4442, w_015_4445, w_015_4447, w_015_4448, w_015_4449, w_015_4454, w_015_4455, w_015_4456, w_015_4457, w_015_4458, w_015_4459, w_015_4460, w_015_4464, w_015_4465, w_015_4466, w_015_4469, w_015_4470, w_015_4472, w_015_4473, w_015_4474, w_015_4475, w_015_4476, w_015_4477, w_015_4478, w_015_4479, w_015_4481, w_015_4482, w_015_4483, w_015_4484, w_015_4485, w_015_4488, w_015_4489, w_015_4490, w_015_4491, w_015_4493, w_015_4494, w_015_4496, w_015_4498, w_015_4499, w_015_4501, w_015_4504, w_015_4505, w_015_4506, w_015_4507, w_015_4509, w_015_4510, w_015_4512, w_015_4513, w_015_4516, w_015_4518, w_015_4519, w_015_4520, w_015_4522, w_015_4523, w_015_4524, w_015_4525, w_015_4526, w_015_4527, w_015_4529, w_015_4530, w_015_4532, w_015_4534, w_015_4535, w_015_4536, w_015_4537, w_015_4538, w_015_4539, w_015_4540, w_015_4542, w_015_4544, w_015_4545, w_015_4547, w_015_4548, w_015_4549, w_015_4550, w_015_4551, w_015_4552, w_015_4554, w_015_4555, w_015_4558, w_015_4559, w_015_4560, w_015_4561, w_015_4563, w_015_4564, w_015_4566, w_015_4567, w_015_4568, w_015_4569, w_015_4571, w_015_4572, w_015_4573, w_015_4574, w_015_4575, w_015_4576, w_015_4578, w_015_4579, w_015_4583, w_015_4584, w_015_4588, w_015_4589, w_015_4590, w_015_4591, w_015_4592, w_015_4593, w_015_4594, w_015_4595, w_015_4598, w_015_4600, w_015_4601, w_015_4602, w_015_4603, w_015_4604, w_015_4605, w_015_4607, w_015_4608, w_015_4609, w_015_4610, w_015_4611, w_015_4612, w_015_4613, w_015_4614, w_015_4615, w_015_4616, w_015_4618, w_015_4619, w_015_4620, w_015_4621, w_015_4622, w_015_4623, w_015_4624, w_015_4625, w_015_4627, w_015_4628, w_015_4629, w_015_4630, w_015_4631, w_015_4632, w_015_4633, w_015_4635, w_015_4636, w_015_4637, w_015_4638, w_015_4639, w_015_4641, w_015_4643, w_015_4644, w_015_4645, w_015_4646, w_015_4649, w_015_4650, w_015_4651, w_015_4652, w_015_4653, w_015_4656, w_015_4660, w_015_4661, w_015_4662, w_015_4665, w_015_4666, w_015_4667, w_015_4668, w_015_4669, w_015_4670, w_015_4672, w_015_4673, w_015_4675, w_015_4676, w_015_4677, w_015_4678, w_015_4679, w_015_4680, w_015_4681, w_015_4685, w_015_4687, w_015_4688, w_015_4689, w_015_4690, w_015_4691, w_015_4693, w_015_4694, w_015_4695, w_015_4696, w_015_4699, w_015_4700, w_015_4701, w_015_4703, w_015_4704, w_015_4705, w_015_4706, w_015_4707, w_015_4708, w_015_4709, w_015_4711, w_015_4712, w_015_4715, w_015_4716, w_015_4718, w_015_4719, w_015_4720, w_015_4721, w_015_4722, w_015_4723, w_015_4725, w_015_4726, w_015_4728, w_015_4730, w_015_4731, w_015_4732, w_015_4734, w_015_4735, w_015_4737, w_015_4738, w_015_4739, w_015_4740, w_015_4741, w_015_4742, w_015_4743, w_015_4744, w_015_4745, w_015_4747, w_015_4748, w_015_4749, w_015_4750, w_015_4751, w_015_4752, w_015_4753, w_015_4755, w_015_4756, w_015_4757, w_015_4758, w_015_4759, w_015_4760, w_015_4761, w_015_4762, w_015_4763, w_015_4765, w_015_4766, w_015_4767, w_015_4770, w_015_4771, w_015_4772, w_015_4774, w_015_4775, w_015_4776, w_015_4777, w_015_4779, w_015_4780, w_015_4781, w_015_4782, w_015_4783, w_015_4784, w_015_4785, w_015_4787, w_015_4788, w_015_4789, w_015_4790, w_015_4792, w_015_4798, w_015_4799, w_015_4800, w_015_4801, w_015_4802, w_015_4803, w_015_4805, w_015_4806, w_015_4808, w_015_4809, w_015_4810, w_015_4811, w_015_4812, w_015_4813, w_015_4814, w_015_4816, w_015_4817, w_015_4821, w_015_4822, w_015_4823, w_015_4825, w_015_4826, w_015_4830, w_015_4831, w_015_4832, w_015_4834, w_015_4835, w_015_4836, w_015_4837, w_015_4839, w_015_4841, w_015_4842, w_015_4844, w_015_4845, w_015_4846, w_015_4848, w_015_4849, w_015_4850, w_015_4851, w_015_4852, w_015_4853, w_015_4855, w_015_4857, w_015_4858, w_015_4859, w_015_4860, w_015_4861, w_015_4862, w_015_4865, w_015_4867, w_015_4868, w_015_4870, w_015_4871, w_015_4873, w_015_4874, w_015_4875, w_015_4876, w_015_4877, w_015_4878, w_015_4880, w_015_4881, w_015_4882, w_015_4883, w_015_4884, w_015_4886, w_015_4888, w_015_4889, w_015_4890, w_015_4891, w_015_4893, w_015_4895, w_015_4896, w_015_4897, w_015_4898, w_015_4899, w_015_4900, w_015_4901, w_015_4902, w_015_4903, w_015_4904, w_015_4905, w_015_4906, w_015_4907, w_015_4909, w_015_4910, w_015_4911, w_015_4912, w_015_4914, w_015_4915, w_015_4916, w_015_4919, w_015_4920, w_015_4922, w_015_4923, w_015_4924, w_015_4925, w_015_4926, w_015_4928, w_015_4929, w_015_4931, w_015_4932, w_015_4933, w_015_4934, w_015_4936, w_015_4937, w_015_4938, w_015_4940, w_015_4941, w_015_4943, w_015_4945, w_015_4946, w_015_4947, w_015_4948, w_015_4949, w_015_4950, w_015_4951, w_015_4952, w_015_4953, w_015_4954, w_015_4955, w_015_4956;
  wire w_016_001, w_016_002, w_016_003, w_016_004, w_016_005, w_016_006, w_016_007, w_016_008, w_016_009, w_016_010, w_016_011, w_016_012, w_016_013, w_016_014, w_016_015, w_016_016, w_016_017, w_016_018, w_016_019, w_016_020, w_016_022, w_016_023, w_016_024, w_016_025, w_016_026, w_016_027, w_016_028, w_016_029, w_016_030, w_016_031, w_016_032, w_016_033, w_016_034, w_016_035, w_016_036, w_016_037, w_016_038, w_016_039, w_016_040, w_016_041, w_016_042, w_016_043, w_016_044, w_016_045, w_016_046, w_016_047, w_016_048, w_016_049, w_016_050, w_016_051, w_016_052, w_016_053, w_016_055, w_016_056, w_016_057, w_016_058, w_016_059, w_016_060, w_016_061, w_016_062, w_016_063, w_016_064, w_016_065, w_016_066, w_016_067, w_016_068, w_016_069, w_016_071, w_016_072, w_016_073, w_016_074, w_016_075, w_016_076, w_016_077, w_016_078, w_016_080, w_016_081, w_016_082, w_016_083, w_016_084, w_016_086, w_016_087, w_016_088, w_016_090, w_016_091, w_016_092, w_016_093, w_016_095, w_016_096, w_016_097, w_016_098, w_016_099, w_016_100, w_016_101, w_016_102, w_016_103, w_016_104, w_016_105, w_016_106, w_016_107, w_016_109, w_016_110, w_016_111, w_016_112, w_016_113, w_016_114, w_016_115, w_016_116, w_016_117, w_016_118, w_016_120, w_016_121, w_016_122, w_016_123, w_016_124, w_016_125, w_016_126, w_016_127, w_016_128, w_016_130, w_016_131, w_016_132, w_016_133, w_016_134, w_016_135, w_016_136, w_016_137, w_016_138, w_016_139, w_016_140, w_016_141, w_016_142, w_016_143, w_016_146, w_016_147, w_016_148, w_016_149, w_016_150, w_016_151, w_016_154, w_016_155, w_016_156, w_016_157, w_016_158, w_016_159, w_016_160, w_016_161, w_016_162, w_016_163, w_016_164, w_016_165, w_016_166, w_016_167, w_016_168, w_016_169, w_016_170, w_016_173, w_016_174, w_016_175, w_016_176, w_016_177, w_016_178, w_016_179, w_016_180, w_016_181, w_016_182, w_016_183, w_016_184, w_016_185, w_016_186, w_016_187, w_016_188, w_016_189, w_016_190, w_016_191, w_016_192, w_016_193, w_016_194, w_016_195, w_016_196, w_016_197, w_016_198, w_016_199, w_016_200, w_016_201, w_016_202, w_016_203, w_016_204, w_016_205, w_016_206, w_016_207, w_016_208, w_016_209, w_016_210, w_016_211, w_016_213, w_016_214, w_016_215, w_016_216, w_016_217, w_016_218, w_016_219, w_016_220, w_016_221, w_016_222, w_016_223, w_016_224, w_016_225, w_016_226, w_016_227, w_016_228, w_016_229, w_016_230, w_016_232, w_016_233, w_016_234, w_016_235, w_016_236, w_016_237, w_016_238, w_016_239, w_016_240, w_016_241, w_016_242, w_016_243, w_016_244, w_016_246, w_016_247, w_016_248, w_016_249, w_016_250, w_016_251, w_016_252, w_016_253, w_016_254, w_016_255, w_016_256, w_016_257, w_016_258, w_016_259, w_016_260, w_016_261, w_016_262, w_016_264, w_016_265, w_016_266, w_016_267, w_016_268, w_016_269, w_016_270, w_016_271, w_016_272, w_016_273, w_016_274, w_016_275, w_016_276, w_016_278, w_016_279, w_016_280, w_016_281, w_016_282, w_016_283, w_016_284, w_016_285, w_016_286, w_016_287, w_016_288, w_016_289, w_016_290, w_016_291, w_016_292, w_016_293, w_016_295, w_016_296, w_016_297, w_016_298, w_016_299, w_016_300, w_016_301, w_016_302, w_016_303, w_016_304, w_016_305, w_016_306, w_016_307, w_016_308, w_016_309, w_016_310, w_016_311, w_016_312, w_016_313, w_016_315, w_016_316, w_016_317, w_016_319, w_016_320, w_016_321, w_016_322, w_016_323, w_016_325, w_016_326, w_016_327, w_016_328, w_016_329, w_016_330, w_016_331, w_016_332, w_016_333, w_016_334, w_016_335, w_016_336, w_016_337, w_016_338, w_016_339, w_016_340, w_016_341, w_016_342, w_016_343, w_016_344, w_016_345, w_016_346, w_016_347, w_016_348, w_016_349, w_016_350, w_016_351, w_016_353, w_016_355, w_016_356, w_016_357, w_016_358, w_016_359, w_016_360, w_016_361, w_016_362, w_016_363, w_016_364, w_016_365, w_016_366, w_016_367, w_016_368, w_016_369, w_016_370, w_016_371, w_016_372, w_016_373, w_016_374, w_016_375, w_016_376, w_016_377, w_016_378, w_016_379, w_016_380, w_016_381, w_016_382, w_016_383, w_016_384, w_016_385, w_016_387, w_016_388, w_016_389, w_016_390, w_016_391, w_016_392, w_016_393, w_016_394, w_016_395, w_016_396, w_016_397, w_016_398, w_016_399, w_016_400, w_016_402, w_016_403, w_016_404, w_016_405, w_016_406, w_016_407, w_016_408, w_016_409, w_016_410, w_016_411, w_016_412, w_016_413, w_016_414, w_016_415, w_016_416, w_016_417, w_016_418, w_016_419, w_016_420, w_016_421, w_016_422, w_016_423, w_016_424, w_016_425, w_016_426, w_016_427, w_016_428, w_016_429, w_016_431, w_016_432, w_016_433, w_016_434, w_016_435, w_016_436, w_016_437, w_016_438, w_016_439, w_016_440, w_016_441, w_016_442, w_016_443, w_016_444, w_016_445, w_016_446, w_016_447, w_016_448, w_016_449, w_016_450, w_016_451, w_016_452, w_016_454, w_016_455, w_016_456, w_016_458, w_016_459, w_016_460, w_016_461, w_016_463, w_016_464, w_016_465, w_016_466, w_016_467, w_016_468, w_016_469, w_016_470, w_016_471, w_016_472, w_016_473, w_016_474, w_016_475, w_016_476, w_016_477, w_016_478, w_016_479, w_016_480, w_016_481, w_016_482, w_016_483, w_016_484, w_016_485, w_016_486, w_016_487, w_016_488, w_016_489, w_016_490, w_016_491, w_016_492, w_016_493, w_016_494, w_016_495, w_016_496, w_016_497, w_016_498, w_016_499, w_016_500, w_016_501, w_016_502, w_016_504, w_016_505, w_016_506, w_016_507, w_016_508, w_016_509, w_016_510, w_016_511, w_016_512, w_016_513, w_016_514, w_016_515, w_016_516, w_016_517, w_016_518, w_016_519, w_016_520, w_016_521, w_016_523, w_016_524, w_016_525, w_016_526, w_016_527, w_016_528, w_016_529, w_016_530, w_016_531, w_016_532, w_016_533, w_016_534, w_016_535, w_016_536, w_016_537, w_016_538, w_016_539, w_016_540, w_016_541, w_016_542, w_016_543, w_016_544, w_016_545, w_016_546, w_016_547, w_016_548, w_016_549, w_016_550, w_016_551, w_016_552, w_016_553, w_016_554, w_016_555, w_016_557, w_016_558, w_016_559, w_016_560, w_016_561, w_016_562, w_016_563, w_016_564, w_016_565, w_016_566, w_016_567, w_016_568, w_016_569, w_016_570, w_016_571, w_016_573, w_016_574, w_016_575, w_016_576, w_016_577, w_016_578, w_016_579, w_016_580, w_016_581, w_016_582, w_016_583, w_016_584, w_016_585, w_016_586, w_016_587, w_016_588, w_016_589, w_016_591, w_016_592, w_016_593, w_016_594, w_016_595, w_016_596, w_016_597, w_016_599, w_016_600, w_016_601, w_016_602, w_016_603, w_016_604, w_016_605, w_016_607, w_016_608, w_016_609, w_016_610, w_016_611, w_016_612, w_016_614, w_016_615, w_016_616, w_016_617, w_016_618, w_016_619, w_016_620, w_016_621, w_016_622, w_016_623, w_016_624, w_016_625, w_016_626, w_016_628, w_016_629, w_016_630, w_016_631, w_016_632, w_016_633, w_016_635, w_016_637, w_016_639, w_016_640, w_016_641, w_016_642, w_016_643, w_016_644, w_016_645, w_016_646, w_016_647, w_016_648, w_016_649, w_016_650, w_016_651, w_016_652, w_016_653, w_016_654, w_016_655, w_016_656, w_016_657, w_016_658, w_016_659, w_016_660, w_016_661, w_016_662, w_016_663, w_016_664, w_016_665, w_016_666, w_016_667, w_016_668, w_016_671, w_016_672, w_016_673, w_016_676, w_016_678, w_016_679, w_016_680, w_016_681, w_016_682, w_016_683, w_016_684, w_016_685, w_016_686, w_016_687, w_016_689, w_016_690, w_016_691, w_016_692, w_016_693, w_016_694, w_016_695, w_016_696, w_016_697, w_016_698, w_016_699, w_016_700, w_016_701, w_016_702, w_016_703, w_016_704, w_016_705, w_016_706, w_016_707, w_016_708, w_016_709, w_016_710, w_016_711, w_016_712, w_016_714, w_016_715, w_016_716, w_016_717, w_016_718, w_016_719, w_016_720, w_016_722, w_016_723, w_016_724, w_016_725, w_016_728, w_016_729, w_016_730, w_016_731, w_016_732, w_016_733, w_016_734, w_016_735, w_016_736, w_016_737, w_016_738, w_016_739, w_016_740, w_016_741, w_016_742, w_016_743, w_016_744, w_016_745, w_016_746, w_016_747, w_016_748, w_016_749, w_016_750, w_016_751, w_016_752, w_016_753, w_016_754, w_016_755, w_016_756, w_016_757, w_016_759, w_016_760, w_016_761, w_016_762, w_016_763, w_016_764, w_016_765, w_016_766, w_016_767, w_016_768, w_016_769, w_016_770, w_016_771, w_016_772, w_016_773, w_016_774, w_016_775, w_016_776, w_016_777, w_016_778, w_016_779, w_016_780, w_016_781, w_016_782, w_016_783, w_016_784, w_016_785, w_016_786, w_016_787, w_016_788, w_016_789, w_016_790, w_016_791, w_016_792, w_016_794, w_016_795, w_016_796, w_016_797, w_016_798, w_016_800, w_016_801, w_016_802, w_016_803, w_016_804, w_016_805, w_016_806, w_016_807, w_016_808, w_016_809, w_016_810, w_016_811, w_016_812, w_016_813, w_016_814, w_016_815, w_016_816, w_016_817, w_016_818, w_016_819, w_016_820, w_016_821, w_016_822, w_016_823, w_016_824, w_016_825, w_016_826, w_016_827, w_016_828, w_016_829, w_016_830, w_016_831, w_016_832, w_016_833, w_016_834, w_016_835, w_016_837, w_016_838, w_016_839, w_016_840, w_016_841, w_016_842, w_016_843, w_016_844, w_016_845, w_016_846, w_016_847, w_016_848, w_016_850, w_016_851, w_016_852, w_016_853, w_016_854, w_016_855, w_016_856, w_016_857, w_016_858, w_016_859, w_016_860, w_016_861, w_016_862, w_016_863, w_016_864, w_016_865, w_016_866, w_016_867, w_016_868, w_016_869, w_016_870, w_016_871, w_016_872, w_016_873, w_016_875, w_016_876, w_016_877, w_016_878, w_016_879, w_016_880, w_016_881, w_016_882, w_016_884, w_016_885, w_016_887, w_016_888, w_016_889, w_016_890, w_016_891, w_016_892, w_016_893, w_016_894, w_016_895, w_016_896, w_016_897, w_016_898, w_016_899, w_016_900, w_016_901, w_016_902, w_016_903, w_016_904, w_016_905, w_016_906, w_016_907, w_016_908, w_016_909, w_016_910, w_016_912, w_016_913, w_016_914, w_016_915, w_016_917, w_016_918, w_016_919, w_016_920, w_016_921, w_016_922, w_016_923, w_016_924, w_016_925, w_016_926, w_016_927, w_016_928, w_016_929, w_016_930, w_016_931, w_016_932, w_016_933, w_016_934, w_016_935, w_016_936, w_016_937, w_016_938, w_016_939, w_016_940, w_016_941, w_016_942, w_016_943, w_016_944, w_016_945, w_016_946, w_016_947, w_016_948, w_016_949, w_016_950, w_016_951, w_016_952, w_016_954, w_016_955, w_016_956, w_016_958, w_016_959, w_016_960, w_016_961, w_016_962, w_016_963, w_016_964, w_016_965, w_016_966, w_016_967, w_016_968, w_016_969, w_016_970, w_016_971, w_016_972, w_016_973, w_016_974, w_016_975, w_016_976, w_016_978, w_016_979, w_016_980, w_016_981, w_016_982, w_016_983, w_016_984, w_016_985, w_016_986, w_016_987, w_016_988, w_016_989, w_016_990, w_016_991, w_016_992, w_016_993, w_016_994, w_016_995, w_016_996, w_016_997, w_016_998, w_016_999, w_016_1000, w_016_1001, w_016_1002, w_016_1003, w_016_1005, w_016_1006, w_016_1007, w_016_1008, w_016_1009, w_016_1010, w_016_1011, w_016_1012, w_016_1013, w_016_1014, w_016_1015, w_016_1016, w_016_1018, w_016_1019, w_016_1020, w_016_1021, w_016_1022, w_016_1023, w_016_1024, w_016_1025, w_016_1026, w_016_1027, w_016_1028, w_016_1029, w_016_1032, w_016_1035, w_016_1036, w_016_1037, w_016_1038, w_016_1039, w_016_1040, w_016_1041, w_016_1042, w_016_1044, w_016_1046, w_016_1047, w_016_1048, w_016_1050, w_016_1051, w_016_1052, w_016_1053, w_016_1054, w_016_1055, w_016_1056, w_016_1057, w_016_1058, w_016_1059, w_016_1060, w_016_1061, w_016_1062, w_016_1063, w_016_1064, w_016_1065, w_016_1066, w_016_1067, w_016_1068, w_016_1069, w_016_1070, w_016_1071, w_016_1072, w_016_1074, w_016_1075, w_016_1076, w_016_1077, w_016_1078, w_016_1079, w_016_1080, w_016_1081, w_016_1082, w_016_1083, w_016_1084, w_016_1085, w_016_1087, w_016_1088, w_016_1091, w_016_1092, w_016_1093, w_016_1094, w_016_1095, w_016_1096, w_016_1097, w_016_1098, w_016_1099, w_016_1100, w_016_1101, w_016_1102, w_016_1103, w_016_1104, w_016_1105, w_016_1106, w_016_1107, w_016_1108, w_016_1109, w_016_1110, w_016_1111, w_016_1112, w_016_1113, w_016_1115, w_016_1116, w_016_1117, w_016_1118, w_016_1120, w_016_1121, w_016_1122, w_016_1123, w_016_1124, w_016_1125, w_016_1126, w_016_1127, w_016_1128, w_016_1129, w_016_1130, w_016_1132, w_016_1133, w_016_1134, w_016_1135, w_016_1136, w_016_1137, w_016_1138, w_016_1139, w_016_1140, w_016_1141, w_016_1142, w_016_1143, w_016_1144, w_016_1145, w_016_1146, w_016_1147, w_016_1148, w_016_1149, w_016_1150, w_016_1151, w_016_1152, w_016_1154, w_016_1155, w_016_1156, w_016_1157, w_016_1158, w_016_1159, w_016_1160, w_016_1161, w_016_1162, w_016_1163, w_016_1164, w_016_1165, w_016_1166, w_016_1168, w_016_1169, w_016_1170, w_016_1173, w_016_1174, w_016_1175, w_016_1176, w_016_1177, w_016_1178, w_016_1179, w_016_1180, w_016_1181, w_016_1182, w_016_1183, w_016_1184, w_016_1185, w_016_1186, w_016_1187, w_016_1188, w_016_1189, w_016_1190, w_016_1191, w_016_1192, w_016_1193, w_016_1194, w_016_1195, w_016_1196, w_016_1197, w_016_1198, w_016_1199, w_016_1201, w_016_1202, w_016_1203, w_016_1204, w_016_1205, w_016_1206, w_016_1207, w_016_1208, w_016_1209, w_016_1210, w_016_1211, w_016_1212, w_016_1213, w_016_1214, w_016_1215, w_016_1216, w_016_1217, w_016_1218, w_016_1219, w_016_1220, w_016_1221, w_016_1222, w_016_1223, w_016_1224, w_016_1225, w_016_1226, w_016_1227, w_016_1228, w_016_1229, w_016_1230, w_016_1231, w_016_1232, w_016_1233, w_016_1234, w_016_1235, w_016_1236, w_016_1237, w_016_1238, w_016_1239, w_016_1240, w_016_1241, w_016_1242, w_016_1243, w_016_1244, w_016_1245, w_016_1246, w_016_1247, w_016_1248, w_016_1249, w_016_1251, w_016_1252, w_016_1253, w_016_1254, w_016_1255, w_016_1256, w_016_1257, w_016_1258, w_016_1259, w_016_1260, w_016_1261, w_016_1262, w_016_1263, w_016_1264, w_016_1265, w_016_1266, w_016_1267, w_016_1268, w_016_1269, w_016_1270, w_016_1271, w_016_1272, w_016_1273, w_016_1274, w_016_1275, w_016_1276, w_016_1277, w_016_1278, w_016_1279, w_016_1280, w_016_1281, w_016_1282, w_016_1283, w_016_1284, w_016_1285, w_016_1286, w_016_1289, w_016_1290, w_016_1291, w_016_1292, w_016_1293, w_016_1294, w_016_1295, w_016_1296, w_016_1298, w_016_1299, w_016_1300, w_016_1302, w_016_1303, w_016_1305, w_016_1306, w_016_1307, w_016_1308, w_016_1309, w_016_1310, w_016_1311, w_016_1312, w_016_1313, w_016_1314, w_016_1315, w_016_1316, w_016_1317, w_016_1318, w_016_1319, w_016_1320, w_016_1321, w_016_1322, w_016_1323, w_016_1324, w_016_1325, w_016_1326, w_016_1327, w_016_1328, w_016_1329, w_016_1330, w_016_1331, w_016_1332, w_016_1333, w_016_1335, w_016_1336, w_016_1338, w_016_1339, w_016_1341, w_016_1342, w_016_1343, w_016_1344, w_016_1345, w_016_1346, w_016_1347, w_016_1348, w_016_1349, w_016_1350, w_016_1351, w_016_1352, w_016_1353, w_016_1354, w_016_1355, w_016_1356, w_016_1357, w_016_1358, w_016_1359, w_016_1360, w_016_1361, w_016_1362, w_016_1363, w_016_1364, w_016_1365, w_016_1366, w_016_1367, w_016_1369, w_016_1371, w_016_1372, w_016_1373, w_016_1374, w_016_1375, w_016_1376, w_016_1377, w_016_1378, w_016_1379, w_016_1380, w_016_1381, w_016_1382, w_016_1383, w_016_1384, w_016_1385, w_016_1386, w_016_1387, w_016_1388, w_016_1389, w_016_1390, w_016_1391, w_016_1392, w_016_1393, w_016_1394, w_016_1395, w_016_1396, w_016_1397, w_016_1398, w_016_1399, w_016_1400, w_016_1401, w_016_1402, w_016_1403, w_016_1404, w_016_1405, w_016_1406, w_016_1407, w_016_1408, w_016_1409, w_016_1410, w_016_1411, w_016_1412, w_016_1413, w_016_1414, w_016_1415, w_016_1416, w_016_1417, w_016_1418, w_016_1419, w_016_1420, w_016_1421, w_016_1422, w_016_1423, w_016_1424, w_016_1425, w_016_1426, w_016_1427, w_016_1428, w_016_1429, w_016_1430, w_016_1431, w_016_1432, w_016_1433, w_016_1434, w_016_1435, w_016_1436, w_016_1437, w_016_1438, w_016_1439, w_016_1441, w_016_1444, w_016_1445, w_016_1446, w_016_1447, w_016_1449, w_016_1450, w_016_1451, w_016_1452, w_016_1455, w_016_1456, w_016_1457, w_016_1458, w_016_1459, w_016_1460, w_016_1461, w_016_1462, w_016_1463, w_016_1464, w_016_1465, w_016_1466, w_016_1467, w_016_1468, w_016_1469, w_016_1470, w_016_1471, w_016_1472, w_016_1474, w_016_1475, w_016_1476, w_016_1477, w_016_1478, w_016_1479, w_016_1480, w_016_1481, w_016_1482, w_016_1483, w_016_1484, w_016_1486, w_016_1487, w_016_1488, w_016_1489, w_016_1490, w_016_1491, w_016_1492, w_016_1493, w_016_1494, w_016_1495, w_016_1496, w_016_1497, w_016_1498, w_016_1499, w_016_1500, w_016_1501, w_016_1504, w_016_1505, w_016_1506, w_016_1509, w_016_1510, w_016_1511, w_016_1512, w_016_1513, w_016_1514, w_016_1515, w_016_1516, w_016_1518, w_016_1519, w_016_1520, w_016_1521, w_016_1522, w_016_1523, w_016_1524, w_016_1525, w_016_1527, w_016_1529, w_016_1530, w_016_1531, w_016_1533, w_016_1534, w_016_1535, w_016_1536, w_016_1537, w_016_1538, w_016_1541, w_016_1542, w_016_1543, w_016_1544, w_016_1545, w_016_1546, w_016_1547, w_016_1548, w_016_1550, w_016_1551, w_016_1553, w_016_1554, w_016_1555, w_016_1556, w_016_1557, w_016_1558, w_016_1559, w_016_1561, w_016_1564, w_016_1566, w_016_1569, w_016_1570, w_016_1571, w_016_1573, w_016_1574, w_016_1575, w_016_1577, w_016_1578, w_016_1579, w_016_1580, w_016_1581, w_016_1582, w_016_1583, w_016_1586, w_016_1588, w_016_1589, w_016_1590, w_016_1591, w_016_1592, w_016_1593, w_016_1594, w_016_1596, w_016_1597, w_016_1598, w_016_1600, w_016_1601, w_016_1602, w_016_1603, w_016_1604, w_016_1605, w_016_1607, w_016_1608, w_016_1609, w_016_1611, w_016_1612, w_016_1615, w_016_1617, w_016_1619, w_016_1620, w_016_1621, w_016_1622, w_016_1623, w_016_1626, w_016_1627, w_016_1628, w_016_1629, w_016_1630, w_016_1631, w_016_1632, w_016_1633, w_016_1634, w_016_1635, w_016_1636, w_016_1637, w_016_1638, w_016_1639, w_016_1640, w_016_1642, w_016_1643, w_016_1644, w_016_1645, w_016_1647, w_016_1648, w_016_1649, w_016_1650, w_016_1651, w_016_1654, w_016_1655, w_016_1656, w_016_1657, w_016_1658, w_016_1661, w_016_1662, w_016_1663, w_016_1664, w_016_1665, w_016_1666, w_016_1667, w_016_1668, w_016_1669, w_016_1670, w_016_1672, w_016_1673, w_016_1674, w_016_1675, w_016_1676, w_016_1678, w_016_1679, w_016_1681, w_016_1682, w_016_1683, w_016_1685, w_016_1686, w_016_1688, w_016_1691, w_016_1692, w_016_1693, w_016_1694, w_016_1696, w_016_1697, w_016_1699, w_016_1700, w_016_1701, w_016_1703, w_016_1704, w_016_1705, w_016_1709, w_016_1711, w_016_1712, w_016_1713, w_016_1714, w_016_1716, w_016_1717, w_016_1718, w_016_1719, w_016_1720, w_016_1721, w_016_1722, w_016_1723, w_016_1724, w_016_1725, w_016_1726, w_016_1728, w_016_1729, w_016_1730, w_016_1731, w_016_1732, w_016_1735, w_016_1736, w_016_1737, w_016_1738, w_016_1739, w_016_1740, w_016_1741, w_016_1742, w_016_1743, w_016_1745, w_016_1747, w_016_1748, w_016_1749, w_016_1751, w_016_1752, w_016_1753, w_016_1755, w_016_1756, w_016_1757, w_016_1758, w_016_1759, w_016_1760, w_016_1761, w_016_1763, w_016_1766, w_016_1768, w_016_1770, w_016_1771, w_016_1773, w_016_1774, w_016_1775, w_016_1776, w_016_1777, w_016_1778, w_016_1780, w_016_1782, w_016_1784, w_016_1786, w_016_1787, w_016_1788, w_016_1789, w_016_1790, w_016_1791, w_016_1793, w_016_1794, w_016_1795, w_016_1796, w_016_1797, w_016_1798, w_016_1799, w_016_1800, w_016_1801, w_016_1802, w_016_1803, w_016_1804, w_016_1806, w_016_1808, w_016_1809, w_016_1810, w_016_1812, w_016_1813, w_016_1815, w_016_1816, w_016_1817, w_016_1818, w_016_1819, w_016_1820, w_016_1821, w_016_1822, w_016_1823, w_016_1824, w_016_1826, w_016_1830, w_016_1831, w_016_1832, w_016_1835, w_016_1838, w_016_1839, w_016_1840, w_016_1841, w_016_1844, w_016_1845, w_016_1846, w_016_1847, w_016_1852, w_016_1853, w_016_1855, w_016_1857, w_016_1858, w_016_1859, w_016_1863, w_016_1864, w_016_1867, w_016_1869, w_016_1870, w_016_1873, w_016_1874, w_016_1875, w_016_1877, w_016_1878, w_016_1880, w_016_1881, w_016_1882, w_016_1883, w_016_1884, w_016_1885, w_016_1886, w_016_1887, w_016_1889, w_016_1891, w_016_1892, w_016_1894, w_016_1896, w_016_1897, w_016_1899, w_016_1901, w_016_1903, w_016_1904, w_016_1905, w_016_1906, w_016_1907, w_016_1909, w_016_1910, w_016_1911, w_016_1912, w_016_1913, w_016_1914, w_016_1915, w_016_1917, w_016_1918, w_016_1919, w_016_1920, w_016_1921, w_016_1922, w_016_1923, w_016_1925, w_016_1926, w_016_1927, w_016_1928, w_016_1929, w_016_1930, w_016_1934, w_016_1935, w_016_1937, w_016_1938, w_016_1939, w_016_1941, w_016_1942, w_016_1944, w_016_1946, w_016_1947, w_016_1948, w_016_1949, w_016_1950, w_016_1951, w_016_1952, w_016_1954, w_016_1955, w_016_1956, w_016_1957, w_016_1958, w_016_1961, w_016_1962, w_016_1963, w_016_1964, w_016_1965, w_016_1966, w_016_1968, w_016_1969, w_016_1970, w_016_1971, w_016_1974, w_016_1975, w_016_1976, w_016_1977, w_016_1982, w_016_1984, w_016_1985, w_016_1986, w_016_1987, w_016_1988, w_016_1990, w_016_1991, w_016_1992, w_016_1994, w_016_1997, w_016_1999, w_016_2002, w_016_2003, w_016_2004, w_016_2006, w_016_2007, w_016_2008, w_016_2009, w_016_2010, w_016_2011, w_016_2012, w_016_2013, w_016_2014, w_016_2016, w_016_2017, w_016_2021, w_016_2022, w_016_2024, w_016_2025, w_016_2026, w_016_2027, w_016_2028, w_016_2029, w_016_2030, w_016_2031, w_016_2033, w_016_2034, w_016_2035, w_016_2036, w_016_2037, w_016_2038, w_016_2039, w_016_2040, w_016_2041, w_016_2043, w_016_2045, w_016_2046, w_016_2048, w_016_2049, w_016_2050, w_016_2051, w_016_2052, w_016_2053, w_016_2054, w_016_2056, w_016_2057, w_016_2059, w_016_2060, w_016_2061, w_016_2062, w_016_2063, w_016_2064, w_016_2065, w_016_2067, w_016_2068, w_016_2071, w_016_2074, w_016_2075, w_016_2077, w_016_2078, w_016_2079, w_016_2082, w_016_2083, w_016_2085, w_016_2086, w_016_2087, w_016_2088, w_016_2089, w_016_2090, w_016_2091, w_016_2092, w_016_2094, w_016_2096, w_016_2097, w_016_2098, w_016_2100, w_016_2101, w_016_2102, w_016_2103, w_016_2105, w_016_2106, w_016_2107, w_016_2108, w_016_2110, w_016_2111, w_016_2112, w_016_2113, w_016_2115, w_016_2118, w_016_2119, w_016_2120, w_016_2122, w_016_2123, w_016_2124, w_016_2126, w_016_2127, w_016_2128, w_016_2130, w_016_2131, w_016_2134, w_016_2135, w_016_2136, w_016_2137, w_016_2138, w_016_2139, w_016_2141, w_016_2142, w_016_2143, w_016_2144, w_016_2146, w_016_2150, w_016_2151, w_016_2152, w_016_2154, w_016_2155, w_016_2157, w_016_2158, w_016_2161, w_016_2163, w_016_2164, w_016_2165, w_016_2166, w_016_2167, w_016_2172, w_016_2173, w_016_2175, w_016_2176, w_016_2177, w_016_2179, w_016_2180, w_016_2181, w_016_2183, w_016_2184, w_016_2185, w_016_2186, w_016_2187, w_016_2189, w_016_2193, w_016_2194, w_016_2195, w_016_2196, w_016_2197, w_016_2198, w_016_2199, w_016_2201, w_016_2202, w_016_2204, w_016_2205, w_016_2206, w_016_2208, w_016_2209, w_016_2210, w_016_2211, w_016_2212, w_016_2213, w_016_2214, w_016_2215, w_016_2216, w_016_2217, w_016_2218, w_016_2220, w_016_2222, w_016_2223, w_016_2224, w_016_2225, w_016_2226, w_016_2227, w_016_2230, w_016_2231, w_016_2235, w_016_2236, w_016_2237, w_016_2240, w_016_2241, w_016_2242, w_016_2244, w_016_2245, w_016_2246, w_016_2248, w_016_2249, w_016_2250, w_016_2253, w_016_2254, w_016_2255, w_016_2258, w_016_2261, w_016_2262, w_016_2265, w_016_2266, w_016_2267, w_016_2268, w_016_2269, w_016_2270, w_016_2272, w_016_2273, w_016_2274, w_016_2275, w_016_2276, w_016_2277, w_016_2279, w_016_2280, w_016_2281, w_016_2282, w_016_2283, w_016_2284, w_016_2285, w_016_2286, w_016_2287, w_016_2288, w_016_2289, w_016_2290, w_016_2293, w_016_2296, w_016_2297, w_016_2298, w_016_2299, w_016_2301, w_016_2302, w_016_2303, w_016_2304, w_016_2305, w_016_2307, w_016_2308, w_016_2310, w_016_2311, w_016_2312, w_016_2313, w_016_2314, w_016_2315, w_016_2317, w_016_2319, w_016_2320, w_016_2321, w_016_2323, w_016_2324, w_016_2326, w_016_2327, w_016_2328, w_016_2329, w_016_2331, w_016_2333, w_016_2334, w_016_2336, w_016_2338, w_016_2339, w_016_2340, w_016_2341, w_016_2342, w_016_2343, w_016_2345, w_016_2346, w_016_2348, w_016_2349, w_016_2350, w_016_2351, w_016_2352, w_016_2355, w_016_2356, w_016_2357, w_016_2358, w_016_2359, w_016_2360, w_016_2361, w_016_2362, w_016_2364, w_016_2365, w_016_2366, w_016_2367, w_016_2368, w_016_2369, w_016_2372, w_016_2373, w_016_2374, w_016_2375, w_016_2376, w_016_2378, w_016_2379, w_016_2380, w_016_2381, w_016_2383, w_016_2384, w_016_2385, w_016_2387, w_016_2389, w_016_2390, w_016_2391, w_016_2392, w_016_2393, w_016_2394, w_016_2397, w_016_2399, w_016_2400, w_016_2401, w_016_2404, w_016_2405, w_016_2406, w_016_2408, w_016_2409, w_016_2411, w_016_2412, w_016_2413, w_016_2414, w_016_2415, w_016_2416, w_016_2417, w_016_2418, w_016_2419, w_016_2420, w_016_2422, w_016_2425, w_016_2427, w_016_2428, w_016_2430, w_016_2431, w_016_2433, w_016_2434, w_016_2436, w_016_2437, w_016_2438, w_016_2439, w_016_2440, w_016_2441, w_016_2442, w_016_2443, w_016_2444, w_016_2445, w_016_2446, w_016_2447, w_016_2448, w_016_2449, w_016_2451, w_016_2452, w_016_2454, w_016_2455, w_016_2456, w_016_2458, w_016_2459, w_016_2460, w_016_2461, w_016_2464, w_016_2465, w_016_2466, w_016_2468, w_016_2470, w_016_2471, w_016_2472, w_016_2474, w_016_2475, w_016_2476, w_016_2477, w_016_2478, w_016_2481, w_016_2482, w_016_2483, w_016_2484, w_016_2485, w_016_2486, w_016_2488, w_016_2490, w_016_2491, w_016_2492, w_016_2493, w_016_2494, w_016_2497, w_016_2501, w_016_2503, w_016_2504, w_016_2505, w_016_2506, w_016_2507, w_016_2508, w_016_2509, w_016_2512, w_016_2513, w_016_2515, w_016_2517, w_016_2519, w_016_2520, w_016_2521, w_016_2524, w_016_2525, w_016_2526, w_016_2528, w_016_2529, w_016_2530, w_016_2531, w_016_2532, w_016_2533, w_016_2534, w_016_2535, w_016_2536, w_016_2537, w_016_2538, w_016_2539, w_016_2540, w_016_2541, w_016_2542, w_016_2543, w_016_2545, w_016_2546, w_016_2548, w_016_2549, w_016_2550, w_016_2551, w_016_2552, w_016_2554, w_016_2556, w_016_2557, w_016_2558, w_016_2559, w_016_2560, w_016_2561, w_016_2562, w_016_2563, w_016_2564, w_016_2566, w_016_2567, w_016_2569, w_016_2570, w_016_2571, w_016_2573, w_016_2574, w_016_2575, w_016_2576, w_016_2577, w_016_2578, w_016_2579, w_016_2580, w_016_2581, w_016_2582, w_016_2583, w_016_2585, w_016_2586, w_016_2587, w_016_2588, w_016_2589, w_016_2590, w_016_2592, w_016_2593, w_016_2594, w_016_2595, w_016_2596, w_016_2597, w_016_2598, w_016_2599, w_016_2600, w_016_2601, w_016_2602, w_016_2603, w_016_2604, w_016_2605, w_016_2606, w_016_2607, w_016_2608, w_016_2609, w_016_2610, w_016_2611, w_016_2613, w_016_2615, w_016_2616, w_016_2617, w_016_2618, w_016_2620, w_016_2621, w_016_2622, w_016_2623, w_016_2624, w_016_2625, w_016_2626, w_016_2629, w_016_2630, w_016_2631, w_016_2632, w_016_2633, w_016_2634, w_016_2635, w_016_2636, w_016_2638, w_016_2639, w_016_2641, w_016_2642, w_016_2644, w_016_2645, w_016_2646, w_016_2647, w_016_2649, w_016_2650, w_016_2652, w_016_2653, w_016_2654, w_016_2656, w_016_2657, w_016_2658, w_016_2659, w_016_2660, w_016_2661, w_016_2662, w_016_2663, w_016_2664, w_016_2666, w_016_2668, w_016_2671, w_016_2672, w_016_2673, w_016_2674, w_016_2676, w_016_2677, w_016_2678, w_016_2680, w_016_2681, w_016_2682, w_016_2683, w_016_2684, w_016_2686, w_016_2687, w_016_2688, w_016_2689, w_016_2690, w_016_2692, w_016_2693, w_016_2694, w_016_2697, w_016_2698, w_016_2699, w_016_2700, w_016_2701, w_016_2704, w_016_2705, w_016_2706, w_016_2707, w_016_2710, w_016_2712, w_016_2713, w_016_2716, w_016_2717, w_016_2719, w_016_2720, w_016_2721, w_016_2722, w_016_2723, w_016_2726, w_016_2727, w_016_2728, w_016_2729, w_016_2730, w_016_2731, w_016_2732, w_016_2734, w_016_2735, w_016_2736, w_016_2737, w_016_2738, w_016_2741, w_016_2742, w_016_2743, w_016_2744, w_016_2745, w_016_2746, w_016_2747, w_016_2748, w_016_2749, w_016_2750, w_016_2753, w_016_2754, w_016_2755, w_016_2757, w_016_2759, w_016_2760, w_016_2761, w_016_2762, w_016_2763, w_016_2764, w_016_2765, w_016_2766, w_016_2767, w_016_2769, w_016_2770, w_016_2771, w_016_2772, w_016_2773, w_016_2774, w_016_2775, w_016_2776, w_016_2777, w_016_2778, w_016_2779, w_016_2780, w_016_2781, w_016_2782, w_016_2783, w_016_2784, w_016_2786, w_016_2787, w_016_2788, w_016_2789, w_016_2790, w_016_2791, w_016_2792, w_016_2793, w_016_2795, w_016_2796, w_016_2799, w_016_2800, w_016_2802, w_016_2803, w_016_2804, w_016_2805, w_016_2807, w_016_2808, w_016_2809, w_016_2810, w_016_2811, w_016_2812, w_016_2813, w_016_2814, w_016_2815, w_016_2816, w_016_2817, w_016_2818, w_016_2820, w_016_2821, w_016_2822, w_016_2824, w_016_2825, w_016_2828, w_016_2829, w_016_2830, w_016_2831, w_016_2832, w_016_2833, w_016_2834, w_016_2835, w_016_2836, w_016_2837, w_016_2838, w_016_2843, w_016_2844, w_016_2845, w_016_2847, w_016_2848, w_016_2849, w_016_2850, w_016_2851, w_016_2852, w_016_2853, w_016_2855, w_016_2856, w_016_2857, w_016_2858, w_016_2859, w_016_2860, w_016_2861, w_016_2862, w_016_2863, w_016_2864, w_016_2865, w_016_2866, w_016_2867, w_016_2868, w_016_2869, w_016_2871, w_016_2873, w_016_2875, w_016_2876, w_016_2878, w_016_2879, w_016_2881, w_016_2882, w_016_2883, w_016_2884, w_016_2886, w_016_2887, w_016_2889, w_016_2890, w_016_2891, w_016_2892, w_016_2893, w_016_2894, w_016_2895, w_016_2896, w_016_2897, w_016_2898, w_016_2900, w_016_2901, w_016_2902, w_016_2903, w_016_2907, w_016_2909, w_016_2911, w_016_2912, w_016_2914, w_016_2915, w_016_2916, w_016_2917, w_016_2918, w_016_2919, w_016_2920, w_016_2921, w_016_2922, w_016_2926, w_016_2927, w_016_2929, w_016_2930, w_016_2931, w_016_2932, w_016_2933, w_016_2934, w_016_2936, w_016_2938, w_016_2939, w_016_2941, w_016_2942, w_016_2944, w_016_2945, w_016_2946, w_016_2947, w_016_2948, w_016_2949, w_016_2950, w_016_2951, w_016_2952, w_016_2953, w_016_2955, w_016_2956, w_016_2958, w_016_2959, w_016_2960, w_016_2961, w_016_2962, w_016_2965, w_016_2967, w_016_2968, w_016_2970, w_016_2972, w_016_2975, w_016_2976, w_016_2978, w_016_2979, w_016_2980, w_016_2981, w_016_2982, w_016_2984, w_016_2986, w_016_2987, w_016_2988, w_016_2990, w_016_2991, w_016_2992, w_016_2994, w_016_2995, w_016_2996, w_016_2998, w_016_3000, w_016_3002, w_016_3004, w_016_3005, w_016_3006, w_016_3007, w_016_3009, w_016_3010, w_016_3011, w_016_3014, w_016_3017, w_016_3018, w_016_3020, w_016_3021, w_016_3022, w_016_3024, w_016_3025, w_016_3027, w_016_3029, w_016_3030, w_016_3031, w_016_3032, w_016_3033, w_016_3034, w_016_3035, w_016_3036, w_016_3037, w_016_3038, w_016_3040, w_016_3041, w_016_3042, w_016_3044, w_016_3045, w_016_3046, w_016_3047, w_016_3050, w_016_3052, w_016_3054, w_016_3055, w_016_3056, w_016_3057, w_016_3060, w_016_3061, w_016_3064, w_016_3066, w_016_3069, w_016_3071, w_016_3072, w_016_3073, w_016_3074, w_016_3075, w_016_3076, w_016_3077, w_016_3079, w_016_3081, w_016_3082, w_016_3083, w_016_3084, w_016_3085, w_016_3086, w_016_3087, w_016_3088, w_016_3090, w_016_3091, w_016_3092, w_016_3094, w_016_3095, w_016_3096, w_016_3098, w_016_3099, w_016_3100, w_016_3101, w_016_3102, w_016_3104, w_016_3105, w_016_3106, w_016_3107, w_016_3110, w_016_3111, w_016_3112, w_016_3113, w_016_3114, w_016_3115, w_016_3116, w_016_3118, w_016_3119, w_016_3121, w_016_3122, w_016_3124, w_016_3125, w_016_3126, w_016_3127, w_016_3128, w_016_3129, w_016_3130, w_016_3131, w_016_3132, w_016_3133, w_016_3134, w_016_3135, w_016_3138, w_016_3139, w_016_3140, w_016_3141, w_016_3142, w_016_3144, w_016_3146, w_016_3147, w_016_3148, w_016_3149, w_016_3150, w_016_3151, w_016_3152, w_016_3153, w_016_3155, w_016_3156, w_016_3157, w_016_3158, w_016_3160, w_016_3161, w_016_3162, w_016_3165, w_016_3167, w_016_3169, w_016_3170, w_016_3171, w_016_3172, w_016_3175, w_016_3176, w_016_3177, w_016_3179, w_016_3181, w_016_3184, w_016_3185, w_016_3186, w_016_3187, w_016_3188, w_016_3189, w_016_3191, w_016_3193, w_016_3194, w_016_3197, w_016_3199, w_016_3200, w_016_3202, w_016_3204, w_016_3205, w_016_3206, w_016_3207, w_016_3209, w_016_3210, w_016_3211, w_016_3212, w_016_3213, w_016_3215, w_016_3216, w_016_3217, w_016_3218, w_016_3219, w_016_3221, w_016_3223, w_016_3225, w_016_3226, w_016_3227, w_016_3228, w_016_3229, w_016_3230, w_016_3231, w_016_3233, w_016_3236, w_016_3237, w_016_3238, w_016_3240, w_016_3241, w_016_3242, w_016_3244, w_016_3245, w_016_3246, w_016_3247, w_016_3248, w_016_3250, w_016_3253, w_016_3255, w_016_3259, w_016_3260, w_016_3261, w_016_3262, w_016_3263, w_016_3264, w_016_3265, w_016_3266, w_016_3267, w_016_3268, w_016_3269, w_016_3270, w_016_3272, w_016_3273, w_016_3274, w_016_3275, w_016_3276, w_016_3277, w_016_3279, w_016_3283, w_016_3285, w_016_3286, w_016_3288, w_016_3289, w_016_3290, w_016_3292, w_016_3293, w_016_3294, w_016_3297, w_016_3299, w_016_3301, w_016_3302, w_016_3303, w_016_3304, w_016_3305, w_016_3306, w_016_3307, w_016_3308, w_016_3309, w_016_3310, w_016_3311, w_016_3312, w_016_3313, w_016_3317, w_016_3318, w_016_3319, w_016_3320, w_016_3321, w_016_3322, w_016_3323, w_016_3325, w_016_3326, w_016_3327, w_016_3328, w_016_3329, w_016_3330, w_016_3333, w_016_3334, w_016_3335, w_016_3336, w_016_3338, w_016_3339, w_016_3341, w_016_3342, w_016_3343, w_016_3345, w_016_3346, w_016_3347, w_016_3349, w_016_3351, w_016_3352, w_016_3353, w_016_3356, w_016_3357, w_016_3358, w_016_3359, w_016_3361, w_016_3362, w_016_3364, w_016_3365, w_016_3367, w_016_3368, w_016_3369, w_016_3371, w_016_3372, w_016_3373, w_016_3375, w_016_3376, w_016_3377, w_016_3381, w_016_3384, w_016_3385, w_016_3386, w_016_3387, w_016_3388, w_016_3390, w_016_3391, w_016_3392, w_016_3393, w_016_3395, w_016_3396, w_016_3397, w_016_3398, w_016_3399, w_016_3401, w_016_3403, w_016_3404, w_016_3406, w_016_3407, w_016_3408, w_016_3409, w_016_3411, w_016_3415, w_016_3416, w_016_3417, w_016_3418, w_016_3419, w_016_3421, w_016_3422, w_016_3423, w_016_3424, w_016_3425, w_016_3426, w_016_3427, w_016_3428, w_016_3429, w_016_3430, w_016_3434, w_016_3435, w_016_3436, w_016_3437, w_016_3438, w_016_3440, w_016_3441, w_016_3442, w_016_3443, w_016_3444, w_016_3445, w_016_3446, w_016_3447, w_016_3448, w_016_3449, w_016_3450, w_016_3451, w_016_3452, w_016_3453, w_016_3456, w_016_3457, w_016_3461, w_016_3462, w_016_3463, w_016_3466, w_016_3467, w_016_3468, w_016_3470, w_016_3471, w_016_3472, w_016_3473, w_016_3474, w_016_3475, w_016_3477, w_016_3478, w_016_3480, w_016_3482, w_016_3483, w_016_3485, w_016_3486, w_016_3487, w_016_3488, w_016_3489, w_016_3490, w_016_3491, w_016_3492, w_016_3493, w_016_3494, w_016_3495, w_016_3496;
  wire w_017_000, w_017_001, w_017_002, w_017_003, w_017_004, w_017_005, w_017_006, w_017_007, w_017_008, w_017_009, w_017_010, w_017_011, w_017_012, w_017_013, w_017_014, w_017_015, w_017_016, w_017_017, w_017_018, w_017_019, w_017_020, w_017_021, w_017_022, w_017_023, w_017_024, w_017_025, w_017_026, w_017_027, w_017_028, w_017_029, w_017_030, w_017_031, w_017_032, w_017_033, w_017_034, w_017_035, w_017_036, w_017_037, w_017_038, w_017_039, w_017_040, w_017_041, w_017_042, w_017_043, w_017_044, w_017_045, w_017_046, w_017_047, w_017_048, w_017_049, w_017_050, w_017_051, w_017_052, w_017_053, w_017_054, w_017_055, w_017_056, w_017_057, w_017_058, w_017_059, w_017_060, w_017_062, w_017_063, w_017_064, w_017_065, w_017_066, w_017_067, w_017_068, w_017_069, w_017_070, w_017_071, w_017_072, w_017_073, w_017_074, w_017_075, w_017_076, w_017_077, w_017_078, w_017_079, w_017_080, w_017_081, w_017_082, w_017_083, w_017_084, w_017_085, w_017_086, w_017_087, w_017_088, w_017_089, w_017_090, w_017_091, w_017_092, w_017_093, w_017_094, w_017_095, w_017_096, w_017_097, w_017_098, w_017_099, w_017_100, w_017_101, w_017_102, w_017_104, w_017_105, w_017_106, w_017_107, w_017_108, w_017_109, w_017_110, w_017_111, w_017_112, w_017_113, w_017_114, w_017_115, w_017_116, w_017_117, w_017_118, w_017_119, w_017_120, w_017_121, w_017_122, w_017_123, w_017_124, w_017_125, w_017_126, w_017_127, w_017_128, w_017_129, w_017_130, w_017_131, w_017_132, w_017_133, w_017_134, w_017_135, w_017_136, w_017_137, w_017_138, w_017_139, w_017_140, w_017_141, w_017_142, w_017_143, w_017_144, w_017_145, w_017_146, w_017_147, w_017_148, w_017_149, w_017_150, w_017_151, w_017_152, w_017_153, w_017_154, w_017_155, w_017_156, w_017_157, w_017_158, w_017_159, w_017_160, w_017_161, w_017_162, w_017_163, w_017_164, w_017_165, w_017_166, w_017_167, w_017_168, w_017_169, w_017_170, w_017_171, w_017_172, w_017_173, w_017_174, w_017_175, w_017_176, w_017_177, w_017_178, w_017_179, w_017_180, w_017_181, w_017_182, w_017_183, w_017_184, w_017_185, w_017_186, w_017_187, w_017_188, w_017_189, w_017_190, w_017_191, w_017_192, w_017_193, w_017_194, w_017_195, w_017_196, w_017_198, w_017_199, w_017_200, w_017_201, w_017_202, w_017_203, w_017_204, w_017_205, w_017_206, w_017_207, w_017_208, w_017_209, w_017_210, w_017_211, w_017_212, w_017_213, w_017_214, w_017_215, w_017_216, w_017_217, w_017_218, w_017_219, w_017_220, w_017_221, w_017_222, w_017_223, w_017_224, w_017_225, w_017_226, w_017_227, w_017_228, w_017_229, w_017_230, w_017_231, w_017_232, w_017_233, w_017_234, w_017_235, w_017_236, w_017_237, w_017_238, w_017_239, w_017_240, w_017_241, w_017_242, w_017_243, w_017_244, w_017_245, w_017_246, w_017_247, w_017_248, w_017_249, w_017_250, w_017_251, w_017_252, w_017_253, w_017_254, w_017_255, w_017_256, w_017_257, w_017_258, w_017_259, w_017_260, w_017_261, w_017_262, w_017_263, w_017_264, w_017_265, w_017_266, w_017_267, w_017_268, w_017_269, w_017_270, w_017_271, w_017_272, w_017_273, w_017_274, w_017_275, w_017_276, w_017_277, w_017_278, w_017_279, w_017_280, w_017_281, w_017_282, w_017_283, w_017_284, w_017_285, w_017_286, w_017_287, w_017_288, w_017_289, w_017_290, w_017_291, w_017_292, w_017_293, w_017_294, w_017_296, w_017_297, w_017_298, w_017_299, w_017_300, w_017_301, w_017_302, w_017_303, w_017_304, w_017_305, w_017_306, w_017_307, w_017_308, w_017_309, w_017_311, w_017_312, w_017_313, w_017_314, w_017_315, w_017_316, w_017_317, w_017_318, w_017_319, w_017_320, w_017_321, w_017_322, w_017_323, w_017_324, w_017_325, w_017_326, w_017_327, w_017_328, w_017_329, w_017_331, w_017_332, w_017_333, w_017_334, w_017_336, w_017_337, w_017_338, w_017_339, w_017_340, w_017_341, w_017_342, w_017_343, w_017_344, w_017_345, w_017_346, w_017_347, w_017_348, w_017_349, w_017_350, w_017_351, w_017_352, w_017_353, w_017_354, w_017_355, w_017_356, w_017_358, w_017_360, w_017_361, w_017_362, w_017_363, w_017_364, w_017_365, w_017_366, w_017_367, w_017_368, w_017_369, w_017_370, w_017_371, w_017_372, w_017_373, w_017_374, w_017_375, w_017_376, w_017_377, w_017_378, w_017_379, w_017_380, w_017_381, w_017_382, w_017_383, w_017_384, w_017_385, w_017_386, w_017_387, w_017_388, w_017_389, w_017_390, w_017_391, w_017_392, w_017_393, w_017_395, w_017_396, w_017_397, w_017_398, w_017_399, w_017_400, w_017_401, w_017_402, w_017_403, w_017_404, w_017_405, w_017_406, w_017_407, w_017_408, w_017_409, w_017_410, w_017_411, w_017_412, w_017_413, w_017_414, w_017_415, w_017_416, w_017_417, w_017_418, w_017_419, w_017_420, w_017_421, w_017_422, w_017_423, w_017_424, w_017_425, w_017_426, w_017_427, w_017_428, w_017_429, w_017_430, w_017_431, w_017_432, w_017_434, w_017_435, w_017_436, w_017_437, w_017_438, w_017_439, w_017_440, w_017_441, w_017_442, w_017_443, w_017_444, w_017_445, w_017_446, w_017_447, w_017_448, w_017_449, w_017_450, w_017_451, w_017_452, w_017_453, w_017_454, w_017_455, w_017_456, w_017_457, w_017_458, w_017_459, w_017_460, w_017_461, w_017_462, w_017_463, w_017_464, w_017_465, w_017_466, w_017_467, w_017_468, w_017_469, w_017_470, w_017_471, w_017_472, w_017_474, w_017_475, w_017_476, w_017_477, w_017_479, w_017_480, w_017_481, w_017_482, w_017_483, w_017_485, w_017_486, w_017_487, w_017_488, w_017_489, w_017_490, w_017_491, w_017_492, w_017_493, w_017_494, w_017_495, w_017_496, w_017_497, w_017_498, w_017_499, w_017_501, w_017_502, w_017_503, w_017_504, w_017_506, w_017_507, w_017_508, w_017_509, w_017_510, w_017_512, w_017_514, w_017_515, w_017_516, w_017_517, w_017_518, w_017_519, w_017_520, w_017_521, w_017_522, w_017_523, w_017_524, w_017_525, w_017_527, w_017_528, w_017_529, w_017_530, w_017_531, w_017_532, w_017_533, w_017_534, w_017_535, w_017_536, w_017_537, w_017_538, w_017_539, w_017_540, w_017_541, w_017_542, w_017_543, w_017_544, w_017_545, w_017_546, w_017_547, w_017_548, w_017_549, w_017_551, w_017_552, w_017_553, w_017_554, w_017_555, w_017_556, w_017_557, w_017_558, w_017_559, w_017_560, w_017_562, w_017_563, w_017_564, w_017_565, w_017_566, w_017_567, w_017_570, w_017_571, w_017_572, w_017_573, w_017_574, w_017_575, w_017_576, w_017_577, w_017_578, w_017_579, w_017_580, w_017_581, w_017_582, w_017_583, w_017_584, w_017_585, w_017_586, w_017_587, w_017_588, w_017_589, w_017_590, w_017_591, w_017_592, w_017_593, w_017_594, w_017_595, w_017_596, w_017_597, w_017_598, w_017_599, w_017_600, w_017_601, w_017_602, w_017_603, w_017_604, w_017_605, w_017_606, w_017_607, w_017_608, w_017_609, w_017_610, w_017_611, w_017_613, w_017_614, w_017_615, w_017_616, w_017_617, w_017_618, w_017_619, w_017_620, w_017_621, w_017_622, w_017_623, w_017_624, w_017_625, w_017_627, w_017_628, w_017_629, w_017_630, w_017_631, w_017_632, w_017_633, w_017_634, w_017_635, w_017_636, w_017_637, w_017_638, w_017_639, w_017_641, w_017_643, w_017_644, w_017_645, w_017_646, w_017_647, w_017_649, w_017_650, w_017_651, w_017_652, w_017_653, w_017_654, w_017_656, w_017_657, w_017_658, w_017_659, w_017_660, w_017_661, w_017_662, w_017_663, w_017_664, w_017_665, w_017_666, w_017_668, w_017_669, w_017_670, w_017_671, w_017_672, w_017_673, w_017_674, w_017_675, w_017_676, w_017_677, w_017_678, w_017_679, w_017_680, w_017_681, w_017_682, w_017_683, w_017_684, w_017_685, w_017_686, w_017_688, w_017_689, w_017_690, w_017_691, w_017_692, w_017_693, w_017_694, w_017_695, w_017_696, w_017_697, w_017_698, w_017_699, w_017_700, w_017_701, w_017_702, w_017_703, w_017_704, w_017_705, w_017_706, w_017_707, w_017_708, w_017_709, w_017_710, w_017_711, w_017_713, w_017_714, w_017_715, w_017_716, w_017_717, w_017_718, w_017_719, w_017_720, w_017_721, w_017_722, w_017_723, w_017_724, w_017_725, w_017_726, w_017_727, w_017_728, w_017_729, w_017_731, w_017_732, w_017_733, w_017_734, w_017_735, w_017_736, w_017_737, w_017_738, w_017_739, w_017_741, w_017_742, w_017_743, w_017_744, w_017_746, w_017_747, w_017_748, w_017_749, w_017_750, w_017_751, w_017_753, w_017_755, w_017_756, w_017_757, w_017_758, w_017_760, w_017_761, w_017_762, w_017_763, w_017_764, w_017_765, w_017_766, w_017_767, w_017_768, w_017_769, w_017_770, w_017_771, w_017_772, w_017_773, w_017_774, w_017_775, w_017_776, w_017_778, w_017_780, w_017_781, w_017_782, w_017_783, w_017_784, w_017_785, w_017_786, w_017_787, w_017_788, w_017_789, w_017_791, w_017_792, w_017_793, w_017_794, w_017_795, w_017_796, w_017_797, w_017_798, w_017_800, w_017_801, w_017_802, w_017_803, w_017_804, w_017_805, w_017_806, w_017_807, w_017_808, w_017_809, w_017_810, w_017_811, w_017_813, w_017_814, w_017_815, w_017_816, w_017_817, w_017_818, w_017_819, w_017_820, w_017_821, w_017_822, w_017_823, w_017_824, w_017_825, w_017_826, w_017_827, w_017_828, w_017_829, w_017_830, w_017_831, w_017_832, w_017_833, w_017_834, w_017_835, w_017_836, w_017_837, w_017_838, w_017_839, w_017_841, w_017_842, w_017_843, w_017_844, w_017_845, w_017_846, w_017_847, w_017_848, w_017_849, w_017_850, w_017_851, w_017_852, w_017_853, w_017_854, w_017_855, w_017_856, w_017_857, w_017_859, w_017_860, w_017_861, w_017_862, w_017_863, w_017_864, w_017_865, w_017_866, w_017_867, w_017_868, w_017_869, w_017_870, w_017_871, w_017_872, w_017_873, w_017_874, w_017_875, w_017_876, w_017_877, w_017_879, w_017_880, w_017_881, w_017_882, w_017_883, w_017_884, w_017_885, w_017_886, w_017_887, w_017_888, w_017_889, w_017_891, w_017_892, w_017_893, w_017_894, w_017_895, w_017_896, w_017_897, w_017_898, w_017_899, w_017_900, w_017_901, w_017_902, w_017_903, w_017_904, w_017_905, w_017_906, w_017_907, w_017_908, w_017_909, w_017_910, w_017_911, w_017_912, w_017_913, w_017_914, w_017_915, w_017_916, w_017_917, w_017_918, w_017_919, w_017_920, w_017_921, w_017_922, w_017_923, w_017_924, w_017_925, w_017_926, w_017_927, w_017_928, w_017_929, w_017_930, w_017_931, w_017_932, w_017_933, w_017_934, w_017_935, w_017_936, w_017_937, w_017_938, w_017_939, w_017_940, w_017_941, w_017_942, w_017_943, w_017_944, w_017_945, w_017_946, w_017_948, w_017_949, w_017_950, w_017_952, w_017_953, w_017_954, w_017_955, w_017_956, w_017_958, w_017_959, w_017_960, w_017_961, w_017_962, w_017_963, w_017_964, w_017_965, w_017_966, w_017_967, w_017_969, w_017_970, w_017_971, w_017_972, w_017_973, w_017_974, w_017_975, w_017_976, w_017_977, w_017_978, w_017_979, w_017_980, w_017_981, w_017_982, w_017_983, w_017_984, w_017_985, w_017_986, w_017_987, w_017_988, w_017_989, w_017_990, w_017_991, w_017_992, w_017_993, w_017_994, w_017_996, w_017_997, w_017_998, w_017_999, w_017_1000, w_017_1002, w_017_1003, w_017_1004, w_017_1005, w_017_1007, w_017_1008, w_017_1009, w_017_1010, w_017_1011, w_017_1012, w_017_1013, w_017_1014, w_017_1015, w_017_1016, w_017_1017, w_017_1018, w_017_1019, w_017_1020, w_017_1021, w_017_1022, w_017_1023, w_017_1024, w_017_1025, w_017_1026, w_017_1027, w_017_1028, w_017_1029, w_017_1030, w_017_1031, w_017_1032, w_017_1033, w_017_1034, w_017_1035, w_017_1036, w_017_1037, w_017_1038, w_017_1039, w_017_1040, w_017_1042, w_017_1043, w_017_1044, w_017_1045, w_017_1046, w_017_1047, w_017_1048, w_017_1049, w_017_1050, w_017_1051, w_017_1052, w_017_1053, w_017_1054, w_017_1055, w_017_1057, w_017_1058, w_017_1059, w_017_1060, w_017_1061, w_017_1062, w_017_1063, w_017_1064, w_017_1065, w_017_1066, w_017_1067, w_017_1068, w_017_1069, w_017_1070, w_017_1071, w_017_1072, w_017_1073, w_017_1075, w_017_1076, w_017_1077, w_017_1078, w_017_1079, w_017_1080, w_017_1081, w_017_1082, w_017_1083, w_017_1084, w_017_1085, w_017_1086, w_017_1087, w_017_1088, w_017_1089, w_017_1092, w_017_1093, w_017_1096, w_017_1097, w_017_1098, w_017_1099, w_017_1100, w_017_1101, w_017_1102, w_017_1103, w_017_1104, w_017_1105, w_017_1106, w_017_1107, w_017_1108, w_017_1109, w_017_1110, w_017_1111, w_017_1112, w_017_1113, w_017_1114, w_017_1115, w_017_1116, w_017_1117, w_017_1118, w_017_1119, w_017_1120, w_017_1121, w_017_1122, w_017_1123, w_017_1124, w_017_1125, w_017_1127, w_017_1128, w_017_1129, w_017_1130, w_017_1131, w_017_1132, w_017_1135, w_017_1136, w_017_1137, w_017_1138, w_017_1140, w_017_1141, w_017_1142, w_017_1144, w_017_1145, w_017_1146, w_017_1147, w_017_1148, w_017_1149, w_017_1150, w_017_1151, w_017_1152, w_017_1154, w_017_1155, w_017_1156, w_017_1157, w_017_1158, w_017_1159, w_017_1160, w_017_1161, w_017_1162, w_017_1163, w_017_1164, w_017_1165, w_017_1166, w_017_1167, w_017_1168, w_017_1169, w_017_1170, w_017_1171, w_017_1172, w_017_1173, w_017_1174, w_017_1175, w_017_1176, w_017_1177, w_017_1178, w_017_1179, w_017_1180, w_017_1181, w_017_1182, w_017_1183, w_017_1185, w_017_1186, w_017_1187, w_017_1188, w_017_1189, w_017_1190, w_017_1192, w_017_1193, w_017_1194, w_017_1195, w_017_1196, w_017_1197, w_017_1198, w_017_1199, w_017_1200, w_017_1201, w_017_1202, w_017_1203, w_017_1204, w_017_1207, w_017_1208, w_017_1209, w_017_1210, w_017_1211, w_017_1212, w_017_1213, w_017_1214, w_017_1215, w_017_1216, w_017_1217, w_017_1218, w_017_1219, w_017_1220, w_017_1221, w_017_1222, w_017_1223, w_017_1224, w_017_1225, w_017_1226, w_017_1227, w_017_1228, w_017_1229, w_017_1231, w_017_1232, w_017_1233, w_017_1234, w_017_1235, w_017_1236, w_017_1237, w_017_1238, w_017_1239, w_017_1240, w_017_1241, w_017_1242, w_017_1243, w_017_1244, w_017_1245, w_017_1246, w_017_1247, w_017_1248, w_017_1249, w_017_1250, w_017_1251, w_017_1252, w_017_1253, w_017_1254, w_017_1255, w_017_1256, w_017_1257, w_017_1258, w_017_1259, w_017_1260, w_017_1261, w_017_1262, w_017_1263, w_017_1264, w_017_1265, w_017_1266, w_017_1267, w_017_1268, w_017_1269, w_017_1270, w_017_1271, w_017_1273, w_017_1274, w_017_1276, w_017_1277, w_017_1278, w_017_1279, w_017_1280, w_017_1282, w_017_1283, w_017_1284, w_017_1285, w_017_1286, w_017_1287, w_017_1288, w_017_1289, w_017_1290, w_017_1294, w_017_1295, w_017_1296, w_017_1297, w_017_1298, w_017_1299, w_017_1300, w_017_1301, w_017_1302, w_017_1303, w_017_1305, w_017_1306, w_017_1307, w_017_1308, w_017_1309, w_017_1311, w_017_1312, w_017_1313, w_017_1314, w_017_1315, w_017_1316, w_017_1317, w_017_1318, w_017_1319, w_017_1320, w_017_1321, w_017_1322, w_017_1323, w_017_1324, w_017_1325, w_017_1326, w_017_1327, w_017_1329, w_017_1330, w_017_1331, w_017_1332, w_017_1333, w_017_1334, w_017_1335, w_017_1336, w_017_1337, w_017_1338, w_017_1339, w_017_1340, w_017_1341, w_017_1342, w_017_1343, w_017_1344, w_017_1345, w_017_1346, w_017_1347, w_017_1348, w_017_1349, w_017_1350, w_017_1351, w_017_1352, w_017_1353, w_017_1354, w_017_1355, w_017_1356, w_017_1357, w_017_1358, w_017_1360, w_017_1361, w_017_1362, w_017_1363, w_017_1364, w_017_1365, w_017_1366, w_017_1367, w_017_1368, w_017_1369, w_017_1370, w_017_1371, w_017_1372, w_017_1373, w_017_1374, w_017_1375, w_017_1376, w_017_1377, w_017_1379, w_017_1380, w_017_1382, w_017_1383, w_017_1384, w_017_1385, w_017_1387, w_017_1388, w_017_1389, w_017_1390, w_017_1391, w_017_1392, w_017_1393, w_017_1394, w_017_1395, w_017_1396, w_017_1397, w_017_1398, w_017_1399, w_017_1400, w_017_1401, w_017_1402, w_017_1403, w_017_1404, w_017_1405, w_017_1406, w_017_1407, w_017_1408, w_017_1410, w_017_1411, w_017_1412, w_017_1413, w_017_1414, w_017_1415, w_017_1416, w_017_1417, w_017_1418, w_017_1419, w_017_1420, w_017_1421, w_017_1422, w_017_1423, w_017_1424, w_017_1425, w_017_1426, w_017_1427, w_017_1428, w_017_1429, w_017_1431, w_017_1432, w_017_1433, w_017_1434, w_017_1435, w_017_1436, w_017_1437, w_017_1438, w_017_1439, w_017_1440, w_017_1441, w_017_1442, w_017_1443, w_017_1444, w_017_1445, w_017_1446, w_017_1447, w_017_1448, w_017_1449, w_017_1450, w_017_1452, w_017_1454, w_017_1455, w_017_1456, w_017_1457, w_017_1458, w_017_1459, w_017_1460, w_017_1462, w_017_1463, w_017_1464, w_017_1465, w_017_1466, w_017_1467, w_017_1469, w_017_1470, w_017_1471, w_017_1472, w_017_1473, w_017_1474, w_017_1475, w_017_1476, w_017_1477, w_017_1478, w_017_1479, w_017_1480, w_017_1481, w_017_1482, w_017_1483, w_017_1484, w_017_1485, w_017_1486, w_017_1487, w_017_1488, w_017_1490, w_017_1491, w_017_1492, w_017_1493, w_017_1494, w_017_1495, w_017_1497, w_017_1498, w_017_1499, w_017_1500, w_017_1501, w_017_1502, w_017_1503, w_017_1504, w_017_1505, w_017_1506, w_017_1507, w_017_1508, w_017_1510, w_017_1511, w_017_1512, w_017_1513, w_017_1514, w_017_1515, w_017_1516, w_017_1517, w_017_1518, w_017_1519, w_017_1520, w_017_1521, w_017_1522, w_017_1523, w_017_1525, w_017_1526, w_017_1527, w_017_1528, w_017_1529, w_017_1530, w_017_1531, w_017_1532, w_017_1533, w_017_1534, w_017_1535, w_017_1536, w_017_1537, w_017_1538, w_017_1539, w_017_1540, w_017_1541, w_017_1542, w_017_1543, w_017_1544, w_017_1545, w_017_1546, w_017_1547, w_017_1548, w_017_1549, w_017_1550, w_017_1551, w_017_1552, w_017_1553, w_017_1554, w_017_1555, w_017_1557, w_017_1558, w_017_1559, w_017_1560, w_017_1561, w_017_1562, w_017_1563, w_017_1564, w_017_1565, w_017_1566, w_017_1567, w_017_1568, w_017_1570, w_017_1571, w_017_1573, w_017_1574, w_017_1575, w_017_1576, w_017_1577, w_017_1578, w_017_1579, w_017_1580, w_017_1581, w_017_1582, w_017_1583, w_017_1584, w_017_1585, w_017_1586, w_017_1587, w_017_1588, w_017_1589, w_017_1590, w_017_1591, w_017_1592, w_017_1593, w_017_1594, w_017_1595, w_017_1596, w_017_1597, w_017_1598, w_017_1599, w_017_1600, w_017_1601, w_017_1602, w_017_1603, w_017_1604, w_017_1605, w_017_1606, w_017_1607, w_017_1608, w_017_1609, w_017_1610, w_017_1611, w_017_1612, w_017_1613, w_017_1614, w_017_1615, w_017_1616, w_017_1617, w_017_1618, w_017_1619, w_017_1620, w_017_1621, w_017_1622, w_017_1623, w_017_1624, w_017_1625, w_017_1626, w_017_1627, w_017_1629, w_017_1630, w_017_1631, w_017_1632, w_017_1633, w_017_1635, w_017_1636, w_017_1637, w_017_1638, w_017_1639, w_017_1640, w_017_1641, w_017_1642, w_017_1643, w_017_1644, w_017_1645, w_017_1646, w_017_1647, w_017_1648, w_017_1649, w_017_1650, w_017_1651, w_017_1652, w_017_1653, w_017_1654, w_017_1655, w_017_1656, w_017_1657, w_017_1659, w_017_1660, w_017_1661, w_017_1662, w_017_1664, w_017_1665, w_017_1666, w_017_1667, w_017_1668, w_017_1669, w_017_1670, w_017_1671, w_017_1672, w_017_1673, w_017_1674, w_017_1675, w_017_1676, w_017_1677, w_017_1679, w_017_1680, w_017_1681, w_017_1682, w_017_1683, w_017_1684, w_017_1685, w_017_1686, w_017_1687, w_017_1689, w_017_1690, w_017_1691, w_017_1692, w_017_1693, w_017_1694, w_017_1695, w_017_1696, w_017_1697, w_017_1698, w_017_1699, w_017_1700, w_017_1701, w_017_1702, w_017_1703, w_017_1705, w_017_1706, w_017_1707, w_017_1709, w_017_1710, w_017_1711, w_017_1712, w_017_1713, w_017_1714, w_017_1715, w_017_1716, w_017_1718, w_017_1719, w_017_1720, w_017_1721, w_017_1722, w_017_1723, w_017_1725, w_017_1726, w_017_1727, w_017_1728, w_017_1729, w_017_1730, w_017_1731, w_017_1732, w_017_1733, w_017_1734, w_017_1735, w_017_1736, w_017_1737, w_017_1738, w_017_1739, w_017_1740, w_017_1741, w_017_1742, w_017_1743, w_017_1744, w_017_1745, w_017_1746, w_017_1747, w_017_1748, w_017_1749, w_017_1750, w_017_1751, w_017_1752, w_017_1753, w_017_1754, w_017_1755, w_017_1756, w_017_1757, w_017_1758, w_017_1759, w_017_1760, w_017_1761, w_017_1762, w_017_1763, w_017_1764, w_017_1765, w_017_1766, w_017_1767, w_017_1768, w_017_1769, w_017_1770, w_017_1771, w_017_1772, w_017_1773, w_017_1774, w_017_1775, w_017_1777, w_017_1778, w_017_1779, w_017_1780, w_017_1781, w_017_1782, w_017_1783, w_017_1785, w_017_1786, w_017_1787, w_017_1788, w_017_1789, w_017_1790, w_017_1791, w_017_1792, w_017_1794, w_017_1795, w_017_1800, w_017_1801, w_017_1802, w_017_1803, w_017_1804, w_017_1805, w_017_1806, w_017_1807, w_017_1808, w_017_1809, w_017_1810, w_017_1811, w_017_1812, w_017_1813, w_017_1814, w_017_1815, w_017_1816, w_017_1817, w_017_1818, w_017_1819, w_017_1820, w_017_1821, w_017_1822, w_017_1823, w_017_1824, w_017_1825, w_017_1826, w_017_1828, w_017_1829, w_017_1830, w_017_1831, w_017_1832, w_017_1833, w_017_1834, w_017_1835, w_017_1836, w_017_1837, w_017_1838, w_017_1839, w_017_1840, w_017_1841, w_017_1843, w_017_1844, w_017_1846, w_017_1847, w_017_1848, w_017_1849, w_017_1850, w_017_1851, w_017_1852, w_017_1853, w_017_1854, w_017_1855, w_017_1856, w_017_1857, w_017_1858, w_017_1859, w_017_1861, w_017_1862, w_017_1864, w_017_1865, w_017_1866, w_017_1867, w_017_1868, w_017_1869, w_017_1870, w_017_1871, w_017_1872, w_017_1874, w_017_1875, w_017_1877, w_017_1878, w_017_1879, w_017_1881, w_017_1882, w_017_1883, w_017_1884, w_017_1885, w_017_1886, w_017_1887, w_017_1888, w_017_1889, w_017_1890, w_017_1891, w_017_1892, w_017_1893, w_017_1894, w_017_1895, w_017_1896, w_017_1897, w_017_1898, w_017_1899, w_017_1900, w_017_1901, w_017_1902, w_017_1903, w_017_1904, w_017_1905, w_017_1907, w_017_1908, w_017_1909, w_017_1910, w_017_1911, w_017_1912, w_017_1913, w_017_1915, w_017_1916, w_017_1917, w_017_1918, w_017_1919, w_017_1920, w_017_1921, w_017_1922, w_017_1923, w_017_1924, w_017_1925, w_017_1926, w_017_1927, w_017_1929, w_017_1930, w_017_1931, w_017_1932, w_017_1933, w_017_1934, w_017_1935, w_017_1936, w_017_1937, w_017_1938, w_017_1939, w_017_1940, w_017_1941, w_017_1942, w_017_1943, w_017_1945, w_017_1946, w_017_1947, w_017_1948, w_017_1949, w_017_1951, w_017_1952, w_017_1954, w_017_1955, w_017_1956, w_017_1957, w_017_1958, w_017_1959, w_017_1960, w_017_1961, w_017_1962, w_017_1963, w_017_1964, w_017_1965, w_017_1966, w_017_1967, w_017_1968, w_017_1969, w_017_1970, w_017_1971, w_017_1972, w_017_1973, w_017_1974, w_017_1975, w_017_1976, w_017_1977, w_017_1978, w_017_1980, w_017_1981, w_017_1982, w_017_1983, w_017_1984, w_017_1985, w_017_1986, w_017_1987, w_017_1988, w_017_1989, w_017_1991, w_017_1992, w_017_1993, w_017_1994, w_017_1995, w_017_1996, w_017_1997, w_017_1998, w_017_1999, w_017_2001, w_017_2002, w_017_2003, w_017_2004, w_017_2005, w_017_2006, w_017_2007, w_017_2008, w_017_2009, w_017_2010, w_017_2011, w_017_2012, w_017_2013, w_017_2014, w_017_2015, w_017_2016, w_017_2017, w_017_2018, w_017_2019, w_017_2020, w_017_2021, w_017_2022, w_017_2023, w_017_2024, w_017_2025, w_017_2026, w_017_2027, w_017_2028, w_017_2029, w_017_2030, w_017_2031, w_017_2032, w_017_2033, w_017_2034, w_017_2035, w_017_2036, w_017_2037, w_017_2038, w_017_2039, w_017_2040, w_017_2041, w_017_2042, w_017_2043, w_017_2044, w_017_2045, w_017_2046, w_017_2047, w_017_2048, w_017_2049, w_017_2050, w_017_2052, w_017_2053, w_017_2054, w_017_2055, w_017_2056, w_017_2057, w_017_2058, w_017_2059, w_017_2060, w_017_2061, w_017_2062, w_017_2063, w_017_2064, w_017_2065, w_017_2067, w_017_2068, w_017_2069, w_017_2070, w_017_2071, w_017_2072, w_017_2073, w_017_2074, w_017_2075, w_017_2076, w_017_2077, w_017_2078, w_017_2079, w_017_2081, w_017_2082, w_017_2084, w_017_2085, w_017_2086, w_017_2087, w_017_2088, w_017_2089, w_017_2090, w_017_2091, w_017_2092, w_017_2093, w_017_2094, w_017_2095, w_017_2096, w_017_2097, w_017_2098, w_017_2099, w_017_2100, w_017_2101, w_017_2102, w_017_2103, w_017_2104, w_017_2105, w_017_2106, w_017_2107, w_017_2108, w_017_2109, w_017_2110, w_017_2111, w_017_2112, w_017_2113, w_017_2114, w_017_2115, w_017_2116, w_017_2117, w_017_2118, w_017_2119, w_017_2120, w_017_2121, w_017_2122, w_017_2124, w_017_2125, w_017_2126, w_017_2127, w_017_2128, w_017_2129, w_017_2130, w_017_2131, w_017_2132, w_017_2133, w_017_2134, w_017_2136, w_017_2137, w_017_2139, w_017_2140, w_017_2141, w_017_2142, w_017_2143, w_017_2144, w_017_2145, w_017_2146, w_017_2147, w_017_2148, w_017_2149, w_017_2150, w_017_2151, w_017_2152, w_017_2153, w_017_2154, w_017_2156, w_017_2157, w_017_2158, w_017_2159, w_017_2160, w_017_2161, w_017_2162, w_017_2163, w_017_2164, w_017_2165, w_017_2166, w_017_2167, w_017_2168, w_017_2169, w_017_2170, w_017_2171, w_017_2172, w_017_2173, w_017_2174, w_017_2175, w_017_2176, w_017_2177, w_017_2178, w_017_2179, w_017_2181, w_017_2182, w_017_2183, w_017_2184, w_017_2185, w_017_2186, w_017_2187, w_017_2188, w_017_2189, w_017_2190, w_017_2191, w_017_2192, w_017_2193, w_017_2194, w_017_2195, w_017_2196, w_017_2197, w_017_2198, w_017_2199, w_017_2200, w_017_2201, w_017_2202, w_017_2203, w_017_2204, w_017_2205, w_017_2206, w_017_2207, w_017_2208, w_017_2209, w_017_2210, w_017_2211, w_017_2212, w_017_2213, w_017_2214, w_017_2215, w_017_2216, w_017_2217, w_017_2218, w_017_2219, w_017_2220, w_017_2221, w_017_2222, w_017_2223, w_017_2224, w_017_2225, w_017_2227, w_017_2228, w_017_2229, w_017_2230, w_017_2231, w_017_2232, w_017_2233, w_017_2234, w_017_2235, w_017_2236, w_017_2237, w_017_2238, w_017_2239, w_017_2240, w_017_2241, w_017_2242, w_017_2243, w_017_2244, w_017_2245, w_017_2246, w_017_2247, w_017_2248, w_017_2249, w_017_2250, w_017_2251, w_017_2252, w_017_2253, w_017_2254, w_017_2255, w_017_2256, w_017_2257, w_017_2258, w_017_2260, w_017_2261, w_017_2262, w_017_2264, w_017_2265, w_017_2266, w_017_2267, w_017_2268, w_017_2269, w_017_2270, w_017_2271, w_017_2272, w_017_2273, w_017_2274, w_017_2275, w_017_2276, w_017_2277, w_017_2278, w_017_2280, w_017_2281, w_017_2282, w_017_2283, w_017_2284, w_017_2285, w_017_2286, w_017_2287, w_017_2288, w_017_2289, w_017_2291, w_017_2292, w_017_2293, w_017_2295, w_017_2296, w_017_2297, w_017_2298, w_017_2299, w_017_2300, w_017_2301, w_017_2302, w_017_2303, w_017_2304, w_017_2306, w_017_2307, w_017_2309, w_017_2310, w_017_2311, w_017_2312, w_017_2313, w_017_2314, w_017_2315, w_017_2317, w_017_2318, w_017_2319, w_017_2321, w_017_2322, w_017_2325, w_017_2326, w_017_2327, w_017_2328, w_017_2329, w_017_2330, w_017_2331, w_017_2332, w_017_2333, w_017_2334, w_017_2335, w_017_2336, w_017_2337, w_017_2338, w_017_2339, w_017_2340, w_017_2341, w_017_2342, w_017_2343, w_017_2344, w_017_2345, w_017_2346, w_017_2348, w_017_2350, w_017_2351, w_017_2352, w_017_2353, w_017_2354, w_017_2356, w_017_2358, w_017_2359, w_017_2360, w_017_2361, w_017_2362;
  wire w_018_000, w_018_001, w_018_002, w_018_003, w_018_004, w_018_005, w_018_006, w_018_007, w_018_008, w_018_009, w_018_010, w_018_011, w_018_012, w_018_013, w_018_014, w_018_015, w_018_016, w_018_017, w_018_018, w_018_019, w_018_020, w_018_021, w_018_022, w_018_023, w_018_024, w_018_025, w_018_026, w_018_027, w_018_028, w_018_029, w_018_030, w_018_031, w_018_032, w_018_033, w_018_034, w_018_035, w_018_036, w_018_037, w_018_038, w_018_039, w_018_040, w_018_041, w_018_042, w_018_043, w_018_044, w_018_045, w_018_046, w_018_047, w_018_048, w_018_049, w_018_050, w_018_051, w_018_052, w_018_053, w_018_054, w_018_055, w_018_056, w_018_057, w_018_058, w_018_059, w_018_060, w_018_061, w_018_062, w_018_063, w_018_064, w_018_065, w_018_066, w_018_067, w_018_068, w_018_069, w_018_070, w_018_071, w_018_072, w_018_073, w_018_074, w_018_075, w_018_076, w_018_077, w_018_078, w_018_079, w_018_080, w_018_081, w_018_082, w_018_083, w_018_084, w_018_085, w_018_086, w_018_087, w_018_088, w_018_089, w_018_090, w_018_091, w_018_092, w_018_093, w_018_094, w_018_095, w_018_096, w_018_097, w_018_098, w_018_099, w_018_100, w_018_101, w_018_102, w_018_103, w_018_104, w_018_105, w_018_106, w_018_107, w_018_108, w_018_109, w_018_110, w_018_111, w_018_112, w_018_113, w_018_114, w_018_115, w_018_116, w_018_117, w_018_118, w_018_119, w_018_120, w_018_121, w_018_122, w_018_123, w_018_124, w_018_125, w_018_126, w_018_127, w_018_128, w_018_129, w_018_130, w_018_131, w_018_132, w_018_133, w_018_134, w_018_135, w_018_136, w_018_137, w_018_138, w_018_139, w_018_140, w_018_141, w_018_142, w_018_143, w_018_144, w_018_145, w_018_146, w_018_147, w_018_148, w_018_149, w_018_150, w_018_151, w_018_152, w_018_153, w_018_154, w_018_155, w_018_156, w_018_157, w_018_158, w_018_159, w_018_160, w_018_161, w_018_162, w_018_163, w_018_164, w_018_165, w_018_166, w_018_167, w_018_168, w_018_169, w_018_170, w_018_171, w_018_172, w_018_173, w_018_174, w_018_175, w_018_176, w_018_177, w_018_178, w_018_179, w_018_180, w_018_181, w_018_182, w_018_183, w_018_184, w_018_185, w_018_186, w_018_187, w_018_188, w_018_189, w_018_190, w_018_191, w_018_192, w_018_193, w_018_194, w_018_195, w_018_196, w_018_197, w_018_198, w_018_199, w_018_200, w_018_201, w_018_202, w_018_203, w_018_204, w_018_205, w_018_206, w_018_207, w_018_208, w_018_209, w_018_210, w_018_211, w_018_212, w_018_213, w_018_214, w_018_215, w_018_216, w_018_217, w_018_218, w_018_219, w_018_220, w_018_221, w_018_222, w_018_223, w_018_224, w_018_225, w_018_226, w_018_227, w_018_228, w_018_229, w_018_230, w_018_231, w_018_232, w_018_233, w_018_234, w_018_235, w_018_236, w_018_237, w_018_238, w_018_239, w_018_240, w_018_241, w_018_242, w_018_243, w_018_244, w_018_245, w_018_246, w_018_247, w_018_248, w_018_250, w_018_251, w_018_252, w_018_253, w_018_254, w_018_255, w_018_256, w_018_257, w_018_258, w_018_259, w_018_261, w_018_263, w_018_264, w_018_265, w_018_267;
  wire w_019_000, w_019_001, w_019_002, w_019_003, w_019_004, w_019_005, w_019_006, w_019_007, w_019_008, w_019_009, w_019_010, w_019_011, w_019_012, w_019_013, w_019_014, w_019_015, w_019_016, w_019_017, w_019_018, w_019_019, w_019_020, w_019_021, w_019_022, w_019_023, w_019_024, w_019_025, w_019_026, w_019_027, w_019_028, w_019_029, w_019_030, w_019_031, w_019_032, w_019_033, w_019_034, w_019_035, w_019_036, w_019_037, w_019_038, w_019_039, w_019_040, w_019_041, w_019_042, w_019_043, w_019_044, w_019_045, w_019_046, w_019_047, w_019_048, w_019_049, w_019_050, w_019_051, w_019_052, w_019_053, w_019_054, w_019_055, w_019_056, w_019_057, w_019_058, w_019_059, w_019_060, w_019_061, w_019_062, w_019_063, w_019_064, w_019_065, w_019_066, w_019_067, w_019_068, w_019_069, w_019_070, w_019_071, w_019_072, w_019_073, w_019_074, w_019_075, w_019_076, w_019_077, w_019_078, w_019_079, w_019_080, w_019_081, w_019_082, w_019_083, w_019_084, w_019_085, w_019_086, w_019_087, w_019_088, w_019_089, w_019_090, w_019_091, w_019_092, w_019_093, w_019_094, w_019_095, w_019_096, w_019_097, w_019_098, w_019_099, w_019_100, w_019_101, w_019_102, w_019_103, w_019_104, w_019_105, w_019_106, w_019_107, w_019_108, w_019_109, w_019_110, w_019_111, w_019_112, w_019_113, w_019_114, w_019_115, w_019_116, w_019_117, w_019_118, w_019_119, w_019_120, w_019_121, w_019_122, w_019_123, w_019_124, w_019_125, w_019_126, w_019_127, w_019_128, w_019_129, w_019_130, w_019_131, w_019_132, w_019_133, w_019_134, w_019_135, w_019_136, w_019_137, w_019_138, w_019_139, w_019_140, w_019_141, w_019_142, w_019_143, w_019_144, w_019_145, w_019_146, w_019_147, w_019_148, w_019_149, w_019_150, w_019_151, w_019_152, w_019_153, w_019_154, w_019_155, w_019_156, w_019_157, w_019_158, w_019_159, w_019_160, w_019_161, w_019_162, w_019_163, w_019_164, w_019_165, w_019_166, w_019_167, w_019_168, w_019_169, w_019_170, w_019_171, w_019_172, w_019_173, w_019_174, w_019_175, w_019_176, w_019_177, w_019_178, w_019_179, w_019_180, w_019_181, w_019_182, w_019_183, w_019_184, w_019_185, w_019_186, w_019_187, w_019_188, w_019_189, w_019_190, w_019_191, w_019_192, w_019_193, w_019_194, w_019_195, w_019_196, w_019_197, w_019_198, w_019_199, w_019_200, w_019_201, w_019_202, w_019_203, w_019_204, w_019_205, w_019_206, w_019_207, w_019_208, w_019_209, w_019_210, w_019_211, w_019_212, w_019_213, w_019_214, w_019_215, w_019_216, w_019_217, w_019_218, w_019_219, w_019_220, w_019_221, w_019_222, w_019_223, w_019_224, w_019_225, w_019_226, w_019_227, w_019_228, w_019_229, w_019_230, w_019_231, w_019_232, w_019_233, w_019_234, w_019_235, w_019_236, w_019_237, w_019_238, w_019_239, w_019_240, w_019_241, w_019_242, w_019_243, w_019_244, w_019_245, w_019_246, w_019_247, w_019_248, w_019_249, w_019_250, w_019_251, w_019_252, w_019_253, w_019_254, w_019_255, w_019_256, w_019_257, w_019_258, w_019_259, w_019_260, w_019_261, w_019_262, w_019_263, w_019_264, w_019_265, w_019_266, w_019_267, w_019_268, w_019_269, w_019_270, w_019_271, w_019_272, w_019_273, w_019_274, w_019_275, w_019_276, w_019_277, w_019_278, w_019_279, w_019_280, w_019_281, w_019_282, w_019_283, w_019_284, w_019_285, w_019_286, w_019_287, w_019_288, w_019_289, w_019_290, w_019_291, w_019_292, w_019_293, w_019_294, w_019_295, w_019_296, w_019_297, w_019_298, w_019_299, w_019_300, w_019_301, w_019_302, w_019_303, w_019_304, w_019_305, w_019_306, w_019_307, w_019_308, w_019_309, w_019_310, w_019_311, w_019_312, w_019_313, w_019_314, w_019_315, w_019_316, w_019_317, w_019_318, w_019_319, w_019_320, w_019_321, w_019_322, w_019_323, w_019_324, w_019_325, w_019_326, w_019_327, w_019_328, w_019_329, w_019_330, w_019_331, w_019_332, w_019_333, w_019_334, w_019_335, w_019_336, w_019_337, w_019_338, w_019_339, w_019_340, w_019_341, w_019_342, w_019_343, w_019_344, w_019_345, w_019_346, w_019_347, w_019_348, w_019_349, w_019_350, w_019_351, w_019_352, w_019_353, w_019_354, w_019_355, w_019_356, w_019_357, w_019_358, w_019_359, w_019_360, w_019_361, w_019_362, w_019_363, w_019_364, w_019_365, w_019_366, w_019_367, w_019_368, w_019_369, w_019_370, w_019_371, w_019_372, w_019_373, w_019_374, w_019_375, w_019_376, w_019_377, w_019_378, w_019_379, w_019_380, w_019_381, w_019_382, w_019_383, w_019_384, w_019_385, w_019_386, w_019_387, w_019_388, w_019_389, w_019_390, w_019_391, w_019_392, w_019_393, w_019_394, w_019_395, w_019_396, w_019_397, w_019_398, w_019_399, w_019_400, w_019_401, w_019_402, w_019_403, w_019_404, w_019_405, w_019_406, w_019_407, w_019_408, w_019_409, w_019_410, w_019_411, w_019_412, w_019_413, w_019_414, w_019_415, w_019_417, w_019_418, w_019_419, w_019_420, w_019_421, w_019_422, w_019_423, w_019_424, w_019_425, w_019_426, w_019_427, w_019_428, w_019_429, w_019_430, w_019_431, w_019_432, w_019_433, w_019_434, w_019_435, w_019_436, w_019_437, w_019_438, w_019_439, w_019_440, w_019_441, w_019_442, w_019_443, w_019_444, w_019_445, w_019_446, w_019_447, w_019_448, w_019_449, w_019_450, w_019_451, w_019_452, w_019_453, w_019_454, w_019_455, w_019_456, w_019_457, w_019_458, w_019_459, w_019_460, w_019_461, w_019_462, w_019_463, w_019_464, w_019_465, w_019_466, w_019_467, w_019_468, w_019_469, w_019_470, w_019_471, w_019_472, w_019_473, w_019_474, w_019_475, w_019_476, w_019_477, w_019_478, w_019_479, w_019_480, w_019_481, w_019_482, w_019_483, w_019_484, w_019_485, w_019_486, w_019_487, w_019_488, w_019_489, w_019_490, w_019_491, w_019_492, w_019_493, w_019_494, w_019_495, w_019_496, w_019_497, w_019_498, w_019_499, w_019_500, w_019_501, w_019_502, w_019_503, w_019_504, w_019_505, w_019_506, w_019_507, w_019_508, w_019_509, w_019_510, w_019_511, w_019_512, w_019_513, w_019_514, w_019_515, w_019_516, w_019_517, w_019_518, w_019_519, w_019_520, w_019_521, w_019_522, w_019_523, w_019_524, w_019_525, w_019_526, w_019_527, w_019_528, w_019_529, w_019_530, w_019_531, w_019_532, w_019_533, w_019_534, w_019_535, w_019_536, w_019_537, w_019_538, w_019_539, w_019_540, w_019_541, w_019_542, w_019_543, w_019_544, w_019_545, w_019_546, w_019_547, w_019_548, w_019_549, w_019_550, w_019_551, w_019_552, w_019_553, w_019_554, w_019_555, w_019_556, w_019_558, w_019_559, w_019_560, w_019_561, w_019_562, w_019_563, w_019_564, w_019_565, w_019_566, w_019_567, w_019_568, w_019_569, w_019_570, w_019_571, w_019_572, w_019_573, w_019_574, w_019_575, w_019_576, w_019_577, w_019_578, w_019_579, w_019_580, w_019_581, w_019_582, w_019_583, w_019_584, w_019_585, w_019_586, w_019_587, w_019_588, w_019_589, w_019_590, w_019_591, w_019_592, w_019_593, w_019_594, w_019_595, w_019_596, w_019_597, w_019_598, w_019_599, w_019_600, w_019_601, w_019_602, w_019_603, w_019_604, w_019_605, w_019_606, w_019_607, w_019_608, w_019_609, w_019_610, w_019_611, w_019_612, w_019_613, w_019_614, w_019_615, w_019_616, w_019_617, w_019_618, w_019_619, w_019_620, w_019_621, w_019_622, w_019_623, w_019_624, w_019_625, w_019_626, w_019_627, w_019_628, w_019_629, w_019_630, w_019_631, w_019_632, w_019_633, w_019_634, w_019_635, w_019_636, w_019_637, w_019_638, w_019_639, w_019_640, w_019_641, w_019_642, w_019_643, w_019_644, w_019_645, w_019_646, w_019_647, w_019_648, w_019_649, w_019_650, w_019_651, w_019_652, w_019_653, w_019_654, w_019_655, w_019_656, w_019_657, w_019_658, w_019_659, w_019_660, w_019_661, w_019_662, w_019_663, w_019_664, w_019_665, w_019_666, w_019_667, w_019_668, w_019_669, w_019_670, w_019_671, w_019_672, w_019_673, w_019_674, w_019_675, w_019_676, w_019_677, w_019_678, w_019_679, w_019_680, w_019_681, w_019_682, w_019_683, w_019_684, w_019_685, w_019_686, w_019_687, w_019_688, w_019_689, w_019_690, w_019_691, w_019_692, w_019_693, w_019_694, w_019_695, w_019_696, w_019_697, w_019_698, w_019_699, w_019_700, w_019_701, w_019_702, w_019_703, w_019_704, w_019_705, w_019_706, w_019_707, w_019_708, w_019_709, w_019_710, w_019_711, w_019_712, w_019_713, w_019_714, w_019_715, w_019_716, w_019_717, w_019_718, w_019_719, w_019_720, w_019_721, w_019_722, w_019_723, w_019_724, w_019_725, w_019_726, w_019_727, w_019_728, w_019_729, w_019_730, w_019_731, w_019_732, w_019_733, w_019_734, w_019_735, w_019_736, w_019_737, w_019_738, w_019_739, w_019_740, w_019_741, w_019_742, w_019_743, w_019_744, w_019_745, w_019_746, w_019_747, w_019_748, w_019_749, w_019_750, w_019_751, w_019_752, w_019_753, w_019_754, w_019_755, w_019_756, w_019_757, w_019_758, w_019_759, w_019_760, w_019_761, w_019_762, w_019_763, w_019_764, w_019_765, w_019_766, w_019_767, w_019_768, w_019_769, w_019_770, w_019_771, w_019_772, w_019_773, w_019_774, w_019_775, w_019_776, w_019_777, w_019_778, w_019_779, w_019_780, w_019_781, w_019_782, w_019_783, w_019_784, w_019_785, w_019_786, w_019_787, w_019_788, w_019_789, w_019_790, w_019_791, w_019_792, w_019_793, w_019_794, w_019_795, w_019_796, w_019_797, w_019_798, w_019_799, w_019_800, w_019_801, w_019_802, w_019_803, w_019_804, w_019_805, w_019_806, w_019_807, w_019_808, w_019_809, w_019_810, w_019_811, w_019_812, w_019_813, w_019_814, w_019_815, w_019_816, w_019_817, w_019_818, w_019_819, w_019_820, w_019_821, w_019_822, w_019_823, w_019_824, w_019_825, w_019_826, w_019_827, w_019_828, w_019_829, w_019_830, w_019_831, w_019_832, w_019_833, w_019_834, w_019_835, w_019_836, w_019_837, w_019_838, w_019_839, w_019_840, w_019_841, w_019_842, w_019_843, w_019_844, w_019_845, w_019_846, w_019_847, w_019_848, w_019_849, w_019_850, w_019_851, w_019_852, w_019_853, w_019_854, w_019_855, w_019_856, w_019_857, w_019_858, w_019_859, w_019_860, w_019_861, w_019_862, w_019_863, w_019_864, w_019_865, w_019_866, w_019_867, w_019_868, w_019_869, w_019_870, w_019_871, w_019_872, w_019_873, w_019_874, w_019_875, w_019_876, w_019_877, w_019_878, w_019_879, w_019_880, w_019_881, w_019_882, w_019_883, w_019_884, w_019_885, w_019_886, w_019_887, w_019_888, w_019_889, w_019_890, w_019_891, w_019_892, w_019_893, w_019_894, w_019_895, w_019_896, w_019_897, w_019_898, w_019_899, w_019_900, w_019_901, w_019_902, w_019_903, w_019_904, w_019_905, w_019_906, w_019_907, w_019_908, w_019_909, w_019_910, w_019_911, w_019_912, w_019_913, w_019_914, w_019_915, w_019_916, w_019_917, w_019_918, w_019_919, w_019_920, w_019_921, w_019_922, w_019_923, w_019_924, w_019_925, w_019_926, w_019_927, w_019_928, w_019_929, w_019_930, w_019_931, w_019_932, w_019_933, w_019_934, w_019_935, w_019_936, w_019_937, w_019_938, w_019_939, w_019_940, w_019_941, w_019_942, w_019_943, w_019_944, w_019_945, w_019_946, w_019_947, w_019_948, w_019_949, w_019_950, w_019_951, w_019_952, w_019_953, w_019_954, w_019_955, w_019_956, w_019_957, w_019_958, w_019_959, w_019_960, w_019_961, w_019_962, w_019_963, w_019_964, w_019_965, w_019_966, w_019_967, w_019_968, w_019_969, w_019_970, w_019_971, w_019_972, w_019_973, w_019_974, w_019_975, w_019_976, w_019_977, w_019_978, w_019_979, w_019_980, w_019_981, w_019_982, w_019_983, w_019_984, w_019_985, w_019_986, w_019_987, w_019_988, w_019_989, w_019_990, w_019_991, w_019_992, w_019_993, w_019_994, w_019_995, w_019_996, w_019_997, w_019_998, w_019_999, w_019_1000, w_019_1001, w_019_1002, w_019_1003, w_019_1004, w_019_1005, w_019_1006, w_019_1007, w_019_1008, w_019_1009, w_019_1010, w_019_1011, w_019_1012, w_019_1013, w_019_1014, w_019_1015, w_019_1016, w_019_1017, w_019_1018, w_019_1019, w_019_1020, w_019_1021, w_019_1022, w_019_1023, w_019_1024, w_019_1025, w_019_1026, w_019_1027, w_019_1028, w_019_1029, w_019_1030, w_019_1031, w_019_1032, w_019_1033, w_019_1034, w_019_1035, w_019_1036, w_019_1037, w_019_1038, w_019_1039, w_019_1040, w_019_1041, w_019_1042, w_019_1043, w_019_1044, w_019_1045, w_019_1046, w_019_1047, w_019_1048, w_019_1049, w_019_1050, w_019_1051, w_019_1052, w_019_1053, w_019_1054, w_019_1055, w_019_1056, w_019_1057, w_019_1058, w_019_1059, w_019_1060, w_019_1061, w_019_1062, w_019_1063, w_019_1064, w_019_1065, w_019_1066, w_019_1067, w_019_1068, w_019_1069, w_019_1070, w_019_1071, w_019_1072, w_019_1073, w_019_1074, w_019_1075, w_019_1076, w_019_1077, w_019_1078, w_019_1079, w_019_1080, w_019_1081, w_019_1082;
  wire w_020_000, w_020_001, w_020_002, w_020_003, w_020_004, w_020_005, w_020_006, w_020_007, w_020_008, w_020_009, w_020_010, w_020_011, w_020_012, w_020_013, w_020_014, w_020_015, w_020_016, w_020_017, w_020_018, w_020_019, w_020_020, w_020_021, w_020_022, w_020_023, w_020_024, w_020_025, w_020_026, w_020_027, w_020_028, w_020_029, w_020_030, w_020_031, w_020_032, w_020_033, w_020_034, w_020_035, w_020_036, w_020_037, w_020_038, w_020_039, w_020_040, w_020_041, w_020_042, w_020_043, w_020_044, w_020_045, w_020_046, w_020_047, w_020_048, w_020_049, w_020_050, w_020_051, w_020_052, w_020_053, w_020_054, w_020_055, w_020_056, w_020_057, w_020_058, w_020_059, w_020_060, w_020_061, w_020_062, w_020_063, w_020_064, w_020_065, w_020_066, w_020_067, w_020_068, w_020_069, w_020_070, w_020_071, w_020_072, w_020_073, w_020_074, w_020_075, w_020_076, w_020_077, w_020_078, w_020_079, w_020_080, w_020_081, w_020_082, w_020_083, w_020_084, w_020_085, w_020_086, w_020_087, w_020_088, w_020_089, w_020_090, w_020_091, w_020_092, w_020_093, w_020_094, w_020_095, w_020_096, w_020_097, w_020_098, w_020_099, w_020_100, w_020_101, w_020_102, w_020_103, w_020_104, w_020_105, w_020_106, w_020_107, w_020_108, w_020_109, w_020_110, w_020_111, w_020_112, w_020_113, w_020_114, w_020_115, w_020_116, w_020_117, w_020_118, w_020_119, w_020_120, w_020_121, w_020_122, w_020_123, w_020_124, w_020_125, w_020_126, w_020_127, w_020_128, w_020_129, w_020_130, w_020_131, w_020_132, w_020_133, w_020_134, w_020_135, w_020_136, w_020_137, w_020_138, w_020_139, w_020_140, w_020_141, w_020_142, w_020_143, w_020_144, w_020_145, w_020_146, w_020_147, w_020_148, w_020_149, w_020_150, w_020_151, w_020_152, w_020_153, w_020_154, w_020_155, w_020_156, w_020_157, w_020_158, w_020_159, w_020_160, w_020_161, w_020_162, w_020_163, w_020_164, w_020_165, w_020_166, w_020_167, w_020_168, w_020_169, w_020_170, w_020_171, w_020_172, w_020_173, w_020_174, w_020_175, w_020_176, w_020_177, w_020_178, w_020_179, w_020_180, w_020_181, w_020_182, w_020_183, w_020_184, w_020_185, w_020_186, w_020_187, w_020_188, w_020_189, w_020_190, w_020_191, w_020_192, w_020_193, w_020_194, w_020_195, w_020_196, w_020_197, w_020_198, w_020_199, w_020_200, w_020_201, w_020_202, w_020_203, w_020_204, w_020_205, w_020_206, w_020_207, w_020_208, w_020_209, w_020_210, w_020_211, w_020_212, w_020_213, w_020_214, w_020_215, w_020_216, w_020_217, w_020_218, w_020_219, w_020_220, w_020_221, w_020_222, w_020_223, w_020_224, w_020_225, w_020_226, w_020_227, w_020_228, w_020_229, w_020_230, w_020_231, w_020_232, w_020_233, w_020_234, w_020_235, w_020_236, w_020_237, w_020_238, w_020_239, w_020_240, w_020_241, w_020_242, w_020_243, w_020_244, w_020_245, w_020_246, w_020_247, w_020_248, w_020_249, w_020_250, w_020_251, w_020_252, w_020_253, w_020_254, w_020_255, w_020_256, w_020_257, w_020_258, w_020_259, w_020_260, w_020_261, w_020_262, w_020_263, w_020_264, w_020_265, w_020_266, w_020_267, w_020_268, w_020_269, w_020_270, w_020_271, w_020_272, w_020_273, w_020_274, w_020_275, w_020_276, w_020_277, w_020_278, w_020_279, w_020_280, w_020_281, w_020_282, w_020_283, w_020_284, w_020_285, w_020_286, w_020_287, w_020_288, w_020_289, w_020_290, w_020_291, w_020_292, w_020_293, w_020_294, w_020_295, w_020_296, w_020_297, w_020_298, w_020_299, w_020_300, w_020_301, w_020_302, w_020_303, w_020_304, w_020_305, w_020_306, w_020_307, w_020_308, w_020_309, w_020_310, w_020_311, w_020_312, w_020_313, w_020_314, w_020_315, w_020_316, w_020_317, w_020_318, w_020_319, w_020_320, w_020_321, w_020_322, w_020_323, w_020_324, w_020_325, w_020_326, w_020_327, w_020_328, w_020_329, w_020_330, w_020_331, w_020_332, w_020_333, w_020_334, w_020_335, w_020_336, w_020_337, w_020_338, w_020_339, w_020_340, w_020_341, w_020_342, w_020_343, w_020_344, w_020_345, w_020_346, w_020_347, w_020_348, w_020_349, w_020_350, w_020_351, w_020_352, w_020_353, w_020_354, w_020_355, w_020_356, w_020_357, w_020_358, w_020_359, w_020_360, w_020_361, w_020_362, w_020_363, w_020_364, w_020_365, w_020_366, w_020_367, w_020_368, w_020_369, w_020_370, w_020_371, w_020_372, w_020_373, w_020_374, w_020_375, w_020_376, w_020_377, w_020_378, w_020_379, w_020_380, w_020_381, w_020_382, w_020_383, w_020_384, w_020_385, w_020_386, w_020_387, w_020_388, w_020_389, w_020_390, w_020_391, w_020_392, w_020_393, w_020_394, w_020_395, w_020_396, w_020_397, w_020_398, w_020_399, w_020_400, w_020_401, w_020_402, w_020_403, w_020_404, w_020_405, w_020_406, w_020_407, w_020_408, w_020_409, w_020_410, w_020_411, w_020_412, w_020_413, w_020_414, w_020_415, w_020_416, w_020_417, w_020_418, w_020_419, w_020_420, w_020_421, w_020_422, w_020_423, w_020_424, w_020_425, w_020_426, w_020_427, w_020_428, w_020_429, w_020_430, w_020_431, w_020_432, w_020_433, w_020_434, w_020_435, w_020_436, w_020_437, w_020_438, w_020_439, w_020_440, w_020_441, w_020_442, w_020_443, w_020_444, w_020_445, w_020_446, w_020_447, w_020_448, w_020_449, w_020_450, w_020_451, w_020_452, w_020_453, w_020_454, w_020_455, w_020_456, w_020_457, w_020_458, w_020_459, w_020_460, w_020_461, w_020_462, w_020_463, w_020_464, w_020_465, w_020_466, w_020_467, w_020_468, w_020_469, w_020_470, w_020_471, w_020_472, w_020_473, w_020_474, w_020_475, w_020_476, w_020_477, w_020_478, w_020_479, w_020_480, w_020_481, w_020_482, w_020_483, w_020_484, w_020_485, w_020_486, w_020_487, w_020_488, w_020_489, w_020_490, w_020_491, w_020_492, w_020_493, w_020_494, w_020_495, w_020_496, w_020_497, w_020_498, w_020_499, w_020_500, w_020_501, w_020_502, w_020_503, w_020_504, w_020_505, w_020_506, w_020_507, w_020_508, w_020_509, w_020_510, w_020_511, w_020_512, w_020_513, w_020_514, w_020_515, w_020_516, w_020_517, w_020_518, w_020_519, w_020_520, w_020_521, w_020_522, w_020_523, w_020_524, w_020_525, w_020_526, w_020_527, w_020_528, w_020_529, w_020_530, w_020_531, w_020_532, w_020_533, w_020_534, w_020_535, w_020_536, w_020_537, w_020_538, w_020_539, w_020_540, w_020_541, w_020_542, w_020_543, w_020_544, w_020_545, w_020_546, w_020_547, w_020_548, w_020_549, w_020_550, w_020_551, w_020_552, w_020_553, w_020_554, w_020_555, w_020_556, w_020_557, w_020_558, w_020_559, w_020_560, w_020_561, w_020_562, w_020_563, w_020_564, w_020_565, w_020_566, w_020_567, w_020_568, w_020_569, w_020_570, w_020_571, w_020_572, w_020_573, w_020_574, w_020_575, w_020_576, w_020_577, w_020_578, w_020_579, w_020_580, w_020_581, w_020_582, w_020_583, w_020_584, w_020_585, w_020_586, w_020_587, w_020_588, w_020_589, w_020_590, w_020_591, w_020_592, w_020_593, w_020_594, w_020_595, w_020_596, w_020_597, w_020_598, w_020_599, w_020_600, w_020_601, w_020_602, w_020_603, w_020_604, w_020_605, w_020_606, w_020_607, w_020_608, w_020_609, w_020_610, w_020_611, w_020_612, w_020_613, w_020_614, w_020_615, w_020_616, w_020_617, w_020_618, w_020_619, w_020_620, w_020_621, w_020_622, w_020_623, w_020_624, w_020_625, w_020_626, w_020_627, w_020_628, w_020_629, w_020_630, w_020_631, w_020_632, w_020_633, w_020_634, w_020_635, w_020_636, w_020_637, w_020_638, w_020_639, w_020_640, w_020_641, w_020_642, w_020_643, w_020_644, w_020_645, w_020_646, w_020_647, w_020_648, w_020_649, w_020_650, w_020_651, w_020_652, w_020_653, w_020_654, w_020_655, w_020_656, w_020_657, w_020_658, w_020_659, w_020_660, w_020_661, w_020_662, w_020_663, w_020_664, w_020_665, w_020_666, w_020_667, w_020_668, w_020_669, w_020_670, w_020_671, w_020_672, w_020_673, w_020_674, w_020_675, w_020_676, w_020_677, w_020_678, w_020_679, w_020_680, w_020_681, w_020_682, w_020_683, w_020_684, w_020_685, w_020_686, w_020_687, w_020_688, w_020_689, w_020_690, w_020_691, w_020_692, w_020_693, w_020_694, w_020_695, w_020_696, w_020_697, w_020_698, w_020_699, w_020_700, w_020_701, w_020_702, w_020_703, w_020_704, w_020_705, w_020_706, w_020_707, w_020_708, w_020_709, w_020_710, w_020_711, w_020_712, w_020_713, w_020_714, w_020_715, w_020_716, w_020_717, w_020_718, w_020_719, w_020_720, w_020_721, w_020_722, w_020_723, w_020_724, w_020_725, w_020_726, w_020_727, w_020_728, w_020_729, w_020_730, w_020_731, w_020_732, w_020_733, w_020_734, w_020_735, w_020_736, w_020_737, w_020_738, w_020_739, w_020_740, w_020_741, w_020_742, w_020_743, w_020_744, w_020_745, w_020_746, w_020_747, w_020_748, w_020_749, w_020_750, w_020_751, w_020_752, w_020_753, w_020_754, w_020_755, w_020_756, w_020_757, w_020_758, w_020_759, w_020_760, w_020_761, w_020_762, w_020_763, w_020_764, w_020_765, w_020_766, w_020_767, w_020_768, w_020_769, w_020_770, w_020_771, w_020_772, w_020_773, w_020_774, w_020_775, w_020_776, w_020_777, w_020_778, w_020_779, w_020_780, w_020_781, w_020_782, w_020_783, w_020_784, w_020_785, w_020_786, w_020_787, w_020_788, w_020_789, w_020_790, w_020_791, w_020_792, w_020_793, w_020_794, w_020_795, w_020_796, w_020_797, w_020_798, w_020_799, w_020_800, w_020_801, w_020_802, w_020_803, w_020_804, w_020_805, w_020_806, w_020_807, w_020_808, w_020_809, w_020_810, w_020_811, w_020_812, w_020_813, w_020_814, w_020_815, w_020_816, w_020_817, w_020_818, w_020_819, w_020_820, w_020_821, w_020_822, w_020_823, w_020_824, w_020_825, w_020_826, w_020_827, w_020_828, w_020_829, w_020_830, w_020_831, w_020_832, w_020_833, w_020_834, w_020_835, w_020_836, w_020_837, w_020_838, w_020_839, w_020_840, w_020_841, w_020_842, w_020_844, w_020_845, w_020_846, w_020_847, w_020_848, w_020_849, w_020_850, w_020_851, w_020_852, w_020_853, w_020_854, w_020_855, w_020_856, w_020_857, w_020_858, w_020_859, w_020_860, w_020_861, w_020_862, w_020_863, w_020_864, w_020_865, w_020_866, w_020_867, w_020_868, w_020_869, w_020_870, w_020_871, w_020_872, w_020_873, w_020_874, w_020_875, w_020_876, w_020_877, w_020_878, w_020_879, w_020_880, w_020_881, w_020_882, w_020_883, w_020_884, w_020_885, w_020_886, w_020_887, w_020_888, w_020_889, w_020_890, w_020_891, w_020_892, w_020_893, w_020_894, w_020_895, w_020_896, w_020_897, w_020_898, w_020_899, w_020_900, w_020_901, w_020_902, w_020_903, w_020_904, w_020_905, w_020_906, w_020_907, w_020_908, w_020_909, w_020_910, w_020_911, w_020_912, w_020_913, w_020_914, w_020_915, w_020_916, w_020_917, w_020_918, w_020_919, w_020_920, w_020_921, w_020_922, w_020_923, w_020_924, w_020_925, w_020_926, w_020_927, w_020_928, w_020_929, w_020_930, w_020_931, w_020_932, w_020_933, w_020_934, w_020_935, w_020_936;
  wire w_021_000, w_021_001, w_021_002, w_021_003, w_021_004, w_021_005, w_021_006, w_021_007, w_021_008, w_021_009, w_021_010, w_021_011, w_021_012, w_021_013, w_021_014, w_021_015, w_021_016, w_021_017, w_021_018, w_021_019, w_021_020, w_021_021, w_021_022, w_021_023, w_021_024, w_021_025, w_021_026, w_021_027, w_021_028, w_021_029, w_021_030, w_021_031, w_021_032, w_021_033, w_021_034, w_021_035, w_021_036, w_021_037, w_021_038, w_021_039, w_021_040, w_021_041, w_021_042, w_021_043, w_021_044, w_021_045, w_021_046, w_021_047, w_021_048, w_021_049, w_021_050, w_021_051, w_021_052, w_021_053, w_021_054, w_021_055, w_021_056, w_021_057, w_021_058, w_021_059, w_021_060, w_021_061, w_021_062, w_021_063, w_021_064, w_021_065, w_021_066, w_021_067, w_021_068, w_021_069, w_021_070, w_021_071, w_021_072, w_021_073, w_021_074, w_021_075, w_021_076, w_021_077, w_021_078, w_021_079, w_021_080, w_021_081, w_021_082, w_021_083, w_021_084, w_021_085, w_021_086, w_021_087, w_021_088, w_021_089, w_021_090, w_021_091, w_021_092, w_021_093, w_021_094, w_021_095, w_021_096, w_021_097, w_021_098, w_021_099, w_021_100, w_021_101, w_021_102, w_021_103, w_021_104, w_021_105, w_021_106, w_021_107, w_021_108, w_021_109, w_021_110, w_021_111, w_021_112, w_021_113, w_021_114, w_021_115, w_021_116, w_021_117, w_021_118, w_021_119, w_021_120, w_021_121, w_021_122, w_021_123, w_021_124, w_021_125, w_021_126, w_021_127, w_021_128, w_021_129, w_021_130, w_021_131, w_021_132, w_021_133, w_021_134, w_021_135, w_021_136, w_021_137, w_021_138, w_021_139, w_021_140, w_021_141, w_021_142, w_021_143, w_021_144, w_021_145, w_021_146, w_021_147, w_021_148, w_021_149, w_021_150, w_021_151, w_021_152, w_021_153, w_021_154, w_021_155, w_021_156, w_021_157, w_021_158, w_021_159, w_021_160, w_021_161, w_021_162, w_021_163, w_021_164, w_021_165, w_021_166, w_021_167, w_021_168, w_021_169, w_021_170, w_021_171, w_021_172, w_021_173, w_021_174, w_021_175, w_021_176, w_021_177, w_021_178, w_021_179, w_021_180, w_021_181, w_021_182, w_021_183, w_021_184, w_021_185, w_021_186, w_021_187, w_021_188, w_021_189, w_021_190, w_021_191, w_021_192, w_021_193, w_021_194, w_021_195, w_021_196, w_021_197, w_021_198, w_021_199, w_021_200, w_021_201, w_021_202, w_021_203, w_021_204, w_021_205, w_021_206, w_021_207, w_021_208, w_021_209, w_021_210, w_021_211, w_021_212, w_021_213, w_021_214, w_021_215, w_021_216, w_021_217, w_021_218, w_021_219, w_021_220, w_021_221, w_021_222, w_021_223, w_021_224, w_021_225, w_021_226, w_021_227, w_021_228, w_021_229, w_021_230, w_021_231, w_021_232, w_021_233, w_021_234, w_021_235, w_021_236, w_021_237, w_021_238, w_021_239, w_021_240, w_021_241, w_021_242, w_021_243, w_021_244, w_021_245, w_021_246, w_021_247, w_021_248, w_021_249, w_021_250, w_021_251, w_021_252, w_021_253, w_021_254, w_021_255, w_021_256, w_021_257, w_021_258, w_021_259, w_021_260, w_021_261, w_021_262, w_021_263, w_021_264, w_021_265, w_021_266, w_021_267, w_021_268, w_021_269, w_021_270, w_021_271, w_021_272, w_021_273, w_021_274, w_021_275, w_021_276, w_021_277, w_021_278, w_021_279, w_021_280, w_021_281, w_021_282, w_021_283, w_021_284, w_021_285, w_021_286, w_021_287, w_021_288, w_021_289, w_021_290, w_021_291, w_021_292, w_021_293, w_021_294, w_021_295, w_021_296, w_021_297, w_021_298, w_021_299, w_021_300, w_021_301, w_021_302, w_021_303, w_021_304, w_021_305, w_021_306, w_021_307, w_021_308, w_021_309, w_021_310, w_021_311, w_021_312, w_021_313, w_021_314, w_021_315, w_021_316, w_021_317, w_021_318, w_021_319, w_021_320, w_021_321, w_021_322, w_021_323, w_021_324, w_021_325, w_021_326, w_021_327, w_021_328, w_021_329, w_021_330, w_021_331, w_021_332, w_021_333, w_021_334, w_021_335, w_021_336, w_021_337, w_021_338, w_021_339, w_021_340, w_021_341, w_021_342, w_021_343, w_021_344, w_021_345, w_021_346, w_021_347, w_021_348, w_021_349, w_021_350, w_021_351, w_021_352, w_021_353, w_021_354, w_021_355, w_021_356, w_021_357, w_021_358, w_021_359, w_021_360, w_021_361, w_021_362, w_021_363, w_021_364, w_021_365, w_021_366, w_021_367, w_021_368, w_021_369, w_021_370, w_021_371, w_021_372, w_021_373, w_021_374, w_021_375, w_021_376, w_021_377, w_021_378, w_021_379, w_021_380, w_021_381, w_021_382, w_021_383, w_021_384, w_021_385, w_021_386, w_021_387, w_021_388, w_021_389, w_021_390, w_021_391, w_021_392, w_021_393, w_021_394, w_021_395, w_021_396, w_021_397, w_021_398, w_021_399, w_021_400, w_021_401, w_021_402, w_021_403, w_021_404, w_021_405, w_021_406, w_021_407, w_021_408, w_021_409, w_021_410, w_021_411, w_021_412, w_021_413, w_021_414, w_021_415, w_021_416, w_021_417, w_021_418, w_021_419, w_021_420, w_021_421, w_021_422, w_021_423, w_021_424, w_021_425, w_021_426, w_021_427, w_021_428, w_021_429, w_021_430, w_021_431, w_021_432, w_021_433, w_021_434, w_021_435, w_021_436, w_021_437, w_021_438, w_021_439, w_021_440, w_021_441, w_021_442, w_021_443, w_021_444, w_021_445, w_021_446, w_021_447, w_021_448, w_021_449, w_021_450, w_021_451, w_021_452, w_021_453, w_021_454, w_021_455, w_021_456, w_021_457, w_021_458, w_021_459, w_021_460, w_021_461, w_021_462, w_021_463, w_021_464, w_021_465, w_021_466, w_021_467, w_021_468, w_021_469, w_021_470, w_021_471, w_021_472, w_021_473, w_021_474, w_021_475, w_021_476, w_021_477, w_021_478, w_021_479, w_021_480, w_021_481, w_021_482, w_021_483, w_021_484, w_021_485, w_021_486, w_021_487, w_021_488, w_021_489, w_021_490, w_021_491, w_021_492, w_021_493, w_021_494, w_021_495, w_021_496, w_021_497, w_021_498, w_021_499, w_021_500, w_021_501, w_021_502, w_021_503, w_021_504, w_021_505, w_021_506, w_021_507, w_021_508, w_021_509, w_021_510, w_021_511, w_021_512, w_021_513, w_021_514, w_021_515, w_021_516, w_021_517, w_021_518, w_021_519, w_021_520, w_021_521, w_021_522, w_021_523, w_021_524, w_021_525, w_021_526, w_021_527, w_021_528, w_021_529, w_021_530, w_021_531, w_021_532, w_021_533, w_021_534, w_021_535, w_021_536, w_021_537, w_021_538, w_021_539, w_021_540, w_021_541, w_021_542, w_021_543, w_021_544, w_021_545, w_021_546, w_021_547, w_021_548, w_021_549, w_021_550, w_021_551, w_021_552, w_021_553, w_021_554, w_021_555, w_021_556, w_021_557, w_021_558, w_021_559, w_021_560, w_021_561, w_021_562, w_021_563, w_021_564, w_021_565, w_021_566, w_021_567, w_021_568, w_021_569, w_021_570, w_021_571, w_021_572, w_021_573, w_021_574, w_021_575, w_021_576, w_021_577, w_021_578, w_021_579, w_021_580, w_021_581, w_021_582, w_021_583, w_021_584, w_021_585, w_021_586, w_021_587, w_021_588, w_021_589, w_021_590, w_021_591, w_021_592, w_021_593, w_021_594, w_021_595, w_021_596, w_021_597, w_021_598, w_021_599, w_021_600, w_021_601, w_021_602, w_021_603, w_021_604, w_021_605, w_021_606, w_021_607, w_021_608, w_021_609, w_021_610, w_021_611, w_021_612, w_021_613, w_021_614, w_021_615, w_021_616, w_021_617, w_021_618, w_021_619, w_021_620, w_021_621, w_021_622, w_021_623, w_021_624, w_021_625, w_021_626, w_021_627, w_021_628, w_021_629, w_021_630, w_021_631, w_021_632, w_021_633, w_021_634, w_021_635, w_021_636, w_021_637, w_021_638, w_021_639, w_021_640, w_021_641, w_021_642, w_021_643, w_021_644, w_021_645, w_021_646, w_021_647, w_021_648, w_021_649, w_021_650, w_021_651, w_021_652, w_021_653, w_021_654, w_021_655, w_021_656, w_021_657, w_021_658, w_021_659, w_021_660, w_021_661, w_021_662, w_021_663, w_021_664, w_021_665, w_021_666, w_021_667, w_021_668, w_021_669, w_021_670, w_021_671, w_021_672, w_021_673, w_021_674, w_021_675, w_021_676, w_021_678, w_021_679, w_021_680, w_021_681, w_021_682, w_021_683, w_021_684, w_021_686;
  wire w_022_000, w_022_001, w_022_002, w_022_003, w_022_004, w_022_005, w_022_006, w_022_007, w_022_008, w_022_009, w_022_010, w_022_011, w_022_012, w_022_013, w_022_014, w_022_015, w_022_017, w_022_018, w_022_020, w_022_022, w_022_023, w_022_024, w_022_027, w_022_028, w_022_029, w_022_030, w_022_031, w_022_032, w_022_033, w_022_034, w_022_036, w_022_037, w_022_038, w_022_039, w_022_040, w_022_041, w_022_043, w_022_046, w_022_047, w_022_048, w_022_049, w_022_050, w_022_051, w_022_052, w_022_053, w_022_054, w_022_055, w_022_056, w_022_057, w_022_058, w_022_059, w_022_060, w_022_061, w_022_062, w_022_063, w_022_064, w_022_065, w_022_067, w_022_068, w_022_069, w_022_070, w_022_071, w_022_072, w_022_073, w_022_074, w_022_075, w_022_076, w_022_077, w_022_079, w_022_081, w_022_082, w_022_083, w_022_084, w_022_085, w_022_086, w_022_087, w_022_088, w_022_090, w_022_091, w_022_092, w_022_093, w_022_094, w_022_095, w_022_096, w_022_097, w_022_098, w_022_099, w_022_100, w_022_101, w_022_102, w_022_103, w_022_104, w_022_105, w_022_106, w_022_107, w_022_108, w_022_109, w_022_110, w_022_112, w_022_113, w_022_114, w_022_115, w_022_116, w_022_117, w_022_118, w_022_119, w_022_120, w_022_121, w_022_122, w_022_123, w_022_124, w_022_125, w_022_126, w_022_127, w_022_129, w_022_130, w_022_131, w_022_132, w_022_133, w_022_134, w_022_136, w_022_137, w_022_139, w_022_140, w_022_141, w_022_142, w_022_143, w_022_144, w_022_145, w_022_146, w_022_147, w_022_148, w_022_149, w_022_150, w_022_151, w_022_152, w_022_153, w_022_154, w_022_155, w_022_156, w_022_158, w_022_159, w_022_160, w_022_161, w_022_162, w_022_163, w_022_164, w_022_165, w_022_166, w_022_167, w_022_169, w_022_170, w_022_171, w_022_172, w_022_173, w_022_174, w_022_175, w_022_176, w_022_177, w_022_178, w_022_179, w_022_180, w_022_181, w_022_182, w_022_183, w_022_184, w_022_185, w_022_186, w_022_187, w_022_188, w_022_189, w_022_191, w_022_192, w_022_193, w_022_194, w_022_195, w_022_196, w_022_198, w_022_199, w_022_200, w_022_201, w_022_202, w_022_203, w_022_204, w_022_205, w_022_206, w_022_207, w_022_208, w_022_209, w_022_210, w_022_212, w_022_213, w_022_214, w_022_215, w_022_216, w_022_217, w_022_218, w_022_219, w_022_220, w_022_221, w_022_222, w_022_223, w_022_224, w_022_225, w_022_226, w_022_227, w_022_228, w_022_229, w_022_230, w_022_232, w_022_233, w_022_234, w_022_235, w_022_236, w_022_237, w_022_238, w_022_239, w_022_240, w_022_241, w_022_242, w_022_243, w_022_244, w_022_245, w_022_246, w_022_247, w_022_248, w_022_250, w_022_251, w_022_252, w_022_253, w_022_254, w_022_255, w_022_256, w_022_257, w_022_258, w_022_259, w_022_260, w_022_261, w_022_262, w_022_263, w_022_264, w_022_265, w_022_266, w_022_267, w_022_268, w_022_269, w_022_270, w_022_271, w_022_272, w_022_273, w_022_274, w_022_275, w_022_276, w_022_277, w_022_278, w_022_279, w_022_281, w_022_282, w_022_283, w_022_284, w_022_285, w_022_286, w_022_287, w_022_288, w_022_289, w_022_290, w_022_291, w_022_293, w_022_294, w_022_295, w_022_296, w_022_297, w_022_298, w_022_299, w_022_300, w_022_301, w_022_302, w_022_303, w_022_304, w_022_305, w_022_306, w_022_307, w_022_308, w_022_309, w_022_310, w_022_312, w_022_313, w_022_314, w_022_315, w_022_316, w_022_317, w_022_318, w_022_319, w_022_320, w_022_321, w_022_323, w_022_324, w_022_325, w_022_327, w_022_328, w_022_329, w_022_330, w_022_331, w_022_332, w_022_333, w_022_334, w_022_335, w_022_336, w_022_337, w_022_338, w_022_339, w_022_340, w_022_341, w_022_342, w_022_343, w_022_344, w_022_346, w_022_347, w_022_348, w_022_349, w_022_351, w_022_352, w_022_353, w_022_354, w_022_355, w_022_356, w_022_357, w_022_358, w_022_359, w_022_361, w_022_362, w_022_363, w_022_364, w_022_365, w_022_366, w_022_367, w_022_369, w_022_370, w_022_371, w_022_372, w_022_373, w_022_374, w_022_375, w_022_376, w_022_377, w_022_378, w_022_379, w_022_380, w_022_381, w_022_382, w_022_383, w_022_384, w_022_385, w_022_386, w_022_387, w_022_388, w_022_389, w_022_390, w_022_391, w_022_392, w_022_393, w_022_394, w_022_395, w_022_396, w_022_397, w_022_398, w_022_399, w_022_400, w_022_401, w_022_402, w_022_403, w_022_405, w_022_406, w_022_407, w_022_408, w_022_411, w_022_412, w_022_413, w_022_414, w_022_415, w_022_417, w_022_418, w_022_419, w_022_420, w_022_422, w_022_423, w_022_424, w_022_425, w_022_426, w_022_427, w_022_428, w_022_429, w_022_430, w_022_431, w_022_433, w_022_434, w_022_435, w_022_436, w_022_437, w_022_438, w_022_439, w_022_441, w_022_442, w_022_443, w_022_444, w_022_445, w_022_446, w_022_447, w_022_448, w_022_449, w_022_450, w_022_451, w_022_452, w_022_453, w_022_454, w_022_455, w_022_456, w_022_457, w_022_458, w_022_459, w_022_460, w_022_461, w_022_462, w_022_463, w_022_464, w_022_465, w_022_466, w_022_467, w_022_468, w_022_469, w_022_470, w_022_471, w_022_472, w_022_473, w_022_474, w_022_475, w_022_476, w_022_477, w_022_478, w_022_479, w_022_480, w_022_481, w_022_482, w_022_483, w_022_484, w_022_485, w_022_486, w_022_488, w_022_489, w_022_490, w_022_491, w_022_492, w_022_494, w_022_495, w_022_496, w_022_498, w_022_499, w_022_500, w_022_501, w_022_502, w_022_503, w_022_504, w_022_505, w_022_506, w_022_507, w_022_508, w_022_509, w_022_511, w_022_512, w_022_513, w_022_514, w_022_517, w_022_518, w_022_519, w_022_522, w_022_523, w_022_524, w_022_525, w_022_526, w_022_528, w_022_529, w_022_530, w_022_531, w_022_532, w_022_533, w_022_534, w_022_535, w_022_536, w_022_537, w_022_539, w_022_540, w_022_541, w_022_542, w_022_543, w_022_544, w_022_546, w_022_547, w_022_548, w_022_549, w_022_550, w_022_551, w_022_553, w_022_554, w_022_555, w_022_556, w_022_557, w_022_558, w_022_559, w_022_560, w_022_561, w_022_562, w_022_563, w_022_564, w_022_565, w_022_566, w_022_567, w_022_568, w_022_569, w_022_570, w_022_572, w_022_573, w_022_574, w_022_575, w_022_576, w_022_577, w_022_579, w_022_580, w_022_582, w_022_583, w_022_584, w_022_585, w_022_586, w_022_587, w_022_588, w_022_589, w_022_590, w_022_591, w_022_592, w_022_594, w_022_595, w_022_596, w_022_597, w_022_598, w_022_599, w_022_600, w_022_602, w_022_603, w_022_604, w_022_605, w_022_606, w_022_607, w_022_608, w_022_609, w_022_610, w_022_611, w_022_612, w_022_613, w_022_614, w_022_615, w_022_616, w_022_617, w_022_618, w_022_619, w_022_620, w_022_621, w_022_622, w_022_623, w_022_624, w_022_625, w_022_626, w_022_627, w_022_628, w_022_629, w_022_630, w_022_631, w_022_632, w_022_633, w_022_634, w_022_635, w_022_637, w_022_638, w_022_639, w_022_640, w_022_641, w_022_642, w_022_644, w_022_645, w_022_646, w_022_648, w_022_649, w_022_650, w_022_652, w_022_653, w_022_654, w_022_655, w_022_656, w_022_657, w_022_658, w_022_659, w_022_660, w_022_661, w_022_662, w_022_663, w_022_664, w_022_665, w_022_666, w_022_667, w_022_668, w_022_669, w_022_670, w_022_671, w_022_672, w_022_673, w_022_674, w_022_676, w_022_677, w_022_678, w_022_679, w_022_680, w_022_681, w_022_684, w_022_685, w_022_686, w_022_687, w_022_688, w_022_689, w_022_690, w_022_691, w_022_692, w_022_693, w_022_694, w_022_695, w_022_696, w_022_697, w_022_698, w_022_699, w_022_700, w_022_701, w_022_702, w_022_703, w_022_704, w_022_705, w_022_706, w_022_708, w_022_709, w_022_710, w_022_711, w_022_712, w_022_713, w_022_714, w_022_715, w_022_716, w_022_717, w_022_718, w_022_719, w_022_720, w_022_721, w_022_722, w_022_723, w_022_724, w_022_725, w_022_726, w_022_728, w_022_729, w_022_730, w_022_731, w_022_732, w_022_733, w_022_734, w_022_735, w_022_738, w_022_740, w_022_741, w_022_742, w_022_743, w_022_745, w_022_746, w_022_747, w_022_748, w_022_749, w_022_751, w_022_752, w_022_753, w_022_755, w_022_756, w_022_757, w_022_758, w_022_759, w_022_760, w_022_761, w_022_762, w_022_763, w_022_764, w_022_765, w_022_766, w_022_767, w_022_768, w_022_769, w_022_770, w_022_771, w_022_772, w_022_773, w_022_774, w_022_776, w_022_777, w_022_778, w_022_779, w_022_780, w_022_781, w_022_782, w_022_783, w_022_784, w_022_785, w_022_786, w_022_787, w_022_788, w_022_789, w_022_790, w_022_791, w_022_792, w_022_793, w_022_794, w_022_795, w_022_796, w_022_797, w_022_798, w_022_799, w_022_801, w_022_802, w_022_803, w_022_804, w_022_805, w_022_806, w_022_807, w_022_808, w_022_809, w_022_812, w_022_813, w_022_814, w_022_815, w_022_817, w_022_818, w_022_820, w_022_821, w_022_822, w_022_823, w_022_824, w_022_825, w_022_826, w_022_827, w_022_828, w_022_829, w_022_830, w_022_831, w_022_832, w_022_833, w_022_834, w_022_835, w_022_836, w_022_838, w_022_839, w_022_840, w_022_841, w_022_842, w_022_845, w_022_846, w_022_847, w_022_848, w_022_849, w_022_850, w_022_851, w_022_852, w_022_853, w_022_854, w_022_855, w_022_856, w_022_857, w_022_858, w_022_859, w_022_860, w_022_861, w_022_862, w_022_863, w_022_864, w_022_866, w_022_867, w_022_870, w_022_871, w_022_872, w_022_873, w_022_874, w_022_875, w_022_876, w_022_877, w_022_878, w_022_879, w_022_880, w_022_881, w_022_882, w_022_883, w_022_884, w_022_885, w_022_886, w_022_887, w_022_888, w_022_889, w_022_890, w_022_891, w_022_892, w_022_893, w_022_894, w_022_895, w_022_896, w_022_897, w_022_898, w_022_899, w_022_900, w_022_901, w_022_902, w_022_903, w_022_904, w_022_905, w_022_906, w_022_907, w_022_908, w_022_909, w_022_910, w_022_911, w_022_912, w_022_913, w_022_914, w_022_915, w_022_916, w_022_917, w_022_918, w_022_919, w_022_920, w_022_921, w_022_922, w_022_923, w_022_924, w_022_925, w_022_926, w_022_927, w_022_928, w_022_929, w_022_931, w_022_932, w_022_933, w_022_934, w_022_935, w_022_936, w_022_937, w_022_938, w_022_939, w_022_941, w_022_942, w_022_943, w_022_944, w_022_945, w_022_946, w_022_947, w_022_948, w_022_949, w_022_950, w_022_951, w_022_952, w_022_953, w_022_954, w_022_955, w_022_956, w_022_957, w_022_958, w_022_959, w_022_960, w_022_961, w_022_962, w_022_963, w_022_964, w_022_965, w_022_966, w_022_967, w_022_970, w_022_971, w_022_972, w_022_975, w_022_976, w_022_977, w_022_978, w_022_979, w_022_982, w_022_984, w_022_985, w_022_986, w_022_987, w_022_988, w_022_989, w_022_990, w_022_991, w_022_992, w_022_993, w_022_994, w_022_995, w_022_996, w_022_997, w_022_998, w_022_999, w_022_1000, w_022_1001, w_022_1002, w_022_1003, w_022_1004, w_022_1005, w_022_1006, w_022_1007, w_022_1008, w_022_1009, w_022_1010, w_022_1014, w_022_1015, w_022_1016, w_022_1019, w_022_1020, w_022_1021, w_022_1022, w_022_1023, w_022_1024, w_022_1025, w_022_1026, w_022_1027, w_022_1028, w_022_1029, w_022_1030, w_022_1032, w_022_1033, w_022_1034, w_022_1038, w_022_1039, w_022_1040, w_022_1041, w_022_1042, w_022_1043, w_022_1044, w_022_1045, w_022_1046, w_022_1047, w_022_1048, w_022_1049, w_022_1050, w_022_1051, w_022_1052, w_022_1053, w_022_1054, w_022_1055, w_022_1056, w_022_1057, w_022_1058, w_022_1059, w_022_1060, w_022_1061, w_022_1062, w_022_1063, w_022_1064, w_022_1065, w_022_1066, w_022_1067, w_022_1068, w_022_1069, w_022_1070, w_022_1071, w_022_1072, w_022_1073, w_022_1074, w_022_1076, w_022_1077, w_022_1078, w_022_1079, w_022_1080, w_022_1081, w_022_1082, w_022_1083, w_022_1085, w_022_1086, w_022_1087, w_022_1088, w_022_1089, w_022_1090, w_022_1091, w_022_1092, w_022_1093, w_022_1094, w_022_1095, w_022_1096, w_022_1097, w_022_1098, w_022_1099, w_022_1100, w_022_1101, w_022_1103, w_022_1104, w_022_1105, w_022_1106, w_022_1107, w_022_1108, w_022_1109, w_022_1110, w_022_1111, w_022_1112, w_022_1113, w_022_1115, w_022_1116, w_022_1118, w_022_1119, w_022_1120, w_022_1122, w_022_1123, w_022_1124, w_022_1125, w_022_1126, w_022_1127, w_022_1128, w_022_1129, w_022_1130, w_022_1131, w_022_1132, w_022_1133, w_022_1135, w_022_1136, w_022_1138, w_022_1139, w_022_1140, w_022_1143, w_022_1144, w_022_1145, w_022_1146, w_022_1147, w_022_1148, w_022_1149, w_022_1150, w_022_1151, w_022_1152, w_022_1153, w_022_1154, w_022_1155, w_022_1156, w_022_1157, w_022_1159, w_022_1161, w_022_1162, w_022_1163, w_022_1164, w_022_1166, w_022_1167, w_022_1168, w_022_1170, w_022_1171, w_022_1172, w_022_1173, w_022_1174, w_022_1175, w_022_1176, w_022_1177, w_022_1178, w_022_1179, w_022_1180, w_022_1181, w_022_1182, w_022_1183, w_022_1184, w_022_1185, w_022_1186, w_022_1187, w_022_1188, w_022_1189, w_022_1190, w_022_1191, w_022_1192, w_022_1193, w_022_1194, w_022_1195, w_022_1196, w_022_1197, w_022_1198, w_022_1199, w_022_1200, w_022_1201, w_022_1203, w_022_1204, w_022_1205, w_022_1206, w_022_1207, w_022_1208, w_022_1209, w_022_1210, w_022_1211, w_022_1212, w_022_1213, w_022_1214, w_022_1215, w_022_1216, w_022_1217, w_022_1218, w_022_1219, w_022_1221, w_022_1222, w_022_1223, w_022_1224, w_022_1225, w_022_1227, w_022_1228, w_022_1229, w_022_1230, w_022_1231, w_022_1232, w_022_1233, w_022_1234, w_022_1236, w_022_1237, w_022_1238, w_022_1240, w_022_1241, w_022_1242, w_022_1243, w_022_1244, w_022_1245, w_022_1246, w_022_1247, w_022_1248, w_022_1249, w_022_1250, w_022_1251, w_022_1252, w_022_1253, w_022_1254, w_022_1256, w_022_1257, w_022_1258, w_022_1259, w_022_1260, w_022_1261, w_022_1262, w_022_1263, w_022_1264, w_022_1265, w_022_1266, w_022_1267, w_022_1268, w_022_1269, w_022_1270, w_022_1271, w_022_1272, w_022_1273, w_022_1274, w_022_1275, w_022_1276, w_022_1277, w_022_1278, w_022_1279, w_022_1281, w_022_1282, w_022_1283, w_022_1284, w_022_1285, w_022_1286, w_022_1287, w_022_1288, w_022_1289, w_022_1290, w_022_1292, w_022_1293, w_022_1294, w_022_1295, w_022_1296, w_022_1297, w_022_1298, w_022_1299, w_022_1300, w_022_1301, w_022_1302, w_022_1303, w_022_1304, w_022_1305, w_022_1306, w_022_1307, w_022_1308, w_022_1309, w_022_1311, w_022_1312, w_022_1313, w_022_1314, w_022_1315, w_022_1316, w_022_1317, w_022_1318, w_022_1319, w_022_1320, w_022_1321, w_022_1322, w_022_1323, w_022_1324, w_022_1325, w_022_1326, w_022_1327, w_022_1328, w_022_1329, w_022_1330, w_022_1331, w_022_1332, w_022_1333, w_022_1334, w_022_1335, w_022_1338, w_022_1339, w_022_1340, w_022_1341, w_022_1342, w_022_1343, w_022_1344, w_022_1345, w_022_1346, w_022_1347, w_022_1348, w_022_1349, w_022_1350, w_022_1351, w_022_1352, w_022_1353, w_022_1354, w_022_1357, w_022_1359, w_022_1360, w_022_1361, w_022_1362, w_022_1363, w_022_1364, w_022_1365, w_022_1366, w_022_1367, w_022_1368, w_022_1369, w_022_1370, w_022_1371, w_022_1372, w_022_1373, w_022_1374, w_022_1375, w_022_1376, w_022_1377, w_022_1378, w_022_1379, w_022_1380, w_022_1381, w_022_1382, w_022_1383, w_022_1384, w_022_1385, w_022_1386, w_022_1387, w_022_1388, w_022_1389, w_022_1390, w_022_1391, w_022_1392, w_022_1393, w_022_1394, w_022_1395, w_022_1396, w_022_1397, w_022_1398, w_022_1399, w_022_1400, w_022_1401, w_022_1402, w_022_1403, w_022_1404, w_022_1405, w_022_1406, w_022_1407, w_022_1408, w_022_1409, w_022_1410, w_022_1411, w_022_1412, w_022_1413, w_022_1414, w_022_1415, w_022_1416, w_022_1417, w_022_1418, w_022_1419, w_022_1420, w_022_1421, w_022_1422, w_022_1423, w_022_1424, w_022_1425, w_022_1426, w_022_1427, w_022_1428, w_022_1429, w_022_1431, w_022_1432, w_022_1433, w_022_1434, w_022_1435, w_022_1436, w_022_1437, w_022_1438, w_022_1439, w_022_1440, w_022_1441, w_022_1442, w_022_1443, w_022_1444, w_022_1445, w_022_1446, w_022_1447, w_022_1448, w_022_1449, w_022_1450, w_022_1451, w_022_1452, w_022_1453, w_022_1454, w_022_1455, w_022_1456, w_022_1457, w_022_1458, w_022_1459, w_022_1460, w_022_1461, w_022_1462, w_022_1463, w_022_1464, w_022_1466, w_022_1467, w_022_1468, w_022_1469, w_022_1470, w_022_1471, w_022_1472, w_022_1473, w_022_1474, w_022_1475, w_022_1476, w_022_1477, w_022_1478, w_022_1479, w_022_1480, w_022_1481, w_022_1482, w_022_1483, w_022_1484, w_022_1485, w_022_1486, w_022_1487, w_022_1488, w_022_1491, w_022_1492, w_022_1493, w_022_1494, w_022_1495, w_022_1496, w_022_1498, w_022_1499, w_022_1500, w_022_1501, w_022_1502, w_022_1503, w_022_1504, w_022_1505, w_022_1506, w_022_1508, w_022_1509, w_022_1510, w_022_1511, w_022_1512, w_022_1513, w_022_1514, w_022_1515, w_022_1516, w_022_1518, w_022_1520, w_022_1521, w_022_1522, w_022_1523, w_022_1524, w_022_1525, w_022_1526, w_022_1527, w_022_1528, w_022_1530, w_022_1531, w_022_1532, w_022_1534, w_022_1536, w_022_1538, w_022_1539, w_022_1540, w_022_1541, w_022_1542, w_022_1543, w_022_1544, w_022_1545, w_022_1546, w_022_1547, w_022_1548, w_022_1549, w_022_1550, w_022_1551, w_022_1552, w_022_1553, w_022_1555, w_022_1556, w_022_1558, w_022_1560, w_022_1561, w_022_1562, w_022_1564, w_022_1565, w_022_1566, w_022_1567, w_022_1568, w_022_1569, w_022_1570, w_022_1571, w_022_1572, w_022_1573, w_022_1574, w_022_1575, w_022_1576, w_022_1577, w_022_1578, w_022_1579, w_022_1580, w_022_1581, w_022_1582, w_022_1583, w_022_1584, w_022_1585, w_022_1586, w_022_1588, w_022_1589, w_022_1590, w_022_1591, w_022_1592, w_022_1593, w_022_1594, w_022_1595, w_022_1596, w_022_1597, w_022_1598, w_022_1600, w_022_1601, w_022_1602, w_022_1603, w_022_1604, w_022_1605, w_022_1606, w_022_1607, w_022_1608, w_022_1609, w_022_1610, w_022_1611, w_022_1612, w_022_1613, w_022_1614, w_022_1615, w_022_1616, w_022_1617, w_022_1618, w_022_1619, w_022_1620, w_022_1621, w_022_1622, w_022_1623, w_022_1624, w_022_1625, w_022_1626, w_022_1627, w_022_1628, w_022_1629, w_022_1630, w_022_1631, w_022_1632, w_022_1633, w_022_1634, w_022_1635, w_022_1636, w_022_1637, w_022_1638, w_022_1639, w_022_1640, w_022_1641, w_022_1642, w_022_1643, w_022_1644, w_022_1646, w_022_1647, w_022_1648, w_022_1649, w_022_1651, w_022_1652, w_022_1653, w_022_1654, w_022_1655, w_022_1656, w_022_1657, w_022_1659, w_022_1660, w_022_1661, w_022_1662, w_022_1663, w_022_1664, w_022_1665, w_022_1667, w_022_1669, w_022_1670, w_022_1671, w_022_1672, w_022_1673, w_022_1674, w_022_1675, w_022_1676, w_022_1677, w_022_1678, w_022_1679, w_022_1680, w_022_1681, w_022_1682, w_022_1683, w_022_1684, w_022_1685, w_022_1686, w_022_1687, w_022_1688, w_022_1689, w_022_1690, w_022_1691, w_022_1692, w_022_1693, w_022_1694, w_022_1695, w_022_1696, w_022_1697, w_022_1698, w_022_1699, w_022_1700, w_022_1701, w_022_1702, w_022_1703, w_022_1704, w_022_1705, w_022_1706, w_022_1707, w_022_1708, w_022_1710, w_022_1711, w_022_1712, w_022_1713, w_022_1714, w_022_1715, w_022_1716, w_022_1717, w_022_1718, w_022_1719, w_022_1720, w_022_1721, w_022_1722, w_022_1723, w_022_1724, w_022_1725, w_022_1726, w_022_1727, w_022_1728, w_022_1729, w_022_1730, w_022_1731, w_022_1732, w_022_1733, w_022_1734, w_022_1735, w_022_1736, w_022_1737, w_022_1738, w_022_1739, w_022_1740, w_022_1741, w_022_1742, w_022_1743, w_022_1744, w_022_1745, w_022_1746, w_022_1747, w_022_1748, w_022_1749, w_022_1750, w_022_1751, w_022_1752, w_022_1753, w_022_1754, w_022_1755, w_022_1756, w_022_1757, w_022_1758, w_022_1759, w_022_1760, w_022_1761, w_022_1762, w_022_1763, w_022_1764, w_022_1765, w_022_1766, w_022_1767, w_022_1768, w_022_1770, w_022_1771, w_022_1772, w_022_1773, w_022_1774, w_022_1775, w_022_1776, w_022_1778, w_022_1779, w_022_1780, w_022_1781, w_022_1782, w_022_1783, w_022_1784, w_022_1785, w_022_1786, w_022_1787, w_022_1788, w_022_1789, w_022_1790, w_022_1791, w_022_1792, w_022_1793, w_022_1794, w_022_1795, w_022_1796, w_022_1797, w_022_1798, w_022_1799, w_022_1801, w_022_1802, w_022_1803, w_022_1804, w_022_1805, w_022_1806, w_022_1807, w_022_1808, w_022_1809, w_022_1810, w_022_1811, w_022_1812, w_022_1813, w_022_1814, w_022_1815, w_022_1816, w_022_1817, w_022_1818, w_022_1819, w_022_1820, w_022_1821, w_022_1822, w_022_1823, w_022_1824, w_022_1825, w_022_1826, w_022_1827, w_022_1828, w_022_1829, w_022_1830, w_022_1831, w_022_1832, w_022_1833, w_022_1834, w_022_1835, w_022_1836, w_022_1837, w_022_1838, w_022_1839, w_022_1840, w_022_1841, w_022_1842, w_022_1843, w_022_1845, w_022_1846, w_022_1847, w_022_1848, w_022_1849, w_022_1850, w_022_1851, w_022_1852, w_022_1854, w_022_1855, w_022_1856, w_022_1857, w_022_1858, w_022_1859, w_022_1860, w_022_1861, w_022_1862, w_022_1863, w_022_1864, w_022_1865, w_022_1866, w_022_1867, w_022_1868, w_022_1869, w_022_1870, w_022_1871, w_022_1872, w_022_1873, w_022_1874, w_022_1875, w_022_1876, w_022_1877, w_022_1878, w_022_1879, w_022_1880, w_022_1881, w_022_1882, w_022_1883, w_022_1884, w_022_1885, w_022_1886, w_022_1888, w_022_1890, w_022_1891, w_022_1892, w_022_1893, w_022_1894, w_022_1895, w_022_1897, w_022_1899, w_022_1902, w_022_1903, w_022_1908, w_022_1910, w_022_1911, w_022_1913, w_022_1914, w_022_1915, w_022_1917, w_022_1920, w_022_1923, w_022_1924, w_022_1925, w_022_1926, w_022_1927, w_022_1928, w_022_1929, w_022_1930, w_022_1931, w_022_1932, w_022_1935, w_022_1936, w_022_1937, w_022_1938, w_022_1939, w_022_1940, w_022_1941, w_022_1944, w_022_1945, w_022_1946, w_022_1948, w_022_1951, w_022_1953, w_022_1954, w_022_1956, w_022_1958, w_022_1960, w_022_1961, w_022_1962, w_022_1963, w_022_1964, w_022_1965, w_022_1966, w_022_1967, w_022_1969, w_022_1970, w_022_1971, w_022_1974, w_022_1975, w_022_1976, w_022_1977, w_022_1978, w_022_1979, w_022_1980, w_022_1981, w_022_1982, w_022_1983, w_022_1985, w_022_1986, w_022_1987, w_022_1988, w_022_1989, w_022_1990, w_022_1992, w_022_1993, w_022_1994, w_022_1996, w_022_1998, w_022_1999, w_022_2000, w_022_2001, w_022_2002, w_022_2003, w_022_2004, w_022_2005, w_022_2006, w_022_2007, w_022_2009, w_022_2010, w_022_2012, w_022_2013, w_022_2015, w_022_2016, w_022_2018, w_022_2019, w_022_2020, w_022_2021, w_022_2022, w_022_2023, w_022_2024, w_022_2025, w_022_2026, w_022_2027, w_022_2029, w_022_2031, w_022_2033, w_022_2034, w_022_2035, w_022_2036, w_022_2037, w_022_2038, w_022_2040, w_022_2044, w_022_2045, w_022_2046, w_022_2048, w_022_2049, w_022_2050, w_022_2051, w_022_2052, w_022_2054, w_022_2055, w_022_2056, w_022_2057, w_022_2058, w_022_2060, w_022_2063, w_022_2064, w_022_2065, w_022_2067, w_022_2070, w_022_2071, w_022_2072, w_022_2073, w_022_2074, w_022_2075, w_022_2076, w_022_2077, w_022_2078, w_022_2079, w_022_2080, w_022_2084, w_022_2085, w_022_2086, w_022_2087, w_022_2089, w_022_2091, w_022_2093, w_022_2094, w_022_2095, w_022_2096, w_022_2098, w_022_2099, w_022_2102, w_022_2103, w_022_2104, w_022_2105, w_022_2107, w_022_2109, w_022_2110, w_022_2114, w_022_2116, w_022_2117, w_022_2120, w_022_2121, w_022_2122, w_022_2123, w_022_2124, w_022_2127, w_022_2128, w_022_2129, w_022_2130, w_022_2131, w_022_2132, w_022_2133, w_022_2134, w_022_2138, w_022_2139, w_022_2140, w_022_2141, w_022_2142, w_022_2143, w_022_2144, w_022_2145, w_022_2146, w_022_2147, w_022_2148, w_022_2149, w_022_2150, w_022_2151, w_022_2152, w_022_2153, w_022_2154, w_022_2155, w_022_2156, w_022_2157, w_022_2158, w_022_2159, w_022_2160, w_022_2163, w_022_2164, w_022_2167, w_022_2168, w_022_2169, w_022_2170, w_022_2171, w_022_2172, w_022_2174, w_022_2176, w_022_2177, w_022_2178, w_022_2180, w_022_2181, w_022_2182, w_022_2183, w_022_2184, w_022_2185, w_022_2186, w_022_2190, w_022_2191, w_022_2192, w_022_2193, w_022_2194, w_022_2195, w_022_2198, w_022_2199, w_022_2200, w_022_2201, w_022_2202, w_022_2204, w_022_2205, w_022_2206, w_022_2209, w_022_2210, w_022_2211, w_022_2212, w_022_2216, w_022_2218, w_022_2221, w_022_2222, w_022_2224, w_022_2225, w_022_2226, w_022_2227, w_022_2228, w_022_2230, w_022_2231, w_022_2232, w_022_2233, w_022_2234, w_022_2235, w_022_2236, w_022_2237, w_022_2238, w_022_2241, w_022_2243, w_022_2244, w_022_2246, w_022_2251, w_022_2253, w_022_2254, w_022_2257, w_022_2258, w_022_2259, w_022_2260, w_022_2261, w_022_2262, w_022_2264, w_022_2265, w_022_2266, w_022_2267, w_022_2268, w_022_2269, w_022_2270, w_022_2271, w_022_2273, w_022_2274, w_022_2275, w_022_2276, w_022_2277, w_022_2279, w_022_2280, w_022_2281, w_022_2282, w_022_2284, w_022_2285, w_022_2287, w_022_2288, w_022_2289, w_022_2290, w_022_2291, w_022_2292, w_022_2293, w_022_2294, w_022_2296, w_022_2299, w_022_2301, w_022_2302, w_022_2303, w_022_2305, w_022_2306, w_022_2307, w_022_2308, w_022_2309, w_022_2310, w_022_2311, w_022_2312, w_022_2315, w_022_2316, w_022_2319, w_022_2320, w_022_2322, w_022_2324, w_022_2326, w_022_2328, w_022_2329, w_022_2330, w_022_2332, w_022_2334, w_022_2335, w_022_2336, w_022_2339, w_022_2341, w_022_2343, w_022_2344, w_022_2346, w_022_2347, w_022_2348, w_022_2350, w_022_2352, w_022_2355, w_022_2356, w_022_2358, w_022_2359, w_022_2362, w_022_2363, w_022_2364, w_022_2365, w_022_2366, w_022_2367, w_022_2369, w_022_2371, w_022_2372, w_022_2373, w_022_2375, w_022_2376, w_022_2377, w_022_2379, w_022_2380, w_022_2381, w_022_2382, w_022_2383, w_022_2384, w_022_2385, w_022_2386, w_022_2388, w_022_2389, w_022_2390, w_022_2391, w_022_2392, w_022_2393, w_022_2394, w_022_2395, w_022_2396, w_022_2397, w_022_2398, w_022_2400, w_022_2402, w_022_2403, w_022_2408, w_022_2409, w_022_2413, w_022_2414, w_022_2415, w_022_2416, w_022_2417, w_022_2418, w_022_2419, w_022_2421, w_022_2422, w_022_2423, w_022_2426, w_022_2427, w_022_2429, w_022_2431, w_022_2436, w_022_2438, w_022_2441, w_022_2442, w_022_2444, w_022_2445, w_022_2447, w_022_2448, w_022_2449, w_022_2450, w_022_2452, w_022_2454, w_022_2457, w_022_2459, w_022_2460, w_022_2461, w_022_2463, w_022_2464, w_022_2466, w_022_2468, w_022_2471, w_022_2472, w_022_2473, w_022_2474, w_022_2476, w_022_2479, w_022_2480, w_022_2481, w_022_2483, w_022_2485, w_022_2489, w_022_2490, w_022_2491, w_022_2493, w_022_2494, w_022_2495, w_022_2496, w_022_2499, w_022_2500, w_022_2501, w_022_2503, w_022_2506, w_022_2507, w_022_2508, w_022_2509, w_022_2510, w_022_2511, w_022_2512, w_022_2514, w_022_2518, w_022_2519, w_022_2520, w_022_2521, w_022_2522, w_022_2524, w_022_2526, w_022_2527, w_022_2528, w_022_2532, w_022_2533, w_022_2534, w_022_2535, w_022_2536, w_022_2537, w_022_2538, w_022_2539, w_022_2542, w_022_2543, w_022_2544, w_022_2545, w_022_2546, w_022_2547, w_022_2548, w_022_2549, w_022_2551, w_022_2553, w_022_2554, w_022_2555, w_022_2556, w_022_2557, w_022_2558, w_022_2559, w_022_2560, w_022_2561, w_022_2562, w_022_2563, w_022_2566, w_022_2567, w_022_2568, w_022_2570, w_022_2571, w_022_2572, w_022_2573, w_022_2575, w_022_2576, w_022_2578, w_022_2579, w_022_2580, w_022_2581, w_022_2583, w_022_2584, w_022_2585, w_022_2586, w_022_2587, w_022_2588, w_022_2589, w_022_2590, w_022_2592, w_022_2593, w_022_2595, w_022_2596, w_022_2597, w_022_2598, w_022_2600, w_022_2601, w_022_2602, w_022_2603, w_022_2605, w_022_2606, w_022_2608, w_022_2609, w_022_2610, w_022_2611, w_022_2612, w_022_2613, w_022_2615, w_022_2616, w_022_2617, w_022_2620, w_022_2621, w_022_2623, w_022_2624, w_022_2625, w_022_2626, w_022_2628, w_022_2631, w_022_2632, w_022_2633, w_022_2634, w_022_2635, w_022_2636, w_022_2637, w_022_2639, w_022_2640, w_022_2644, w_022_2645, w_022_2646, w_022_2648, w_022_2649, w_022_2652, w_022_2653, w_022_2654, w_022_2655, w_022_2656, w_022_2657, w_022_2658, w_022_2660, w_022_2661, w_022_2662, w_022_2663, w_022_2665, w_022_2669, w_022_2671, w_022_2672, w_022_2673, w_022_2675, w_022_2676, w_022_2677, w_022_2678, w_022_2679, w_022_2680, w_022_2681, w_022_2682, w_022_2684, w_022_2686, w_022_2688, w_022_2689, w_022_2691, w_022_2692, w_022_2694, w_022_2695, w_022_2696, w_022_2697, w_022_2700, w_022_2701, w_022_2702, w_022_2704, w_022_2707, w_022_2708, w_022_2710, w_022_2711, w_022_2713, w_022_2714, w_022_2715, w_022_2716, w_022_2717, w_022_2718, w_022_2719, w_022_2721, w_022_2722, w_022_2725, w_022_2728, w_022_2729, w_022_2730, w_022_2731, w_022_2732, w_022_2733, w_022_2734, w_022_2735, w_022_2736, w_022_2737, w_022_2738, w_022_2740, w_022_2741, w_022_2742, w_022_2743, w_022_2744, w_022_2745, w_022_2746, w_022_2748, w_022_2751, w_022_2754, w_022_2755, w_022_2756, w_022_2760, w_022_2761, w_022_2762, w_022_2763, w_022_2765, w_022_2768, w_022_2769, w_022_2772, w_022_2773, w_022_2774, w_022_2775, w_022_2776, w_022_2777, w_022_2781, w_022_2782, w_022_2783, w_022_2784, w_022_2785, w_022_2786, w_022_2787, w_022_2788, w_022_2789, w_022_2790, w_022_2791, w_022_2792, w_022_2793, w_022_2795, w_022_2796, w_022_2798, w_022_2799, w_022_2800, w_022_2801, w_022_2803, w_022_2805, w_022_2806, w_022_2807, w_022_2808, w_022_2809, w_022_2810, w_022_2812, w_022_2815, w_022_2816, w_022_2822, w_022_2823, w_022_2825, w_022_2826, w_022_2828, w_022_2830, w_022_2832, w_022_2833, w_022_2834, w_022_2835, w_022_2838, w_022_2840, w_022_2842, w_022_2843, w_022_2844, w_022_2845, w_022_2846, w_022_2847, w_022_2850, w_022_2851, w_022_2852, w_022_2854, w_022_2855, w_022_2856, w_022_2857, w_022_2858, w_022_2859, w_022_2860, w_022_2861, w_022_2862, w_022_2863, w_022_2864, w_022_2865, w_022_2866, w_022_2869, w_022_2872, w_022_2876, w_022_2877, w_022_2878, w_022_2879, w_022_2880, w_022_2882, w_022_2883, w_022_2885, w_022_2886, w_022_2887, w_022_2893, w_022_2894, w_022_2895, w_022_2896, w_022_2897, w_022_2898, w_022_2899, w_022_2900, w_022_2901, w_022_2902, w_022_2903, w_022_2904, w_022_2905, w_022_2907, w_022_2909, w_022_2911, w_022_2914, w_022_2915, w_022_2916, w_022_2917, w_022_2918, w_022_2919, w_022_2920, w_022_2922, w_022_2923, w_022_2924, w_022_2925, w_022_2927, w_022_2928, w_022_2929, w_022_2930, w_022_2933, w_022_2934, w_022_2935, w_022_2936, w_022_2937, w_022_2939, w_022_2941, w_022_2942, w_022_2943, w_022_2946, w_022_2947, w_022_2949, w_022_2950, w_022_2951, w_022_2954, w_022_2955, w_022_2956, w_022_2957, w_022_2959, w_022_2961, w_022_2962, w_022_2963, w_022_2966, w_022_2967, w_022_2968, w_022_2969, w_022_2971, w_022_2973, w_022_2974, w_022_2975, w_022_2980, w_022_2981, w_022_2982, w_022_2984, w_022_2986, w_022_2990, w_022_2991, w_022_2992, w_022_2993, w_022_2995, w_022_2998, w_022_3001, w_022_3003, w_022_3004, w_022_3005, w_022_3006, w_022_3007, w_022_3010, w_022_3012, w_022_3014, w_022_3015, w_022_3016, w_022_3017, w_022_3019, w_022_3020, w_022_3021, w_022_3022, w_022_3024, w_022_3025, w_022_3026, w_022_3027, w_022_3028, w_022_3029, w_022_3030, w_022_3034, w_022_3035, w_022_3036, w_022_3039, w_022_3040, w_022_3044, w_022_3045, w_022_3046, w_022_3048, w_022_3049, w_022_3050, w_022_3051, w_022_3052, w_022_3053, w_022_3055, w_022_3056, w_022_3057, w_022_3059, w_022_3060, w_022_3061, w_022_3062, w_022_3064, w_022_3065, w_022_3066, w_022_3067, w_022_3068, w_022_3069, w_022_3071, w_022_3072, w_022_3073, w_022_3074, w_022_3075, w_022_3077, w_022_3078, w_022_3079, w_022_3082, w_022_3085, w_022_3087, w_022_3088, w_022_3089, w_022_3090, w_022_3092, w_022_3094, w_022_3097, w_022_3098, w_022_3099, w_022_3101, w_022_3102, w_022_3103, w_022_3104;
  wire w_023_000, w_023_001, w_023_002, w_023_003, w_023_004, w_023_005, w_023_006, w_023_007, w_023_008, w_023_009, w_023_010, w_023_011, w_023_012, w_023_013, w_023_014, w_023_015, w_023_016, w_023_017, w_023_018, w_023_019, w_023_020, w_023_021, w_023_022, w_023_023, w_023_024, w_023_025, w_023_026, w_023_027, w_023_028, w_023_029, w_023_030, w_023_031, w_023_032, w_023_033, w_023_034, w_023_035, w_023_036, w_023_037, w_023_038, w_023_039, w_023_040, w_023_041, w_023_042, w_023_043, w_023_044, w_023_045, w_023_046, w_023_047, w_023_048, w_023_049, w_023_050, w_023_051, w_023_052, w_023_053, w_023_054, w_023_055, w_023_056, w_023_057, w_023_058, w_023_059, w_023_060, w_023_061, w_023_062, w_023_063, w_023_064, w_023_065, w_023_066, w_023_067, w_023_068, w_023_069, w_023_070, w_023_071, w_023_072, w_023_073, w_023_074, w_023_075, w_023_076, w_023_077, w_023_078, w_023_079, w_023_080, w_023_081, w_023_082, w_023_083, w_023_084, w_023_085, w_023_086, w_023_087, w_023_088, w_023_089, w_023_090, w_023_091, w_023_092, w_023_093, w_023_094, w_023_095, w_023_096, w_023_097, w_023_098, w_023_099, w_023_100, w_023_101, w_023_102, w_023_103, w_023_104, w_023_105, w_023_106, w_023_107, w_023_108, w_023_109, w_023_110, w_023_111, w_023_112, w_023_113, w_023_114, w_023_115, w_023_116, w_023_117, w_023_118, w_023_119, w_023_120, w_023_121, w_023_122, w_023_123, w_023_124, w_023_125, w_023_126, w_023_127, w_023_128, w_023_129, w_023_130, w_023_131, w_023_132, w_023_133, w_023_134, w_023_135, w_023_136, w_023_137, w_023_138, w_023_139, w_023_140, w_023_141, w_023_142, w_023_143, w_023_144, w_023_145, w_023_146, w_023_147, w_023_148, w_023_149, w_023_150, w_023_151, w_023_152, w_023_153, w_023_154, w_023_155, w_023_156, w_023_157, w_023_158, w_023_159, w_023_160, w_023_161, w_023_162, w_023_163, w_023_164, w_023_165, w_023_166, w_023_167, w_023_168, w_023_169, w_023_170, w_023_171, w_023_172, w_023_173, w_023_174, w_023_175, w_023_176, w_023_177, w_023_178, w_023_179, w_023_180, w_023_181, w_023_182, w_023_183, w_023_184, w_023_185, w_023_186, w_023_187, w_023_188, w_023_189, w_023_190, w_023_191, w_023_192, w_023_193, w_023_194, w_023_195, w_023_196, w_023_197, w_023_198, w_023_199, w_023_200, w_023_201, w_023_202, w_023_203, w_023_204, w_023_205, w_023_206, w_023_207, w_023_208, w_023_209, w_023_210, w_023_211, w_023_212, w_023_213, w_023_214, w_023_215, w_023_216, w_023_217, w_023_218, w_023_219, w_023_220, w_023_221, w_023_222, w_023_223, w_023_224, w_023_225, w_023_226, w_023_227, w_023_228, w_023_229, w_023_230, w_023_231, w_023_232, w_023_233, w_023_234, w_023_235, w_023_236, w_023_237, w_023_238, w_023_239, w_023_240, w_023_241, w_023_242, w_023_243, w_023_244, w_023_245, w_023_246, w_023_247, w_023_248, w_023_249, w_023_250, w_023_251, w_023_252, w_023_253, w_023_254, w_023_255, w_023_256, w_023_257, w_023_258, w_023_259, w_023_260, w_023_261, w_023_262, w_023_263, w_023_264, w_023_265, w_023_266, w_023_267, w_023_268, w_023_269, w_023_270, w_023_271, w_023_272, w_023_273, w_023_274, w_023_275, w_023_276, w_023_277, w_023_278, w_023_279, w_023_280, w_023_281, w_023_282, w_023_283, w_023_284, w_023_285, w_023_286, w_023_287, w_023_288, w_023_289, w_023_290, w_023_291, w_023_292, w_023_293, w_023_294, w_023_295, w_023_296, w_023_297, w_023_298, w_023_299, w_023_300, w_023_301, w_023_302, w_023_303, w_023_304, w_023_305, w_023_306, w_023_307, w_023_308, w_023_309, w_023_310, w_023_311, w_023_312, w_023_313, w_023_314, w_023_315, w_023_316, w_023_317, w_023_318, w_023_319, w_023_320, w_023_321, w_023_322, w_023_323, w_023_324, w_023_325, w_023_326, w_023_327, w_023_328, w_023_329, w_023_330, w_023_331, w_023_332, w_023_333, w_023_334, w_023_335, w_023_336, w_023_337, w_023_338, w_023_339, w_023_340, w_023_341, w_023_342, w_023_343, w_023_344, w_023_345, w_023_346, w_023_347, w_023_348, w_023_349, w_023_350, w_023_351, w_023_352, w_023_353, w_023_354, w_023_355, w_023_356, w_023_357, w_023_358, w_023_359, w_023_360, w_023_361, w_023_362, w_023_363, w_023_364, w_023_365, w_023_366, w_023_367, w_023_368, w_023_369, w_023_370, w_023_371, w_023_372, w_023_373, w_023_374, w_023_375, w_023_376, w_023_377, w_023_378, w_023_379, w_023_380, w_023_381, w_023_382, w_023_383, w_023_384, w_023_385, w_023_386, w_023_387, w_023_388, w_023_389, w_023_390, w_023_391, w_023_392, w_023_393, w_023_394, w_023_395, w_023_396, w_023_397, w_023_398, w_023_399, w_023_400, w_023_401, w_023_402, w_023_403, w_023_404, w_023_405, w_023_406, w_023_407, w_023_408, w_023_409, w_023_410, w_023_411, w_023_412, w_023_413, w_023_414, w_023_415, w_023_416, w_023_417, w_023_418, w_023_419, w_023_420, w_023_421, w_023_422, w_023_423, w_023_424, w_023_425, w_023_426, w_023_427, w_023_428, w_023_429, w_023_430, w_023_431, w_023_432, w_023_433, w_023_434, w_023_435, w_023_436, w_023_437, w_023_438, w_023_439, w_023_440, w_023_441, w_023_442, w_023_443, w_023_444, w_023_445, w_023_446, w_023_447, w_023_448, w_023_449, w_023_450, w_023_451, w_023_452, w_023_453, w_023_454, w_023_455, w_023_456, w_023_457, w_023_458, w_023_459, w_023_460, w_023_461, w_023_462, w_023_463, w_023_464, w_023_465, w_023_466, w_023_467, w_023_468, w_023_469, w_023_470, w_023_471, w_023_472, w_023_473, w_023_474, w_023_475, w_023_476, w_023_477, w_023_478, w_023_479, w_023_480, w_023_481, w_023_482, w_023_483, w_023_484, w_023_485, w_023_486, w_023_487, w_023_488, w_023_489, w_023_490, w_023_491, w_023_492, w_023_493, w_023_494, w_023_495, w_023_496, w_023_497, w_023_498, w_023_499, w_023_500, w_023_501, w_023_502, w_023_503, w_023_504, w_023_505, w_023_506, w_023_507, w_023_508, w_023_509, w_023_510, w_023_511, w_023_512, w_023_513, w_023_514, w_023_515, w_023_516, w_023_517, w_023_518, w_023_519, w_023_520, w_023_521, w_023_522, w_023_523, w_023_524, w_023_525, w_023_526, w_023_527, w_023_528, w_023_529, w_023_530, w_023_531, w_023_532, w_023_533, w_023_534, w_023_535, w_023_536, w_023_537, w_023_538, w_023_539, w_023_540, w_023_541, w_023_542, w_023_543, w_023_544, w_023_545, w_023_546, w_023_547, w_023_548, w_023_549, w_023_550, w_023_551, w_023_552, w_023_553, w_023_554, w_023_555, w_023_556, w_023_557, w_023_558, w_023_559, w_023_560, w_023_561, w_023_562, w_023_563, w_023_564, w_023_565, w_023_566, w_023_567, w_023_568, w_023_569, w_023_570, w_023_571, w_023_572, w_023_573, w_023_574, w_023_575, w_023_576, w_023_577, w_023_578, w_023_579, w_023_580, w_023_581, w_023_583, w_023_584, w_023_585, w_023_586, w_023_587, w_023_588, w_023_589, w_023_591;
  wire w_024_000, w_024_001, w_024_002, w_024_005, w_024_006, w_024_007, w_024_008, w_024_010, w_024_011, w_024_012, w_024_013, w_024_014, w_024_015, w_024_016, w_024_017, w_024_018, w_024_019, w_024_020, w_024_021, w_024_022, w_024_023, w_024_024, w_024_025, w_024_026, w_024_027, w_024_028, w_024_030, w_024_031, w_024_032, w_024_033, w_024_034, w_024_035, w_024_037, w_024_038, w_024_039, w_024_040, w_024_041, w_024_043, w_024_044, w_024_045, w_024_046, w_024_047, w_024_048, w_024_049, w_024_050, w_024_051, w_024_052, w_024_053, w_024_054, w_024_055, w_024_056, w_024_057, w_024_058, w_024_059, w_024_060, w_024_061, w_024_063, w_024_064, w_024_065, w_024_066, w_024_067, w_024_068, w_024_069, w_024_070, w_024_071, w_024_072, w_024_073, w_024_074, w_024_075, w_024_077, w_024_078, w_024_079, w_024_080, w_024_081, w_024_082, w_024_083, w_024_084, w_024_085, w_024_087, w_024_088, w_024_089, w_024_090, w_024_091, w_024_092, w_024_093, w_024_094, w_024_095, w_024_096, w_024_097, w_024_099, w_024_101, w_024_102, w_024_103, w_024_104, w_024_105, w_024_106, w_024_107, w_024_108, w_024_109, w_024_111, w_024_112, w_024_113, w_024_115, w_024_116, w_024_117, w_024_118, w_024_119, w_024_120, w_024_122, w_024_123, w_024_124, w_024_125, w_024_126, w_024_127, w_024_128, w_024_129, w_024_130, w_024_131, w_024_132, w_024_133, w_024_135, w_024_136, w_024_137, w_024_138, w_024_139, w_024_140, w_024_141, w_024_142, w_024_143, w_024_144, w_024_145, w_024_146, w_024_147, w_024_148, w_024_149, w_024_150, w_024_151, w_024_152, w_024_153, w_024_154, w_024_155, w_024_156, w_024_157, w_024_158, w_024_159, w_024_160, w_024_161, w_024_162, w_024_163, w_024_164, w_024_165, w_024_166, w_024_167, w_024_169, w_024_170, w_024_171, w_024_172, w_024_173, w_024_174, w_024_175, w_024_176, w_024_177, w_024_178, w_024_179, w_024_180, w_024_181, w_024_182, w_024_183, w_024_184, w_024_185, w_024_186, w_024_187, w_024_188, w_024_189, w_024_190, w_024_191, w_024_193, w_024_194, w_024_195, w_024_196, w_024_197, w_024_198, w_024_199, w_024_200, w_024_201, w_024_202, w_024_203, w_024_205, w_024_206, w_024_207, w_024_208, w_024_209, w_024_210, w_024_211, w_024_212, w_024_213, w_024_214, w_024_215, w_024_216, w_024_217, w_024_218, w_024_219, w_024_220, w_024_222, w_024_223, w_024_224, w_024_225, w_024_226, w_024_227, w_024_229, w_024_230, w_024_231, w_024_232, w_024_233, w_024_234, w_024_235, w_024_236, w_024_237, w_024_238, w_024_239, w_024_240, w_024_241, w_024_242, w_024_243, w_024_244, w_024_245, w_024_246, w_024_247, w_024_248, w_024_249, w_024_250, w_024_251, w_024_252, w_024_253, w_024_254, w_024_255, w_024_256, w_024_257, w_024_258, w_024_259, w_024_260, w_024_261, w_024_262, w_024_263, w_024_265, w_024_266, w_024_267, w_024_268, w_024_269, w_024_270, w_024_271, w_024_272, w_024_273, w_024_274, w_024_275, w_024_276, w_024_277, w_024_278, w_024_279, w_024_280, w_024_281, w_024_282, w_024_283, w_024_284, w_024_285, w_024_286, w_024_288, w_024_290, w_024_291, w_024_292, w_024_293, w_024_294, w_024_296, w_024_297, w_024_298, w_024_299, w_024_300, w_024_301, w_024_303, w_024_305, w_024_306, w_024_308, w_024_309, w_024_310, w_024_313, w_024_314, w_024_315, w_024_318, w_024_320, w_024_321, w_024_322, w_024_323, w_024_324, w_024_325, w_024_326, w_024_327, w_024_328, w_024_329, w_024_330, w_024_331, w_024_334, w_024_335, w_024_337, w_024_338, w_024_340, w_024_341, w_024_342, w_024_344, w_024_345, w_024_348, w_024_349, w_024_350, w_024_351, w_024_352, w_024_354, w_024_356, w_024_357, w_024_359, w_024_360, w_024_362, w_024_363, w_024_364, w_024_365, w_024_366, w_024_367, w_024_369, w_024_371, w_024_372, w_024_373, w_024_374, w_024_375, w_024_376, w_024_380, w_024_382, w_024_383, w_024_384, w_024_385, w_024_386, w_024_388, w_024_390, w_024_391, w_024_392, w_024_393, w_024_394, w_024_397, w_024_398, w_024_399, w_024_400, w_024_402, w_024_403, w_024_405, w_024_406, w_024_409, w_024_414, w_024_415, w_024_416, w_024_418, w_024_421, w_024_422, w_024_423, w_024_424, w_024_427, w_024_428, w_024_430, w_024_431, w_024_433, w_024_434, w_024_435, w_024_436, w_024_437, w_024_438, w_024_439, w_024_440, w_024_442, w_024_443, w_024_445, w_024_446, w_024_447, w_024_448, w_024_452, w_024_453, w_024_455, w_024_457, w_024_459, w_024_460, w_024_462, w_024_463, w_024_464, w_024_465, w_024_466, w_024_467, w_024_470, w_024_471, w_024_472, w_024_474, w_024_475, w_024_476, w_024_478, w_024_479, w_024_480, w_024_481, w_024_482, w_024_485, w_024_486, w_024_487, w_024_488, w_024_489, w_024_490, w_024_492, w_024_495, w_024_496, w_024_499, w_024_500, w_024_501, w_024_503, w_024_506, w_024_507, w_024_508, w_024_510, w_024_511, w_024_513, w_024_515, w_024_516, w_024_517, w_024_518, w_024_519, w_024_520, w_024_521, w_024_522, w_024_523, w_024_524, w_024_525, w_024_526, w_024_529, w_024_531, w_024_532, w_024_534, w_024_535, w_024_537, w_024_538, w_024_539, w_024_541, w_024_542, w_024_543, w_024_544, w_024_545, w_024_547, w_024_550, w_024_551, w_024_553, w_024_555, w_024_556, w_024_559, w_024_562, w_024_563, w_024_567, w_024_568, w_024_571, w_024_572, w_024_574, w_024_575, w_024_577, w_024_578, w_024_579, w_024_580, w_024_581, w_024_582, w_024_585, w_024_586, w_024_590, w_024_591, w_024_592, w_024_593, w_024_594, w_024_596, w_024_597, w_024_603, w_024_604, w_024_607, w_024_608, w_024_609, w_024_610, w_024_612, w_024_613, w_024_615, w_024_616, w_024_618, w_024_619, w_024_622, w_024_625, w_024_626, w_024_627, w_024_630, w_024_631, w_024_632, w_024_634, w_024_635, w_024_638, w_024_639, w_024_640, w_024_645, w_024_646, w_024_648, w_024_650, w_024_651, w_024_652, w_024_655, w_024_657, w_024_661, w_024_662, w_024_663, w_024_664, w_024_665, w_024_668, w_024_670, w_024_671, w_024_672, w_024_674, w_024_675, w_024_676, w_024_677, w_024_678, w_024_679, w_024_680, w_024_682, w_024_683, w_024_684, w_024_685, w_024_686, w_024_687, w_024_688, w_024_689, w_024_691, w_024_692, w_024_693, w_024_694, w_024_697, w_024_698, w_024_699, w_024_700, w_024_701, w_024_702, w_024_703, w_024_704, w_024_705, w_024_706, w_024_707, w_024_708, w_024_710, w_024_711, w_024_712, w_024_713, w_024_715, w_024_716, w_024_717, w_024_719, w_024_720, w_024_722, w_024_724, w_024_725, w_024_727, w_024_729, w_024_730, w_024_733, w_024_734, w_024_736, w_024_738, w_024_739, w_024_740, w_024_741, w_024_742, w_024_743, w_024_744, w_024_745, w_024_748, w_024_749, w_024_750, w_024_751, w_024_753, w_024_754, w_024_756, w_024_757, w_024_759, w_024_762, w_024_764, w_024_765, w_024_768, w_024_770, w_024_771, w_024_772, w_024_773, w_024_774, w_024_775, w_024_776, w_024_778, w_024_779, w_024_781, w_024_782, w_024_783, w_024_785, w_024_788, w_024_790, w_024_791, w_024_793, w_024_794, w_024_797, w_024_798, w_024_799, w_024_800, w_024_801, w_024_804, w_024_806, w_024_807, w_024_808, w_024_809, w_024_810, w_024_811, w_024_814, w_024_816, w_024_817, w_024_818, w_024_819, w_024_820, w_024_821, w_024_822, w_024_823, w_024_825, w_024_826, w_024_828, w_024_829, w_024_830, w_024_831, w_024_833, w_024_835, w_024_837, w_024_840, w_024_841, w_024_842, w_024_845, w_024_846, w_024_847, w_024_848, w_024_851, w_024_852, w_024_853, w_024_855, w_024_857, w_024_860, w_024_862, w_024_863, w_024_865, w_024_866, w_024_867, w_024_868, w_024_869, w_024_870, w_024_871, w_024_872, w_024_873, w_024_875, w_024_876, w_024_877, w_024_878, w_024_879, w_024_880, w_024_881, w_024_882, w_024_884, w_024_885, w_024_886, w_024_888, w_024_889, w_024_890, w_024_891, w_024_893, w_024_896, w_024_898, w_024_899, w_024_901, w_024_902, w_024_903, w_024_904, w_024_905, w_024_907, w_024_908, w_024_909, w_024_910, w_024_913, w_024_914, w_024_917, w_024_919, w_024_920, w_024_921, w_024_922, w_024_923, w_024_924, w_024_927, w_024_929, w_024_930, w_024_933, w_024_934, w_024_935, w_024_938, w_024_940, w_024_943, w_024_944, w_024_945, w_024_946, w_024_948, w_024_950, w_024_954, w_024_956, w_024_957, w_024_958, w_024_959, w_024_961, w_024_962, w_024_964, w_024_965, w_024_966, w_024_968, w_024_969, w_024_971, w_024_972, w_024_973, w_024_974, w_024_977, w_024_978, w_024_979, w_024_980, w_024_982, w_024_983, w_024_984, w_024_985, w_024_986, w_024_987, w_024_989, w_024_990, w_024_991, w_024_994, w_024_995, w_024_996, w_024_997, w_024_998, w_024_999, w_024_1000, w_024_1001, w_024_1002, w_024_1003, w_024_1005, w_024_1008, w_024_1009, w_024_1010, w_024_1012, w_024_1013, w_024_1014, w_024_1015, w_024_1016, w_024_1018, w_024_1020, w_024_1022, w_024_1023, w_024_1024, w_024_1025, w_024_1028, w_024_1031, w_024_1034, w_024_1036, w_024_1038, w_024_1040, w_024_1041, w_024_1042, w_024_1043, w_024_1045, w_024_1048, w_024_1049, w_024_1050, w_024_1051, w_024_1052, w_024_1053, w_024_1055, w_024_1056, w_024_1057, w_024_1058, w_024_1060, w_024_1062, w_024_1063, w_024_1064, w_024_1065, w_024_1067, w_024_1069, w_024_1071, w_024_1072, w_024_1074, w_024_1075, w_024_1076, w_024_1077, w_024_1078, w_024_1079, w_024_1080, w_024_1081, w_024_1082, w_024_1085, w_024_1086, w_024_1087, w_024_1088, w_024_1090, w_024_1091, w_024_1094, w_024_1096, w_024_1099, w_024_1100, w_024_1101, w_024_1102, w_024_1106, w_024_1107, w_024_1109, w_024_1110, w_024_1112, w_024_1113, w_024_1114, w_024_1116, w_024_1117, w_024_1119, w_024_1121, w_024_1122, w_024_1123, w_024_1124, w_024_1126, w_024_1127, w_024_1128, w_024_1129, w_024_1130, w_024_1131, w_024_1132, w_024_1133, w_024_1134, w_024_1135, w_024_1136, w_024_1139, w_024_1140, w_024_1145, w_024_1147, w_024_1149, w_024_1150, w_024_1151, w_024_1153, w_024_1154, w_024_1155, w_024_1156, w_024_1158, w_024_1159, w_024_1160, w_024_1161, w_024_1162, w_024_1164, w_024_1166, w_024_1169, w_024_1170, w_024_1171, w_024_1172, w_024_1173, w_024_1174, w_024_1175, w_024_1177, w_024_1180, w_024_1181, w_024_1182, w_024_1184, w_024_1185, w_024_1186, w_024_1190, w_024_1194, w_024_1196, w_024_1197, w_024_1198, w_024_1199, w_024_1200, w_024_1201, w_024_1202, w_024_1203, w_024_1204, w_024_1205, w_024_1207, w_024_1208, w_024_1210, w_024_1211, w_024_1212, w_024_1213, w_024_1214, w_024_1216, w_024_1217, w_024_1219, w_024_1221, w_024_1222, w_024_1223, w_024_1224, w_024_1226, w_024_1227, w_024_1228, w_024_1229, w_024_1230, w_024_1231, w_024_1232, w_024_1233, w_024_1235, w_024_1236, w_024_1237, w_024_1238, w_024_1240, w_024_1241, w_024_1242, w_024_1246, w_024_1247, w_024_1249, w_024_1250, w_024_1252, w_024_1253, w_024_1254, w_024_1256, w_024_1257, w_024_1258, w_024_1260, w_024_1261, w_024_1262, w_024_1263, w_024_1267, w_024_1268, w_024_1269, w_024_1270, w_024_1272, w_024_1275, w_024_1277, w_024_1278, w_024_1279, w_024_1283, w_024_1284, w_024_1287, w_024_1288, w_024_1289, w_024_1290, w_024_1292, w_024_1293, w_024_1294, w_024_1295, w_024_1297, w_024_1298, w_024_1299, w_024_1302, w_024_1303, w_024_1304, w_024_1305, w_024_1307, w_024_1309, w_024_1311, w_024_1312, w_024_1313, w_024_1314, w_024_1315, w_024_1317, w_024_1318, w_024_1319, w_024_1320, w_024_1321, w_024_1322, w_024_1323, w_024_1324, w_024_1325, w_024_1328, w_024_1329, w_024_1332, w_024_1334, w_024_1336, w_024_1337, w_024_1338, w_024_1339, w_024_1342, w_024_1344, w_024_1347, w_024_1348, w_024_1349, w_024_1350, w_024_1355, w_024_1356, w_024_1357, w_024_1358, w_024_1359, w_024_1361, w_024_1362, w_024_1363, w_024_1366, w_024_1369, w_024_1370, w_024_1371, w_024_1372, w_024_1374, w_024_1378, w_024_1379, w_024_1380, w_024_1381, w_024_1383, w_024_1384, w_024_1385, w_024_1386, w_024_1387, w_024_1388, w_024_1389, w_024_1390, w_024_1391, w_024_1394, w_024_1395, w_024_1397, w_024_1398, w_024_1399, w_024_1402, w_024_1403, w_024_1404, w_024_1406, w_024_1407, w_024_1408, w_024_1409, w_024_1410, w_024_1411, w_024_1412, w_024_1413, w_024_1415, w_024_1417, w_024_1419, w_024_1420, w_024_1421, w_024_1422, w_024_1423, w_024_1426, w_024_1429, w_024_1430, w_024_1431, w_024_1432, w_024_1434, w_024_1435, w_024_1436, w_024_1437, w_024_1438, w_024_1441, w_024_1443, w_024_1444, w_024_1445, w_024_1448, w_024_1450, w_024_1451, w_024_1452, w_024_1454, w_024_1456, w_024_1457, w_024_1461, w_024_1463, w_024_1464, w_024_1467, w_024_1468, w_024_1470, w_024_1471, w_024_1472, w_024_1473, w_024_1474, w_024_1475, w_024_1476, w_024_1478, w_024_1479, w_024_1480, w_024_1481, w_024_1482, w_024_1483, w_024_1485, w_024_1488, w_024_1489, w_024_1493, w_024_1494, w_024_1495, w_024_1496, w_024_1497, w_024_1501, w_024_1502, w_024_1504, w_024_1505, w_024_1506, w_024_1512, w_024_1514, w_024_1515, w_024_1518, w_024_1519, w_024_1521, w_024_1523, w_024_1524, w_024_1525, w_024_1526, w_024_1527, w_024_1529, w_024_1531, w_024_1532, w_024_1534, w_024_1535, w_024_1536, w_024_1537, w_024_1541, w_024_1542, w_024_1544, w_024_1545, w_024_1546, w_024_1547, w_024_1548, w_024_1550, w_024_1552, w_024_1553, w_024_1554, w_024_1556, w_024_1557, w_024_1558, w_024_1559, w_024_1561, w_024_1562, w_024_1563, w_024_1566, w_024_1567, w_024_1568, w_024_1569, w_024_1573, w_024_1574, w_024_1575, w_024_1577, w_024_1578, w_024_1579, w_024_1580, w_024_1581, w_024_1582, w_024_1583, w_024_1584, w_024_1585, w_024_1586, w_024_1587, w_024_1588, w_024_1589, w_024_1590, w_024_1591, w_024_1592, w_024_1593, w_024_1594, w_024_1596, w_024_1601, w_024_1602, w_024_1605, w_024_1606, w_024_1609, w_024_1615, w_024_1617, w_024_1618, w_024_1623, w_024_1626, w_024_1627, w_024_1628, w_024_1631, w_024_1632, w_024_1633, w_024_1634, w_024_1636, w_024_1637, w_024_1640, w_024_1641, w_024_1642, w_024_1643, w_024_1645, w_024_1647, w_024_1648, w_024_1651, w_024_1652, w_024_1653, w_024_1656, w_024_1658, w_024_1659, w_024_1660, w_024_1662, w_024_1663, w_024_1664, w_024_1665, w_024_1669, w_024_1670, w_024_1671, w_024_1672, w_024_1673, w_024_1674, w_024_1676, w_024_1677, w_024_1678, w_024_1679, w_024_1681, w_024_1684, w_024_1685, w_024_1687, w_024_1688, w_024_1689, w_024_1690, w_024_1691, w_024_1692, w_024_1696, w_024_1697, w_024_1699, w_024_1700, w_024_1701, w_024_1702, w_024_1704, w_024_1706, w_024_1707, w_024_1708, w_024_1709, w_024_1714, w_024_1715, w_024_1716, w_024_1719, w_024_1722, w_024_1724, w_024_1725, w_024_1726, w_024_1727, w_024_1728, w_024_1729, w_024_1730, w_024_1731, w_024_1732, w_024_1734, w_024_1735, w_024_1737, w_024_1738, w_024_1739, w_024_1740, w_024_1742, w_024_1743, w_024_1746, w_024_1747, w_024_1748, w_024_1749, w_024_1750, w_024_1751, w_024_1752, w_024_1754, w_024_1757, w_024_1759, w_024_1760, w_024_1763, w_024_1764, w_024_1766, w_024_1767, w_024_1768, w_024_1769, w_024_1770, w_024_1771, w_024_1773, w_024_1777, w_024_1781, w_024_1782, w_024_1783, w_024_1784, w_024_1786, w_024_1787, w_024_1788, w_024_1789, w_024_1790, w_024_1791, w_024_1792, w_024_1793, w_024_1794, w_024_1795, w_024_1796, w_024_1797, w_024_1798, w_024_1800, w_024_1804, w_024_1806, w_024_1808, w_024_1810, w_024_1812, w_024_1813, w_024_1814, w_024_1815, w_024_1817, w_024_1818, w_024_1819, w_024_1821, w_024_1824, w_024_1825, w_024_1826, w_024_1827, w_024_1828, w_024_1829, w_024_1832, w_024_1833, w_024_1834, w_024_1836, w_024_1838, w_024_1839, w_024_1840, w_024_1841, w_024_1842, w_024_1843, w_024_1845, w_024_1846, w_024_1848, w_024_1849, w_024_1851, w_024_1852, w_024_1853, w_024_1855, w_024_1856, w_024_1857, w_024_1858, w_024_1862, w_024_1863, w_024_1864, w_024_1866, w_024_1867, w_024_1868, w_024_1869, w_024_1870, w_024_1871, w_024_1872, w_024_1875, w_024_1877, w_024_1878, w_024_1879, w_024_1881, w_024_1882, w_024_1884, w_024_1885, w_024_1886, w_024_1887, w_024_1888, w_024_1890, w_024_1892, w_024_1893, w_024_1894, w_024_1896, w_024_1898, w_024_1899, w_024_1900, w_024_1901, w_024_1902, w_024_1904, w_024_1906, w_024_1907, w_024_1908, w_024_1910, w_024_1913, w_024_1915, w_024_1917, w_024_1918, w_024_1919, w_024_1920, w_024_1921, w_024_1922, w_024_1924, w_024_1925, w_024_1926, w_024_1928, w_024_1929, w_024_1930, w_024_1931, w_024_1932, w_024_1933, w_024_1938, w_024_1941, w_024_1942, w_024_1943, w_024_1944, w_024_1945, w_024_1947, w_024_1948, w_024_1949, w_024_1951, w_024_1952, w_024_1953, w_024_1954, w_024_1956, w_024_1957, w_024_1958, w_024_1961, w_024_1963, w_024_1966, w_024_1968, w_024_1969, w_024_1970, w_024_1971, w_024_1974, w_024_1975, w_024_1976, w_024_1979, w_024_1981, w_024_1982, w_024_1983, w_024_1985, w_024_1987, w_024_1988, w_024_1990, w_024_1992, w_024_1993, w_024_1994, w_024_1997, w_024_1998, w_024_1999, w_024_2001, w_024_2003, w_024_2004, w_024_2006, w_024_2007, w_024_2008, w_024_2009, w_024_2010, w_024_2011, w_024_2014, w_024_2015, w_024_2016, w_024_2018, w_024_2020, w_024_2022, w_024_2023, w_024_2024, w_024_2025, w_024_2026, w_024_2029, w_024_2030, w_024_2031, w_024_2032, w_024_2033, w_024_2035, w_024_2036, w_024_2037, w_024_2040, w_024_2041, w_024_2042, w_024_2045, w_024_2048, w_024_2050, w_024_2051, w_024_2052, w_024_2053, w_024_2054, w_024_2056, w_024_2057, w_024_2061, w_024_2062, w_024_2064, w_024_2065, w_024_2068, w_024_2069, w_024_2071, w_024_2073, w_024_2074, w_024_2077, w_024_2078, w_024_2079, w_024_2082, w_024_2084, w_024_2085, w_024_2086, w_024_2089, w_024_2090, w_024_2091, w_024_2092, w_024_2093, w_024_2096, w_024_2097, w_024_2099, w_024_2100, w_024_2101, w_024_2104, w_024_2106, w_024_2107, w_024_2108, w_024_2110, w_024_2111, w_024_2113, w_024_2114, w_024_2115, w_024_2116, w_024_2119, w_024_2120, w_024_2121, w_024_2125, w_024_2126, w_024_2127, w_024_2129, w_024_2130, w_024_2132, w_024_2134, w_024_2135, w_024_2136, w_024_2137, w_024_2138, w_024_2140, w_024_2141, w_024_2142, w_024_2143, w_024_2144, w_024_2145, w_024_2146, w_024_2147, w_024_2148, w_024_2149, w_024_2150, w_024_2151, w_024_2152, w_024_2153, w_024_2154, w_024_2156, w_024_2157, w_024_2160, w_024_2162, w_024_2163, w_024_2164, w_024_2168, w_024_2169, w_024_2170, w_024_2172, w_024_2173, w_024_2175, w_024_2177, w_024_2178, w_024_2180, w_024_2182, w_024_2185, w_024_2187, w_024_2188, w_024_2189, w_024_2191, w_024_2192, w_024_2193, w_024_2194, w_024_2196, w_024_2197, w_024_2199, w_024_2200, w_024_2202, w_024_2203, w_024_2204, w_024_2205, w_024_2206, w_024_2207, w_024_2208, w_024_2209, w_024_2210, w_024_2211, w_024_2212, w_024_2213, w_024_2215, w_024_2216, w_024_2218, w_024_2219, w_024_2220, w_024_2221, w_024_2222, w_024_2223, w_024_2224, w_024_2225, w_024_2229, w_024_2230, w_024_2231, w_024_2233, w_024_2234, w_024_2235, w_024_2237, w_024_2239, w_024_2242, w_024_2244, w_024_2245, w_024_2246, w_024_2250, w_024_2251, w_024_2252, w_024_2253, w_024_2254, w_024_2257, w_024_2260, w_024_2261, w_024_2262, w_024_2263, w_024_2264, w_024_2265, w_024_2266, w_024_2267, w_024_2269, w_024_2272, w_024_2273, w_024_2274, w_024_2276, w_024_2278, w_024_2279, w_024_2280, w_024_2282, w_024_2283, w_024_2285, w_024_2286, w_024_2287, w_024_2288, w_024_2290, w_024_2291, w_024_2292, w_024_2293, w_024_2296, w_024_2297, w_024_2299, w_024_2300, w_024_2301, w_024_2302, w_024_2303, w_024_2304, w_024_2307, w_024_2309, w_024_2310, w_024_2311, w_024_2312, w_024_2313, w_024_2314, w_024_2315, w_024_2316, w_024_2317, w_024_2318, w_024_2319, w_024_2320, w_024_2322, w_024_2323, w_024_2324, w_024_2326, w_024_2327, w_024_2329, w_024_2330, w_024_2331, w_024_2332, w_024_2333, w_024_2334, w_024_2335, w_024_2336, w_024_2338, w_024_2339, w_024_2340, w_024_2342, w_024_2345, w_024_2346, w_024_2347, w_024_2349, w_024_2350, w_024_2351, w_024_2353, w_024_2354, w_024_2355, w_024_2356, w_024_2357, w_024_2358, w_024_2359, w_024_2360, w_024_2363, w_024_2365, w_024_2366, w_024_2369, w_024_2370, w_024_2371, w_024_2372, w_024_2374, w_024_2375, w_024_2377, w_024_2380, w_024_2381, w_024_2382, w_024_2384, w_024_2386, w_024_2389, w_024_2390, w_024_2391, w_024_2395, w_024_2396, w_024_2399, w_024_2400, w_024_2401, w_024_2402, w_024_2403, w_024_2406, w_024_2407, w_024_2408, w_024_2409, w_024_2410, w_024_2412, w_024_2416, w_024_2417, w_024_2418, w_024_2419, w_024_2420, w_024_2421, w_024_2422, w_024_2423, w_024_2424, w_024_2426, w_024_2427, w_024_2428, w_024_2429, w_024_2431, w_024_2432, w_024_2435, w_024_2437, w_024_2439, w_024_2440, w_024_2441, w_024_2442, w_024_2444, w_024_2445, w_024_2446, w_024_2449, w_024_2450, w_024_2451, w_024_2452, w_024_2453, w_024_2454, w_024_2456, w_024_2457, w_024_2458, w_024_2459, w_024_2460, w_024_2461, w_024_2462, w_024_2464, w_024_2465, w_024_2466, w_024_2467, w_024_2471, w_024_2472, w_024_2474, w_024_2475, w_024_2476, w_024_2477, w_024_2479, w_024_2480, w_024_2481, w_024_2484, w_024_2487, w_024_2488, w_024_2490, w_024_2491, w_024_2492, w_024_2493, w_024_2494, w_024_2496, w_024_2497, w_024_2498, w_024_2499, w_024_2500, w_024_2501, w_024_2503, w_024_2504, w_024_2508, w_024_2509, w_024_2510, w_024_2512, w_024_2513, w_024_2514, w_024_2515, w_024_2516, w_024_2518, w_024_2519, w_024_2520, w_024_2521, w_024_2522, w_024_2523, w_024_2525, w_024_2526, w_024_2527, w_024_2528, w_024_2529, w_024_2530, w_024_2532, w_024_2533, w_024_2534, w_024_2535, w_024_2536, w_024_2537, w_024_2538, w_024_2539, w_024_2540, w_024_2541, w_024_2542, w_024_2545, w_024_2546, w_024_2548, w_024_2549, w_024_2550, w_024_2551, w_024_2552, w_024_2553, w_024_2554, w_024_2555, w_024_2556, w_024_2557, w_024_2558, w_024_2559, w_024_2560, w_024_2561, w_024_2562, w_024_2563, w_024_2565, w_024_2566, w_024_2569, w_024_2570, w_024_2571, w_024_2573, w_024_2575, w_024_2576, w_024_2578, w_024_2580, w_024_2581, w_024_2582, w_024_2583, w_024_2584, w_024_2585, w_024_2587, w_024_2592, w_024_2593, w_024_2594, w_024_2595, w_024_2596, w_024_2597, w_024_2598, w_024_2599, w_024_2600, w_024_2601, w_024_2602, w_024_2604, w_024_2606, w_024_2607, w_024_2609, w_024_2610, w_024_2613, w_024_2614, w_024_2616, w_024_2617, w_024_2618, w_024_2619, w_024_2621, w_024_2622, w_024_2623, w_024_2625, w_024_2627, w_024_2629, w_024_2630, w_024_2631, w_024_2632, w_024_2635, w_024_2636, w_024_2638, w_024_2639, w_024_2640, w_024_2641, w_024_2642, w_024_2647, w_024_2649, w_024_2650, w_024_2651, w_024_2652, w_024_2653, w_024_2658, w_024_2660, w_024_2663, w_024_2664, w_024_2667, w_024_2670, w_024_2672, w_024_2673, w_024_2675, w_024_2676, w_024_2677, w_024_2678, w_024_2679, w_024_2680, w_024_2682, w_024_2684, w_024_2685, w_024_2686, w_024_2687, w_024_2688, w_024_2689, w_024_2691, w_024_2694, w_024_2696, w_024_2697, w_024_2699, w_024_2700, w_024_2701, w_024_2702, w_024_2704, w_024_2705, w_024_2706, w_024_2708, w_024_2710, w_024_2711, w_024_2712, w_024_2713, w_024_2714, w_024_2716, w_024_2717, w_024_2718, w_024_2719, w_024_2720, w_024_2721, w_024_2722, w_024_2723, w_024_2724, w_024_2725, w_024_2726, w_024_2727, w_024_2731, w_024_2732, w_024_2733, w_024_2735, w_024_2736, w_024_2737, w_024_2739, w_024_2740, w_024_2741, w_024_2742, w_024_2743, w_024_2744, w_024_2745, w_024_2746, w_024_2747, w_024_2750, w_024_2751, w_024_2752, w_024_2753, w_024_2754, w_024_2755, w_024_2759, w_024_2760, w_024_2762, w_024_2763, w_024_2765, w_024_2766, w_024_2767, w_024_2768, w_024_2769, w_024_2770, w_024_2771, w_024_2773, w_024_2775, w_024_2776, w_024_2779, w_024_2780, w_024_2781, w_024_2782, w_024_2783, w_024_2784, w_024_2785, w_024_2786, w_024_2788, w_024_2789, w_024_2790, w_024_2792, w_024_2794, w_024_2795, w_024_2796, w_024_2797, w_024_2798, w_024_2799, w_024_2800, w_024_2801, w_024_2802, w_024_2804, w_024_2805, w_024_2806, w_024_2808, w_024_2810, w_024_2812, w_024_2813, w_024_2814, w_024_2815, w_024_2818, w_024_2819, w_024_2821, w_024_2824, w_024_2827, w_024_2829, w_024_2830, w_024_2831, w_024_2832, w_024_2833, w_024_2834, w_024_2835, w_024_2837, w_024_2839, w_024_2840, w_024_2841, w_024_2843, w_024_2844, w_024_2845, w_024_2846, w_024_2848, w_024_2850, w_024_2851, w_024_2852, w_024_2853, w_024_2854, w_024_2857, w_024_2859, w_024_2860, w_024_2861, w_024_2862, w_024_2863, w_024_2864, w_024_2867, w_024_2868, w_024_2869, w_024_2870, w_024_2871, w_024_2872, w_024_2873, w_024_2874, w_024_2875, w_024_2879, w_024_2880, w_024_2881, w_024_2882, w_024_2883, w_024_2884, w_024_2886, w_024_2888, w_024_2889, w_024_2890, w_024_2891, w_024_2893, w_024_2895, w_024_2896, w_024_2897, w_024_2898, w_024_2899, w_024_2900, w_024_2902, w_024_2904, w_024_2905, w_024_2906, w_024_2907, w_024_2910, w_024_2912, w_024_2913, w_024_2914, w_024_2917, w_024_2919, w_024_2920, w_024_2921, w_024_2923, w_024_2925, w_024_2926, w_024_2932, w_024_2933, w_024_2936, w_024_2937, w_024_2940, w_024_2943, w_024_2944, w_024_2945, w_024_2947, w_024_2948, w_024_2950, w_024_2952, w_024_2953, w_024_2958, w_024_2959, w_024_2960, w_024_2961, w_024_2963, w_024_2965, w_024_2967, w_024_2968, w_024_2970, w_024_2972, w_024_2973, w_024_2974, w_024_2975, w_024_2976, w_024_2977, w_024_2978, w_024_2979, w_024_2981, w_024_2982, w_024_2983, w_024_2984, w_024_2985, w_024_2986, w_024_2987, w_024_2989, w_024_2990, w_024_2991, w_024_2994, w_024_2995, w_024_2996, w_024_2997, w_024_2998, w_024_3000, w_024_3001, w_024_3004, w_024_3006, w_024_3008, w_024_3009, w_024_3010, w_024_3011, w_024_3012, w_024_3013, w_024_3014, w_024_3016, w_024_3017, w_024_3019, w_024_3020, w_024_3021, w_024_3022, w_024_3024, w_024_3026, w_024_3027, w_024_3028, w_024_3032, w_024_3033, w_024_3035, w_024_3036, w_024_3037, w_024_3038, w_024_3039, w_024_3040, w_024_3041, w_024_3042, w_024_3045, w_024_3046, w_024_3048, w_024_3050, w_024_3051, w_024_3052, w_024_3053, w_024_3054, w_024_3055, w_024_3056, w_024_3057, w_024_3058, w_024_3059, w_024_3060, w_024_3061, w_024_3063, w_024_3064, w_024_3066, w_024_3068, w_024_3071, w_024_3072, w_024_3074, w_024_3075, w_024_3076, w_024_3077, w_024_3079, w_024_3082, w_024_3083, w_024_3084, w_024_3087, w_024_3088, w_024_3089, w_024_3090, w_024_3091, w_024_3092, w_024_3094, w_024_3098, w_024_3099, w_024_3100, w_024_3101, w_024_3103, w_024_3104, w_024_3105, w_024_3106, w_024_3107, w_024_3108, w_024_3112, w_024_3113, w_024_3115, w_024_3116, w_024_3119, w_024_3120, w_024_3121, w_024_3122, w_024_3124, w_024_3125, w_024_3126, w_024_3127, w_024_3128, w_024_3129, w_024_3130, w_024_3131, w_024_3132, w_024_3133, w_024_3135, w_024_3136, w_024_3137, w_024_3138, w_024_3139, w_024_3146, w_024_3147, w_024_3149, w_024_3150, w_024_3151, w_024_3154, w_024_3155, w_024_3157, w_024_3158, w_024_3162, w_024_3163, w_024_3164, w_024_3165, w_024_3166, w_024_3168, w_024_3169, w_024_3173, w_024_3175, w_024_3177, w_024_3178, w_024_3179, w_024_3180, w_024_3181, w_024_3182, w_024_3183, w_024_3188, w_024_3189, w_024_3190, w_024_3191, w_024_3192, w_024_3193, w_024_3195, w_024_3196, w_024_3197, w_024_3198, w_024_3199, w_024_3202, w_024_3204, w_024_3205, w_024_3207, w_024_3208, w_024_3209, w_024_3210, w_024_3212, w_024_3214, w_024_3215, w_024_3216, w_024_3217, w_024_3218, w_024_3219, w_024_3220, w_024_3221, w_024_3223, w_024_3224, w_024_3230, w_024_3232, w_024_3233, w_024_3235, w_024_3237, w_024_3238, w_024_3239, w_024_3240, w_024_3242, w_024_3243, w_024_3244, w_024_3245, w_024_3246, w_024_3250, w_024_3251, w_024_3252, w_024_3253, w_024_3254, w_024_3256, w_024_3257, w_024_3259, w_024_3260, w_024_3262, w_024_3263, w_024_3265, w_024_3266, w_024_3267, w_024_3269, w_024_3270, w_024_3271, w_024_3276, w_024_3278, w_024_3279, w_024_3280, w_024_3281, w_024_3288, w_024_3289, w_024_3290, w_024_3291, w_024_3293, w_024_3294, w_024_3295, w_024_3296, w_024_3298, w_024_3299, w_024_3300, w_024_3301, w_024_3303, w_024_3304, w_024_3306, w_024_3307, w_024_3308, w_024_3312, w_024_3313, w_024_3315, w_024_3316, w_024_3317, w_024_3318, w_024_3319, w_024_3321, w_024_3322, w_024_3324, w_024_3325, w_024_3328, w_024_3330, w_024_3331, w_024_3336, w_024_3339, w_024_3340, w_024_3341, w_024_3342, w_024_3343, w_024_3348, w_024_3349, w_024_3350, w_024_3351, w_024_3352, w_024_3353, w_024_3354, w_024_3358, w_024_3359, w_024_3360, w_024_3361, w_024_3363, w_024_3364, w_024_3365, w_024_3366, w_024_3368, w_024_3369, w_024_3371, w_024_3372, w_024_3373, w_024_3375, w_024_3376, w_024_3377, w_024_3378, w_024_3380, w_024_3383, w_024_3384, w_024_3385, w_024_3387, w_024_3388, w_024_3391, w_024_3392, w_024_3393, w_024_3394, w_024_3398, w_024_3402, w_024_3403, w_024_3404, w_024_3405, w_024_3406, w_024_3407, w_024_3409, w_024_3410, w_024_3414, w_024_3415, w_024_3418, w_024_3420, w_024_3424, w_024_3425, w_024_3427, w_024_3430, w_024_3433, w_024_3434, w_024_3435, w_024_3436, w_024_3437, w_024_3439, w_024_3440, w_024_3441, w_024_3443, w_024_3444, w_024_3445, w_024_3446, w_024_3447, w_024_3449, w_024_3453, w_024_3454, w_024_3457, w_024_3458, w_024_3459, w_024_3461, w_024_3462, w_024_3464, w_024_3465, w_024_3466, w_024_3467, w_024_3468, w_024_3469, w_024_3470, w_024_3472, w_024_3473, w_024_3475, w_024_3477, w_024_3478, w_024_3479, w_024_3480, w_024_3481, w_024_3482, w_024_3483, w_024_3485, w_024_3487, w_024_3488, w_024_3489, w_024_3492, w_024_3493, w_024_3494, w_024_3495, w_024_3496, w_024_3497, w_024_3498, w_024_3499, w_024_3501, w_024_3504, w_024_3505, w_024_3506, w_024_3507, w_024_3509, w_024_3511, w_024_3513, w_024_3519, w_024_3522, w_024_3523, w_024_3526, w_024_3528, w_024_3529, w_024_3530, w_024_3531, w_024_3532, w_024_3533, w_024_3534, w_024_3535, w_024_3538, w_024_3539, w_024_3540, w_024_3541, w_024_3542, w_024_3543, w_024_3545, w_024_3546, w_024_3547, w_024_3548, w_024_3550, w_024_3551, w_024_3553, w_024_3554, w_024_3556, w_024_3557, w_024_3558, w_024_3559, w_024_3560, w_024_3561, w_024_3562, w_024_3564, w_024_3567, w_024_3571, w_024_3572, w_024_3573, w_024_3575, w_024_3577, w_024_3579, w_024_3580, w_024_3581, w_024_3582, w_024_3583, w_024_3584, w_024_3585, w_024_3588, w_024_3591, w_024_3592, w_024_3594, w_024_3595, w_024_3596, w_024_3598, w_024_3600, w_024_3602, w_024_3603, w_024_3604, w_024_3605, w_024_3606, w_024_3607, w_024_3608, w_024_3609, w_024_3611, w_024_3612, w_024_3613, w_024_3616, w_024_3617, w_024_3618, w_024_3619, w_024_3620, w_024_3621, w_024_3622, w_024_3623, w_024_3624, w_024_3625, w_024_3626, w_024_3629, w_024_3630, w_024_3631, w_024_3633, w_024_3635, w_024_3636, w_024_3638, w_024_3639, w_024_3640, w_024_3641, w_024_3642, w_024_3644, w_024_3645, w_024_3646, w_024_3647, w_024_3650, w_024_3651, w_024_3652, w_024_3653, w_024_3654, w_024_3655, w_024_3656, w_024_3657, w_024_3658, w_024_3659, w_024_3665, w_024_3667, w_024_3668, w_024_3669, w_024_3670, w_024_3671, w_024_3672, w_024_3673, w_024_3674, w_024_3675, w_024_3676, w_024_3677, w_024_3678, w_024_3679, w_024_3681, w_024_3683, w_024_3689, w_024_3690, w_024_3691, w_024_3692, w_024_3693, w_024_3694, w_024_3695, w_024_3696, w_024_3697, w_024_3701, w_024_3702, w_024_3703, w_024_3704, w_024_3705, w_024_3706, w_024_3707, w_024_3711, w_024_3712, w_024_3713, w_024_3714, w_024_3717, w_024_3718, w_024_3719, w_024_3720, w_024_3726, w_024_3727, w_024_3728, w_024_3729, w_024_3730, w_024_3731, w_024_3732, w_024_3733, w_024_3734, w_024_3735, w_024_3740, w_024_3741, w_024_3743, w_024_3745, w_024_3746, w_024_3748, w_024_3749, w_024_3750, w_024_3751, w_024_3752, w_024_3755, w_024_3757, w_024_3759, w_024_3760, w_024_3762, w_024_3763, w_024_3764, w_024_3765, w_024_3767, w_024_3768, w_024_3771, w_024_3772, w_024_3773, w_024_3774, w_024_3775, w_024_3776, w_024_3778, w_024_3779, w_024_3782, w_024_3783, w_024_3784, w_024_3786, w_024_3787, w_024_3790, w_024_3791, w_024_3792, w_024_3793, w_024_3796, w_024_3797, w_024_3798, w_024_3800, w_024_3801, w_024_3803, w_024_3804, w_024_3805, w_024_3806, w_024_3807, w_024_3809, w_024_3811, w_024_3813, w_024_3814, w_024_3816, w_024_3817, w_024_3818, w_024_3820, w_024_3822, w_024_3824, w_024_3825, w_024_3826, w_024_3827, w_024_3828, w_024_3829, w_024_3830, w_024_3831, w_024_3832, w_024_3833, w_024_3835, w_024_3836, w_024_3839, w_024_3840, w_024_3841, w_024_3842, w_024_3843, w_024_3844, w_024_3845, w_024_3846, w_024_3847, w_024_3852, w_024_3853, w_024_3858, w_024_3861, w_024_3862, w_024_3863, w_024_3864, w_024_3865, w_024_3866, w_024_3867, w_024_3868, w_024_3869, w_024_3871, w_024_3874, w_024_3875, w_024_3876, w_024_3877, w_024_3878, w_024_3879, w_024_3880, w_024_3882, w_024_3885, w_024_3886, w_024_3888, w_024_3890, w_024_3892, w_024_3893, w_024_3896, w_024_3897, w_024_3898, w_024_3899, w_024_3900, w_024_3902, w_024_3905, w_024_3906, w_024_3907, w_024_3908, w_024_3911, w_024_3912, w_024_3914, w_024_3916, w_024_3917, w_024_3918, w_024_3922, w_024_3925, w_024_3927, w_024_3929, w_024_3932, w_024_3933, w_024_3935, w_024_3937, w_024_3938, w_024_3939, w_024_3941, w_024_3945, w_024_3946, w_024_3948, w_024_3951, w_024_3952, w_024_3953, w_024_3955, w_024_3957, w_024_3958, w_024_3961, w_024_3962, w_024_3963, w_024_3964, w_024_3965, w_024_3967, w_024_3968, w_024_3970, w_024_3971, w_024_3972, w_024_3973, w_024_3974, w_024_3975, w_024_3976, w_024_3978, w_024_3981, w_024_3982, w_024_3983, w_024_3986, w_024_3987, w_024_3988, w_024_3989, w_024_3992, w_024_3997, w_024_3998, w_024_4000, w_024_4001, w_024_4002, w_024_4003, w_024_4005, w_024_4006, w_024_4009, w_024_4011, w_024_4013, w_024_4014, w_024_4015, w_024_4017, w_024_4019, w_024_4020, w_024_4021, w_024_4022, w_024_4023, w_024_4025, w_024_4027, w_024_4028, w_024_4030, w_024_4033, w_024_4034, w_024_4035, w_024_4037, w_024_4038, w_024_4039, w_024_4040, w_024_4041, w_024_4042, w_024_4043, w_024_4044, w_024_4045, w_024_4046, w_024_4047, w_024_4048, w_024_4051, w_024_4052, w_024_4055, w_024_4059, w_024_4060, w_024_4061, w_024_4062, w_024_4063, w_024_4064, w_024_4067, w_024_4068, w_024_4069, w_024_4070, w_024_4071, w_024_4072, w_024_4073, w_024_4074, w_024_4075, w_024_4077, w_024_4079, w_024_4081, w_024_4082, w_024_4083, w_024_4084, w_024_4085, w_024_4086, w_024_4087, w_024_4088, w_024_4089, w_024_4091, w_024_4092, w_024_4094, w_024_4095, w_024_4097, w_024_4100, w_024_4101, w_024_4103, w_024_4104, w_024_4105, w_024_4106, w_024_4107, w_024_4109, w_024_4111, w_024_4112, w_024_4113, w_024_4115, w_024_4116, w_024_4119, w_024_4121, w_024_4122, w_024_4123, w_024_4124, w_024_4125, w_024_4126, w_024_4127, w_024_4128, w_024_4129, w_024_4130, w_024_4131, w_024_4132, w_024_4135, w_024_4136, w_024_4137, w_024_4140, w_024_4141, w_024_4142, w_024_4143, w_024_4145, w_024_4147, w_024_4148, w_024_4149, w_024_4150, w_024_4153, w_024_4154, w_024_4155, w_024_4160, w_024_4161, w_024_4162, w_024_4163, w_024_4164, w_024_4165, w_024_4167, w_024_4168, w_024_4169, w_024_4171, w_024_4172, w_024_4173, w_024_4177, w_024_4178, w_024_4179, w_024_4180, w_024_4182, w_024_4183, w_024_4185, w_024_4186, w_024_4188, w_024_4189, w_024_4190, w_024_4193, w_024_4194, w_024_4195, w_024_4196, w_024_4197, w_024_4198, w_024_4199, w_024_4200, w_024_4201, w_024_4202, w_024_4203, w_024_4204, w_024_4205, w_024_4207, w_024_4208, w_024_4209, w_024_4211, w_024_4212, w_024_4215, w_024_4217, w_024_4220, w_024_4222, w_024_4223, w_024_4225, w_024_4226, w_024_4228, w_024_4229, w_024_4230, w_024_4231, w_024_4232, w_024_4234, w_024_4236, w_024_4237, w_024_4244, w_024_4245, w_024_4246, w_024_4247, w_024_4248, w_024_4251, w_024_4254, w_024_4255, w_024_4256, w_024_4257, w_024_4258, w_024_4259, w_024_4261, w_024_4262, w_024_4263, w_024_4264, w_024_4268, w_024_4270, w_024_4271, w_024_4273, w_024_4275, w_024_4276, w_024_4277, w_024_4278, w_024_4279, w_024_4282, w_024_4283, w_024_4284, w_024_4286, w_024_4287, w_024_4289, w_024_4291, w_024_4292, w_024_4294, w_024_4295, w_024_4296, w_024_4297, w_024_4299, w_024_4300, w_024_4302, w_024_4303, w_024_4304, w_024_4306, w_024_4307, w_024_4308, w_024_4309, w_024_4310, w_024_4311, w_024_4312, w_024_4313, w_024_4314, w_024_4315, w_024_4316, w_024_4317, w_024_4318, w_024_4320, w_024_4321, w_024_4322, w_024_4325, w_024_4326, w_024_4327, w_024_4331, w_024_4332, w_024_4333, w_024_4336, w_024_4338, w_024_4339, w_024_4342, w_024_4343, w_024_4344, w_024_4345, w_024_4346, w_024_4347, w_024_4348, w_024_4349, w_024_4350, w_024_4353, w_024_4356, w_024_4357, w_024_4359, w_024_4360, w_024_4361, w_024_4363, w_024_4365, w_024_4366, w_024_4367, w_024_4368, w_024_4369, w_024_4371, w_024_4373, w_024_4374, w_024_4375, w_024_4377, w_024_4378, w_024_4379, w_024_4380, w_024_4382, w_024_4383, w_024_4384, w_024_4385, w_024_4387, w_024_4389, w_024_4391, w_024_4392, w_024_4393, w_024_4395, w_024_4400, w_024_4402, w_024_4403, w_024_4404, w_024_4405, w_024_4406, w_024_4407, w_024_4408, w_024_4411, w_024_4412, w_024_4415, w_024_4416, w_024_4417, w_024_4418, w_024_4424, w_024_4425, w_024_4426, w_024_4427, w_024_4428, w_024_4429, w_024_4430, w_024_4433, w_024_4434, w_024_4435, w_024_4436, w_024_4439, w_024_4442, w_024_4443, w_024_4444, w_024_4445, w_024_4446, w_024_4447, w_024_4448, w_024_4449, w_024_4451, w_024_4454, w_024_4456, w_024_4458, w_024_4460, w_024_4461, w_024_4462, w_024_4464, w_024_4466, w_024_4467, w_024_4471, w_024_4472, w_024_4474, w_024_4475, w_024_4476, w_024_4477, w_024_4479, w_024_4480, w_024_4482, w_024_4483, w_024_4485, w_024_4486, w_024_4488, w_024_4489, w_024_4490, w_024_4491, w_024_4492, w_024_4493, w_024_4496, w_024_4497, w_024_4498, w_024_4499, w_024_4500, w_024_4501, w_024_4503, w_024_4504, w_024_4505, w_024_4506, w_024_4507, w_024_4508, w_024_4509, w_024_4512, w_024_4513, w_024_4514, w_024_4516, w_024_4517, w_024_4518, w_024_4521, w_024_4523, w_024_4524, w_024_4525, w_024_4526, w_024_4527, w_024_4529, w_024_4531, w_024_4533, w_024_4534, w_024_4536, w_024_4537, w_024_4538, w_024_4539, w_024_4542, w_024_4543, w_024_4544, w_024_4545, w_024_4546, w_024_4547, w_024_4548, w_024_4549, w_024_4550, w_024_4551, w_024_4554, w_024_4556, w_024_4557, w_024_4558, w_024_4559, w_024_4568, w_024_4569, w_024_4570, w_024_4571, w_024_4572, w_024_4573, w_024_4574, w_024_4577, w_024_4578, w_024_4582, w_024_4583, w_024_4585, w_024_4586, w_024_4587, w_024_4588, w_024_4589, w_024_4591, w_024_4594, w_024_4595, w_024_4596, w_024_4600, w_024_4601, w_024_4602, w_024_4604, w_024_4605, w_024_4606, w_024_4609, w_024_4610, w_024_4611, w_024_4613, w_024_4617, w_024_4618, w_024_4619, w_024_4620, w_024_4621, w_024_4622, w_024_4623, w_024_4624, w_024_4625, w_024_4627, w_024_4628, w_024_4629, w_024_4630, w_024_4631, w_024_4633, w_024_4635, w_024_4636, w_024_4639, w_024_4640, w_024_4641, w_024_4642, w_024_4643, w_024_4644, w_024_4646, w_024_4647, w_024_4648, w_024_4650, w_024_4651, w_024_4652, w_024_4654, w_024_4655, w_024_4657, w_024_4660, w_024_4662, w_024_4663, w_024_4664, w_024_4665, w_024_4667, w_024_4669, w_024_4671, w_024_4672, w_024_4673, w_024_4675, w_024_4676, w_024_4677, w_024_4679, w_024_4681, w_024_4684, w_024_4687, w_024_4690, w_024_4692, w_024_4696, w_024_4697, w_024_4700;
  wire w_025_000, w_025_001, w_025_002, w_025_003, w_025_004, w_025_005, w_025_006, w_025_008, w_025_009, w_025_010, w_025_011, w_025_012, w_025_013, w_025_014, w_025_015, w_025_016, w_025_017, w_025_018, w_025_019, w_025_020, w_025_022, w_025_024, w_025_025, w_025_026, w_025_027, w_025_028, w_025_029, w_025_030, w_025_031, w_025_032, w_025_033, w_025_034, w_025_035, w_025_036, w_025_037, w_025_038, w_025_039, w_025_040, w_025_041, w_025_042, w_025_043, w_025_044, w_025_045, w_025_046, w_025_047, w_025_048, w_025_049, w_025_050, w_025_051, w_025_052, w_025_053, w_025_054, w_025_055, w_025_056, w_025_057, w_025_058, w_025_059, w_025_060, w_025_061, w_025_062, w_025_063, w_025_064, w_025_065, w_025_066, w_025_067, w_025_068, w_025_069, w_025_070, w_025_071, w_025_072, w_025_073, w_025_074, w_025_075, w_025_076, w_025_077, w_025_078, w_025_079, w_025_080, w_025_081, w_025_082, w_025_083, w_025_084, w_025_085, w_025_086, w_025_087, w_025_088, w_025_089, w_025_091, w_025_092, w_025_093, w_025_094, w_025_096, w_025_097, w_025_098, w_025_099, w_025_100, w_025_101, w_025_102, w_025_103, w_025_104, w_025_105, w_025_106, w_025_107, w_025_108, w_025_109, w_025_110, w_025_111, w_025_112, w_025_113, w_025_114, w_025_115, w_025_116, w_025_117, w_025_118, w_025_119, w_025_120, w_025_121, w_025_122, w_025_123, w_025_124, w_025_125, w_025_126, w_025_127, w_025_128, w_025_129, w_025_130, w_025_131, w_025_132, w_025_133, w_025_134, w_025_135, w_025_136, w_025_137, w_025_138, w_025_139, w_025_140, w_025_141, w_025_142, w_025_143, w_025_144, w_025_145, w_025_146, w_025_147, w_025_148, w_025_149, w_025_150, w_025_152, w_025_153, w_025_154, w_025_155, w_025_156, w_025_157, w_025_158, w_025_159, w_025_160, w_025_161, w_025_162, w_025_163, w_025_164, w_025_165, w_025_166, w_025_167, w_025_168, w_025_169, w_025_170, w_025_171, w_025_172, w_025_173, w_025_174, w_025_175, w_025_176, w_025_177, w_025_178, w_025_179, w_025_180, w_025_181, w_025_182, w_025_183, w_025_184, w_025_185, w_025_186, w_025_187, w_025_188, w_025_189, w_025_190, w_025_191, w_025_192, w_025_193, w_025_194, w_025_195, w_025_196, w_025_197, w_025_198, w_025_199, w_025_200, w_025_201, w_025_202, w_025_203, w_025_204, w_025_205, w_025_206, w_025_207, w_025_208, w_025_209, w_025_210, w_025_212, w_025_213, w_025_214, w_025_215, w_025_216, w_025_217, w_025_218, w_025_219, w_025_220, w_025_221, w_025_222, w_025_223, w_025_224, w_025_225, w_025_226, w_025_227, w_025_228, w_025_229, w_025_230, w_025_231, w_025_232, w_025_233, w_025_234, w_025_235, w_025_236, w_025_237, w_025_238, w_025_239, w_025_240, w_025_241, w_025_242, w_025_243, w_025_244, w_025_245, w_025_246, w_025_247, w_025_248, w_025_249, w_025_250, w_025_251, w_025_252, w_025_253, w_025_254, w_025_255, w_025_256, w_025_257, w_025_258, w_025_259, w_025_260, w_025_261, w_025_262, w_025_263, w_025_264, w_025_265, w_025_266, w_025_267, w_025_268, w_025_269, w_025_270, w_025_271, w_025_272, w_025_273, w_025_274, w_025_275, w_025_276, w_025_277, w_025_278, w_025_279, w_025_282, w_025_283, w_025_284, w_025_285, w_025_286, w_025_287, w_025_288, w_025_289, w_025_290, w_025_291, w_025_292, w_025_293, w_025_295, w_025_296, w_025_297, w_025_298, w_025_299, w_025_300, w_025_301, w_025_302, w_025_303, w_025_304, w_025_305, w_025_306, w_025_307, w_025_308, w_025_309, w_025_310, w_025_311, w_025_312, w_025_313, w_025_314, w_025_315, w_025_316, w_025_317, w_025_318, w_025_319, w_025_320, w_025_321, w_025_322, w_025_323, w_025_324, w_025_325, w_025_326, w_025_327, w_025_328, w_025_329, w_025_330, w_025_331, w_025_333, w_025_334, w_025_335, w_025_336, w_025_337, w_025_338, w_025_339, w_025_340, w_025_341, w_025_342, w_025_343, w_025_344, w_025_345, w_025_346, w_025_347, w_025_348, w_025_349, w_025_350, w_025_351, w_025_352, w_025_353, w_025_354, w_025_355, w_025_356, w_025_357, w_025_358, w_025_359, w_025_360, w_025_361, w_025_362, w_025_363, w_025_364, w_025_365, w_025_366, w_025_367, w_025_368, w_025_369, w_025_370, w_025_371, w_025_372, w_025_373, w_025_374, w_025_375, w_025_376, w_025_377, w_025_378, w_025_379, w_025_381, w_025_382, w_025_383, w_025_384, w_025_385, w_025_386, w_025_387, w_025_388, w_025_389, w_025_390, w_025_391, w_025_392, w_025_393, w_025_394, w_025_395, w_025_396, w_025_397, w_025_398, w_025_399, w_025_400, w_025_401, w_025_402, w_025_403, w_025_404, w_025_405, w_025_406, w_025_407, w_025_408, w_025_409, w_025_410, w_025_411, w_025_412, w_025_413, w_025_415, w_025_416, w_025_417, w_025_418, w_025_419, w_025_420, w_025_421, w_025_422, w_025_423, w_025_424, w_025_425, w_025_426, w_025_427, w_025_428, w_025_429, w_025_430, w_025_431, w_025_432, w_025_433, w_025_434, w_025_435, w_025_436, w_025_437, w_025_438, w_025_439, w_025_440, w_025_441, w_025_442, w_025_443, w_025_444, w_025_445, w_025_446, w_025_447, w_025_448, w_025_449, w_025_450, w_025_451, w_025_452, w_025_454, w_025_455, w_025_456, w_025_457, w_025_458, w_025_459, w_025_460, w_025_462, w_025_463, w_025_464, w_025_465, w_025_466, w_025_467, w_025_468, w_025_469, w_025_470, w_025_471, w_025_472, w_025_473, w_025_474, w_025_475, w_025_476, w_025_477, w_025_478, w_025_479, w_025_480, w_025_481, w_025_482, w_025_483, w_025_484, w_025_485, w_025_486, w_025_487, w_025_488, w_025_489, w_025_490, w_025_491, w_025_492, w_025_493, w_025_494, w_025_495, w_025_496, w_025_497, w_025_498, w_025_499, w_025_500, w_025_501, w_025_502, w_025_503, w_025_504, w_025_505, w_025_506, w_025_507, w_025_508, w_025_509, w_025_510, w_025_511, w_025_512, w_025_513, w_025_514, w_025_515, w_025_516, w_025_517, w_025_518, w_025_519, w_025_520, w_025_521, w_025_522, w_025_523, w_025_525, w_025_526, w_025_527, w_025_528, w_025_529, w_025_530, w_025_531, w_025_532, w_025_533, w_025_534, w_025_535, w_025_536, w_025_537, w_025_538, w_025_539, w_025_540, w_025_541, w_025_542, w_025_543, w_025_544, w_025_546, w_025_547, w_025_548, w_025_549, w_025_550, w_025_551, w_025_552, w_025_553, w_025_554, w_025_555, w_025_556, w_025_557, w_025_558, w_025_559, w_025_560, w_025_561, w_025_563, w_025_564, w_025_565, w_025_566, w_025_567, w_025_568, w_025_569, w_025_570, w_025_571, w_025_572, w_025_573, w_025_574, w_025_575, w_025_576, w_025_577, w_025_578, w_025_579, w_025_580, w_025_581, w_025_582, w_025_583, w_025_584, w_025_585, w_025_586, w_025_588, w_025_589, w_025_590, w_025_592, w_025_593, w_025_594, w_025_595, w_025_596, w_025_597, w_025_598, w_025_599, w_025_600, w_025_601, w_025_602, w_025_603, w_025_604, w_025_605, w_025_606, w_025_607, w_025_608, w_025_609, w_025_610, w_025_611, w_025_612, w_025_613, w_025_614, w_025_615, w_025_616, w_025_617, w_025_618, w_025_619, w_025_620, w_025_621, w_025_622, w_025_623, w_025_624, w_025_625, w_025_626, w_025_627, w_025_628, w_025_629, w_025_630, w_025_631, w_025_632, w_025_633, w_025_634, w_025_635, w_025_636, w_025_637, w_025_638, w_025_639, w_025_640, w_025_641, w_025_642, w_025_643, w_025_644, w_025_645, w_025_646, w_025_647, w_025_648, w_025_649, w_025_650, w_025_651, w_025_652, w_025_654, w_025_655, w_025_656, w_025_657, w_025_658, w_025_659, w_025_660, w_025_661, w_025_662, w_025_664, w_025_665, w_025_666, w_025_667, w_025_668, w_025_669, w_025_670, w_025_671, w_025_672, w_025_673, w_025_674, w_025_675, w_025_676, w_025_677, w_025_678, w_025_679, w_025_681, w_025_682, w_025_684, w_025_685, w_025_686, w_025_687, w_025_688, w_025_689, w_025_690, w_025_691, w_025_692, w_025_693, w_025_694, w_025_695, w_025_696, w_025_697, w_025_698, w_025_699, w_025_700, w_025_701, w_025_702, w_025_703, w_025_704, w_025_705, w_025_706, w_025_707, w_025_708, w_025_709, w_025_710, w_025_711, w_025_712, w_025_713, w_025_715, w_025_716, w_025_717, w_025_718, w_025_719, w_025_720, w_025_721, w_025_722, w_025_723, w_025_724, w_025_725, w_025_726, w_025_727, w_025_728, w_025_729, w_025_730, w_025_731, w_025_732, w_025_733, w_025_734, w_025_735, w_025_736, w_025_737, w_025_738, w_025_739, w_025_740, w_025_741, w_025_742, w_025_743, w_025_744, w_025_745, w_025_746, w_025_747, w_025_748, w_025_749, w_025_751, w_025_752, w_025_753, w_025_754, w_025_755, w_025_756, w_025_757, w_025_758, w_025_759, w_025_760, w_025_761, w_025_762, w_025_763, w_025_764, w_025_765, w_025_766, w_025_767, w_025_768, w_025_769, w_025_770, w_025_771, w_025_772, w_025_773, w_025_774, w_025_775, w_025_776, w_025_777, w_025_778, w_025_779, w_025_780, w_025_781, w_025_782, w_025_783, w_025_784, w_025_785, w_025_786, w_025_787, w_025_788, w_025_789, w_025_791, w_025_792, w_025_793, w_025_794, w_025_795, w_025_796, w_025_797, w_025_798, w_025_800, w_025_801, w_025_802, w_025_803, w_025_804, w_025_805, w_025_806, w_025_807, w_025_808, w_025_809, w_025_810, w_025_811, w_025_812, w_025_813, w_025_814, w_025_815, w_025_816, w_025_817, w_025_819, w_025_820, w_025_821, w_025_822, w_025_823, w_025_824, w_025_825, w_025_826, w_025_827, w_025_828, w_025_829, w_025_830, w_025_831, w_025_832, w_025_833, w_025_834, w_025_835, w_025_836, w_025_837, w_025_838, w_025_839, w_025_840, w_025_841, w_025_842, w_025_843, w_025_844, w_025_845, w_025_846, w_025_847, w_025_848, w_025_849, w_025_850, w_025_851, w_025_852, w_025_853, w_025_854, w_025_855, w_025_856, w_025_857, w_025_858, w_025_859, w_025_860, w_025_861, w_025_862, w_025_863, w_025_864, w_025_865, w_025_867, w_025_868, w_025_869, w_025_870, w_025_871, w_025_872, w_025_873, w_025_874, w_025_875, w_025_876, w_025_877, w_025_878, w_025_879, w_025_880, w_025_881, w_025_882, w_025_883, w_025_884, w_025_885, w_025_886, w_025_887, w_025_888, w_025_889, w_025_890, w_025_891, w_025_892, w_025_893, w_025_894, w_025_895, w_025_896, w_025_897, w_025_898, w_025_899, w_025_900, w_025_901, w_025_903, w_025_904, w_025_905, w_025_906, w_025_907, w_025_908, w_025_909, w_025_910, w_025_912, w_025_913, w_025_914, w_025_915, w_025_916, w_025_917, w_025_918, w_025_919, w_025_920, w_025_921, w_025_922, w_025_924, w_025_925, w_025_926, w_025_927, w_025_928, w_025_929, w_025_930, w_025_931, w_025_932, w_025_933, w_025_934, w_025_935, w_025_936, w_025_937, w_025_938, w_025_939, w_025_940, w_025_941, w_025_942, w_025_943, w_025_944, w_025_945, w_025_946, w_025_947, w_025_948, w_025_949, w_025_950, w_025_951, w_025_952, w_025_953, w_025_955, w_025_956, w_025_957, w_025_958, w_025_959, w_025_960, w_025_961, w_025_962, w_025_963, w_025_964, w_025_965, w_025_966, w_025_967, w_025_968, w_025_969, w_025_970, w_025_971, w_025_972, w_025_973, w_025_974, w_025_975, w_025_977, w_025_978, w_025_979, w_025_980, w_025_981, w_025_982, w_025_983, w_025_984, w_025_985, w_025_986, w_025_987, w_025_988, w_025_989, w_025_990, w_025_992, w_025_993, w_025_994, w_025_995, w_025_996, w_025_997, w_025_998, w_025_999, w_025_1000, w_025_1001, w_025_1002, w_025_1003, w_025_1005, w_025_1006, w_025_1007, w_025_1008, w_025_1009, w_025_1010, w_025_1011, w_025_1012, w_025_1013, w_025_1014, w_025_1015, w_025_1016, w_025_1018, w_025_1019, w_025_1020, w_025_1021, w_025_1022, w_025_1023, w_025_1024, w_025_1025, w_025_1026, w_025_1027, w_025_1028, w_025_1029, w_025_1030, w_025_1031, w_025_1032, w_025_1033, w_025_1034, w_025_1035, w_025_1036, w_025_1037, w_025_1038, w_025_1039, w_025_1040, w_025_1041, w_025_1042, w_025_1043, w_025_1044, w_025_1045, w_025_1046, w_025_1047, w_025_1048, w_025_1049, w_025_1050, w_025_1051, w_025_1052, w_025_1053, w_025_1054, w_025_1055, w_025_1056, w_025_1057, w_025_1058, w_025_1059, w_025_1060, w_025_1061, w_025_1062, w_025_1063, w_025_1064, w_025_1066, w_025_1067, w_025_1068, w_025_1069, w_025_1070, w_025_1071, w_025_1072, w_025_1073, w_025_1074, w_025_1075, w_025_1076, w_025_1077, w_025_1078, w_025_1079, w_025_1080, w_025_1081, w_025_1082, w_025_1083, w_025_1084, w_025_1085, w_025_1086, w_025_1087, w_025_1088, w_025_1089, w_025_1090, w_025_1091, w_025_1092, w_025_1093, w_025_1094, w_025_1095, w_025_1096, w_025_1097, w_025_1098, w_025_1099, w_025_1100, w_025_1101, w_025_1102, w_025_1103, w_025_1104, w_025_1105, w_025_1106, w_025_1107, w_025_1108, w_025_1109, w_025_1110, w_025_1111, w_025_1112, w_025_1113, w_025_1114, w_025_1115, w_025_1116, w_025_1117, w_025_1118, w_025_1119, w_025_1120, w_025_1121, w_025_1122, w_025_1123, w_025_1124, w_025_1125, w_025_1126, w_025_1127, w_025_1128, w_025_1129, w_025_1130, w_025_1131, w_025_1132, w_025_1133, w_025_1134, w_025_1135, w_025_1136, w_025_1137, w_025_1138, w_025_1139, w_025_1140, w_025_1141, w_025_1142, w_025_1143, w_025_1144, w_025_1145, w_025_1146, w_025_1147, w_025_1148, w_025_1149, w_025_1150, w_025_1151, w_025_1152, w_025_1153, w_025_1154, w_025_1155, w_025_1156, w_025_1157, w_025_1158, w_025_1159, w_025_1160, w_025_1161, w_025_1162, w_025_1163, w_025_1164, w_025_1165, w_025_1166, w_025_1167, w_025_1168, w_025_1169, w_025_1170, w_025_1171, w_025_1172, w_025_1173, w_025_1174, w_025_1175, w_025_1176, w_025_1177, w_025_1178, w_025_1179, w_025_1180, w_025_1181, w_025_1182, w_025_1183, w_025_1184, w_025_1186, w_025_1187, w_025_1188, w_025_1189, w_025_1190, w_025_1191, w_025_1192, w_025_1193, w_025_1194, w_025_1195, w_025_1196, w_025_1197, w_025_1198, w_025_1200, w_025_1201, w_025_1202, w_025_1203, w_025_1204, w_025_1206, w_025_1207, w_025_1208, w_025_1209, w_025_1210, w_025_1211, w_025_1212, w_025_1213, w_025_1214, w_025_1215, w_025_1216, w_025_1217, w_025_1218, w_025_1219, w_025_1220, w_025_1221, w_025_1222, w_025_1223, w_025_1224, w_025_1225, w_025_1226, w_025_1227, w_025_1228, w_025_1229, w_025_1231, w_025_1232, w_025_1233, w_025_1234, w_025_1235, w_025_1236, w_025_1237, w_025_1238, w_025_1239, w_025_1240, w_025_1241, w_025_1242, w_025_1243, w_025_1244, w_025_1245, w_025_1246, w_025_1247, w_025_1248, w_025_1249, w_025_1250, w_025_1251, w_025_1252, w_025_1253, w_025_1254, w_025_1255, w_025_1256, w_025_1257, w_025_1258, w_025_1259, w_025_1260, w_025_1261, w_025_1262, w_025_1263, w_025_1264, w_025_1265, w_025_1266, w_025_1267, w_025_1268, w_025_1269, w_025_1270, w_025_1271, w_025_1272, w_025_1273, w_025_1274, w_025_1275, w_025_1276, w_025_1277, w_025_1278, w_025_1279, w_025_1280, w_025_1281, w_025_1282, w_025_1283, w_025_1284, w_025_1285, w_025_1286, w_025_1287, w_025_1288, w_025_1289, w_025_1290, w_025_1291, w_025_1292, w_025_1293, w_025_1294, w_025_1295, w_025_1296, w_025_1297, w_025_1298, w_025_1299, w_025_1300, w_025_1302, w_025_1303, w_025_1304, w_025_1305, w_025_1306, w_025_1307, w_025_1308, w_025_1309, w_025_1310, w_025_1311, w_025_1312, w_025_1313, w_025_1314, w_025_1315, w_025_1316, w_025_1317, w_025_1318, w_025_1319, w_025_1320, w_025_1321, w_025_1322, w_025_1323, w_025_1324, w_025_1325, w_025_1326, w_025_1327, w_025_1328, w_025_1329, w_025_1331, w_025_1332, w_025_1333, w_025_1334, w_025_1335, w_025_1336, w_025_1337, w_025_1338, w_025_1339, w_025_1340, w_025_1341, w_025_1342, w_025_1343, w_025_1344, w_025_1345, w_025_1346, w_025_1347, w_025_1348, w_025_1349, w_025_1350, w_025_1351, w_025_1352, w_025_1353, w_025_1354, w_025_1355, w_025_1356, w_025_1357, w_025_1358, w_025_1359, w_025_1360, w_025_1361, w_025_1362, w_025_1363, w_025_1364, w_025_1365, w_025_1366, w_025_1367, w_025_1368, w_025_1369, w_025_1370, w_025_1371, w_025_1372, w_025_1373, w_025_1374, w_025_1375, w_025_1376, w_025_1377, w_025_1379, w_025_1380, w_025_1381, w_025_1382, w_025_1383, w_025_1384, w_025_1386, w_025_1387, w_025_1390, w_025_1391, w_025_1392, w_025_1393, w_025_1394, w_025_1395, w_025_1396, w_025_1397, w_025_1398, w_025_1399, w_025_1400, w_025_1402, w_025_1403, w_025_1404, w_025_1405, w_025_1406, w_025_1407, w_025_1409, w_025_1410, w_025_1411, w_025_1412, w_025_1413, w_025_1414, w_025_1415, w_025_1417, w_025_1418, w_025_1419, w_025_1420, w_025_1421, w_025_1423, w_025_1424, w_025_1425, w_025_1426, w_025_1427, w_025_1428, w_025_1429, w_025_1430, w_025_1431, w_025_1432, w_025_1433, w_025_1434, w_025_1435, w_025_1436, w_025_1437, w_025_1438, w_025_1439, w_025_1440, w_025_1441, w_025_1442, w_025_1443, w_025_1444, w_025_1445, w_025_1446, w_025_1447, w_025_1448, w_025_1449, w_025_1450, w_025_1451, w_025_1452, w_025_1453, w_025_1454, w_025_1455, w_025_1456, w_025_1457, w_025_1458, w_025_1459, w_025_1460, w_025_1461, w_025_1462, w_025_1463, w_025_1464, w_025_1465, w_025_1466, w_025_1467, w_025_1468, w_025_1469, w_025_1470, w_025_1471, w_025_1472, w_025_1473, w_025_1474, w_025_1477, w_025_1478, w_025_1479, w_025_1480, w_025_1481, w_025_1483, w_025_1484, w_025_1486, w_025_1487, w_025_1488, w_025_1489, w_025_1490, w_025_1491, w_025_1492, w_025_1494, w_025_1495, w_025_1497, w_025_1498, w_025_1499, w_025_1500, w_025_1501, w_025_1502, w_025_1504, w_025_1505, w_025_1506, w_025_1508, w_025_1509, w_025_1510, w_025_1511, w_025_1512, w_025_1513, w_025_1514, w_025_1515, w_025_1516, w_025_1517, w_025_1518, w_025_1519, w_025_1520, w_025_1521, w_025_1522, w_025_1523, w_025_1524, w_025_1525, w_025_1526, w_025_1527, w_025_1528, w_025_1530, w_025_1531, w_025_1532, w_025_1533, w_025_1534, w_025_1535, w_025_1538, w_025_1539, w_025_1540, w_025_1541, w_025_1543, w_025_1544, w_025_1546, w_025_1547, w_025_1548, w_025_1549, w_025_1550, w_025_1551, w_025_1553, w_025_1554, w_025_1555, w_025_1556, w_025_1557, w_025_1558, w_025_1559, w_025_1560, w_025_1561, w_025_1562, w_025_1563, w_025_1565, w_025_1566, w_025_1568, w_025_1569, w_025_1570, w_025_1571, w_025_1572, w_025_1573, w_025_1574, w_025_1575, w_025_1576, w_025_1577, w_025_1578, w_025_1579, w_025_1580, w_025_1582, w_025_1584, w_025_1585, w_025_1586, w_025_1587, w_025_1588, w_025_1589, w_025_1590, w_025_1592, w_025_1593, w_025_1594, w_025_1595, w_025_1597, w_025_1598, w_025_1599, w_025_1600, w_025_1601, w_025_1602, w_025_1603, w_025_1604, w_025_1605, w_025_1606, w_025_1607, w_025_1609, w_025_1610, w_025_1611, w_025_1612, w_025_1613, w_025_1614, w_025_1615, w_025_1616, w_025_1617, w_025_1618, w_025_1619, w_025_1620, w_025_1621, w_025_1622, w_025_1623, w_025_1624, w_025_1625, w_025_1626, w_025_1627, w_025_1628, w_025_1629, w_025_1630, w_025_1632, w_025_1633, w_025_1634, w_025_1635, w_025_1636, w_025_1637, w_025_1638, w_025_1640, w_025_1641, w_025_1642, w_025_1643, w_025_1644, w_025_1645, w_025_1646, w_025_1647, w_025_1648, w_025_1649, w_025_1650, w_025_1651, w_025_1652, w_025_1653, w_025_1654, w_025_1657, w_025_1659, w_025_1660, w_025_1661, w_025_1662, w_025_1663, w_025_1664, w_025_1665, w_025_1666, w_025_1667, w_025_1668, w_025_1669, w_025_1670, w_025_1671, w_025_1672, w_025_1673, w_025_1674, w_025_1675, w_025_1676, w_025_1677, w_025_1678, w_025_1679, w_025_1680, w_025_1681, w_025_1682, w_025_1683, w_025_1686, w_025_1687, w_025_1688, w_025_1689, w_025_1690, w_025_1691, w_025_1692, w_025_1693, w_025_1694, w_025_1695, w_025_1696, w_025_1698, w_025_1699, w_025_1700, w_025_1701, w_025_1702, w_025_1703, w_025_1704, w_025_1706, w_025_1707, w_025_1708, w_025_1709, w_025_1710, w_025_1711, w_025_1712, w_025_1713, w_025_1714, w_025_1715, w_025_1716, w_025_1717, w_025_1718, w_025_1719, w_025_1720, w_025_1721, w_025_1722, w_025_1723, w_025_1724, w_025_1725, w_025_1726, w_025_1727, w_025_1728, w_025_1729, w_025_1730, w_025_1732, w_025_1733, w_025_1735, w_025_1736, w_025_1737, w_025_1738, w_025_1739, w_025_1741, w_025_1742, w_025_1743, w_025_1745, w_025_1746, w_025_1747, w_025_1748, w_025_1749, w_025_1750, w_025_1751, w_025_1752, w_025_1753, w_025_1754, w_025_1755, w_025_1756, w_025_1757, w_025_1758, w_025_1759, w_025_1760, w_025_1761, w_025_1762, w_025_1764, w_025_1765, w_025_1766, w_025_1767, w_025_1768, w_025_1769, w_025_1770, w_025_1771, w_025_1772, w_025_1773, w_025_1774, w_025_1775, w_025_1776, w_025_1777, w_025_1778, w_025_1779, w_025_1780, w_025_1781, w_025_1783, w_025_1784, w_025_1785, w_025_1786, w_025_1787, w_025_1788, w_025_1790, w_025_1791, w_025_1792, w_025_1794, w_025_1795, w_025_1796, w_025_1797, w_025_1798, w_025_1800, w_025_1801, w_025_1802, w_025_1804, w_025_1805, w_025_1806, w_025_1807, w_025_1808, w_025_1809, w_025_1810, w_025_1811, w_025_1812, w_025_1813, w_025_1814, w_025_1815, w_025_1816, w_025_1817;
  wire w_026_000, w_026_001, w_026_002, w_026_003, w_026_004, w_026_005, w_026_006, w_026_007, w_026_008, w_026_009, w_026_010, w_026_012, w_026_013, w_026_014, w_026_015, w_026_016, w_026_017, w_026_018, w_026_019, w_026_020, w_026_021, w_026_022, w_026_023, w_026_024, w_026_025, w_026_026, w_026_027, w_026_028, w_026_029, w_026_030, w_026_031, w_026_032, w_026_033, w_026_034, w_026_035, w_026_036, w_026_037, w_026_039, w_026_040, w_026_041, w_026_042, w_026_043, w_026_044, w_026_045, w_026_046, w_026_047, w_026_049, w_026_050, w_026_051, w_026_052, w_026_053, w_026_054, w_026_055, w_026_056, w_026_057, w_026_059, w_026_060, w_026_061, w_026_062, w_026_063, w_026_064, w_026_065, w_026_066, w_026_067, w_026_068, w_026_069, w_026_070, w_026_071, w_026_072, w_026_073, w_026_075, w_026_076, w_026_077, w_026_078, w_026_079, w_026_080, w_026_081, w_026_082, w_026_083, w_026_084, w_026_085, w_026_086, w_026_087, w_026_088, w_026_089, w_026_090, w_026_091, w_026_092, w_026_093, w_026_094, w_026_095, w_026_096, w_026_097, w_026_098, w_026_100, w_026_101, w_026_102, w_026_103, w_026_104, w_026_105, w_026_106, w_026_107, w_026_108, w_026_109, w_026_111, w_026_112, w_026_113, w_026_114, w_026_115, w_026_116, w_026_117, w_026_118, w_026_119, w_026_120, w_026_122, w_026_123, w_026_124, w_026_125, w_026_126, w_026_127, w_026_128, w_026_129, w_026_130, w_026_131, w_026_132, w_026_133, w_026_135, w_026_136, w_026_137, w_026_138, w_026_139, w_026_140, w_026_141, w_026_142, w_026_143, w_026_144, w_026_145, w_026_146, w_026_147, w_026_148, w_026_149, w_026_150, w_026_151, w_026_152, w_026_153, w_026_154, w_026_156, w_026_157, w_026_158, w_026_159, w_026_160, w_026_161, w_026_162, w_026_163, w_026_164, w_026_165, w_026_166, w_026_167, w_026_168, w_026_169, w_026_170, w_026_171, w_026_172, w_026_173, w_026_174, w_026_175, w_026_176, w_026_177, w_026_178, w_026_179, w_026_180, w_026_181, w_026_182, w_026_183, w_026_184, w_026_185, w_026_186, w_026_187, w_026_188, w_026_189, w_026_190, w_026_191, w_026_192, w_026_193, w_026_194, w_026_195, w_026_196, w_026_197, w_026_198, w_026_199, w_026_200, w_026_201, w_026_202, w_026_203, w_026_204, w_026_205, w_026_206, w_026_207, w_026_208, w_026_209, w_026_210, w_026_211, w_026_212, w_026_213, w_026_214, w_026_215, w_026_216, w_026_217, w_026_218, w_026_219, w_026_220, w_026_221, w_026_222, w_026_223, w_026_224, w_026_225, w_026_226, w_026_227, w_026_228, w_026_229, w_026_230, w_026_231, w_026_232, w_026_233, w_026_234, w_026_235, w_026_236, w_026_237, w_026_238, w_026_239, w_026_240, w_026_241, w_026_242, w_026_243, w_026_244, w_026_245, w_026_246, w_026_247, w_026_248, w_026_249, w_026_250, w_026_251, w_026_252, w_026_253, w_026_254, w_026_255, w_026_256, w_026_257, w_026_258, w_026_259, w_026_260, w_026_261, w_026_262, w_026_263, w_026_264, w_026_265, w_026_266, w_026_267, w_026_268, w_026_269, w_026_270, w_026_271, w_026_272, w_026_273, w_026_274, w_026_275, w_026_276, w_026_277, w_026_278, w_026_279, w_026_280, w_026_281, w_026_282, w_026_283, w_026_284, w_026_285, w_026_286, w_026_287, w_026_288, w_026_290, w_026_291, w_026_292, w_026_293, w_026_294, w_026_295, w_026_297, w_026_298, w_026_299, w_026_300, w_026_301, w_026_302, w_026_303, w_026_304, w_026_305, w_026_306, w_026_307, w_026_308, w_026_309, w_026_310, w_026_311, w_026_312, w_026_313, w_026_314, w_026_315, w_026_316, w_026_317, w_026_318, w_026_319, w_026_320, w_026_321, w_026_323, w_026_325, w_026_326, w_026_327, w_026_328, w_026_329, w_026_330, w_026_331, w_026_332, w_026_333, w_026_334, w_026_335, w_026_336, w_026_337, w_026_339, w_026_340, w_026_341, w_026_343, w_026_345, w_026_346, w_026_347, w_026_348, w_026_349, w_026_350, w_026_351, w_026_352, w_026_353, w_026_354, w_026_355, w_026_356, w_026_357, w_026_358, w_026_359, w_026_360, w_026_361, w_026_362, w_026_364, w_026_365, w_026_366, w_026_367, w_026_368, w_026_369, w_026_370, w_026_371, w_026_372, w_026_373, w_026_374, w_026_375, w_026_376, w_026_377, w_026_378, w_026_380, w_026_381, w_026_382, w_026_383, w_026_384, w_026_385, w_026_386, w_026_387, w_026_388, w_026_389, w_026_390, w_026_391, w_026_392, w_026_393, w_026_394, w_026_395, w_026_396, w_026_397, w_026_399, w_026_400, w_026_401, w_026_402, w_026_403, w_026_404, w_026_405, w_026_406, w_026_407, w_026_408, w_026_409, w_026_410, w_026_411, w_026_412, w_026_413, w_026_414, w_026_415, w_026_416, w_026_417, w_026_418, w_026_419, w_026_420, w_026_421, w_026_423, w_026_424, w_026_425, w_026_426, w_026_427, w_026_428, w_026_429, w_026_430, w_026_431, w_026_432, w_026_433, w_026_434, w_026_436, w_026_438, w_026_439, w_026_440, w_026_441, w_026_442, w_026_443, w_026_444, w_026_445, w_026_446, w_026_447, w_026_448, w_026_449, w_026_450, w_026_451, w_026_452, w_026_453, w_026_454, w_026_455, w_026_456, w_026_457, w_026_458, w_026_459, w_026_460, w_026_461, w_026_463, w_026_464, w_026_465, w_026_466, w_026_467, w_026_468, w_026_469, w_026_470, w_026_471, w_026_472, w_026_473, w_026_474, w_026_475, w_026_476, w_026_477, w_026_478, w_026_480, w_026_481, w_026_482, w_026_483, w_026_484, w_026_485, w_026_486, w_026_487, w_026_489, w_026_490, w_026_491, w_026_493, w_026_494, w_026_495, w_026_496, w_026_497, w_026_498, w_026_499, w_026_500, w_026_501, w_026_503, w_026_504, w_026_505, w_026_506, w_026_507, w_026_508, w_026_510, w_026_511, w_026_512, w_026_514, w_026_515, w_026_516, w_026_517, w_026_518, w_026_519, w_026_520, w_026_521, w_026_522, w_026_523, w_026_525, w_026_526, w_026_527, w_026_528, w_026_529, w_026_530, w_026_531, w_026_532, w_026_533, w_026_534, w_026_535, w_026_536, w_026_538, w_026_539, w_026_540, w_026_542, w_026_543, w_026_544, w_026_546, w_026_547, w_026_549, w_026_550, w_026_551, w_026_552, w_026_553, w_026_554, w_026_556, w_026_557, w_026_558, w_026_559, w_026_560, w_026_561, w_026_562, w_026_563, w_026_564, w_026_565, w_026_566, w_026_567, w_026_568, w_026_569, w_026_570, w_026_571, w_026_572, w_026_573, w_026_574, w_026_575, w_026_576, w_026_577, w_026_578, w_026_579, w_026_580, w_026_581, w_026_582, w_026_583, w_026_584, w_026_585, w_026_586, w_026_587, w_026_588, w_026_589, w_026_590, w_026_591, w_026_592, w_026_593, w_026_594, w_026_595, w_026_596, w_026_597, w_026_598, w_026_599, w_026_600, w_026_601, w_026_602, w_026_603, w_026_605, w_026_606, w_026_607, w_026_608, w_026_609, w_026_610, w_026_611, w_026_612, w_026_613, w_026_615, w_026_616, w_026_617, w_026_618, w_026_619, w_026_620, w_026_621, w_026_622, w_026_623, w_026_624, w_026_625, w_026_626, w_026_627, w_026_629, w_026_630, w_026_631, w_026_632, w_026_633, w_026_634, w_026_636, w_026_638, w_026_639, w_026_640, w_026_641, w_026_642, w_026_643, w_026_644, w_026_645, w_026_646, w_026_647, w_026_648, w_026_649, w_026_650, w_026_652, w_026_653, w_026_654, w_026_655, w_026_656, w_026_657, w_026_658, w_026_659, w_026_660, w_026_661, w_026_662, w_026_663, w_026_664, w_026_665, w_026_666, w_026_667, w_026_668, w_026_669, w_026_670, w_026_671, w_026_672, w_026_674, w_026_675, w_026_676, w_026_677, w_026_678, w_026_679, w_026_680, w_026_681, w_026_682, w_026_683, w_026_684, w_026_685, w_026_686, w_026_687, w_026_688, w_026_689, w_026_690, w_026_691, w_026_692, w_026_693, w_026_694, w_026_695, w_026_697, w_026_698, w_026_699, w_026_700, w_026_701, w_026_702, w_026_703, w_026_704, w_026_706, w_026_707, w_026_708, w_026_709, w_026_710, w_026_711, w_026_712, w_026_714, w_026_715, w_026_716, w_026_717, w_026_718, w_026_719, w_026_720, w_026_721, w_026_722, w_026_723, w_026_724, w_026_725, w_026_726, w_026_727, w_026_728, w_026_729, w_026_730, w_026_731, w_026_732, w_026_733, w_026_734, w_026_736, w_026_737, w_026_738, w_026_740, w_026_741, w_026_742, w_026_743, w_026_744, w_026_745, w_026_746, w_026_747, w_026_748, w_026_749, w_026_750, w_026_751, w_026_752, w_026_755, w_026_756, w_026_757, w_026_759, w_026_760, w_026_761, w_026_762, w_026_763, w_026_764, w_026_766, w_026_767, w_026_768, w_026_769, w_026_770, w_026_771, w_026_772, w_026_773, w_026_774, w_026_775, w_026_776, w_026_777, w_026_778, w_026_779, w_026_780, w_026_781, w_026_783, w_026_784, w_026_785, w_026_786, w_026_787, w_026_788, w_026_789, w_026_790, w_026_792, w_026_793, w_026_794, w_026_795, w_026_798, w_026_799, w_026_800, w_026_801, w_026_802, w_026_803, w_026_804, w_026_805, w_026_806, w_026_807, w_026_808, w_026_809, w_026_811, w_026_812, w_026_813, w_026_814, w_026_815, w_026_816, w_026_817, w_026_818, w_026_819, w_026_820, w_026_821, w_026_822, w_026_823, w_026_824, w_026_825, w_026_826, w_026_827, w_026_830, w_026_831, w_026_832, w_026_833, w_026_834, w_026_835, w_026_836, w_026_837, w_026_838, w_026_839, w_026_840, w_026_841, w_026_842, w_026_843, w_026_844, w_026_845, w_026_847, w_026_848, w_026_849, w_026_850, w_026_851, w_026_852, w_026_854, w_026_855, w_026_856, w_026_857, w_026_858, w_026_859, w_026_861, w_026_862, w_026_863, w_026_864, w_026_865, w_026_866, w_026_867, w_026_868, w_026_869, w_026_870, w_026_871, w_026_872, w_026_873, w_026_874, w_026_875, w_026_876, w_026_877, w_026_878, w_026_879, w_026_880, w_026_881, w_026_882, w_026_883, w_026_884, w_026_885, w_026_886, w_026_888, w_026_889, w_026_890, w_026_891, w_026_892, w_026_893, w_026_894, w_026_895, w_026_897, w_026_898, w_026_899, w_026_900, w_026_901, w_026_902, w_026_904, w_026_905, w_026_906, w_026_907, w_026_909, w_026_910, w_026_911, w_026_912, w_026_913, w_026_914, w_026_915, w_026_916, w_026_918, w_026_919, w_026_920, w_026_922, w_026_923, w_026_925, w_026_926, w_026_927, w_026_928, w_026_929, w_026_930, w_026_931, w_026_932, w_026_933, w_026_934, w_026_935, w_026_936, w_026_937, w_026_938, w_026_939, w_026_940, w_026_941, w_026_942, w_026_943, w_026_944, w_026_945, w_026_946, w_026_947, w_026_948, w_026_949, w_026_950, w_026_952, w_026_953, w_026_954, w_026_956, w_026_957, w_026_958, w_026_959, w_026_960, w_026_961, w_026_962, w_026_963, w_026_964, w_026_965, w_026_966, w_026_967, w_026_968, w_026_969, w_026_970, w_026_971, w_026_972, w_026_973, w_026_974, w_026_975, w_026_976, w_026_977, w_026_978, w_026_979, w_026_980, w_026_981, w_026_982, w_026_983, w_026_984, w_026_985, w_026_986, w_026_988, w_026_989, w_026_990, w_026_992, w_026_993, w_026_994, w_026_995, w_026_996, w_026_997, w_026_998, w_026_999, w_026_1000, w_026_1001, w_026_1002, w_026_1003, w_026_1004, w_026_1005, w_026_1007, w_026_1008, w_026_1009, w_026_1010, w_026_1011, w_026_1013, w_026_1015, w_026_1016, w_026_1017, w_026_1018, w_026_1020, w_026_1021, w_026_1022, w_026_1023, w_026_1025, w_026_1026, w_026_1027, w_026_1029, w_026_1031, w_026_1032, w_026_1033, w_026_1034, w_026_1035, w_026_1038, w_026_1039, w_026_1040, w_026_1041, w_026_1042, w_026_1043, w_026_1044, w_026_1045, w_026_1046, w_026_1047, w_026_1048, w_026_1049, w_026_1050, w_026_1051, w_026_1052, w_026_1053, w_026_1054, w_026_1056, w_026_1057, w_026_1058, w_026_1059, w_026_1060, w_026_1061, w_026_1062, w_026_1063, w_026_1064, w_026_1065, w_026_1066, w_026_1067, w_026_1068, w_026_1069, w_026_1070, w_026_1071, w_026_1072, w_026_1073, w_026_1074, w_026_1075, w_026_1076, w_026_1077, w_026_1078, w_026_1079, w_026_1080, w_026_1081, w_026_1082, w_026_1083, w_026_1084, w_026_1085, w_026_1087, w_026_1088, w_026_1089, w_026_1090, w_026_1091, w_026_1092, w_026_1093, w_026_1095, w_026_1097, w_026_1098, w_026_1100, w_026_1101, w_026_1102, w_026_1103, w_026_1104, w_026_1105, w_026_1106, w_026_1107, w_026_1108, w_026_1109, w_026_1110, w_026_1111, w_026_1112, w_026_1114, w_026_1115, w_026_1116, w_026_1117, w_026_1118, w_026_1119, w_026_1120, w_026_1121, w_026_1124, w_026_1125, w_026_1126, w_026_1127, w_026_1128, w_026_1129, w_026_1130, w_026_1131, w_026_1133, w_026_1134, w_026_1135, w_026_1136, w_026_1137, w_026_1138, w_026_1139, w_026_1140, w_026_1141, w_026_1142, w_026_1143, w_026_1144, w_026_1145, w_026_1146, w_026_1147, w_026_1148, w_026_1149, w_026_1150, w_026_1151, w_026_1152, w_026_1153, w_026_1154, w_026_1156, w_026_1157, w_026_1158, w_026_1159, w_026_1160, w_026_1162, w_026_1163, w_026_1164, w_026_1165, w_026_1167, w_026_1168, w_026_1169, w_026_1170, w_026_1172, w_026_1173, w_026_1174, w_026_1175, w_026_1176, w_026_1177, w_026_1178, w_026_1179, w_026_1180, w_026_1181, w_026_1182, w_026_1183, w_026_1184, w_026_1185, w_026_1186, w_026_1187, w_026_1188, w_026_1189, w_026_1192, w_026_1193, w_026_1194, w_026_1195, w_026_1197, w_026_1198, w_026_1199, w_026_1200, w_026_1202, w_026_1204, w_026_1205, w_026_1206, w_026_1208, w_026_1209, w_026_1210, w_026_1213, w_026_1214, w_026_1215, w_026_1216, w_026_1218, w_026_1219, w_026_1220, w_026_1221, w_026_1222, w_026_1223, w_026_1224, w_026_1225, w_026_1226, w_026_1227, w_026_1228, w_026_1230, w_026_1231, w_026_1232, w_026_1233, w_026_1234, w_026_1235, w_026_1236, w_026_1237, w_026_1238, w_026_1239, w_026_1240, w_026_1241, w_026_1242, w_026_1243, w_026_1244, w_026_1245, w_026_1246, w_026_1247, w_026_1248, w_026_1249, w_026_1250, w_026_1251, w_026_1253, w_026_1254, w_026_1255, w_026_1256, w_026_1257, w_026_1258, w_026_1259, w_026_1260, w_026_1261, w_026_1262, w_026_1263, w_026_1264, w_026_1265, w_026_1266, w_026_1267, w_026_1268, w_026_1269, w_026_1270, w_026_1271, w_026_1272, w_026_1273, w_026_1274, w_026_1275, w_026_1276, w_026_1277, w_026_1280, w_026_1281, w_026_1282, w_026_1283, w_026_1285, w_026_1286, w_026_1287, w_026_1289, w_026_1290, w_026_1291, w_026_1292, w_026_1294, w_026_1295, w_026_1296, w_026_1297, w_026_1299, w_026_1300, w_026_1301, w_026_1302, w_026_1303, w_026_1304, w_026_1305, w_026_1306, w_026_1307, w_026_1308, w_026_1310, w_026_1311, w_026_1312, w_026_1313, w_026_1314, w_026_1315, w_026_1316, w_026_1317, w_026_1318, w_026_1319, w_026_1320, w_026_1321, w_026_1322, w_026_1323, w_026_1324, w_026_1325, w_026_1326, w_026_1328, w_026_1329, w_026_1330, w_026_1331, w_026_1332, w_026_1333, w_026_1334, w_026_1335, w_026_1336, w_026_1337, w_026_1338, w_026_1339, w_026_1340, w_026_1341, w_026_1342, w_026_1344, w_026_1345, w_026_1346, w_026_1347, w_026_1348, w_026_1349, w_026_1350, w_026_1352, w_026_1353, w_026_1354, w_026_1355, w_026_1357, w_026_1359, w_026_1360, w_026_1361, w_026_1362, w_026_1363, w_026_1364, w_026_1365, w_026_1367, w_026_1368, w_026_1369, w_026_1371, w_026_1372, w_026_1373, w_026_1374, w_026_1375, w_026_1376, w_026_1377, w_026_1378, w_026_1379, w_026_1380, w_026_1381, w_026_1382, w_026_1383, w_026_1384, w_026_1385, w_026_1386, w_026_1387, w_026_1388, w_026_1390, w_026_1391, w_026_1392, w_026_1394, w_026_1395, w_026_1396, w_026_1397, w_026_1398, w_026_1399, w_026_1401, w_026_1403, w_026_1404, w_026_1405, w_026_1407, w_026_1408, w_026_1409, w_026_1410, w_026_1411, w_026_1412, w_026_1413, w_026_1414, w_026_1415, w_026_1416, w_026_1417, w_026_1418, w_026_1419, w_026_1420, w_026_1421, w_026_1422, w_026_1424, w_026_1425, w_026_1427, w_026_1428, w_026_1429, w_026_1430, w_026_1431, w_026_1432, w_026_1433, w_026_1434, w_026_1435, w_026_1436, w_026_1437, w_026_1438, w_026_1439, w_026_1441, w_026_1442, w_026_1443, w_026_1444, w_026_1445, w_026_1446, w_026_1447, w_026_1448, w_026_1449, w_026_1450, w_026_1451, w_026_1452, w_026_1453, w_026_1455, w_026_1456, w_026_1457, w_026_1458, w_026_1459, w_026_1460, w_026_1461, w_026_1462, w_026_1463, w_026_1465, w_026_1466, w_026_1467, w_026_1468, w_026_1470, w_026_1471, w_026_1472, w_026_1473, w_026_1474, w_026_1476, w_026_1477, w_026_1478, w_026_1479, w_026_1480, w_026_1481, w_026_1482, w_026_1483, w_026_1484, w_026_1485, w_026_1486, w_026_1487, w_026_1489, w_026_1490, w_026_1491, w_026_1492, w_026_1495, w_026_1496, w_026_1497, w_026_1498, w_026_1499, w_026_1500, w_026_1502, w_026_1503, w_026_1504, w_026_1505, w_026_1506, w_026_1507, w_026_1508, w_026_1509, w_026_1510, w_026_1511, w_026_1513, w_026_1514, w_026_1515, w_026_1516, w_026_1517, w_026_1518, w_026_1519, w_026_1520, w_026_1521, w_026_1522, w_026_1523, w_026_1524, w_026_1525, w_026_1526, w_026_1527, w_026_1528, w_026_1529, w_026_1530, w_026_1531, w_026_1532, w_026_1533, w_026_1534, w_026_1535, w_026_1536, w_026_1537, w_026_1539, w_026_1540, w_026_1541, w_026_1542, w_026_1544, w_026_1545, w_026_1546, w_026_1548, w_026_1549, w_026_1551, w_026_1552, w_026_1553, w_026_1555, w_026_1556, w_026_1557, w_026_1558, w_026_1559, w_026_1560, w_026_1561, w_026_1562, w_026_1563, w_026_1564, w_026_1566, w_026_1567, w_026_1568, w_026_1569, w_026_1570, w_026_1571, w_026_1573, w_026_1574, w_026_1575, w_026_1576, w_026_1577, w_026_1578, w_026_1579, w_026_1580, w_026_1581, w_026_1582, w_026_1583, w_026_1584, w_026_1585, w_026_1587, w_026_1588, w_026_1590, w_026_1592, w_026_1593, w_026_1594, w_026_1595, w_026_1598, w_026_1599, w_026_1600, w_026_1601, w_026_1602, w_026_1604, w_026_1605, w_026_1606, w_026_1607, w_026_1608, w_026_1609, w_026_1610, w_026_1611, w_026_1612, w_026_1613, w_026_1614, w_026_1616, w_026_1617, w_026_1618, w_026_1619, w_026_1620, w_026_1621, w_026_1622, w_026_1623, w_026_1624, w_026_1625, w_026_1626, w_026_1627, w_026_1628, w_026_1629, w_026_1630, w_026_1632, w_026_1633, w_026_1634, w_026_1635, w_026_1636, w_026_1637, w_026_1638, w_026_1639, w_026_1640, w_026_1641, w_026_1642, w_026_1643, w_026_1644, w_026_1645, w_026_1646, w_026_1648, w_026_1649, w_026_1650, w_026_1652, w_026_1653, w_026_1654, w_026_1655, w_026_1656, w_026_1657, w_026_1658, w_026_1659, w_026_1660, w_026_1661, w_026_1662, w_026_1663, w_026_1665, w_026_1666, w_026_1667, w_026_1668, w_026_1669, w_026_1670, w_026_1671, w_026_1672, w_026_1673, w_026_1674, w_026_1675, w_026_1676, w_026_1677, w_026_1678, w_026_1679, w_026_1680, w_026_1681, w_026_1682, w_026_1683, w_026_1686, w_026_1687, w_026_1688, w_026_1689, w_026_1690, w_026_1691, w_026_1692, w_026_1693, w_026_1696, w_026_1697, w_026_1698, w_026_1699, w_026_1701, w_026_1703, w_026_1704, w_026_1705, w_026_1706, w_026_1707, w_026_1708, w_026_1709, w_026_1710, w_026_1711, w_026_1713, w_026_1714, w_026_1715, w_026_1718, w_026_1719, w_026_1720, w_026_1721, w_026_1722, w_026_1723, w_026_1724, w_026_1725, w_026_1726, w_026_1727, w_026_1728, w_026_1730, w_026_1731, w_026_1732, w_026_1733, w_026_1734, w_026_1735, w_026_1736, w_026_1737, w_026_1738, w_026_1739, w_026_1740, w_026_1741, w_026_1743, w_026_1744, w_026_1745, w_026_1746, w_026_1747, w_026_1748, w_026_1750, w_026_1751, w_026_1752, w_026_1754, w_026_1755, w_026_1756, w_026_1757, w_026_1758, w_026_1759, w_026_1760, w_026_1761, w_026_1763, w_026_1765, w_026_1766, w_026_1768, w_026_1769, w_026_1770, w_026_1771, w_026_1772, w_026_1773, w_026_1774, w_026_1776, w_026_1777, w_026_1778, w_026_1779, w_026_1780, w_026_1781, w_026_1782, w_026_1783, w_026_1784, w_026_1785, w_026_1786, w_026_1787, w_026_1788, w_026_1790, w_026_1791, w_026_1792, w_026_1793, w_026_1794, w_026_1795, w_026_1797, w_026_1798, w_026_1799, w_026_1800, w_026_1801, w_026_1802, w_026_1803, w_026_1804, w_026_1806, w_026_1807, w_026_1808, w_026_1809, w_026_1812, w_026_1813, w_026_1814, w_026_1815, w_026_1816, w_026_1817, w_026_1818, w_026_1819, w_026_1820, w_026_1821, w_026_1822, w_026_1823, w_026_1824, w_026_1825, w_026_1827, w_026_1828, w_026_1829, w_026_1830, w_026_1831, w_026_1832, w_026_1833, w_026_1834, w_026_1835, w_026_1836, w_026_1837, w_026_1838, w_026_1839, w_026_1840, w_026_1841, w_026_1842, w_026_1843, w_026_1845, w_026_1846, w_026_1847, w_026_1848, w_026_1849, w_026_1850, w_026_1851, w_026_1852, w_026_1853, w_026_1854, w_026_1855, w_026_1856, w_026_1857, w_026_1858, w_026_1859, w_026_1860, w_026_1861, w_026_1862, w_026_1863, w_026_1864, w_026_1865, w_026_1866, w_026_1867, w_026_1869, w_026_1870, w_026_1871, w_026_1872, w_026_1873, w_026_1874, w_026_1875, w_026_1877, w_026_1878, w_026_1879, w_026_1881, w_026_1882, w_026_1883, w_026_1885, w_026_1886, w_026_1888, w_026_1889, w_026_1890, w_026_1891, w_026_1892, w_026_1893, w_026_1894, w_026_1895, w_026_1896, w_026_1898, w_026_1899, w_026_1900, w_026_1901, w_026_1902, w_026_1903, w_026_1904, w_026_1905, w_026_1906, w_026_1907, w_026_1908, w_026_1909, w_026_1910, w_026_1911, w_026_1912, w_026_1913, w_026_1914, w_026_1915, w_026_1916, w_026_1917, w_026_1918, w_026_1919, w_026_1920, w_026_1922, w_026_1923, w_026_1924, w_026_1925, w_026_1926, w_026_1928, w_026_1929, w_026_1930, w_026_1931, w_026_1932, w_026_1933, w_026_1935, w_026_1937, w_026_1938, w_026_1939, w_026_1940, w_026_1942, w_026_1943, w_026_1944, w_026_1945, w_026_1946, w_026_1947, w_026_1948, w_026_1949, w_026_1950, w_026_1952, w_026_1953, w_026_1954, w_026_1955, w_026_1956, w_026_1957, w_026_1958, w_026_1959, w_026_1960, w_026_1961, w_026_1962, w_026_1963, w_026_1964, w_026_1965, w_026_1966, w_026_1967, w_026_1968, w_026_1969, w_026_1970, w_026_1971, w_026_1972, w_026_1973, w_026_1974, w_026_1975, w_026_1976, w_026_1978, w_026_1979, w_026_1980, w_026_1981, w_026_1982, w_026_1984, w_026_1985, w_026_1986, w_026_1987, w_026_1988, w_026_1989, w_026_1990, w_026_1991, w_026_1993, w_026_1994, w_026_1995, w_026_1996, w_026_1997, w_026_1998, w_026_1999, w_026_2000, w_026_2001, w_026_2002, w_026_2003, w_026_2004, w_026_2005, w_026_2006, w_026_2007, w_026_2008, w_026_2010, w_026_2011, w_026_2012, w_026_2013, w_026_2014, w_026_2015, w_026_2016, w_026_2017, w_026_2018, w_026_2019, w_026_2020, w_026_2021, w_026_2022, w_026_2023, w_026_2025, w_026_2026, w_026_2027, w_026_2028, w_026_2029, w_026_2030, w_026_2031, w_026_2032, w_026_2033, w_026_2034, w_026_2035, w_026_2036, w_026_2037, w_026_2038, w_026_2039, w_026_2040, w_026_2041, w_026_2042, w_026_2043, w_026_2044, w_026_2045, w_026_2046, w_026_2047, w_026_2048, w_026_2049, w_026_2050, w_026_2052, w_026_2053, w_026_2054, w_026_2055, w_026_2056, w_026_2057, w_026_2058, w_026_2059, w_026_2060, w_026_2061, w_026_2062, w_026_2063, w_026_2064, w_026_2066, w_026_2067, w_026_2068, w_026_2069, w_026_2070, w_026_2071, w_026_2072, w_026_2074, w_026_2075, w_026_2076, w_026_2077, w_026_2078, w_026_2079, w_026_2080, w_026_2081, w_026_2082, w_026_2083, w_026_2084, w_026_2085, w_026_2086, w_026_2087, w_026_2089, w_026_2090, w_026_2091, w_026_2092, w_026_2093, w_026_2094, w_026_2095, w_026_2096, w_026_2099, w_026_2101, w_026_2102, w_026_2103, w_026_2104, w_026_2105, w_026_2107, w_026_2108, w_026_2109, w_026_2110, w_026_2111, w_026_2112, w_026_2113, w_026_2114, w_026_2115, w_026_2116, w_026_2117, w_026_2118, w_026_2119, w_026_2121, w_026_2122, w_026_2123, w_026_2125, w_026_2126, w_026_2128, w_026_2129, w_026_2130, w_026_2132, w_026_2133, w_026_2134, w_026_2135, w_026_2136, w_026_2137, w_026_2139, w_026_2140, w_026_2141, w_026_2142, w_026_2143, w_026_2144, w_026_2145, w_026_2146, w_026_2147, w_026_2148, w_026_2149, w_026_2150, w_026_2151, w_026_2152, w_026_2153, w_026_2154, w_026_2156, w_026_2157, w_026_2159, w_026_2160, w_026_2161, w_026_2163, w_026_2164, w_026_2165, w_026_2166, w_026_2167, w_026_2168, w_026_2169, w_026_2170, w_026_2171, w_026_2173, w_026_2175, w_026_2176, w_026_2177, w_026_2178, w_026_2179, w_026_2180, w_026_2181, w_026_2182, w_026_2184, w_026_2185, w_026_2186, w_026_2187, w_026_2188, w_026_2189, w_026_2190, w_026_2191, w_026_2194, w_026_2195, w_026_2196, w_026_2199, w_026_2201, w_026_2203, w_026_2204, w_026_2205, w_026_2206, w_026_2207, w_026_2208, w_026_2210, w_026_2211, w_026_2212, w_026_2213, w_026_2214, w_026_2215, w_026_2216, w_026_2217, w_026_2218, w_026_2219, w_026_2220, w_026_2221, w_026_2222, w_026_2223, w_026_2224, w_026_2225, w_026_2226, w_026_2227, w_026_2228, w_026_2229, w_026_2230, w_026_2231, w_026_2232, w_026_2233, w_026_2235, w_026_2236, w_026_2237, w_026_2238, w_026_2239, w_026_2241, w_026_2242, w_026_2243, w_026_2244, w_026_2245, w_026_2246, w_026_2247, w_026_2248, w_026_2249, w_026_2254, w_026_2255, w_026_2256, w_026_2257, w_026_2258, w_026_2259, w_026_2260, w_026_2261, w_026_2263, w_026_2264, w_026_2265, w_026_2266, w_026_2267, w_026_2272, w_026_2273, w_026_2274, w_026_2275, w_026_2276, w_026_2277, w_026_2278, w_026_2279, w_026_2280, w_026_2281, w_026_2282, w_026_2283, w_026_2284, w_026_2285, w_026_2288, w_026_2289, w_026_2290, w_026_2291, w_026_2292, w_026_2293, w_026_2294, w_026_2296, w_026_2297, w_026_2298, w_026_2299, w_026_2300, w_026_2301, w_026_2302, w_026_2303, w_026_2304, w_026_2305, w_026_2306, w_026_2307, w_026_2308, w_026_2309, w_026_2310, w_026_2311, w_026_2312, w_026_2313, w_026_2314, w_026_2315, w_026_2316, w_026_2317, w_026_2318, w_026_2319, w_026_2320, w_026_2321, w_026_2322, w_026_2323, w_026_2324, w_026_2326, w_026_2327, w_026_2329, w_026_2330, w_026_2331, w_026_2332, w_026_2333, w_026_2334, w_026_2335, w_026_2336, w_026_2337, w_026_2338, w_026_2339, w_026_2340, w_026_2341, w_026_2342, w_026_2343, w_026_2344, w_026_2345, w_026_2346, w_026_2348, w_026_2349, w_026_2350, w_026_2351, w_026_2352, w_026_2354, w_026_2356, w_026_2357, w_026_2358, w_026_2359, w_026_2360, w_026_2361, w_026_2362, w_026_2363, w_026_2364, w_026_2367;
  wire w_027_000, w_027_001, w_027_002, w_027_003, w_027_004, w_027_005, w_027_006, w_027_007, w_027_008, w_027_009, w_027_010, w_027_011, w_027_012, w_027_013, w_027_014, w_027_015, w_027_016, w_027_017, w_027_018, w_027_019, w_027_020, w_027_021, w_027_022, w_027_023, w_027_024, w_027_025, w_027_026, w_027_027, w_027_028, w_027_029, w_027_030, w_027_031, w_027_032, w_027_033, w_027_034, w_027_035, w_027_036, w_027_037, w_027_038, w_027_039, w_027_040, w_027_041, w_027_042, w_027_043, w_027_044, w_027_045, w_027_046, w_027_047, w_027_048, w_027_049, w_027_050, w_027_051, w_027_052, w_027_053, w_027_054, w_027_055, w_027_056, w_027_057, w_027_058, w_027_059, w_027_060, w_027_061, w_027_062, w_027_063, w_027_064, w_027_065, w_027_066, w_027_067, w_027_068, w_027_069, w_027_070, w_027_071, w_027_072, w_027_073, w_027_074, w_027_075, w_027_076, w_027_077, w_027_078, w_027_079, w_027_080, w_027_081, w_027_082, w_027_083, w_027_084, w_027_085, w_027_086, w_027_087, w_027_088, w_027_089, w_027_091, w_027_092, w_027_093, w_027_094, w_027_095, w_027_096, w_027_097, w_027_098, w_027_099, w_027_100, w_027_101, w_027_102, w_027_103, w_027_104, w_027_105, w_027_106, w_027_107, w_027_108, w_027_109, w_027_110, w_027_111, w_027_112, w_027_113, w_027_114, w_027_115, w_027_116, w_027_117, w_027_119, w_027_120, w_027_121, w_027_122, w_027_123, w_027_124, w_027_125, w_027_126, w_027_127, w_027_128, w_027_129, w_027_130, w_027_131, w_027_132, w_027_133, w_027_134, w_027_135, w_027_136, w_027_137, w_027_138, w_027_139, w_027_140, w_027_141, w_027_142, w_027_143, w_027_144, w_027_145, w_027_146, w_027_147, w_027_148, w_027_149, w_027_150, w_027_151, w_027_152, w_027_153, w_027_154, w_027_155, w_027_156, w_027_157, w_027_158, w_027_159, w_027_160, w_027_161, w_027_162, w_027_163, w_027_165, w_027_166, w_027_168, w_027_169, w_027_170, w_027_171, w_027_172, w_027_173, w_027_174, w_027_175, w_027_176, w_027_177, w_027_179, w_027_180, w_027_181, w_027_182, w_027_183, w_027_184, w_027_185, w_027_186, w_027_187, w_027_188, w_027_189, w_027_190, w_027_191, w_027_192, w_027_193, w_027_194, w_027_195, w_027_196, w_027_197, w_027_198, w_027_199, w_027_200, w_027_201, w_027_202, w_027_203, w_027_204, w_027_205, w_027_206, w_027_207, w_027_208, w_027_209, w_027_210, w_027_211, w_027_212, w_027_213, w_027_214, w_027_215, w_027_216, w_027_217, w_027_218, w_027_219, w_027_220, w_027_221, w_027_222, w_027_223, w_027_224, w_027_225, w_027_226, w_027_227, w_027_228, w_027_229, w_027_231, w_027_233, w_027_234, w_027_235, w_027_236, w_027_237, w_027_239, w_027_240, w_027_241, w_027_242, w_027_243, w_027_244, w_027_245, w_027_246, w_027_247, w_027_248, w_027_249, w_027_250, w_027_251, w_027_252, w_027_253, w_027_254, w_027_255, w_027_256, w_027_257, w_027_259, w_027_260, w_027_261, w_027_262, w_027_263, w_027_264, w_027_265, w_027_266, w_027_267, w_027_268, w_027_269, w_027_270, w_027_271, w_027_272, w_027_274, w_027_275, w_027_276, w_027_277, w_027_278, w_027_279, w_027_280, w_027_281, w_027_282, w_027_283, w_027_284, w_027_285, w_027_286, w_027_287, w_027_288, w_027_289, w_027_291, w_027_292, w_027_293, w_027_295, w_027_296, w_027_297, w_027_298, w_027_299, w_027_301, w_027_302, w_027_303, w_027_304, w_027_305, w_027_306, w_027_307, w_027_308, w_027_309, w_027_310, w_027_311, w_027_312, w_027_313, w_027_314, w_027_315, w_027_316, w_027_317, w_027_318, w_027_319, w_027_320, w_027_321, w_027_322, w_027_323, w_027_324, w_027_325, w_027_326, w_027_327, w_027_328, w_027_329, w_027_330, w_027_331, w_027_332, w_027_333, w_027_334, w_027_335, w_027_336, w_027_337, w_027_338, w_027_339, w_027_340, w_027_341, w_027_342, w_027_343, w_027_344, w_027_345, w_027_347, w_027_348, w_027_349, w_027_350, w_027_351, w_027_352, w_027_353, w_027_354, w_027_355, w_027_356, w_027_357, w_027_358, w_027_359, w_027_360, w_027_361, w_027_362, w_027_363, w_027_364, w_027_365, w_027_366, w_027_367, w_027_368, w_027_369, w_027_370, w_027_371, w_027_372, w_027_373, w_027_374, w_027_375, w_027_376, w_027_377, w_027_378, w_027_379, w_027_380, w_027_382, w_027_383, w_027_384, w_027_385, w_027_386, w_027_387, w_027_388, w_027_389, w_027_390, w_027_391, w_027_392, w_027_393, w_027_394, w_027_395, w_027_396, w_027_397, w_027_398, w_027_399, w_027_400, w_027_401, w_027_402, w_027_403, w_027_404, w_027_405, w_027_406, w_027_407, w_027_408, w_027_409, w_027_410, w_027_411, w_027_412, w_027_413, w_027_414, w_027_415, w_027_416, w_027_417, w_027_418, w_027_419, w_027_420, w_027_421, w_027_422, w_027_423, w_027_424, w_027_425, w_027_426, w_027_427, w_027_428, w_027_429, w_027_430, w_027_431, w_027_432, w_027_433, w_027_434, w_027_435, w_027_436, w_027_437, w_027_438, w_027_439, w_027_440, w_027_441, w_027_442, w_027_443, w_027_444, w_027_445, w_027_446, w_027_447, w_027_448, w_027_449, w_027_450, w_027_451, w_027_452, w_027_453, w_027_454, w_027_455, w_027_456, w_027_457, w_027_458, w_027_459, w_027_460, w_027_461, w_027_462, w_027_463, w_027_465, w_027_466, w_027_467, w_027_468, w_027_469, w_027_470, w_027_471, w_027_472, w_027_473, w_027_474, w_027_475, w_027_476, w_027_477, w_027_478, w_027_479, w_027_480, w_027_481, w_027_482, w_027_483, w_027_484, w_027_485, w_027_486, w_027_487, w_027_488, w_027_489, w_027_490, w_027_491, w_027_492, w_027_493, w_027_494, w_027_495, w_027_496, w_027_497, w_027_498, w_027_499, w_027_500, w_027_501, w_027_503, w_027_504, w_027_505, w_027_506, w_027_507, w_027_508, w_027_509, w_027_510, w_027_511, w_027_512, w_027_513, w_027_514, w_027_515, w_027_516, w_027_517, w_027_518, w_027_520, w_027_521, w_027_522, w_027_523, w_027_524, w_027_525, w_027_526, w_027_527, w_027_528, w_027_529, w_027_530, w_027_531, w_027_532, w_027_533, w_027_534, w_027_535, w_027_536, w_027_538, w_027_539, w_027_540, w_027_541, w_027_542, w_027_543, w_027_544, w_027_545, w_027_546, w_027_547, w_027_548, w_027_549, w_027_550, w_027_551, w_027_552, w_027_553, w_027_554, w_027_555, w_027_556, w_027_557, w_027_558, w_027_559, w_027_560, w_027_561, w_027_563, w_027_564, w_027_565, w_027_566, w_027_567, w_027_568, w_027_569, w_027_570, w_027_572, w_027_573, w_027_574, w_027_575, w_027_576, w_027_577, w_027_579, w_027_580, w_027_581, w_027_582, w_027_583, w_027_584, w_027_585, w_027_586, w_027_587, w_027_589, w_027_590, w_027_591, w_027_592, w_027_593, w_027_594, w_027_595, w_027_596, w_027_597, w_027_598, w_027_599, w_027_600, w_027_601, w_027_602, w_027_603, w_027_604, w_027_605, w_027_606, w_027_607, w_027_608, w_027_609, w_027_611, w_027_612, w_027_613, w_027_614, w_027_615, w_027_616, w_027_618, w_027_619, w_027_620, w_027_621, w_027_622, w_027_623, w_027_624, w_027_625, w_027_626, w_027_627, w_027_628, w_027_629, w_027_630, w_027_631, w_027_632, w_027_634, w_027_635, w_027_636, w_027_637, w_027_638, w_027_639, w_027_640, w_027_641, w_027_642, w_027_643, w_027_644, w_027_645, w_027_646, w_027_647, w_027_648, w_027_649, w_027_650, w_027_652, w_027_653, w_027_654, w_027_655, w_027_656, w_027_657, w_027_658, w_027_659, w_027_660, w_027_661, w_027_662, w_027_664, w_027_665, w_027_666, w_027_667, w_027_668, w_027_669, w_027_670, w_027_671, w_027_672, w_027_673, w_027_674, w_027_675, w_027_676, w_027_677, w_027_678, w_027_679, w_027_680, w_027_681, w_027_682, w_027_683, w_027_684, w_027_685, w_027_686, w_027_687, w_027_688, w_027_689, w_027_690, w_027_691, w_027_692, w_027_693, w_027_694, w_027_695, w_027_696, w_027_697, w_027_698, w_027_699, w_027_700, w_027_701, w_027_702, w_027_703, w_027_704, w_027_705, w_027_706, w_027_707, w_027_708, w_027_709, w_027_710, w_027_711, w_027_712, w_027_713, w_027_714, w_027_715, w_027_716, w_027_717, w_027_718, w_027_719, w_027_720, w_027_721, w_027_722, w_027_723, w_027_724, w_027_725, w_027_726, w_027_727, w_027_728, w_027_729, w_027_730, w_027_731, w_027_732, w_027_733, w_027_734, w_027_735, w_027_736, w_027_737, w_027_738, w_027_739, w_027_740, w_027_741, w_027_742, w_027_743, w_027_744, w_027_745, w_027_746, w_027_747, w_027_748, w_027_749, w_027_750, w_027_751, w_027_752, w_027_753, w_027_754, w_027_755, w_027_756, w_027_757, w_027_758, w_027_759, w_027_760, w_027_761, w_027_762, w_027_763, w_027_764, w_027_765, w_027_766, w_027_767, w_027_768, w_027_769, w_027_770, w_027_771, w_027_772, w_027_773, w_027_774, w_027_775, w_027_776, w_027_777, w_027_778, w_027_779, w_027_780, w_027_781, w_027_782, w_027_783, w_027_784, w_027_785, w_027_786, w_027_787, w_027_788, w_027_789, w_027_790, w_027_791, w_027_792, w_027_793, w_027_794, w_027_795, w_027_796, w_027_797, w_027_798, w_027_799, w_027_800, w_027_801, w_027_802, w_027_803, w_027_804, w_027_805, w_027_806, w_027_807, w_027_808, w_027_809, w_027_810, w_027_811, w_027_812, w_027_813, w_027_814, w_027_815, w_027_816, w_027_817, w_027_818, w_027_819, w_027_820, w_027_821, w_027_822, w_027_823, w_027_824, w_027_826, w_027_827, w_027_828, w_027_829, w_027_830, w_027_831, w_027_832, w_027_833, w_027_834, w_027_835, w_027_836, w_027_837, w_027_838, w_027_840, w_027_841, w_027_842, w_027_843, w_027_844, w_027_845, w_027_846, w_027_847, w_027_849, w_027_850, w_027_851, w_027_852, w_027_853, w_027_854, w_027_855, w_027_856, w_027_857, w_027_858, w_027_859, w_027_860, w_027_861, w_027_862, w_027_863, w_027_864, w_027_865, w_027_866, w_027_867, w_027_868, w_027_869, w_027_870, w_027_871, w_027_872, w_027_873, w_027_874, w_027_875, w_027_876, w_027_877, w_027_878, w_027_879, w_027_880, w_027_881, w_027_882, w_027_883, w_027_884, w_027_885, w_027_886, w_027_887, w_027_888, w_027_889, w_027_890, w_027_892, w_027_893, w_027_894, w_027_896, w_027_897, w_027_898, w_027_899, w_027_900, w_027_901, w_027_902, w_027_903, w_027_904, w_027_905, w_027_906, w_027_908, w_027_909, w_027_910, w_027_911, w_027_912, w_027_913, w_027_914, w_027_915, w_027_916, w_027_917, w_027_918, w_027_919, w_027_920, w_027_921, w_027_922, w_027_923, w_027_924, w_027_925, w_027_926, w_027_928, w_027_929, w_027_930, w_027_931, w_027_932, w_027_933, w_027_934, w_027_935, w_027_936, w_027_937, w_027_938, w_027_939, w_027_940, w_027_941, w_027_942, w_027_943, w_027_944, w_027_945, w_027_946, w_027_947, w_027_948, w_027_949, w_027_950, w_027_951, w_027_952, w_027_953, w_027_954, w_027_955, w_027_956, w_027_957, w_027_958, w_027_959, w_027_960, w_027_961, w_027_962, w_027_963, w_027_964, w_027_965, w_027_966, w_027_967, w_027_968, w_027_969, w_027_970, w_027_971, w_027_972, w_027_973, w_027_974, w_027_975, w_027_976, w_027_977, w_027_978, w_027_979, w_027_980, w_027_981, w_027_982, w_027_983, w_027_984, w_027_985, w_027_986, w_027_987, w_027_988, w_027_989, w_027_990, w_027_992, w_027_993, w_027_994, w_027_995, w_027_996, w_027_997, w_027_998, w_027_999, w_027_1000, w_027_1001, w_027_1002, w_027_1003, w_027_1004, w_027_1005, w_027_1006, w_027_1007, w_027_1008, w_027_1009, w_027_1010, w_027_1011, w_027_1012, w_027_1013, w_027_1014, w_027_1015, w_027_1016, w_027_1017, w_027_1018, w_027_1019, w_027_1020, w_027_1021, w_027_1022, w_027_1023, w_027_1024, w_027_1025, w_027_1026, w_027_1027, w_027_1028, w_027_1029, w_027_1030, w_027_1031, w_027_1032, w_027_1033, w_027_1034, w_027_1035, w_027_1036, w_027_1037, w_027_1039, w_027_1040, w_027_1041, w_027_1042, w_027_1043, w_027_1044, w_027_1045, w_027_1046, w_027_1047, w_027_1048, w_027_1049, w_027_1050, w_027_1051, w_027_1052, w_027_1053, w_027_1054, w_027_1055, w_027_1056, w_027_1057, w_027_1058, w_027_1059, w_027_1060, w_027_1061, w_027_1062, w_027_1063, w_027_1064, w_027_1065, w_027_1066, w_027_1067, w_027_1068, w_027_1069, w_027_1070, w_027_1071, w_027_1072, w_027_1073, w_027_1074, w_027_1075, w_027_1076, w_027_1077, w_027_1078, w_027_1079, w_027_1080, w_027_1081, w_027_1082, w_027_1083, w_027_1084, w_027_1085, w_027_1086, w_027_1087, w_027_1088, w_027_1089, w_027_1090, w_027_1091, w_027_1092, w_027_1093, w_027_1094, w_027_1095, w_027_1096, w_027_1097, w_027_1098, w_027_1099, w_027_1100, w_027_1101, w_027_1102, w_027_1103, w_027_1105, w_027_1106, w_027_1107, w_027_1108, w_027_1109, w_027_1110, w_027_1111, w_027_1112, w_027_1113, w_027_1114, w_027_1115, w_027_1116, w_027_1117, w_027_1118, w_027_1119, w_027_1120, w_027_1121, w_027_1122, w_027_1123, w_027_1124, w_027_1125, w_027_1126, w_027_1127, w_027_1128, w_027_1129, w_027_1130, w_027_1131, w_027_1132, w_027_1133, w_027_1134, w_027_1135, w_027_1136, w_027_1137, w_027_1138, w_027_1139, w_027_1140, w_027_1141, w_027_1142, w_027_1143, w_027_1144, w_027_1145, w_027_1146, w_027_1147, w_027_1148, w_027_1149, w_027_1150, w_027_1151, w_027_1152, w_027_1153, w_027_1154, w_027_1155, w_027_1156, w_027_1157, w_027_1158, w_027_1159, w_027_1160, w_027_1161, w_027_1162, w_027_1163, w_027_1164, w_027_1165, w_027_1166, w_027_1167, w_027_1168, w_027_1169, w_027_1170, w_027_1171, w_027_1174, w_027_1175, w_027_1176, w_027_1177, w_027_1178, w_027_1179, w_027_1180, w_027_1181, w_027_1182, w_027_1183, w_027_1184, w_027_1185, w_027_1186, w_027_1187, w_027_1188, w_027_1189, w_027_1190, w_027_1191, w_027_1192, w_027_1193, w_027_1194, w_027_1195, w_027_1196, w_027_1197, w_027_1198, w_027_1199, w_027_1200, w_027_1201, w_027_1202, w_027_1203, w_027_1204, w_027_1205, w_027_1206, w_027_1207, w_027_1208, w_027_1209, w_027_1210, w_027_1211, w_027_1212, w_027_1213, w_027_1214, w_027_1215, w_027_1216, w_027_1217, w_027_1218, w_027_1219, w_027_1220, w_027_1221, w_027_1222, w_027_1223, w_027_1224, w_027_1225, w_027_1226, w_027_1227, w_027_1228, w_027_1229, w_027_1230, w_027_1231, w_027_1232, w_027_1233, w_027_1234, w_027_1235, w_027_1236, w_027_1237, w_027_1238, w_027_1239, w_027_1240, w_027_1241, w_027_1242, w_027_1243, w_027_1244, w_027_1245, w_027_1246, w_027_1247, w_027_1248, w_027_1249, w_027_1250, w_027_1251, w_027_1252, w_027_1254, w_027_1255, w_027_1256, w_027_1257, w_027_1258, w_027_1259, w_027_1260, w_027_1261, w_027_1263, w_027_1264, w_027_1265, w_027_1266, w_027_1267, w_027_1268, w_027_1269, w_027_1270, w_027_1271, w_027_1272, w_027_1273, w_027_1274, w_027_1275, w_027_1276, w_027_1277, w_027_1278, w_027_1279, w_027_1280, w_027_1281, w_027_1282, w_027_1283, w_027_1284, w_027_1285, w_027_1286, w_027_1287, w_027_1288, w_027_1289, w_027_1290, w_027_1291, w_027_1292, w_027_1293, w_027_1294, w_027_1295, w_027_1296, w_027_1297, w_027_1298, w_027_1299, w_027_1300, w_027_1301, w_027_1302, w_027_1304, w_027_1305, w_027_1306, w_027_1307, w_027_1308, w_027_1309, w_027_1310, w_027_1311, w_027_1312, w_027_1313, w_027_1314, w_027_1315, w_027_1316, w_027_1317, w_027_1318, w_027_1319, w_027_1320, w_027_1321, w_027_1322, w_027_1323, w_027_1324, w_027_1325, w_027_1326, w_027_1327, w_027_1328, w_027_1329, w_027_1330, w_027_1331, w_027_1332, w_027_1333, w_027_1334, w_027_1335, w_027_1337, w_027_1340, w_027_1341, w_027_1342, w_027_1343, w_027_1344, w_027_1345, w_027_1346, w_027_1347, w_027_1348, w_027_1349, w_027_1350, w_027_1351, w_027_1352, w_027_1353, w_027_1354, w_027_1355, w_027_1356, w_027_1357, w_027_1358, w_027_1359, w_027_1360, w_027_1361, w_027_1362, w_027_1363, w_027_1364, w_027_1366, w_027_1367, w_027_1368, w_027_1369, w_027_1370, w_027_1371, w_027_1372, w_027_1373, w_027_1374, w_027_1375, w_027_1376, w_027_1377, w_027_1378, w_027_1379, w_027_1380, w_027_1381, w_027_1382, w_027_1383, w_027_1384, w_027_1385, w_027_1386, w_027_1387, w_027_1388, w_027_1389, w_027_1390, w_027_1391, w_027_1392, w_027_1393, w_027_1394, w_027_1395, w_027_1396, w_027_1397, w_027_1398, w_027_1399, w_027_1400, w_027_1401, w_027_1402, w_027_1403, w_027_1404, w_027_1405, w_027_1406, w_027_1407, w_027_1408, w_027_1409, w_027_1410, w_027_1411, w_027_1412, w_027_1413, w_027_1414, w_027_1415, w_027_1416, w_027_1418, w_027_1419, w_027_1420, w_027_1421, w_027_1422, w_027_1424, w_027_1425, w_027_1426, w_027_1427, w_027_1428, w_027_1429, w_027_1430, w_027_1431, w_027_1432, w_027_1433, w_027_1434, w_027_1435, w_027_1436, w_027_1437, w_027_1438, w_027_1439, w_027_1440, w_027_1441, w_027_1442, w_027_1444, w_027_1446, w_027_1447, w_027_1448, w_027_1449, w_027_1450, w_027_1451, w_027_1452, w_027_1453, w_027_1454, w_027_1455, w_027_1456, w_027_1457, w_027_1458, w_027_1459, w_027_1460, w_027_1461, w_027_1462, w_027_1463, w_027_1464, w_027_1465, w_027_1466, w_027_1467, w_027_1468, w_027_1469, w_027_1470, w_027_1471, w_027_1472, w_027_1473, w_027_1474, w_027_1475, w_027_1476, w_027_1477, w_027_1479, w_027_1481, w_027_1482, w_027_1483, w_027_1484, w_027_1485, w_027_1486, w_027_1487, w_027_1488, w_027_1489, w_027_1490, w_027_1491, w_027_1492, w_027_1493, w_027_1494, w_027_1495, w_027_1496, w_027_1497, w_027_1498, w_027_1499, w_027_1500, w_027_1501, w_027_1502, w_027_1505, w_027_1506, w_027_1507, w_027_1508, w_027_1509, w_027_1510, w_027_1511, w_027_1512, w_027_1513, w_027_1514, w_027_1515, w_027_1516, w_027_1517, w_027_1518, w_027_1519, w_027_1520, w_027_1521, w_027_1522, w_027_1523, w_027_1524, w_027_1525, w_027_1526, w_027_1527, w_027_1528, w_027_1529, w_027_1530, w_027_1531, w_027_1532, w_027_1533, w_027_1534, w_027_1535, w_027_1536, w_027_1537, w_027_1538, w_027_1539, w_027_1540, w_027_1541, w_027_1542, w_027_1543, w_027_1544, w_027_1545, w_027_1546, w_027_1547, w_027_1548, w_027_1549, w_027_1550, w_027_1551, w_027_1552, w_027_1553, w_027_1554, w_027_1555, w_027_1556, w_027_1557, w_027_1558, w_027_1559, w_027_1560, w_027_1561, w_027_1562, w_027_1563, w_027_1564, w_027_1565, w_027_1566, w_027_1567, w_027_1568, w_027_1569, w_027_1570, w_027_1571, w_027_1572, w_027_1573, w_027_1574, w_027_1575, w_027_1576, w_027_1577, w_027_1579, w_027_1580, w_027_1581, w_027_1582, w_027_1583, w_027_1584, w_027_1585, w_027_1586, w_027_1587, w_027_1588, w_027_1589, w_027_1590, w_027_1591, w_027_1592, w_027_1593, w_027_1594, w_027_1595, w_027_1596, w_027_1597, w_027_1598, w_027_1599, w_027_1600, w_027_1601, w_027_1602, w_027_1603, w_027_1604, w_027_1605, w_027_1606, w_027_1607, w_027_1608, w_027_1609, w_027_1610, w_027_1611, w_027_1612, w_027_1613, w_027_1614, w_027_1615, w_027_1616, w_027_1617, w_027_1618, w_027_1619, w_027_1620, w_027_1621, w_027_1622, w_027_1623, w_027_1624, w_027_1625, w_027_1626, w_027_1627, w_027_1628, w_027_1629, w_027_1630, w_027_1631, w_027_1632, w_027_1633, w_027_1634, w_027_1635, w_027_1636, w_027_1637, w_027_1638, w_027_1640, w_027_1641, w_027_1642, w_027_1643, w_027_1644, w_027_1645, w_027_1646, w_027_1647, w_027_1649, w_027_1651, w_027_1652, w_027_1653, w_027_1654, w_027_1655, w_027_1656, w_027_1657, w_027_1658, w_027_1659, w_027_1660, w_027_1661, w_027_1663;
  wire w_028_000, w_028_001, w_028_002, w_028_003, w_028_005, w_028_010, w_028_011, w_028_012, w_028_013, w_028_014, w_028_015, w_028_016, w_028_017, w_028_018, w_028_019, w_028_020, w_028_021, w_028_022, w_028_024, w_028_025, w_028_027, w_028_028, w_028_029, w_028_030, w_028_031, w_028_033, w_028_035, w_028_036, w_028_038, w_028_039, w_028_040, w_028_041, w_028_042, w_028_043, w_028_045, w_028_046, w_028_047, w_028_048, w_028_049, w_028_050, w_028_051, w_028_053, w_028_054, w_028_055, w_028_056, w_028_057, w_028_058, w_028_059, w_028_060, w_028_062, w_028_063, w_028_064, w_028_065, w_028_067, w_028_068, w_028_069, w_028_070, w_028_072, w_028_073, w_028_074, w_028_076, w_028_077, w_028_078, w_028_079, w_028_080, w_028_081, w_028_082, w_028_083, w_028_084, w_028_086, w_028_087, w_028_088, w_028_089, w_028_090, w_028_091, w_028_092, w_028_093, w_028_094, w_028_095, w_028_096, w_028_098, w_028_100, w_028_101, w_028_102, w_028_103, w_028_105, w_028_106, w_028_107, w_028_108, w_028_109, w_028_110, w_028_111, w_028_113, w_028_114, w_028_115, w_028_116, w_028_117, w_028_118, w_028_119, w_028_120, w_028_121, w_028_123, w_028_124, w_028_125, w_028_126, w_028_128, w_028_130, w_028_131, w_028_132, w_028_133, w_028_134, w_028_135, w_028_136, w_028_137, w_028_138, w_028_139, w_028_140, w_028_141, w_028_142, w_028_143, w_028_144, w_028_146, w_028_148, w_028_149, w_028_150, w_028_151, w_028_152, w_028_153, w_028_154, w_028_155, w_028_156, w_028_157, w_028_158, w_028_159, w_028_160, w_028_161, w_028_162, w_028_163, w_028_164, w_028_165, w_028_166, w_028_167, w_028_168, w_028_169, w_028_170, w_028_171, w_028_172, w_028_173, w_028_174, w_028_175, w_028_176, w_028_177, w_028_178, w_028_179, w_028_180, w_028_181, w_028_182, w_028_183, w_028_184, w_028_185, w_028_186, w_028_187, w_028_188, w_028_189, w_028_190, w_028_191, w_028_192, w_028_193, w_028_194, w_028_195, w_028_196, w_028_197, w_028_198, w_028_200, w_028_201, w_028_202, w_028_203, w_028_204, w_028_205, w_028_206, w_028_207, w_028_209, w_028_210, w_028_212, w_028_213, w_028_214, w_028_215, w_028_216, w_028_218, w_028_219, w_028_220, w_028_221, w_028_222, w_028_223, w_028_224, w_028_225, w_028_226, w_028_227, w_028_228, w_028_229, w_028_230, w_028_231, w_028_232, w_028_233, w_028_234, w_028_235, w_028_236, w_028_237, w_028_238, w_028_239, w_028_240, w_028_242, w_028_243, w_028_244, w_028_245, w_028_246, w_028_247, w_028_250, w_028_251, w_028_252, w_028_253, w_028_254, w_028_256, w_028_257, w_028_258, w_028_259, w_028_260, w_028_261, w_028_262, w_028_263, w_028_264, w_028_265, w_028_266, w_028_267, w_028_268, w_028_269, w_028_270, w_028_271, w_028_272, w_028_273, w_028_274, w_028_275, w_028_276, w_028_279, w_028_280, w_028_282, w_028_283, w_028_284, w_028_285, w_028_287, w_028_288, w_028_289, w_028_290, w_028_291, w_028_292, w_028_293, w_028_294, w_028_295, w_028_296, w_028_297, w_028_298, w_028_299, w_028_300, w_028_302, w_028_303, w_028_304, w_028_305, w_028_306, w_028_307, w_028_308, w_028_309, w_028_310, w_028_312, w_028_313, w_028_314, w_028_315, w_028_316, w_028_317, w_028_318, w_028_319, w_028_320, w_028_321, w_028_322, w_028_323, w_028_324, w_028_325, w_028_326, w_028_327, w_028_328, w_028_329, w_028_331, w_028_333, w_028_334, w_028_335, w_028_337, w_028_338, w_028_340, w_028_341, w_028_342, w_028_344, w_028_345, w_028_346, w_028_347, w_028_348, w_028_349, w_028_350, w_028_351, w_028_352, w_028_353, w_028_354, w_028_355, w_028_356, w_028_358, w_028_359, w_028_360, w_028_361, w_028_362, w_028_364, w_028_365, w_028_366, w_028_367, w_028_368, w_028_369, w_028_370, w_028_371, w_028_372, w_028_374, w_028_375, w_028_376, w_028_377, w_028_378, w_028_379, w_028_381, w_028_382, w_028_383, w_028_384, w_028_385, w_028_386, w_028_387, w_028_388, w_028_389, w_028_390, w_028_391, w_028_392, w_028_393, w_028_394, w_028_396, w_028_398, w_028_399, w_028_400, w_028_401, w_028_402, w_028_403, w_028_404, w_028_405, w_028_406, w_028_408, w_028_409, w_028_410, w_028_411, w_028_412, w_028_413, w_028_414, w_028_415, w_028_417, w_028_418, w_028_420, w_028_421, w_028_422, w_028_423, w_028_424, w_028_425, w_028_426, w_028_427, w_028_428, w_028_429, w_028_430, w_028_431, w_028_432, w_028_433, w_028_434, w_028_436, w_028_438, w_028_439, w_028_440, w_028_441, w_028_442, w_028_443, w_028_444, w_028_445, w_028_448, w_028_449, w_028_451, w_028_453, w_028_454, w_028_455, w_028_456, w_028_457, w_028_458, w_028_459, w_028_460, w_028_461, w_028_462, w_028_463, w_028_464, w_028_465, w_028_466, w_028_467, w_028_468, w_028_469, w_028_470, w_028_471, w_028_472, w_028_473, w_028_474, w_028_475, w_028_476, w_028_477, w_028_479, w_028_480, w_028_481, w_028_482, w_028_483, w_028_484, w_028_485, w_028_486, w_028_487, w_028_488, w_028_489, w_028_490, w_028_491, w_028_492, w_028_493, w_028_494, w_028_495, w_028_496, w_028_497, w_028_498, w_028_499, w_028_500, w_028_501, w_028_502, w_028_503, w_028_504, w_028_505, w_028_506, w_028_507, w_028_508, w_028_509, w_028_510, w_028_511, w_028_513, w_028_514, w_028_515, w_028_516, w_028_517, w_028_518, w_028_519, w_028_520, w_028_521, w_028_522, w_028_524, w_028_525, w_028_527, w_028_528, w_028_529, w_028_530, w_028_531, w_028_532, w_028_533, w_028_534, w_028_535, w_028_536, w_028_538, w_028_539, w_028_540, w_028_541, w_028_542, w_028_544, w_028_545, w_028_546, w_028_547, w_028_548, w_028_549, w_028_550, w_028_551, w_028_554, w_028_555, w_028_556, w_028_557, w_028_558, w_028_559, w_028_560, w_028_561, w_028_562, w_028_563, w_028_565, w_028_567, w_028_568, w_028_569, w_028_570, w_028_571, w_028_572, w_028_573, w_028_574, w_028_576, w_028_577, w_028_578, w_028_579, w_028_580, w_028_581, w_028_582, w_028_583, w_028_585, w_028_586, w_028_587, w_028_588, w_028_589, w_028_590, w_028_591, w_028_593, w_028_594, w_028_595, w_028_596, w_028_597, w_028_598, w_028_599, w_028_600, w_028_601, w_028_602, w_028_603, w_028_604, w_028_605, w_028_606, w_028_607, w_028_608, w_028_609, w_028_610, w_028_611, w_028_612, w_028_613, w_028_614, w_028_615, w_028_616, w_028_617, w_028_618, w_028_619, w_028_620, w_028_621, w_028_622, w_028_623, w_028_624, w_028_625, w_028_626, w_028_627, w_028_629, w_028_630, w_028_632, w_028_634, w_028_635, w_028_637, w_028_638, w_028_639, w_028_641, w_028_642, w_028_643, w_028_645, w_028_646, w_028_648, w_028_649, w_028_650, w_028_651, w_028_652, w_028_653, w_028_655, w_028_656, w_028_657, w_028_658, w_028_659, w_028_660, w_028_661, w_028_662, w_028_663, w_028_664, w_028_665, w_028_666, w_028_667, w_028_668, w_028_670, w_028_672, w_028_673, w_028_674, w_028_675, w_028_676, w_028_677, w_028_678, w_028_679, w_028_680, w_028_681, w_028_682, w_028_683, w_028_684, w_028_685, w_028_687, w_028_688, w_028_691, w_028_692, w_028_694, w_028_695, w_028_697, w_028_698, w_028_699, w_028_700, w_028_701, w_028_702, w_028_705, w_028_706, w_028_707, w_028_708, w_028_709, w_028_710, w_028_711, w_028_712, w_028_713, w_028_714, w_028_715, w_028_716, w_028_717, w_028_718, w_028_719, w_028_720, w_028_721, w_028_723, w_028_724, w_028_725, w_028_726, w_028_727, w_028_728, w_028_731, w_028_732, w_028_733, w_028_734, w_028_735, w_028_737, w_028_738, w_028_740, w_028_741, w_028_742, w_028_743, w_028_744, w_028_745, w_028_746, w_028_748, w_028_749, w_028_750, w_028_751, w_028_752, w_028_754, w_028_755, w_028_756, w_028_757, w_028_758, w_028_759, w_028_760, w_028_761, w_028_762, w_028_763, w_028_765, w_028_766, w_028_767, w_028_768, w_028_769, w_028_770, w_028_771, w_028_773, w_028_775, w_028_776, w_028_777, w_028_779, w_028_780, w_028_781, w_028_783, w_028_784, w_028_785, w_028_786, w_028_787, w_028_788, w_028_789, w_028_790, w_028_791, w_028_793, w_028_794, w_028_795, w_028_796, w_028_798, w_028_799, w_028_800, w_028_801, w_028_802, w_028_803, w_028_804, w_028_805, w_028_806, w_028_807, w_028_808, w_028_810, w_028_811, w_028_812, w_028_813, w_028_815, w_028_816, w_028_817, w_028_818, w_028_819, w_028_820, w_028_821, w_028_822, w_028_823, w_028_824, w_028_825, w_028_826, w_028_827, w_028_828, w_028_830, w_028_831, w_028_832, w_028_833, w_028_834, w_028_835, w_028_836, w_028_838, w_028_839, w_028_840, w_028_841, w_028_842, w_028_843, w_028_844, w_028_845, w_028_849, w_028_850, w_028_852, w_028_853, w_028_854, w_028_855, w_028_856, w_028_857, w_028_858, w_028_859, w_028_860, w_028_861, w_028_862, w_028_863, w_028_864, w_028_865, w_028_866, w_028_867, w_028_868, w_028_869, w_028_870, w_028_871, w_028_872, w_028_873, w_028_874, w_028_875, w_028_876, w_028_877, w_028_878, w_028_879, w_028_880, w_028_881, w_028_882, w_028_883, w_028_884, w_028_885, w_028_886, w_028_888, w_028_889, w_028_890, w_028_891, w_028_892, w_028_893, w_028_894, w_028_896, w_028_897, w_028_899, w_028_900, w_028_901, w_028_902, w_028_903, w_028_904, w_028_905, w_028_906, w_028_907, w_028_908, w_028_909, w_028_910, w_028_911, w_028_913, w_028_914, w_028_915, w_028_918, w_028_919, w_028_920, w_028_921, w_028_922, w_028_923, w_028_924, w_028_925, w_028_927, w_028_929, w_028_931, w_028_932, w_028_933, w_028_934, w_028_935, w_028_936, w_028_937, w_028_938, w_028_939, w_028_940, w_028_941, w_028_942, w_028_943, w_028_944, w_028_945, w_028_946, w_028_947, w_028_948, w_028_949, w_028_950, w_028_951, w_028_953, w_028_954, w_028_955, w_028_957, w_028_958, w_028_959, w_028_960, w_028_961, w_028_962, w_028_964, w_028_965, w_028_966, w_028_967, w_028_968, w_028_969, w_028_970, w_028_971, w_028_973, w_028_974, w_028_975, w_028_976, w_028_977, w_028_978, w_028_979, w_028_980, w_028_981, w_028_982, w_028_983, w_028_984, w_028_986, w_028_987, w_028_988, w_028_989, w_028_990, w_028_991, w_028_992, w_028_993, w_028_994, w_028_995, w_028_996, w_028_997, w_028_998, w_028_999, w_028_1000, w_028_1001, w_028_1002, w_028_1003, w_028_1004, w_028_1005, w_028_1006, w_028_1007, w_028_1008, w_028_1009, w_028_1010, w_028_1011, w_028_1012, w_028_1013, w_028_1014, w_028_1015, w_028_1016, w_028_1018, w_028_1019, w_028_1020, w_028_1021, w_028_1022, w_028_1024, w_028_1025, w_028_1026, w_028_1027, w_028_1028, w_028_1029, w_028_1030, w_028_1031, w_028_1033, w_028_1034, w_028_1035, w_028_1036, w_028_1037, w_028_1038, w_028_1040, w_028_1041, w_028_1043, w_028_1044, w_028_1046, w_028_1047, w_028_1048, w_028_1049, w_028_1051, w_028_1052, w_028_1053, w_028_1054, w_028_1056, w_028_1057, w_028_1058, w_028_1060, w_028_1062, w_028_1063, w_028_1064, w_028_1065, w_028_1066, w_028_1067, w_028_1068, w_028_1069, w_028_1070, w_028_1071, w_028_1072, w_028_1073, w_028_1074, w_028_1075, w_028_1076, w_028_1077, w_028_1078, w_028_1080, w_028_1081, w_028_1082, w_028_1083, w_028_1084, w_028_1085, w_028_1086, w_028_1087, w_028_1088, w_028_1089, w_028_1091, w_028_1092, w_028_1093, w_028_1094, w_028_1095, w_028_1096, w_028_1097, w_028_1099, w_028_1100, w_028_1101, w_028_1102, w_028_1103, w_028_1104, w_028_1105, w_028_1106, w_028_1107, w_028_1108, w_028_1109, w_028_1110, w_028_1111, w_028_1113, w_028_1114, w_028_1115, w_028_1116, w_028_1117, w_028_1118, w_028_1119, w_028_1120, w_028_1121, w_028_1122, w_028_1124, w_028_1125, w_028_1126, w_028_1127, w_028_1128, w_028_1130, w_028_1131, w_028_1132, w_028_1133, w_028_1134, w_028_1135, w_028_1137, w_028_1138, w_028_1139, w_028_1140, w_028_1141, w_028_1142, w_028_1143, w_028_1144, w_028_1145, w_028_1146, w_028_1147, w_028_1148, w_028_1149, w_028_1150, w_028_1151, w_028_1152, w_028_1153, w_028_1154, w_028_1156, w_028_1157, w_028_1158, w_028_1159, w_028_1160, w_028_1161, w_028_1162, w_028_1163, w_028_1164, w_028_1165, w_028_1166, w_028_1167, w_028_1169, w_028_1170, w_028_1171, w_028_1172, w_028_1173, w_028_1174, w_028_1176, w_028_1177, w_028_1180, w_028_1181, w_028_1182, w_028_1183, w_028_1184, w_028_1185, w_028_1186, w_028_1187, w_028_1189, w_028_1191, w_028_1192, w_028_1193, w_028_1194, w_028_1195, w_028_1196, w_028_1197, w_028_1198, w_028_1200, w_028_1201, w_028_1202, w_028_1203, w_028_1204, w_028_1205, w_028_1206, w_028_1207, w_028_1208, w_028_1213, w_028_1214, w_028_1216, w_028_1217, w_028_1218, w_028_1219, w_028_1220, w_028_1221, w_028_1222, w_028_1223, w_028_1224, w_028_1225, w_028_1226, w_028_1228, w_028_1229, w_028_1230, w_028_1231, w_028_1232, w_028_1234, w_028_1235, w_028_1236, w_028_1237, w_028_1238, w_028_1239, w_028_1240, w_028_1241, w_028_1242, w_028_1243, w_028_1244, w_028_1245, w_028_1246, w_028_1247, w_028_1248, w_028_1249, w_028_1250, w_028_1251, w_028_1252, w_028_1253, w_028_1254, w_028_1255, w_028_1259, w_028_1260, w_028_1261, w_028_1262, w_028_1264, w_028_1265, w_028_1266, w_028_1267, w_028_1268, w_028_1269, w_028_1270, w_028_1271, w_028_1272, w_028_1274, w_028_1275, w_028_1276, w_028_1277, w_028_1278, w_028_1279, w_028_1280, w_028_1281, w_028_1282, w_028_1283, w_028_1285, w_028_1286, w_028_1287, w_028_1288, w_028_1290, w_028_1291, w_028_1292, w_028_1293, w_028_1295, w_028_1296, w_028_1297, w_028_1298, w_028_1299, w_028_1300, w_028_1301, w_028_1302, w_028_1303, w_028_1304, w_028_1305, w_028_1306, w_028_1307, w_028_1309, w_028_1311, w_028_1313, w_028_1314, w_028_1315, w_028_1316, w_028_1317, w_028_1318, w_028_1319, w_028_1320, w_028_1321, w_028_1323, w_028_1324, w_028_1325, w_028_1327, w_028_1328, w_028_1329, w_028_1330, w_028_1331, w_028_1332, w_028_1333, w_028_1334, w_028_1335, w_028_1336, w_028_1337, w_028_1338, w_028_1339, w_028_1340, w_028_1341, w_028_1342, w_028_1343, w_028_1344, w_028_1345, w_028_1347, w_028_1348, w_028_1349, w_028_1350, w_028_1351, w_028_1352, w_028_1353, w_028_1354, w_028_1355, w_028_1356, w_028_1357, w_028_1360, w_028_1361, w_028_1362, w_028_1364, w_028_1365, w_028_1366, w_028_1368, w_028_1369, w_028_1370, w_028_1371, w_028_1372, w_028_1373, w_028_1374, w_028_1376, w_028_1377, w_028_1378, w_028_1379, w_028_1381, w_028_1382, w_028_1383, w_028_1385, w_028_1386, w_028_1387, w_028_1388, w_028_1390, w_028_1391, w_028_1392, w_028_1393, w_028_1395, w_028_1396, w_028_1397, w_028_1398, w_028_1399, w_028_1400, w_028_1401, w_028_1402, w_028_1403, w_028_1404, w_028_1405, w_028_1406, w_028_1407, w_028_1410, w_028_1411, w_028_1412, w_028_1414, w_028_1415, w_028_1416, w_028_1418, w_028_1420, w_028_1421, w_028_1422, w_028_1425, w_028_1427, w_028_1429, w_028_1430, w_028_1431, w_028_1436, w_028_1439, w_028_1440, w_028_1441, w_028_1442, w_028_1445, w_028_1446, w_028_1448, w_028_1450, w_028_1451, w_028_1452, w_028_1453, w_028_1456, w_028_1457, w_028_1458, w_028_1460, w_028_1461, w_028_1462, w_028_1464, w_028_1465, w_028_1466, w_028_1468, w_028_1469, w_028_1470, w_028_1472, w_028_1473, w_028_1474, w_028_1475, w_028_1476, w_028_1477, w_028_1478, w_028_1481, w_028_1482, w_028_1485, w_028_1486, w_028_1487, w_028_1488, w_028_1489, w_028_1490, w_028_1491, w_028_1492, w_028_1493, w_028_1495, w_028_1496, w_028_1498, w_028_1499, w_028_1500, w_028_1502, w_028_1503, w_028_1504, w_028_1505, w_028_1506, w_028_1507, w_028_1509, w_028_1510, w_028_1512, w_028_1519, w_028_1520, w_028_1522, w_028_1523, w_028_1524, w_028_1526, w_028_1528, w_028_1531, w_028_1533, w_028_1538, w_028_1539, w_028_1540, w_028_1542, w_028_1544, w_028_1545, w_028_1546, w_028_1551, w_028_1552, w_028_1553, w_028_1554, w_028_1555, w_028_1556, w_028_1557, w_028_1558, w_028_1559, w_028_1560, w_028_1563, w_028_1564, w_028_1565, w_028_1566, w_028_1567, w_028_1568, w_028_1569, w_028_1572, w_028_1573, w_028_1574, w_028_1576, w_028_1579, w_028_1583, w_028_1584, w_028_1586, w_028_1587, w_028_1588, w_028_1589, w_028_1590, w_028_1592, w_028_1593, w_028_1595, w_028_1596, w_028_1597, w_028_1599, w_028_1602, w_028_1603, w_028_1605, w_028_1606, w_028_1608, w_028_1609, w_028_1610, w_028_1611, w_028_1612, w_028_1613, w_028_1615, w_028_1616, w_028_1619, w_028_1620, w_028_1623, w_028_1626, w_028_1627, w_028_1628, w_028_1631, w_028_1632, w_028_1635, w_028_1636, w_028_1637, w_028_1638, w_028_1639, w_028_1640, w_028_1642, w_028_1644, w_028_1645, w_028_1647, w_028_1648, w_028_1649, w_028_1650, w_028_1651, w_028_1652, w_028_1653, w_028_1655, w_028_1657, w_028_1658, w_028_1659, w_028_1661, w_028_1665, w_028_1666, w_028_1667, w_028_1668, w_028_1670, w_028_1671, w_028_1672, w_028_1673, w_028_1675, w_028_1679, w_028_1680, w_028_1682, w_028_1683, w_028_1684, w_028_1685, w_028_1688, w_028_1689, w_028_1691, w_028_1692, w_028_1693, w_028_1694, w_028_1695, w_028_1697, w_028_1698, w_028_1699, w_028_1701, w_028_1702, w_028_1703, w_028_1705, w_028_1706, w_028_1709, w_028_1715, w_028_1716, w_028_1717, w_028_1718, w_028_1719, w_028_1720, w_028_1721, w_028_1724, w_028_1725, w_028_1726, w_028_1728, w_028_1729, w_028_1730, w_028_1732, w_028_1733, w_028_1734, w_028_1735, w_028_1736, w_028_1738, w_028_1739, w_028_1740, w_028_1741, w_028_1742, w_028_1743, w_028_1744, w_028_1745, w_028_1746, w_028_1747, w_028_1748, w_028_1750, w_028_1752, w_028_1753, w_028_1754, w_028_1755, w_028_1756, w_028_1757, w_028_1759, w_028_1762, w_028_1764, w_028_1765, w_028_1766, w_028_1767, w_028_1768, w_028_1770, w_028_1773, w_028_1774, w_028_1776, w_028_1777, w_028_1778, w_028_1779, w_028_1780, w_028_1781, w_028_1784, w_028_1785, w_028_1788, w_028_1791, w_028_1794, w_028_1795, w_028_1796, w_028_1798, w_028_1799, w_028_1801, w_028_1802, w_028_1803, w_028_1804, w_028_1805, w_028_1806, w_028_1807, w_028_1808, w_028_1809, w_028_1811, w_028_1812, w_028_1813, w_028_1814, w_028_1816, w_028_1817, w_028_1818, w_028_1819, w_028_1821, w_028_1823, w_028_1825, w_028_1828, w_028_1829, w_028_1831, w_028_1832, w_028_1833, w_028_1835, w_028_1836, w_028_1837, w_028_1838, w_028_1840, w_028_1842, w_028_1843, w_028_1844, w_028_1845, w_028_1846, w_028_1847, w_028_1850, w_028_1851, w_028_1852, w_028_1853, w_028_1854, w_028_1855, w_028_1859, w_028_1861, w_028_1862, w_028_1863, w_028_1865, w_028_1868, w_028_1870, w_028_1872, w_028_1873, w_028_1874, w_028_1875, w_028_1876, w_028_1877, w_028_1880, w_028_1882, w_028_1883, w_028_1885, w_028_1886, w_028_1888, w_028_1889, w_028_1890, w_028_1894, w_028_1895, w_028_1896, w_028_1898, w_028_1899, w_028_1900, w_028_1901, w_028_1903, w_028_1904, w_028_1905, w_028_1906, w_028_1908, w_028_1909, w_028_1911, w_028_1912, w_028_1913, w_028_1914, w_028_1916, w_028_1917, w_028_1918, w_028_1919, w_028_1923, w_028_1925, w_028_1926, w_028_1927, w_028_1929, w_028_1931, w_028_1932, w_028_1933, w_028_1934, w_028_1935, w_028_1937, w_028_1941, w_028_1942, w_028_1943, w_028_1944, w_028_1946, w_028_1947, w_028_1948, w_028_1950, w_028_1951, w_028_1952, w_028_1953, w_028_1954, w_028_1955, w_028_1956, w_028_1957, w_028_1959, w_028_1961, w_028_1963, w_028_1964, w_028_1965, w_028_1969, w_028_1971, w_028_1972, w_028_1973, w_028_1974, w_028_1975, w_028_1977, w_028_1978, w_028_1979, w_028_1980, w_028_1985, w_028_1987, w_028_1988, w_028_1989, w_028_1990, w_028_1991, w_028_1992, w_028_1993, w_028_1994, w_028_1996, w_028_1997, w_028_1998, w_028_1999, w_028_2000, w_028_2002, w_028_2003, w_028_2004, w_028_2005, w_028_2006, w_028_2008, w_028_2011, w_028_2014, w_028_2016, w_028_2017, w_028_2018, w_028_2019, w_028_2022, w_028_2023, w_028_2024, w_028_2025, w_028_2026, w_028_2027, w_028_2028, w_028_2030, w_028_2031, w_028_2032, w_028_2033, w_028_2034, w_028_2038, w_028_2040, w_028_2041, w_028_2042, w_028_2043, w_028_2044, w_028_2045, w_028_2047, w_028_2049, w_028_2051, w_028_2053, w_028_2054, w_028_2055, w_028_2058, w_028_2059, w_028_2060, w_028_2061, w_028_2064, w_028_2066, w_028_2067, w_028_2068, w_028_2069, w_028_2070, w_028_2071, w_028_2073, w_028_2075, w_028_2076, w_028_2078, w_028_2080, w_028_2081, w_028_2082, w_028_2088, w_028_2089, w_028_2091, w_028_2093, w_028_2094, w_028_2097, w_028_2101, w_028_2102, w_028_2104, w_028_2106, w_028_2107, w_028_2108, w_028_2110, w_028_2111, w_028_2112, w_028_2114, w_028_2115, w_028_2116, w_028_2117, w_028_2118, w_028_2119, w_028_2121, w_028_2122, w_028_2123, w_028_2124, w_028_2127, w_028_2129, w_028_2130, w_028_2131, w_028_2133, w_028_2135, w_028_2136, w_028_2137, w_028_2138, w_028_2139, w_028_2141, w_028_2142, w_028_2144, w_028_2146, w_028_2147, w_028_2148, w_028_2150, w_028_2151, w_028_2152, w_028_2153, w_028_2154, w_028_2155, w_028_2156, w_028_2158, w_028_2160, w_028_2161, w_028_2162, w_028_2164, w_028_2165, w_028_2167, w_028_2168, w_028_2170, w_028_2171, w_028_2172, w_028_2174, w_028_2177, w_028_2180, w_028_2182, w_028_2184, w_028_2185, w_028_2186, w_028_2187, w_028_2190, w_028_2192, w_028_2195, w_028_2197, w_028_2200, w_028_2201, w_028_2203, w_028_2204, w_028_2206, w_028_2208, w_028_2209, w_028_2210, w_028_2211, w_028_2215, w_028_2217, w_028_2219, w_028_2220, w_028_2221, w_028_2222, w_028_2223, w_028_2224, w_028_2225, w_028_2226, w_028_2230, w_028_2231, w_028_2232, w_028_2234, w_028_2237, w_028_2239, w_028_2243, w_028_2244, w_028_2245, w_028_2246, w_028_2247, w_028_2249, w_028_2252, w_028_2254, w_028_2256, w_028_2257, w_028_2259, w_028_2261, w_028_2262, w_028_2263, w_028_2264, w_028_2266, w_028_2268, w_028_2269, w_028_2270, w_028_2272, w_028_2274, w_028_2275, w_028_2276, w_028_2282, w_028_2283, w_028_2284, w_028_2285, w_028_2286, w_028_2287, w_028_2288, w_028_2291, w_028_2293, w_028_2295, w_028_2298, w_028_2299, w_028_2300, w_028_2301, w_028_2303, w_028_2304, w_028_2305, w_028_2307, w_028_2309, w_028_2310, w_028_2311, w_028_2314, w_028_2315, w_028_2316, w_028_2318, w_028_2321, w_028_2323, w_028_2326, w_028_2327, w_028_2328, w_028_2329, w_028_2330, w_028_2331, w_028_2332, w_028_2333, w_028_2335, w_028_2337, w_028_2338, w_028_2339, w_028_2340, w_028_2342, w_028_2344, w_028_2345, w_028_2346, w_028_2349, w_028_2351, w_028_2353, w_028_2355, w_028_2356, w_028_2358, w_028_2359, w_028_2361, w_028_2362, w_028_2363, w_028_2365, w_028_2366, w_028_2368, w_028_2370, w_028_2372, w_028_2374, w_028_2375, w_028_2376, w_028_2377, w_028_2378, w_028_2379, w_028_2381, w_028_2382, w_028_2383, w_028_2384, w_028_2386, w_028_2389, w_028_2391, w_028_2394, w_028_2396, w_028_2399, w_028_2400, w_028_2401, w_028_2402, w_028_2405, w_028_2406, w_028_2407, w_028_2408, w_028_2410, w_028_2412, w_028_2413, w_028_2414, w_028_2415, w_028_2417, w_028_2418, w_028_2419, w_028_2421, w_028_2422, w_028_2424, w_028_2425, w_028_2426, w_028_2428, w_028_2429, w_028_2430, w_028_2431, w_028_2432, w_028_2434, w_028_2436, w_028_2437, w_028_2439, w_028_2441, w_028_2442, w_028_2443, w_028_2445, w_028_2446, w_028_2447, w_028_2448, w_028_2449, w_028_2451, w_028_2453, w_028_2454, w_028_2456, w_028_2457, w_028_2459, w_028_2460, w_028_2461, w_028_2463, w_028_2464, w_028_2465, w_028_2466, w_028_2468, w_028_2469, w_028_2470, w_028_2472, w_028_2474, w_028_2475, w_028_2480, w_028_2481, w_028_2482, w_028_2483, w_028_2484, w_028_2485, w_028_2487, w_028_2488, w_028_2489, w_028_2491, w_028_2492, w_028_2493, w_028_2494, w_028_2495, w_028_2497, w_028_2498, w_028_2500, w_028_2501, w_028_2502, w_028_2503, w_028_2504, w_028_2506, w_028_2507, w_028_2509, w_028_2510, w_028_2512, w_028_2513, w_028_2517, w_028_2519, w_028_2520, w_028_2521, w_028_2522, w_028_2523, w_028_2524, w_028_2525, w_028_2526, w_028_2528, w_028_2530, w_028_2531, w_028_2533, w_028_2534, w_028_2535, w_028_2536, w_028_2538, w_028_2539, w_028_2540, w_028_2541, w_028_2542, w_028_2544, w_028_2545, w_028_2546, w_028_2548, w_028_2549, w_028_2551, w_028_2552, w_028_2553, w_028_2554, w_028_2555, w_028_2556, w_028_2557, w_028_2559, w_028_2560, w_028_2562, w_028_2563, w_028_2565, w_028_2566, w_028_2568, w_028_2570, w_028_2571, w_028_2573, w_028_2574, w_028_2575, w_028_2576, w_028_2577, w_028_2578, w_028_2579, w_028_2580, w_028_2581, w_028_2582, w_028_2585, w_028_2586, w_028_2587, w_028_2589, w_028_2591, w_028_2593, w_028_2595, w_028_2596, w_028_2597, w_028_2598, w_028_2599, w_028_2600, w_028_2601, w_028_2602, w_028_2603, w_028_2604, w_028_2605, w_028_2608, w_028_2609, w_028_2612, w_028_2613, w_028_2614, w_028_2619, w_028_2620, w_028_2621, w_028_2622, w_028_2624, w_028_2625, w_028_2626, w_028_2627, w_028_2628, w_028_2629, w_028_2630, w_028_2631, w_028_2633, w_028_2634, w_028_2636, w_028_2638, w_028_2639, w_028_2640, w_028_2641, w_028_2644, w_028_2646, w_028_2647, w_028_2650, w_028_2651, w_028_2653, w_028_2654, w_028_2655, w_028_2656, w_028_2657, w_028_2659, w_028_2661, w_028_2663, w_028_2664, w_028_2665, w_028_2666, w_028_2667, w_028_2668, w_028_2669, w_028_2670, w_028_2672, w_028_2673, w_028_2674, w_028_2675, w_028_2677, w_028_2678, w_028_2680, w_028_2681, w_028_2683, w_028_2684, w_028_2685, w_028_2687, w_028_2688, w_028_2689, w_028_2691, w_028_2692, w_028_2693, w_028_2694, w_028_2697, w_028_2698, w_028_2699, w_028_2700, w_028_2701, w_028_2702, w_028_2705, w_028_2706, w_028_2708, w_028_2709, w_028_2711, w_028_2712, w_028_2713, w_028_2714, w_028_2716, w_028_2718, w_028_2719, w_028_2720, w_028_2722, w_028_2723, w_028_2724, w_028_2725, w_028_2728, w_028_2730, w_028_2731, w_028_2738, w_028_2740, w_028_2741, w_028_2742, w_028_2744, w_028_2746, w_028_2747, w_028_2749, w_028_2750, w_028_2752, w_028_2754, w_028_2756, w_028_2758, w_028_2759, w_028_2761, w_028_2763, w_028_2764, w_028_2765, w_028_2767, w_028_2769, w_028_2770, w_028_2771, w_028_2772, w_028_2773, w_028_2774, w_028_2777, w_028_2778, w_028_2781, w_028_2783, w_028_2784, w_028_2785, w_028_2786, w_028_2788, w_028_2789, w_028_2790, w_028_2791, w_028_2792, w_028_2793, w_028_2794, w_028_2797, w_028_2798, w_028_2799, w_028_2801, w_028_2802, w_028_2803, w_028_2804, w_028_2806, w_028_2809, w_028_2810, w_028_2813, w_028_2814, w_028_2815, w_028_2818, w_028_2819, w_028_2820, w_028_2823, w_028_2825, w_028_2826, w_028_2829, w_028_2830, w_028_2832, w_028_2833, w_028_2836, w_028_2837, w_028_2839, w_028_2840, w_028_2841, w_028_2842, w_028_2843, w_028_2846, w_028_2847, w_028_2848, w_028_2849, w_028_2850, w_028_2851, w_028_2852, w_028_2853, w_028_2854, w_028_2856, w_028_2859, w_028_2860, w_028_2862, w_028_2863, w_028_2867, w_028_2868, w_028_2869, w_028_2870, w_028_2871, w_028_2872, w_028_2873, w_028_2875, w_028_2876, w_028_2878, w_028_2879, w_028_2880, w_028_2881, w_028_2882, w_028_2883, w_028_2884, w_028_2885, w_028_2886, w_028_2887, w_028_2889, w_028_2891, w_028_2892, w_028_2893, w_028_2897, w_028_2899, w_028_2900, w_028_2901, w_028_2902, w_028_2904, w_028_2905, w_028_2907, w_028_2908, w_028_2909, w_028_2910, w_028_2911, w_028_2913, w_028_2915, w_028_2917, w_028_2918, w_028_2919, w_028_2921, w_028_2925, w_028_2926, w_028_2927, w_028_2928, w_028_2929, w_028_2930, w_028_2931, w_028_2932, w_028_2933, w_028_2935, w_028_2937, w_028_2939, w_028_2941, w_028_2942, w_028_2944, w_028_2945, w_028_2947, w_028_2948, w_028_2949, w_028_2950, w_028_2951, w_028_2954, w_028_2955, w_028_2956, w_028_2957, w_028_2958, w_028_2959, w_028_2960, w_028_2961, w_028_2962, w_028_2963, w_028_2964, w_028_2965, w_028_2966, w_028_2967, w_028_2968, w_028_2969, w_028_2970, w_028_2971, w_028_2972, w_028_2974, w_028_2976, w_028_2977, w_028_2980, w_028_2981, w_028_2982, w_028_2984, w_028_2985, w_028_2988, w_028_2989, w_028_2990, w_028_2992, w_028_2993, w_028_2995, w_028_2996, w_028_2997, w_028_2999, w_028_3002, w_028_3004, w_028_3005, w_028_3006, w_028_3007, w_028_3009, w_028_3011, w_028_3012, w_028_3017, w_028_3019, w_028_3020, w_028_3021, w_028_3023, w_028_3024, w_028_3026, w_028_3027, w_028_3028, w_028_3029, w_028_3030, w_028_3031, w_028_3032, w_028_3034, w_028_3035, w_028_3036, w_028_3038, w_028_3040, w_028_3041, w_028_3044, w_028_3045, w_028_3046, w_028_3047, w_028_3048, w_028_3049, w_028_3050, w_028_3051, w_028_3052, w_028_3054, w_028_3056, w_028_3057, w_028_3060, w_028_3061, w_028_3063, w_028_3064, w_028_3066, w_028_3067, w_028_3068, w_028_3069, w_028_3071, w_028_3072, w_028_3073, w_028_3074, w_028_3075, w_028_3076, w_028_3077, w_028_3078, w_028_3079, w_028_3080, w_028_3082, w_028_3083, w_028_3085, w_028_3086, w_028_3087, w_028_3089, w_028_3090, w_028_3093, w_028_3096, w_028_3097, w_028_3098, w_028_3099, w_028_3100, w_028_3102, w_028_3103, w_028_3105, w_028_3106, w_028_3107, w_028_3108, w_028_3109, w_028_3111, w_028_3112, w_028_3113, w_028_3114, w_028_3115, w_028_3116, w_028_3117, w_028_3118, w_028_3120, w_028_3121, w_028_3122, w_028_3123, w_028_3124, w_028_3126, w_028_3127, w_028_3128, w_028_3130, w_028_3133, w_028_3134, w_028_3135, w_028_3136, w_028_3137, w_028_3139, w_028_3141, w_028_3142, w_028_3143, w_028_3145, w_028_3146, w_028_3147, w_028_3148, w_028_3149, w_028_3151, w_028_3154, w_028_3156, w_028_3157, w_028_3158, w_028_3160, w_028_3161, w_028_3164, w_028_3167, w_028_3170, w_028_3175, w_028_3176, w_028_3177, w_028_3179, w_028_3180, w_028_3181, w_028_3182, w_028_3183, w_028_3185, w_028_3189, w_028_3193, w_028_3194, w_028_3195, w_028_3196, w_028_3197, w_028_3202, w_028_3203, w_028_3204, w_028_3206, w_028_3207, w_028_3208, w_028_3209, w_028_3212, w_028_3215, w_028_3216, w_028_3217, w_028_3218, w_028_3220, w_028_3221, w_028_3224, w_028_3225, w_028_3226, w_028_3228, w_028_3230, w_028_3231, w_028_3233, w_028_3236, w_028_3237, w_028_3239, w_028_3240, w_028_3242, w_028_3243, w_028_3245, w_028_3247, w_028_3248, w_028_3249, w_028_3251, w_028_3252, w_028_3253, w_028_3254, w_028_3255, w_028_3256, w_028_3258, w_028_3259, w_028_3262, w_028_3265, w_028_3266, w_028_3267, w_028_3268, w_028_3269, w_028_3270, w_028_3271, w_028_3273, w_028_3274, w_028_3275, w_028_3276, w_028_3277, w_028_3278, w_028_3279, w_028_3280, w_028_3282, w_028_3284, w_028_3285, w_028_3286, w_028_3288, w_028_3289, w_028_3291, w_028_3292, w_028_3295, w_028_3296, w_028_3297, w_028_3298, w_028_3299, w_028_3300, w_028_3302, w_028_3303, w_028_3304, w_028_3305, w_028_3306, w_028_3307, w_028_3309, w_028_3310, w_028_3311, w_028_3312, w_028_3314, w_028_3315, w_028_3316, w_028_3317, w_028_3318, w_028_3319, w_028_3320, w_028_3322, w_028_3323, w_028_3324, w_028_3325, w_028_3326, w_028_3328, w_028_3329, w_028_3331, w_028_3332, w_028_3333, w_028_3334, w_028_3336, w_028_3338, w_028_3341, w_028_3342, w_028_3343, w_028_3344, w_028_3345, w_028_3346, w_028_3348, w_028_3349, w_028_3353, w_028_3354, w_028_3355, w_028_3356, w_028_3357, w_028_3359, w_028_3363, w_028_3365, w_028_3366, w_028_3367, w_028_3368, w_028_3369, w_028_3371, w_028_3375, w_028_3376, w_028_3381, w_028_3382, w_028_3383, w_028_3384, w_028_3385, w_028_3387, w_028_3390, w_028_3392, w_028_3394, w_028_3396, w_028_3397, w_028_3398, w_028_3399, w_028_3400, w_028_3402, w_028_3403, w_028_3405, w_028_3406, w_028_3408, w_028_3409, w_028_3410, w_028_3412, w_028_3414, w_028_3416, w_028_3417, w_028_3418, w_028_3422, w_028_3423, w_028_3424, w_028_3425, w_028_3427, w_028_3428, w_028_3429, w_028_3430, w_028_3434, w_028_3435, w_028_3436, w_028_3437, w_028_3441, w_028_3442, w_028_3443, w_028_3444, w_028_3445, w_028_3448, w_028_3452, w_028_3453, w_028_3454, w_028_3455, w_028_3456, w_028_3457, w_028_3458, w_028_3459, w_028_3461, w_028_3465, w_028_3468, w_028_3470, w_028_3471, w_028_3472, w_028_3473, w_028_3474, w_028_3478, w_028_3479, w_028_3480, w_028_3482, w_028_3483, w_028_3484, w_028_3485, w_028_3486, w_028_3487, w_028_3488, w_028_3489, w_028_3490, w_028_3492, w_028_3496, w_028_3499, w_028_3500, w_028_3501, w_028_3503, w_028_3505, w_028_3508, w_028_3509, w_028_3511, w_028_3512, w_028_3514, w_028_3515, w_028_3517, w_028_3518, w_028_3520, w_028_3521, w_028_3522, w_028_3524, w_028_3528, w_028_3529, w_028_3530, w_028_3533, w_028_3534, w_028_3535, w_028_3538, w_028_3540, w_028_3542, w_028_3543, w_028_3544, w_028_3545, w_028_3547, w_028_3549, w_028_3550, w_028_3551, w_028_3552, w_028_3553, w_028_3555, w_028_3556, w_028_3558, w_028_3559, w_028_3560, w_028_3561, w_028_3562, w_028_3565, w_028_3566, w_028_3567, w_028_3568, w_028_3570, w_028_3571, w_028_3573, w_028_3574, w_028_3575, w_028_3576, w_028_3577, w_028_3579, w_028_3580, w_028_3581, w_028_3582, w_028_3583, w_028_3584, w_028_3585, w_028_3586, w_028_3587, w_028_3589, w_028_3591, w_028_3592, w_028_3593, w_028_3594, w_028_3595, w_028_3596, w_028_3597, w_028_3598, w_028_3599, w_028_3600, w_028_3601, w_028_3602, w_028_3604;
  wire w_029_001, w_029_002, w_029_003, w_029_004, w_029_006, w_029_007, w_029_008, w_029_009, w_029_010, w_029_011, w_029_013, w_029_014, w_029_015, w_029_016, w_029_018, w_029_019, w_029_020, w_029_021, w_029_022, w_029_023, w_029_024, w_029_025, w_029_026, w_029_027, w_029_028, w_029_031, w_029_033, w_029_034, w_029_036, w_029_037, w_029_038, w_029_040, w_029_041, w_029_042, w_029_043, w_029_044, w_029_045, w_029_046, w_029_047, w_029_048, w_029_049, w_029_050, w_029_052, w_029_053, w_029_054, w_029_055, w_029_056, w_029_057, w_029_059, w_029_060, w_029_061, w_029_063, w_029_064, w_029_065, w_029_066, w_029_067, w_029_068, w_029_069, w_029_070, w_029_071, w_029_072, w_029_073, w_029_074, w_029_075, w_029_076, w_029_077, w_029_078, w_029_079, w_029_081, w_029_082, w_029_083, w_029_084, w_029_085, w_029_086, w_029_087, w_029_088, w_029_089, w_029_090, w_029_093, w_029_094, w_029_095, w_029_096, w_029_098, w_029_099, w_029_100, w_029_101, w_029_102, w_029_103, w_029_104, w_029_105, w_029_106, w_029_108, w_029_109, w_029_111, w_029_112, w_029_113, w_029_114, w_029_115, w_029_116, w_029_117, w_029_118, w_029_119, w_029_120, w_029_121, w_029_122, w_029_123, w_029_124, w_029_125, w_029_126, w_029_127, w_029_128, w_029_130, w_029_131, w_029_132, w_029_133, w_029_134, w_029_135, w_029_136, w_029_137, w_029_138, w_029_139, w_029_140, w_029_141, w_029_142, w_029_144, w_029_145, w_029_146, w_029_147, w_029_148, w_029_149, w_029_150, w_029_151, w_029_152, w_029_153, w_029_154, w_029_155, w_029_156, w_029_157, w_029_158, w_029_159, w_029_160, w_029_161, w_029_162, w_029_163, w_029_164, w_029_165, w_029_167, w_029_168, w_029_169, w_029_170, w_029_171, w_029_172, w_029_174, w_029_176, w_029_177, w_029_178, w_029_179, w_029_180, w_029_181, w_029_182, w_029_183, w_029_185, w_029_186, w_029_187, w_029_188, w_029_189, w_029_190, w_029_193, w_029_194, w_029_195, w_029_196, w_029_197, w_029_198, w_029_199, w_029_200, w_029_201, w_029_202, w_029_203, w_029_204, w_029_205, w_029_206, w_029_207, w_029_208, w_029_209, w_029_210, w_029_211, w_029_212, w_029_214, w_029_215, w_029_216, w_029_217, w_029_218, w_029_220, w_029_221, w_029_222, w_029_223, w_029_224, w_029_225, w_029_226, w_029_227, w_029_228, w_029_230, w_029_231, w_029_233, w_029_234, w_029_235, w_029_236, w_029_237, w_029_238, w_029_240, w_029_241, w_029_242, w_029_243, w_029_244, w_029_245, w_029_246, w_029_248, w_029_249, w_029_251, w_029_252, w_029_253, w_029_254, w_029_255, w_029_256, w_029_259, w_029_260, w_029_262, w_029_263, w_029_264, w_029_265, w_029_266, w_029_267, w_029_268, w_029_269, w_029_270, w_029_271, w_029_272, w_029_273, w_029_274, w_029_275, w_029_276, w_029_277, w_029_278, w_029_279, w_029_280, w_029_281, w_029_282, w_029_283, w_029_284, w_029_286, w_029_287, w_029_288, w_029_289, w_029_291, w_029_292, w_029_293, w_029_294, w_029_295, w_029_296, w_029_297, w_029_298, w_029_299, w_029_300, w_029_301, w_029_302, w_029_303, w_029_304, w_029_305, w_029_306, w_029_308, w_029_309, w_029_310, w_029_311, w_029_312, w_029_313, w_029_314, w_029_315, w_029_316, w_029_317, w_029_318, w_029_319, w_029_320, w_029_323, w_029_324, w_029_326, w_029_327, w_029_328, w_029_329, w_029_330, w_029_331, w_029_333, w_029_334, w_029_335, w_029_336, w_029_337, w_029_338, w_029_339, w_029_340, w_029_341, w_029_343, w_029_344, w_029_345, w_029_346, w_029_350, w_029_352, w_029_354, w_029_355, w_029_356, w_029_357, w_029_358, w_029_359, w_029_360, w_029_361, w_029_362, w_029_363, w_029_364, w_029_366, w_029_367, w_029_368, w_029_369, w_029_370, w_029_372, w_029_373, w_029_374, w_029_375, w_029_376, w_029_377, w_029_378, w_029_379, w_029_380, w_029_381, w_029_382, w_029_383, w_029_384, w_029_386, w_029_387, w_029_388, w_029_389, w_029_390, w_029_391, w_029_392, w_029_394, w_029_395, w_029_396, w_029_397, w_029_398, w_029_399, w_029_400, w_029_401, w_029_402, w_029_403, w_029_404, w_029_405, w_029_406, w_029_408, w_029_410, w_029_411, w_029_412, w_029_413, w_029_414, w_029_415, w_029_416, w_029_418, w_029_420, w_029_421, w_029_422, w_029_423, w_029_424, w_029_425, w_029_426, w_029_427, w_029_429, w_029_430, w_029_431, w_029_432, w_029_433, w_029_434, w_029_435, w_029_436, w_029_437, w_029_438, w_029_439, w_029_440, w_029_441, w_029_442, w_029_443, w_029_444, w_029_445, w_029_446, w_029_447, w_029_448, w_029_449, w_029_450, w_029_451, w_029_452, w_029_453, w_029_454, w_029_455, w_029_456, w_029_457, w_029_458, w_029_459, w_029_460, w_029_462, w_029_463, w_029_464, w_029_465, w_029_466, w_029_467, w_029_468, w_029_470, w_029_471, w_029_472, w_029_473, w_029_474, w_029_475, w_029_476, w_029_477, w_029_480, w_029_481, w_029_482, w_029_483, w_029_484, w_029_485, w_029_486, w_029_487, w_029_489, w_029_491, w_029_492, w_029_493, w_029_494, w_029_495, w_029_497, w_029_498, w_029_499, w_029_500, w_029_501, w_029_502, w_029_503, w_029_504, w_029_505, w_029_506, w_029_507, w_029_508, w_029_510, w_029_511, w_029_513, w_029_514, w_029_515, w_029_516, w_029_517, w_029_518, w_029_519, w_029_521, w_029_523, w_029_524, w_029_525, w_029_526, w_029_527, w_029_528, w_029_531, w_029_533, w_029_534, w_029_536, w_029_537, w_029_538, w_029_539, w_029_540, w_029_541, w_029_542, w_029_543, w_029_546, w_029_547, w_029_548, w_029_549, w_029_550, w_029_551, w_029_552, w_029_553, w_029_554, w_029_555, w_029_556, w_029_557, w_029_558, w_029_559, w_029_560, w_029_561, w_029_562, w_029_563, w_029_564, w_029_565, w_029_567, w_029_568, w_029_569, w_029_570, w_029_571, w_029_572, w_029_573, w_029_574, w_029_575, w_029_576, w_029_577, w_029_578, w_029_579, w_029_580, w_029_582, w_029_583, w_029_584, w_029_586, w_029_588, w_029_589, w_029_590, w_029_591, w_029_592, w_029_593, w_029_594, w_029_595, w_029_598, w_029_599, w_029_600, w_029_601, w_029_602, w_029_603, w_029_604, w_029_605, w_029_606, w_029_607, w_029_608, w_029_609, w_029_610, w_029_611, w_029_612, w_029_613, w_029_614, w_029_615, w_029_616, w_029_618, w_029_620, w_029_621, w_029_622, w_029_623, w_029_624, w_029_625, w_029_626, w_029_627, w_029_628, w_029_629, w_029_630, w_029_631, w_029_633, w_029_634, w_029_635, w_029_636, w_029_637, w_029_638, w_029_639, w_029_640, w_029_641, w_029_642, w_029_643, w_029_645, w_029_646, w_029_647, w_029_648, w_029_650, w_029_651, w_029_652, w_029_654, w_029_655, w_029_656, w_029_657, w_029_660, w_029_661, w_029_662, w_029_663, w_029_664, w_029_665, w_029_666, w_029_667, w_029_668, w_029_669, w_029_670, w_029_671, w_029_672, w_029_673, w_029_674, w_029_675, w_029_676, w_029_677, w_029_678, w_029_679, w_029_680, w_029_681, w_029_682, w_029_683, w_029_684, w_029_685, w_029_686, w_029_687, w_029_688, w_029_689, w_029_690, w_029_691, w_029_692, w_029_693, w_029_694, w_029_695, w_029_696, w_029_698, w_029_699, w_029_700, w_029_701, w_029_703, w_029_704, w_029_705, w_029_706, w_029_707, w_029_708, w_029_709, w_029_710, w_029_711, w_029_712, w_029_713, w_029_714, w_029_715, w_029_716, w_029_717, w_029_718, w_029_719, w_029_720, w_029_721, w_029_722, w_029_723, w_029_724, w_029_725, w_029_726, w_029_727, w_029_729, w_029_730, w_029_731, w_029_732, w_029_733, w_029_734, w_029_735, w_029_736, w_029_737, w_029_738, w_029_739, w_029_740, w_029_741, w_029_742, w_029_743, w_029_744, w_029_746, w_029_747, w_029_748, w_029_749, w_029_750, w_029_751, w_029_752, w_029_754, w_029_755, w_029_756, w_029_757, w_029_758, w_029_759, w_029_760, w_029_761, w_029_762, w_029_764, w_029_765, w_029_766, w_029_767, w_029_769, w_029_770, w_029_771, w_029_772, w_029_773, w_029_775, w_029_777, w_029_778, w_029_779, w_029_780, w_029_781, w_029_782, w_029_783, w_029_784, w_029_785, w_029_786, w_029_787, w_029_788, w_029_789, w_029_790, w_029_791, w_029_792, w_029_793, w_029_794, w_029_795, w_029_797, w_029_798, w_029_799, w_029_802, w_029_803, w_029_804, w_029_806, w_029_807, w_029_808, w_029_809, w_029_810, w_029_811, w_029_812, w_029_813, w_029_815, w_029_816, w_029_817, w_029_818, w_029_820, w_029_821, w_029_822, w_029_824, w_029_825, w_029_826, w_029_828, w_029_829, w_029_830, w_029_831, w_029_832, w_029_833, w_029_834, w_029_835, w_029_836, w_029_837, w_029_838, w_029_839, w_029_840, w_029_842, w_029_843, w_029_844, w_029_845, w_029_846, w_029_847, w_029_848, w_029_849, w_029_850, w_029_851, w_029_852, w_029_853, w_029_856, w_029_857, w_029_858, w_029_859, w_029_860, w_029_861, w_029_862, w_029_863, w_029_864, w_029_865, w_029_866, w_029_867, w_029_868, w_029_869, w_029_870, w_029_871, w_029_872, w_029_873, w_029_874, w_029_875, w_029_876, w_029_877, w_029_878, w_029_880, w_029_881, w_029_882, w_029_883, w_029_884, w_029_885, w_029_886, w_029_887, w_029_888, w_029_890, w_029_891, w_029_892, w_029_893, w_029_894, w_029_895, w_029_896, w_029_897, w_029_898, w_029_899, w_029_900, w_029_901, w_029_903, w_029_904, w_029_905, w_029_906, w_029_907, w_029_908, w_029_909, w_029_910, w_029_911, w_029_912, w_029_913, w_029_914, w_029_915, w_029_916, w_029_917, w_029_918, w_029_919, w_029_920, w_029_921, w_029_922, w_029_923, w_029_925, w_029_926, w_029_927, w_029_930, w_029_932, w_029_933, w_029_934, w_029_935, w_029_936, w_029_937, w_029_939, w_029_940, w_029_941, w_029_942, w_029_943, w_029_945, w_029_947, w_029_948, w_029_949, w_029_950, w_029_951, w_029_952, w_029_953, w_029_954, w_029_955, w_029_956, w_029_957, w_029_958, w_029_959, w_029_960, w_029_961, w_029_962, w_029_964, w_029_965, w_029_966, w_029_967, w_029_969, w_029_970, w_029_971, w_029_972, w_029_973, w_029_974, w_029_975, w_029_976, w_029_977, w_029_978, w_029_979, w_029_981, w_029_982, w_029_984, w_029_985, w_029_986, w_029_987, w_029_988, w_029_989, w_029_990, w_029_991, w_029_992, w_029_993, w_029_994, w_029_995, w_029_996, w_029_997, w_029_998, w_029_1001, w_029_1002, w_029_1003, w_029_1004, w_029_1005, w_029_1006, w_029_1007, w_029_1008, w_029_1010, w_029_1011, w_029_1013, w_029_1014, w_029_1015, w_029_1016, w_029_1017, w_029_1019, w_029_1020, w_029_1021, w_029_1022, w_029_1023, w_029_1024, w_029_1025, w_029_1027, w_029_1028, w_029_1029, w_029_1030, w_029_1031, w_029_1033, w_029_1034, w_029_1035, w_029_1036, w_029_1037, w_029_1038, w_029_1039, w_029_1040, w_029_1041, w_029_1043, w_029_1044, w_029_1045, w_029_1046, w_029_1047, w_029_1048, w_029_1049, w_029_1050, w_029_1051, w_029_1052, w_029_1053, w_029_1054, w_029_1055, w_029_1058, w_029_1059, w_029_1060, w_029_1061, w_029_1062, w_029_1063, w_029_1066, w_029_1067, w_029_1068, w_029_1070, w_029_1071, w_029_1072, w_029_1074, w_029_1076, w_029_1077, w_029_1078, w_029_1079, w_029_1081, w_029_1082, w_029_1083, w_029_1084, w_029_1085, w_029_1086, w_029_1087, w_029_1088, w_029_1089, w_029_1090, w_029_1091, w_029_1092, w_029_1093, w_029_1094, w_029_1096, w_029_1097, w_029_1098, w_029_1100, w_029_1101, w_029_1102, w_029_1103, w_029_1104, w_029_1105, w_029_1106, w_029_1107, w_029_1108, w_029_1109, w_029_1110, w_029_1111, w_029_1112, w_029_1114, w_029_1115, w_029_1116, w_029_1117, w_029_1118, w_029_1120, w_029_1122, w_029_1123, w_029_1124, w_029_1125, w_029_1126, w_029_1127, w_029_1128, w_029_1129, w_029_1130, w_029_1131, w_029_1132, w_029_1133, w_029_1134, w_029_1135, w_029_1136, w_029_1137, w_029_1138, w_029_1139, w_029_1141, w_029_1142, w_029_1144, w_029_1145, w_029_1146, w_029_1147, w_029_1148, w_029_1149, w_029_1150, w_029_1151, w_029_1153, w_029_1154, w_029_1155, w_029_1156, w_029_1158, w_029_1159, w_029_1160, w_029_1161, w_029_1162, w_029_1163, w_029_1164, w_029_1165, w_029_1166, w_029_1167, w_029_1168, w_029_1169, w_029_1170, w_029_1171, w_029_1172, w_029_1173, w_029_1174, w_029_1175, w_029_1176, w_029_1177, w_029_1178, w_029_1179, w_029_1181, w_029_1182, w_029_1184, w_029_1185, w_029_1186, w_029_1187, w_029_1188, w_029_1189, w_029_1190, w_029_1191, w_029_1192, w_029_1194, w_029_1195, w_029_1196, w_029_1197, w_029_1198, w_029_1199, w_029_1200, w_029_1201, w_029_1202, w_029_1203, w_029_1204, w_029_1205, w_029_1206, w_029_1208, w_029_1210, w_029_1211, w_029_1212, w_029_1214, w_029_1215, w_029_1216, w_029_1217, w_029_1218, w_029_1219, w_029_1220, w_029_1221, w_029_1222, w_029_1223, w_029_1224, w_029_1225, w_029_1226, w_029_1227, w_029_1228, w_029_1229, w_029_1230, w_029_1231, w_029_1232, w_029_1233, w_029_1234, w_029_1235, w_029_1236, w_029_1237, w_029_1238, w_029_1239, w_029_1240, w_029_1241, w_029_1242, w_029_1243, w_029_1244, w_029_1245, w_029_1246, w_029_1247, w_029_1248, w_029_1249, w_029_1251, w_029_1252, w_029_1254, w_029_1256, w_029_1257, w_029_1258, w_029_1259, w_029_1260, w_029_1261, w_029_1263, w_029_1264, w_029_1265, w_029_1266, w_029_1267, w_029_1268, w_029_1270, w_029_1271, w_029_1273, w_029_1274, w_029_1275, w_029_1276, w_029_1278, w_029_1279, w_029_1280, w_029_1281, w_029_1282, w_029_1283, w_029_1284, w_029_1285, w_029_1287, w_029_1288, w_029_1289, w_029_1290, w_029_1291, w_029_1293, w_029_1294, w_029_1295, w_029_1296, w_029_1297, w_029_1298, w_029_1300, w_029_1301, w_029_1302, w_029_1303, w_029_1304, w_029_1305, w_029_1306, w_029_1307, w_029_1308, w_029_1309, w_029_1310, w_029_1312, w_029_1313, w_029_1315, w_029_1316, w_029_1317, w_029_1318, w_029_1319, w_029_1320, w_029_1321, w_029_1322, w_029_1323, w_029_1324, w_029_1325, w_029_1326, w_029_1327, w_029_1328, w_029_1329, w_029_1330, w_029_1331, w_029_1332, w_029_1333, w_029_1334, w_029_1335, w_029_1336, w_029_1337, w_029_1338, w_029_1339, w_029_1340, w_029_1341, w_029_1343, w_029_1345, w_029_1346, w_029_1347, w_029_1348, w_029_1350, w_029_1351, w_029_1352, w_029_1354, w_029_1355, w_029_1356, w_029_1357, w_029_1358, w_029_1359, w_029_1360, w_029_1361, w_029_1362, w_029_1363, w_029_1365, w_029_1366, w_029_1367, w_029_1368, w_029_1369, w_029_1370, w_029_1371, w_029_1372, w_029_1373, w_029_1374, w_029_1375, w_029_1376, w_029_1377, w_029_1379, w_029_1380, w_029_1381, w_029_1382, w_029_1383, w_029_1384, w_029_1385, w_029_1386, w_029_1387, w_029_1388, w_029_1389, w_029_1390, w_029_1391, w_029_1392, w_029_1393, w_029_1394, w_029_1395, w_029_1396, w_029_1397, w_029_1398, w_029_1399, w_029_1402, w_029_1403, w_029_1404, w_029_1406, w_029_1407, w_029_1408, w_029_1409, w_029_1411, w_029_1412, w_029_1413, w_029_1415, w_029_1416, w_029_1417, w_029_1418, w_029_1419, w_029_1420, w_029_1421, w_029_1422, w_029_1423, w_029_1424, w_029_1425, w_029_1426, w_029_1427, w_029_1428, w_029_1429, w_029_1430, w_029_1431, w_029_1432, w_029_1433, w_029_1435, w_029_1436, w_029_1438, w_029_1439, w_029_1440, w_029_1441, w_029_1442, w_029_1443, w_029_1444, w_029_1445, w_029_1446, w_029_1447, w_029_1448, w_029_1449, w_029_1451, w_029_1454, w_029_1455, w_029_1456, w_029_1457, w_029_1458, w_029_1459, w_029_1460, w_029_1461, w_029_1462, w_029_1463, w_029_1464, w_029_1465, w_029_1466, w_029_1467, w_029_1469, w_029_1470, w_029_1471, w_029_1472, w_029_1473, w_029_1474, w_029_1475, w_029_1476, w_029_1477, w_029_1478, w_029_1480, w_029_1481, w_029_1482, w_029_1483, w_029_1484, w_029_1485, w_029_1486, w_029_1487, w_029_1488, w_029_1489, w_029_1490, w_029_1491, w_029_1493, w_029_1494, w_029_1495, w_029_1496, w_029_1497, w_029_1498, w_029_1499, w_029_1500, w_029_1501, w_029_1502, w_029_1503, w_029_1504, w_029_1505, w_029_1507, w_029_1508, w_029_1509, w_029_1510, w_029_1511, w_029_1512, w_029_1513, w_029_1514, w_029_1515, w_029_1516, w_029_1517, w_029_1519, w_029_1520, w_029_1521, w_029_1522, w_029_1523, w_029_1524, w_029_1525, w_029_1526, w_029_1527, w_029_1528, w_029_1529, w_029_1530, w_029_1531, w_029_1533, w_029_1534, w_029_1535, w_029_1536, w_029_1537, w_029_1539, w_029_1540, w_029_1541, w_029_1542, w_029_1543, w_029_1544, w_029_1545, w_029_1546, w_029_1547, w_029_1548, w_029_1549, w_029_1550, w_029_1553, w_029_1554, w_029_1555, w_029_1556, w_029_1557, w_029_1558, w_029_1560, w_029_1561, w_029_1562, w_029_1563, w_029_1564, w_029_1565, w_029_1566, w_029_1567, w_029_1568, w_029_1569, w_029_1570, w_029_1571, w_029_1572, w_029_1574, w_029_1575, w_029_1576, w_029_1578, w_029_1579, w_029_1581, w_029_1582, w_029_1583, w_029_1584, w_029_1585, w_029_1586, w_029_1588, w_029_1589, w_029_1590, w_029_1593, w_029_1594, w_029_1595, w_029_1596, w_029_1597, w_029_1598, w_029_1599, w_029_1600, w_029_1601, w_029_1602, w_029_1603, w_029_1605, w_029_1606, w_029_1607, w_029_1608, w_029_1609, w_029_1610, w_029_1611, w_029_1612, w_029_1613, w_029_1614, w_029_1615, w_029_1616, w_029_1617, w_029_1618, w_029_1619, w_029_1620, w_029_1621, w_029_1622, w_029_1623, w_029_1626, w_029_1627, w_029_1629, w_029_1630, w_029_1631, w_029_1632, w_029_1633, w_029_1634, w_029_1635, w_029_1637, w_029_1638, w_029_1639, w_029_1640, w_029_1641, w_029_1642, w_029_1643, w_029_1644, w_029_1645, w_029_1646, w_029_1648, w_029_1649, w_029_1650, w_029_1651, w_029_1652, w_029_1653, w_029_1654, w_029_1655, w_029_1656, w_029_1657, w_029_1660, w_029_1661, w_029_1662, w_029_1663, w_029_1664, w_029_1665, w_029_1666, w_029_1667, w_029_1668, w_029_1669, w_029_1670, w_029_1671, w_029_1672, w_029_1673, w_029_1674, w_029_1676, w_029_1677, w_029_1678, w_029_1679, w_029_1680, w_029_1681, w_029_1682, w_029_1684, w_029_1685, w_029_1686, w_029_1687, w_029_1690, w_029_1691, w_029_1692, w_029_1693, w_029_1694, w_029_1695, w_029_1696, w_029_1697, w_029_1700, w_029_1701, w_029_1702, w_029_1703, w_029_1705, w_029_1706, w_029_1707, w_029_1708, w_029_1709, w_029_1710, w_029_1711, w_029_1713, w_029_1714, w_029_1715, w_029_1716, w_029_1717, w_029_1718, w_029_1719, w_029_1720, w_029_1723, w_029_1724, w_029_1725, w_029_1726, w_029_1727, w_029_1728, w_029_1729, w_029_1730, w_029_1731, w_029_1732, w_029_1733, w_029_1734, w_029_1736, w_029_1737, w_029_1738, w_029_1739, w_029_1740, w_029_1741, w_029_1742, w_029_1743, w_029_1744, w_029_1745, w_029_1746, w_029_1749, w_029_1750, w_029_1751, w_029_1752, w_029_1753, w_029_1755, w_029_1756, w_029_1758, w_029_1760, w_029_1761, w_029_1762, w_029_1764, w_029_1765, w_029_1766, w_029_1767, w_029_1768, w_029_1769, w_029_1770, w_029_1771, w_029_1772, w_029_1773, w_029_1774, w_029_1775, w_029_1776, w_029_1777, w_029_1779, w_029_1780, w_029_1781, w_029_1782, w_029_1783, w_029_1784, w_029_1785, w_029_1786, w_029_1787, w_029_1788, w_029_1789, w_029_1790, w_029_1791, w_029_1792, w_029_1794, w_029_1795, w_029_1796, w_029_1797, w_029_1799, w_029_1800, w_029_1801, w_029_1802, w_029_1803, w_029_1804, w_029_1806, w_029_1807, w_029_1808, w_029_1809, w_029_1810, w_029_1811, w_029_1812, w_029_1813, w_029_1815, w_029_1816, w_029_1818, w_029_1819, w_029_1821, w_029_1822, w_029_1824, w_029_1825, w_029_1827, w_029_1828, w_029_1829, w_029_1830, w_029_1831, w_029_1833, w_029_1835, w_029_1836, w_029_1837, w_029_1838, w_029_1839, w_029_1841, w_029_1842, w_029_1844, w_029_1845, w_029_1846, w_029_1847, w_029_1848, w_029_1849, w_029_1850, w_029_1851, w_029_1852, w_029_1853, w_029_1854, w_029_1855, w_029_1856, w_029_1857, w_029_1858, w_029_1859, w_029_1860, w_029_1861, w_029_1862, w_029_1863, w_029_1864, w_029_1865, w_029_1866, w_029_1867, w_029_1868, w_029_1869, w_029_1870, w_029_1871, w_029_1872, w_029_1873, w_029_1874, w_029_1875, w_029_1876, w_029_1877, w_029_1878, w_029_1879, w_029_1880, w_029_1881, w_029_1882, w_029_1883, w_029_1884, w_029_1885, w_029_1886, w_029_1887, w_029_1888, w_029_1889, w_029_1890, w_029_1891, w_029_1892, w_029_1893, w_029_1895, w_029_1897, w_029_1898, w_029_1899, w_029_1901, w_029_1903, w_029_1904, w_029_1905, w_029_1907, w_029_1908, w_029_1909, w_029_1910, w_029_1911, w_029_1912, w_029_1914, w_029_1915, w_029_1916, w_029_1917, w_029_1918, w_029_1919, w_029_1921, w_029_1922, w_029_1923, w_029_1924, w_029_1925, w_029_1926, w_029_1927, w_029_1928, w_029_1929, w_029_1930, w_029_1931, w_029_1932, w_029_1934, w_029_1935, w_029_1936, w_029_1938, w_029_1939, w_029_1940, w_029_1942, w_029_1943, w_029_1944, w_029_1945, w_029_1946, w_029_1947, w_029_1948, w_029_1949, w_029_1950, w_029_1951, w_029_1953, w_029_1955, w_029_1956, w_029_1957, w_029_1958, w_029_1959, w_029_1960, w_029_1961, w_029_1963, w_029_1965, w_029_1966, w_029_1967, w_029_1968, w_029_1969, w_029_1970, w_029_1972, w_029_1973, w_029_1974, w_029_1975, w_029_1976, w_029_1977, w_029_1978, w_029_1979, w_029_1980, w_029_1981, w_029_1982, w_029_1983, w_029_1984, w_029_1985, w_029_1986, w_029_1987, w_029_1988, w_029_1989, w_029_1990, w_029_1991, w_029_1992, w_029_1993, w_029_1994, w_029_1995, w_029_1996, w_029_1997, w_029_1999, w_029_2000, w_029_2001, w_029_2002, w_029_2003, w_029_2004, w_029_2005, w_029_2006, w_029_2007, w_029_2008, w_029_2010, w_029_2011, w_029_2012, w_029_2013, w_029_2015, w_029_2016, w_029_2017, w_029_2018, w_029_2019, w_029_2020, w_029_2021, w_029_2022, w_029_2024, w_029_2025, w_029_2026, w_029_2027, w_029_2028, w_029_2029, w_029_2030, w_029_2031, w_029_2032, w_029_2033, w_029_2034, w_029_2035, w_029_2037, w_029_2038, w_029_2039, w_029_2040, w_029_2041, w_029_2042, w_029_2043, w_029_2044, w_029_2045, w_029_2046, w_029_2047, w_029_2048, w_029_2049, w_029_2050, w_029_2051, w_029_2052, w_029_2053, w_029_2054, w_029_2055, w_029_2057, w_029_2059, w_029_2060, w_029_2061, w_029_2062, w_029_2063, w_029_2065, w_029_2066, w_029_2067, w_029_2068, w_029_2069, w_029_2070, w_029_2071, w_029_2072, w_029_2073, w_029_2075, w_029_2076, w_029_2077, w_029_2078, w_029_2079, w_029_2080, w_029_2081, w_029_2082, w_029_2083, w_029_2084, w_029_2085, w_029_2086, w_029_2087, w_029_2088, w_029_2090, w_029_2091, w_029_2092, w_029_2093, w_029_2096, w_029_2097, w_029_2098, w_029_2100, w_029_2101, w_029_2102, w_029_2103, w_029_2104, w_029_2105, w_029_2106, w_029_2107, w_029_2108, w_029_2109, w_029_2110, w_029_2111, w_029_2112, w_029_2113, w_029_2114, w_029_2116, w_029_2117, w_029_2118, w_029_2119, w_029_2120, w_029_2121, w_029_2122, w_029_2123, w_029_2125, w_029_2128, w_029_2129, w_029_2130, w_029_2131, w_029_2132, w_029_2133, w_029_2134, w_029_2135, w_029_2136, w_029_2137, w_029_2138, w_029_2139, w_029_2140, w_029_2141, w_029_2143, w_029_2144, w_029_2145, w_029_2146, w_029_2147, w_029_2149, w_029_2150, w_029_2152, w_029_2153, w_029_2154, w_029_2155, w_029_2156, w_029_2158, w_029_2159, w_029_2160, w_029_2161, w_029_2162, w_029_2163, w_029_2165, w_029_2166, w_029_2167, w_029_2168, w_029_2169, w_029_2170, w_029_2172, w_029_2174, w_029_2176, w_029_2178, w_029_2180, w_029_2181, w_029_2182, w_029_2184, w_029_2185, w_029_2186, w_029_2187, w_029_2188, w_029_2190, w_029_2192, w_029_2194, w_029_2195, w_029_2196, w_029_2197, w_029_2198, w_029_2199, w_029_2200, w_029_2201, w_029_2202, w_029_2203, w_029_2204, w_029_2206, w_029_2207, w_029_2208, w_029_2209, w_029_2210, w_029_2211, w_029_2212, w_029_2213, w_029_2214, w_029_2215, w_029_2216, w_029_2218, w_029_2219, w_029_2221, w_029_2222, w_029_2223, w_029_2224, w_029_2225, w_029_2226, w_029_2227, w_029_2228, w_029_2229, w_029_2230, w_029_2231, w_029_2232, w_029_2233, w_029_2234, w_029_2235, w_029_2236, w_029_2237, w_029_2238, w_029_2239, w_029_2240, w_029_2241, w_029_2242, w_029_2243, w_029_2244, w_029_2245, w_029_2246, w_029_2247, w_029_2248, w_029_2249, w_029_2250, w_029_2253, w_029_2254, w_029_2256, w_029_2257, w_029_2258, w_029_2259, w_029_2260, w_029_2261, w_029_2263, w_029_2264, w_029_2265, w_029_2266, w_029_2268, w_029_2270, w_029_2271, w_029_2272, w_029_2273, w_029_2274, w_029_2275, w_029_2276, w_029_2277, w_029_2278, w_029_2279, w_029_2280, w_029_2281, w_029_2285, w_029_2287, w_029_2288, w_029_2289, w_029_2290, w_029_2291, w_029_2292, w_029_2296, w_029_2299, w_029_2300, w_029_2302, w_029_2303, w_029_2304, w_029_2305, w_029_2306, w_029_2309, w_029_2310, w_029_2313, w_029_2314, w_029_2315, w_029_2316, w_029_2317, w_029_2320, w_029_2321, w_029_2322, w_029_2323, w_029_2325, w_029_2326, w_029_2327, w_029_2329, w_029_2331, w_029_2334, w_029_2335, w_029_2336, w_029_2337, w_029_2338, w_029_2339, w_029_2342, w_029_2344, w_029_2345, w_029_2346, w_029_2348, w_029_2349, w_029_2351, w_029_2353, w_029_2354, w_029_2355, w_029_2356, w_029_2358, w_029_2360, w_029_2361, w_029_2365, w_029_2366, w_029_2367, w_029_2368, w_029_2369, w_029_2370, w_029_2373, w_029_2375, w_029_2376, w_029_2377, w_029_2378, w_029_2385, w_029_2388, w_029_2391, w_029_2393, w_029_2395, w_029_2400, w_029_2401, w_029_2402, w_029_2403, w_029_2405, w_029_2406, w_029_2407, w_029_2408, w_029_2409, w_029_2412, w_029_2414, w_029_2417, w_029_2418, w_029_2419, w_029_2421, w_029_2422, w_029_2423, w_029_2425, w_029_2426, w_029_2428, w_029_2429, w_029_2430, w_029_2431, w_029_2432, w_029_2434, w_029_2436, w_029_2437, w_029_2439, w_029_2440, w_029_2442, w_029_2443, w_029_2446, w_029_2447, w_029_2448, w_029_2450, w_029_2451, w_029_2455, w_029_2456, w_029_2458, w_029_2464, w_029_2465, w_029_2466, w_029_2471, w_029_2473, w_029_2474, w_029_2475, w_029_2477, w_029_2479, w_029_2481, w_029_2485, w_029_2486, w_029_2487, w_029_2488, w_029_2489, w_029_2490, w_029_2493, w_029_2495, w_029_2496, w_029_2498, w_029_2500, w_029_2501, w_029_2502, w_029_2503, w_029_2505, w_029_2506, w_029_2508, w_029_2509, w_029_2510, w_029_2511, w_029_2512, w_029_2513, w_029_2516, w_029_2517, w_029_2518, w_029_2519, w_029_2520, w_029_2521, w_029_2522, w_029_2527, w_029_2528, w_029_2529, w_029_2532, w_029_2533, w_029_2534, w_029_2536, w_029_2538, w_029_2539, w_029_2540, w_029_2542, w_029_2543, w_029_2544, w_029_2545, w_029_2546, w_029_2547, w_029_2548, w_029_2550, w_029_2552, w_029_2553, w_029_2555, w_029_2557, w_029_2558, w_029_2560, w_029_2563, w_029_2564, w_029_2565, w_029_2566, w_029_2568, w_029_2569, w_029_2570, w_029_2571, w_029_2572, w_029_2573, w_029_2574, w_029_2576, w_029_2578, w_029_2579, w_029_2580, w_029_2581, w_029_2583, w_029_2584, w_029_2585, w_029_2586, w_029_2587, w_029_2588, w_029_2589, w_029_2590, w_029_2591, w_029_2592, w_029_2593, w_029_2594, w_029_2595, w_029_2597, w_029_2598, w_029_2599, w_029_2600, w_029_2601, w_029_2603, w_029_2605, w_029_2606, w_029_2607, w_029_2609, w_029_2611, w_029_2612, w_029_2613, w_029_2614, w_029_2615, w_029_2616, w_029_2618, w_029_2619, w_029_2620, w_029_2621, w_029_2622, w_029_2624, w_029_2625, w_029_2626, w_029_2627, w_029_2628, w_029_2629, w_029_2630, w_029_2631, w_029_2632, w_029_2633, w_029_2635, w_029_2636, w_029_2638, w_029_2639, w_029_2640, w_029_2641, w_029_2642, w_029_2646, w_029_2649, w_029_2651, w_029_2652, w_029_2653, w_029_2654, w_029_2655, w_029_2656, w_029_2657, w_029_2658, w_029_2663, w_029_2666, w_029_2669, w_029_2670, w_029_2671, w_029_2673, w_029_2674, w_029_2676, w_029_2677, w_029_2678, w_029_2679, w_029_2680, w_029_2681, w_029_2682, w_029_2683, w_029_2684, w_029_2685, w_029_2686, w_029_2687, w_029_2688, w_029_2689, w_029_2692, w_029_2693, w_029_2694, w_029_2696, w_029_2697, w_029_2701, w_029_2703, w_029_2704, w_029_2705, w_029_2706, w_029_2709, w_029_2711, w_029_2712, w_029_2713, w_029_2715, w_029_2717, w_029_2718, w_029_2719, w_029_2721, w_029_2722, w_029_2723;
  wire w_030_000, w_030_001, w_030_002, w_030_003, w_030_004, w_030_005, w_030_006, w_030_007, w_030_008, w_030_009, w_030_010, w_030_011, w_030_012, w_030_013, w_030_014, w_030_015, w_030_016, w_030_017, w_030_018, w_030_019, w_030_020, w_030_021, w_030_022, w_030_023, w_030_024, w_030_025, w_030_026, w_030_027, w_030_028, w_030_029, w_030_030, w_030_031, w_030_032, w_030_035, w_030_036, w_030_038, w_030_039, w_030_040, w_030_041, w_030_042, w_030_043, w_030_044, w_030_046, w_030_047, w_030_048, w_030_049, w_030_050, w_030_051, w_030_053, w_030_054, w_030_055, w_030_056, w_030_057, w_030_058, w_030_059, w_030_060, w_030_061, w_030_062, w_030_063, w_030_064, w_030_065, w_030_066, w_030_067, w_030_068, w_030_069, w_030_070, w_030_071, w_030_072, w_030_073, w_030_074, w_030_075, w_030_076, w_030_077, w_030_078, w_030_079, w_030_080, w_030_081, w_030_082, w_030_083, w_030_084, w_030_085, w_030_086, w_030_087, w_030_088, w_030_089, w_030_090, w_030_091, w_030_092, w_030_093, w_030_094, w_030_095, w_030_096, w_030_097, w_030_098, w_030_099, w_030_100, w_030_101, w_030_102, w_030_103, w_030_104, w_030_105, w_030_106, w_030_107, w_030_108, w_030_109, w_030_111, w_030_113, w_030_114, w_030_115, w_030_117, w_030_118, w_030_120, w_030_121, w_030_122, w_030_123, w_030_124, w_030_125, w_030_126, w_030_127, w_030_128, w_030_129, w_030_130, w_030_131, w_030_132, w_030_133, w_030_134, w_030_135, w_030_136, w_030_137, w_030_138, w_030_139, w_030_140, w_030_141, w_030_142, w_030_143, w_030_144, w_030_145, w_030_146, w_030_148, w_030_149, w_030_150, w_030_151, w_030_152, w_030_154, w_030_155, w_030_156, w_030_157, w_030_158, w_030_159, w_030_160, w_030_161, w_030_162, w_030_163, w_030_164, w_030_165, w_030_166, w_030_167, w_030_168, w_030_169, w_030_170, w_030_171, w_030_172, w_030_173, w_030_174, w_030_175, w_030_176, w_030_177, w_030_178, w_030_179, w_030_180, w_030_181, w_030_182, w_030_183, w_030_184, w_030_185, w_030_186, w_030_187, w_030_188, w_030_189, w_030_190, w_030_191, w_030_192, w_030_193, w_030_194, w_030_195, w_030_196, w_030_197, w_030_198, w_030_199, w_030_200, w_030_201, w_030_202, w_030_203, w_030_204, w_030_205, w_030_206, w_030_207, w_030_208, w_030_209, w_030_210, w_030_211, w_030_212, w_030_213, w_030_214, w_030_215, w_030_216, w_030_217, w_030_218, w_030_219, w_030_220, w_030_221, w_030_222, w_030_223, w_030_224, w_030_225, w_030_226, w_030_227, w_030_228, w_030_229, w_030_230, w_030_231, w_030_232, w_030_233, w_030_234, w_030_235, w_030_236, w_030_237, w_030_238, w_030_239, w_030_240, w_030_241, w_030_242, w_030_243, w_030_244, w_030_245, w_030_246, w_030_247, w_030_248, w_030_249, w_030_250, w_030_251, w_030_252, w_030_253, w_030_254, w_030_255, w_030_256, w_030_258, w_030_259, w_030_260, w_030_261, w_030_262, w_030_263, w_030_264, w_030_265, w_030_266, w_030_267, w_030_268, w_030_269, w_030_270, w_030_272, w_030_273, w_030_274, w_030_275, w_030_276, w_030_277, w_030_278, w_030_279, w_030_280, w_030_281, w_030_282, w_030_283, w_030_285, w_030_286, w_030_287, w_030_288, w_030_289, w_030_290, w_030_291, w_030_292, w_030_293, w_030_294, w_030_295, w_030_296, w_030_297, w_030_298, w_030_299, w_030_300, w_030_301, w_030_302, w_030_303, w_030_304, w_030_305, w_030_306, w_030_307, w_030_309, w_030_310, w_030_311, w_030_312, w_030_313, w_030_314, w_030_315, w_030_316, w_030_317, w_030_318, w_030_319, w_030_320, w_030_321, w_030_322, w_030_323, w_030_324, w_030_325, w_030_326, w_030_327, w_030_328, w_030_329, w_030_330, w_030_331, w_030_332, w_030_333, w_030_334, w_030_335, w_030_336, w_030_337, w_030_338, w_030_339, w_030_340, w_030_341, w_030_342, w_030_343, w_030_344, w_030_345, w_030_347, w_030_348, w_030_349, w_030_350, w_030_351, w_030_352, w_030_353, w_030_354, w_030_355, w_030_356, w_030_357, w_030_358, w_030_359, w_030_360, w_030_361, w_030_362, w_030_363, w_030_364, w_030_365, w_030_366, w_030_367, w_030_368, w_030_370, w_030_371, w_030_372, w_030_373, w_030_375, w_030_376, w_030_377, w_030_378, w_030_379, w_030_380, w_030_381, w_030_382, w_030_383, w_030_384, w_030_385, w_030_386, w_030_388, w_030_389, w_030_390, w_030_391, w_030_392, w_030_394, w_030_395, w_030_396, w_030_397, w_030_398, w_030_399, w_030_400, w_030_401, w_030_403, w_030_405, w_030_406, w_030_407, w_030_408, w_030_409, w_030_410, w_030_411, w_030_412, w_030_413, w_030_414, w_030_415, w_030_416, w_030_417, w_030_418, w_030_419, w_030_420, w_030_421, w_030_422, w_030_423, w_030_424, w_030_425, w_030_426, w_030_427, w_030_428, w_030_429, w_030_430, w_030_431, w_030_432, w_030_433, w_030_434, w_030_435, w_030_436, w_030_437, w_030_438, w_030_439, w_030_440, w_030_441, w_030_442, w_030_444, w_030_445, w_030_446, w_030_447, w_030_448, w_030_449, w_030_450, w_030_451, w_030_452, w_030_453, w_030_454, w_030_455, w_030_456, w_030_457, w_030_458, w_030_459, w_030_460, w_030_461, w_030_463, w_030_464, w_030_465, w_030_466, w_030_468, w_030_469, w_030_470, w_030_471, w_030_472, w_030_473, w_030_474, w_030_475, w_030_476, w_030_477, w_030_479, w_030_480, w_030_481, w_030_482, w_030_483, w_030_484, w_030_485, w_030_486, w_030_487, w_030_488, w_030_489, w_030_490, w_030_491, w_030_492, w_030_493, w_030_494, w_030_496, w_030_497, w_030_498, w_030_499, w_030_500, w_030_501, w_030_502, w_030_503, w_030_504, w_030_505, w_030_506, w_030_507, w_030_508, w_030_509, w_030_510, w_030_511, w_030_512, w_030_513, w_030_514, w_030_515, w_030_516, w_030_517, w_030_518, w_030_519, w_030_520, w_030_521, w_030_522, w_030_523, w_030_524, w_030_525, w_030_526, w_030_527, w_030_528, w_030_529, w_030_530, w_030_531, w_030_532, w_030_533, w_030_534, w_030_535, w_030_536, w_030_538, w_030_539, w_030_540, w_030_541, w_030_542, w_030_543, w_030_544, w_030_545, w_030_546, w_030_547, w_030_548, w_030_549, w_030_550, w_030_551, w_030_552, w_030_553, w_030_554, w_030_555, w_030_556, w_030_557, w_030_558, w_030_559, w_030_560, w_030_561, w_030_562, w_030_563, w_030_564, w_030_565, w_030_566, w_030_567, w_030_568, w_030_570, w_030_571, w_030_572, w_030_573, w_030_574, w_030_575, w_030_576, w_030_577, w_030_578, w_030_579, w_030_580, w_030_581, w_030_582, w_030_583, w_030_584, w_030_585, w_030_586, w_030_587, w_030_588, w_030_589, w_030_590, w_030_591, w_030_592, w_030_593, w_030_594, w_030_595, w_030_596, w_030_597, w_030_598, w_030_599, w_030_600, w_030_601, w_030_603, w_030_604, w_030_605, w_030_606, w_030_607, w_030_608, w_030_609, w_030_610, w_030_611, w_030_612, w_030_613, w_030_614, w_030_615, w_030_616, w_030_617, w_030_618, w_030_619, w_030_620, w_030_621, w_030_622, w_030_623, w_030_624, w_030_625, w_030_626, w_030_627, w_030_628, w_030_629, w_030_631, w_030_632, w_030_633, w_030_634, w_030_635, w_030_636, w_030_637, w_030_638, w_030_639, w_030_640, w_030_641, w_030_642, w_030_643, w_030_644, w_030_645, w_030_646, w_030_647, w_030_648, w_030_649, w_030_650, w_030_651, w_030_652, w_030_655, w_030_656, w_030_657, w_030_658, w_030_659, w_030_660, w_030_661, w_030_662, w_030_663, w_030_664, w_030_665, w_030_666, w_030_667, w_030_668, w_030_669, w_030_670, w_030_672, w_030_674, w_030_675, w_030_676, w_030_677, w_030_678, w_030_679, w_030_680, w_030_681, w_030_682, w_030_683, w_030_684, w_030_685, w_030_686, w_030_687, w_030_688, w_030_689, w_030_690, w_030_691, w_030_692, w_030_693, w_030_694, w_030_695, w_030_696, w_030_697, w_030_698, w_030_699, w_030_700, w_030_701, w_030_702, w_030_703, w_030_704, w_030_705, w_030_706, w_030_707, w_030_708, w_030_710, w_030_711, w_030_712, w_030_713, w_030_714, w_030_715, w_030_716, w_030_717, w_030_718, w_030_719, w_030_720, w_030_721, w_030_722, w_030_723, w_030_724, w_030_725, w_030_726, w_030_727, w_030_728, w_030_729, w_030_730, w_030_731, w_030_732, w_030_733, w_030_734, w_030_735, w_030_736, w_030_738, w_030_739, w_030_740, w_030_741, w_030_742, w_030_743, w_030_744, w_030_745, w_030_746, w_030_747, w_030_748, w_030_749, w_030_750, w_030_752, w_030_753, w_030_754, w_030_755, w_030_756, w_030_757, w_030_758, w_030_759, w_030_760, w_030_761, w_030_762, w_030_763, w_030_764, w_030_765, w_030_766, w_030_767, w_030_768, w_030_769, w_030_770, w_030_771, w_030_772, w_030_773, w_030_774, w_030_775, w_030_776, w_030_777, w_030_778, w_030_779, w_030_780, w_030_781, w_030_782, w_030_783, w_030_784, w_030_785, w_030_786, w_030_787, w_030_788, w_030_790, w_030_791, w_030_792, w_030_793, w_030_794, w_030_795, w_030_796, w_030_797, w_030_798, w_030_799, w_030_800, w_030_801, w_030_802, w_030_803, w_030_804, w_030_805, w_030_806, w_030_807, w_030_808, w_030_809, w_030_810, w_030_811, w_030_812, w_030_813, w_030_815, w_030_816, w_030_817, w_030_818, w_030_819, w_030_820, w_030_821, w_030_822, w_030_823, w_030_824, w_030_825, w_030_826, w_030_827, w_030_828, w_030_829, w_030_830, w_030_831, w_030_832, w_030_833, w_030_834, w_030_835, w_030_836, w_030_837, w_030_838, w_030_839, w_030_840, w_030_841, w_030_842, w_030_843, w_030_844, w_030_845, w_030_846, w_030_847, w_030_849, w_030_850, w_030_851, w_030_852, w_030_853, w_030_854, w_030_855, w_030_856, w_030_858, w_030_859, w_030_860, w_030_861, w_030_862, w_030_863, w_030_864, w_030_865, w_030_866, w_030_867, w_030_868, w_030_869, w_030_870, w_030_871, w_030_872, w_030_873, w_030_874, w_030_875, w_030_876, w_030_877, w_030_878, w_030_879, w_030_880, w_030_881, w_030_882, w_030_883, w_030_884, w_030_885, w_030_886, w_030_887, w_030_888, w_030_889, w_030_890, w_030_891, w_030_894, w_030_895, w_030_896, w_030_897, w_030_898, w_030_899, w_030_900, w_030_901, w_030_902, w_030_903, w_030_904, w_030_905, w_030_906, w_030_907, w_030_908, w_030_909, w_030_910, w_030_911, w_030_912, w_030_913, w_030_914, w_030_915, w_030_916, w_030_918, w_030_919, w_030_920, w_030_921, w_030_922, w_030_923, w_030_924, w_030_925, w_030_927, w_030_928, w_030_929, w_030_930, w_030_931, w_030_932, w_030_933, w_030_934, w_030_935, w_030_936, w_030_937, w_030_938, w_030_939, w_030_940, w_030_941, w_030_942, w_030_943, w_030_944, w_030_945, w_030_946, w_030_947, w_030_948, w_030_949, w_030_950, w_030_951, w_030_952, w_030_953, w_030_954, w_030_955, w_030_956, w_030_957, w_030_958, w_030_959, w_030_960, w_030_961, w_030_962, w_030_963, w_030_964, w_030_965, w_030_966, w_030_967, w_030_968, w_030_969, w_030_970, w_030_971, w_030_972, w_030_973, w_030_974, w_030_975, w_030_976, w_030_977, w_030_978, w_030_979, w_030_980, w_030_981, w_030_982, w_030_983, w_030_985, w_030_986, w_030_987, w_030_988, w_030_989, w_030_990, w_030_991, w_030_992, w_030_993, w_030_994, w_030_995, w_030_996, w_030_997, w_030_998, w_030_999, w_030_1000, w_030_1001, w_030_1002, w_030_1003, w_030_1005, w_030_1006, w_030_1007, w_030_1008, w_030_1009, w_030_1010, w_030_1011, w_030_1012, w_030_1013, w_030_1014, w_030_1015, w_030_1016, w_030_1017, w_030_1018, w_030_1019, w_030_1020, w_030_1021, w_030_1022, w_030_1023, w_030_1025, w_030_1026, w_030_1027, w_030_1028, w_030_1030, w_030_1032, w_030_1033, w_030_1034, w_030_1035, w_030_1036, w_030_1037, w_030_1038, w_030_1039, w_030_1040, w_030_1041, w_030_1042, w_030_1043, w_030_1044, w_030_1045, w_030_1046, w_030_1047, w_030_1048, w_030_1049, w_030_1050, w_030_1052, w_030_1054, w_030_1055, w_030_1056, w_030_1057, w_030_1059, w_030_1060, w_030_1061, w_030_1062, w_030_1063, w_030_1064, w_030_1065, w_030_1066, w_030_1067, w_030_1068, w_030_1069, w_030_1070, w_030_1071, w_030_1072, w_030_1073, w_030_1074, w_030_1075, w_030_1076, w_030_1077, w_030_1078, w_030_1079, w_030_1080, w_030_1081, w_030_1082, w_030_1083, w_030_1084, w_030_1085, w_030_1086, w_030_1087, w_030_1088, w_030_1089, w_030_1090, w_030_1091, w_030_1092, w_030_1093, w_030_1094, w_030_1095, w_030_1096, w_030_1097, w_030_1098, w_030_1099, w_030_1100, w_030_1101, w_030_1102, w_030_1103, w_030_1105, w_030_1106, w_030_1107, w_030_1108, w_030_1109, w_030_1110, w_030_1111, w_030_1112, w_030_1113, w_030_1114, w_030_1115, w_030_1116, w_030_1117, w_030_1118, w_030_1119, w_030_1120, w_030_1121, w_030_1122, w_030_1123, w_030_1124, w_030_1125, w_030_1126, w_030_1127, w_030_1128, w_030_1129, w_030_1130, w_030_1131, w_030_1132, w_030_1133, w_030_1134, w_030_1135, w_030_1136, w_030_1137, w_030_1138, w_030_1139, w_030_1141, w_030_1142, w_030_1143, w_030_1144, w_030_1145, w_030_1146, w_030_1147, w_030_1148, w_030_1149, w_030_1150, w_030_1151, w_030_1152, w_030_1153, w_030_1154, w_030_1155, w_030_1156, w_030_1157, w_030_1158, w_030_1159, w_030_1160, w_030_1161, w_030_1162, w_030_1163, w_030_1164, w_030_1165, w_030_1166, w_030_1167, w_030_1169, w_030_1170, w_030_1173, w_030_1174, w_030_1175, w_030_1176, w_030_1177, w_030_1178, w_030_1179, w_030_1180, w_030_1182, w_030_1183, w_030_1184, w_030_1185, w_030_1186, w_030_1187, w_030_1188, w_030_1189, w_030_1190, w_030_1191, w_030_1192, w_030_1193, w_030_1195, w_030_1196, w_030_1197, w_030_1198, w_030_1199, w_030_1200, w_030_1201, w_030_1202, w_030_1203, w_030_1204, w_030_1205, w_030_1208, w_030_1209, w_030_1210, w_030_1211, w_030_1212, w_030_1213, w_030_1214, w_030_1215, w_030_1216, w_030_1217, w_030_1218, w_030_1219, w_030_1220, w_030_1221, w_030_1222, w_030_1223, w_030_1225, w_030_1226, w_030_1227, w_030_1228, w_030_1229, w_030_1230, w_030_1231, w_030_1232, w_030_1233, w_030_1234, w_030_1236, w_030_1237, w_030_1238, w_030_1239, w_030_1240, w_030_1241, w_030_1242, w_030_1243, w_030_1244, w_030_1245, w_030_1246, w_030_1247, w_030_1248, w_030_1249, w_030_1250, w_030_1251, w_030_1252, w_030_1253, w_030_1254, w_030_1255, w_030_1256, w_030_1257, w_030_1258, w_030_1259, w_030_1260, w_030_1261, w_030_1262, w_030_1264, w_030_1265, w_030_1266, w_030_1267, w_030_1268, w_030_1269, w_030_1270, w_030_1271, w_030_1272, w_030_1273, w_030_1274, w_030_1275, w_030_1276, w_030_1277, w_030_1278, w_030_1279, w_030_1280, w_030_1281, w_030_1283, w_030_1284, w_030_1285, w_030_1286, w_030_1287, w_030_1288, w_030_1289, w_030_1290, w_030_1291, w_030_1292, w_030_1293, w_030_1294, w_030_1295, w_030_1296, w_030_1297, w_030_1298, w_030_1299, w_030_1300, w_030_1301, w_030_1302, w_030_1303, w_030_1304, w_030_1305, w_030_1306, w_030_1307, w_030_1308, w_030_1309, w_030_1310, w_030_1311, w_030_1312, w_030_1313, w_030_1314, w_030_1315, w_030_1316, w_030_1317, w_030_1318, w_030_1319, w_030_1320, w_030_1321, w_030_1322, w_030_1323, w_030_1324, w_030_1325, w_030_1326, w_030_1327, w_030_1328, w_030_1329, w_030_1330, w_030_1331, w_030_1332, w_030_1333, w_030_1334, w_030_1335, w_030_1336, w_030_1337, w_030_1338, w_030_1339, w_030_1340, w_030_1341, w_030_1342, w_030_1343, w_030_1344, w_030_1345, w_030_1346, w_030_1347, w_030_1349, w_030_1350, w_030_1351, w_030_1352, w_030_1354, w_030_1355, w_030_1356, w_030_1357, w_030_1358, w_030_1359, w_030_1360, w_030_1361, w_030_1362, w_030_1363, w_030_1364, w_030_1365, w_030_1366, w_030_1367, w_030_1368, w_030_1369, w_030_1370, w_030_1371, w_030_1372, w_030_1373, w_030_1374, w_030_1375, w_030_1376, w_030_1377, w_030_1378, w_030_1379, w_030_1380, w_030_1381, w_030_1382, w_030_1383, w_030_1384, w_030_1385, w_030_1386, w_030_1387, w_030_1388, w_030_1389, w_030_1390, w_030_1391, w_030_1393, w_030_1394, w_030_1395, w_030_1396, w_030_1397, w_030_1398, w_030_1399, w_030_1400, w_030_1401, w_030_1402, w_030_1404, w_030_1406, w_030_1407, w_030_1408, w_030_1409, w_030_1410, w_030_1411, w_030_1412, w_030_1414, w_030_1416, w_030_1417, w_030_1418, w_030_1419, w_030_1420, w_030_1421, w_030_1423, w_030_1424, w_030_1425, w_030_1426, w_030_1427, w_030_1428, w_030_1429, w_030_1430, w_030_1431, w_030_1432, w_030_1433, w_030_1434, w_030_1435, w_030_1436, w_030_1437, w_030_1438, w_030_1439, w_030_1440, w_030_1441, w_030_1442, w_030_1443, w_030_1445, w_030_1446, w_030_1448, w_030_1449, w_030_1450, w_030_1451, w_030_1452, w_030_1453, w_030_1454, w_030_1455, w_030_1456, w_030_1457, w_030_1458, w_030_1460, w_030_1461, w_030_1462, w_030_1463, w_030_1464, w_030_1465, w_030_1466, w_030_1467, w_030_1468, w_030_1469, w_030_1470, w_030_1471, w_030_1472, w_030_1473, w_030_1474, w_030_1475, w_030_1476, w_030_1477, w_030_1478, w_030_1479, w_030_1481, w_030_1482, w_030_1484, w_030_1485, w_030_1486, w_030_1487, w_030_1488, w_030_1489, w_030_1490, w_030_1491, w_030_1492, w_030_1493, w_030_1494, w_030_1495, w_030_1496, w_030_1497, w_030_1498, w_030_1499, w_030_1500, w_030_1501, w_030_1502, w_030_1503, w_030_1504, w_030_1505, w_030_1506, w_030_1507, w_030_1508, w_030_1509, w_030_1510, w_030_1511, w_030_1512, w_030_1513, w_030_1514, w_030_1515, w_030_1516, w_030_1517, w_030_1518, w_030_1519, w_030_1520, w_030_1522, w_030_1523, w_030_1524, w_030_1525, w_030_1526, w_030_1527, w_030_1528, w_030_1529, w_030_1530, w_030_1531, w_030_1532, w_030_1533, w_030_1534, w_030_1535, w_030_1536, w_030_1537, w_030_1538, w_030_1540, w_030_1541, w_030_1542, w_030_1543, w_030_1544, w_030_1545, w_030_1547, w_030_1548, w_030_1549, w_030_1550, w_030_1554, w_030_1555, w_030_1556, w_030_1557, w_030_1558, w_030_1559, w_030_1560, w_030_1561, w_030_1562, w_030_1563, w_030_1565, w_030_1566, w_030_1567, w_030_1568, w_030_1570, w_030_1571, w_030_1573, w_030_1574, w_030_1575, w_030_1577, w_030_1578, w_030_1579, w_030_1580, w_030_1581, w_030_1582, w_030_1583, w_030_1584, w_030_1585, w_030_1586, w_030_1587, w_030_1590, w_030_1591, w_030_1592, w_030_1593, w_030_1594, w_030_1595, w_030_1596, w_030_1597, w_030_1598, w_030_1599, w_030_1600, w_030_1601, w_030_1602, w_030_1603, w_030_1604, w_030_1605, w_030_1606, w_030_1607, w_030_1608, w_030_1610, w_030_1611, w_030_1612, w_030_1613, w_030_1614, w_030_1615, w_030_1616, w_030_1617, w_030_1618, w_030_1619, w_030_1620, w_030_1621, w_030_1622, w_030_1623, w_030_1624, w_030_1626, w_030_1627, w_030_1628, w_030_1629, w_030_1630, w_030_1631, w_030_1632, w_030_1633, w_030_1634, w_030_1635, w_030_1636, w_030_1637, w_030_1638, w_030_1640, w_030_1641, w_030_1642, w_030_1643, w_030_1644, w_030_1645, w_030_1646, w_030_1648, w_030_1649, w_030_1650, w_030_1652, w_030_1653, w_030_1654, w_030_1655, w_030_1658, w_030_1659, w_030_1660, w_030_1661, w_030_1662, w_030_1665, w_030_1667, w_030_1668, w_030_1669, w_030_1670, w_030_1671, w_030_1672, w_030_1673, w_030_1676, w_030_1677, w_030_1678, w_030_1679, w_030_1680, w_030_1682, w_030_1683, w_030_1684, w_030_1686, w_030_1687, w_030_1688, w_030_1689, w_030_1691, w_030_1693, w_030_1694, w_030_1695, w_030_1697, w_030_1698, w_030_1699, w_030_1700, w_030_1701, w_030_1702, w_030_1703, w_030_1704, w_030_1705, w_030_1707, w_030_1708, w_030_1709, w_030_1711, w_030_1712, w_030_1713, w_030_1714, w_030_1715, w_030_1716, w_030_1717, w_030_1718, w_030_1719, w_030_1720, w_030_1722, w_030_1724, w_030_1725, w_030_1726, w_030_1727;
  wire w_031_000, w_031_001, w_031_002, w_031_003, w_031_004, w_031_005, w_031_006, w_031_007, w_031_008, w_031_009, w_031_010, w_031_011, w_031_012, w_031_013, w_031_014, w_031_015, w_031_016, w_031_017, w_031_018, w_031_019, w_031_020, w_031_021, w_031_022, w_031_023, w_031_024, w_031_025, w_031_026, w_031_027, w_031_028, w_031_029, w_031_030, w_031_031, w_031_032, w_031_033, w_031_034, w_031_035, w_031_036, w_031_037, w_031_038, w_031_039, w_031_040, w_031_041, w_031_042, w_031_043, w_031_044, w_031_045, w_031_046, w_031_047, w_031_048, w_031_049, w_031_050, w_031_051, w_031_052, w_031_053, w_031_054, w_031_055, w_031_056, w_031_057, w_031_058, w_031_059, w_031_060, w_031_061, w_031_062, w_031_063, w_031_064, w_031_065, w_031_066, w_031_067, w_031_068, w_031_069, w_031_070, w_031_071, w_031_072, w_031_073, w_031_074, w_031_075, w_031_076, w_031_077, w_031_078, w_031_079, w_031_080, w_031_081, w_031_082, w_031_083, w_031_084, w_031_085, w_031_086, w_031_087, w_031_088, w_031_089, w_031_090, w_031_091, w_031_092, w_031_093, w_031_094, w_031_095, w_031_096, w_031_097, w_031_098, w_031_099, w_031_100, w_031_101, w_031_102, w_031_103, w_031_104, w_031_105, w_031_106, w_031_107, w_031_108, w_031_109, w_031_110, w_031_111, w_031_112, w_031_113, w_031_114, w_031_115, w_031_116, w_031_117, w_031_118, w_031_119, w_031_120, w_031_121, w_031_123, w_031_124, w_031_125, w_031_126, w_031_127, w_031_128, w_031_129, w_031_130, w_031_132, w_031_133, w_031_134, w_031_135, w_031_136, w_031_137, w_031_138, w_031_139, w_031_140, w_031_141, w_031_142, w_031_143, w_031_144, w_031_145, w_031_146, w_031_147, w_031_148, w_031_149, w_031_150, w_031_151, w_031_152, w_031_153, w_031_154, w_031_155, w_031_156, w_031_157, w_031_158, w_031_159, w_031_160, w_031_161, w_031_162, w_031_163, w_031_164, w_031_165, w_031_166, w_031_167, w_031_168, w_031_169, w_031_170, w_031_171, w_031_172, w_031_173, w_031_174, w_031_175, w_031_176, w_031_177, w_031_178, w_031_179, w_031_180, w_031_181, w_031_182, w_031_183, w_031_184, w_031_185, w_031_186, w_031_187, w_031_188, w_031_189, w_031_190, w_031_191, w_031_192, w_031_193, w_031_194, w_031_195, w_031_196, w_031_197, w_031_198, w_031_199, w_031_200, w_031_201, w_031_202, w_031_203, w_031_204, w_031_205, w_031_206, w_031_207, w_031_208, w_031_209, w_031_210, w_031_211, w_031_212, w_031_213, w_031_214, w_031_215, w_031_216, w_031_217, w_031_218, w_031_219, w_031_220, w_031_221, w_031_222, w_031_223, w_031_224, w_031_225, w_031_226, w_031_227, w_031_228, w_031_229, w_031_230, w_031_231, w_031_232, w_031_233, w_031_234, w_031_235, w_031_236, w_031_237, w_031_238, w_031_239, w_031_240, w_031_241, w_031_242, w_031_243, w_031_244, w_031_245, w_031_246, w_031_247, w_031_248, w_031_249, w_031_250, w_031_251, w_031_252, w_031_253, w_031_254, w_031_255, w_031_256, w_031_257, w_031_258, w_031_259, w_031_260, w_031_261, w_031_262, w_031_263, w_031_264, w_031_265, w_031_266, w_031_267, w_031_268, w_031_269, w_031_270, w_031_271, w_031_272, w_031_273, w_031_274, w_031_275, w_031_276, w_031_277, w_031_278, w_031_279, w_031_280, w_031_281, w_031_282, w_031_283, w_031_284, w_031_285, w_031_286, w_031_287, w_031_288, w_031_289, w_031_290, w_031_291, w_031_292, w_031_293, w_031_294, w_031_295, w_031_296, w_031_297, w_031_298, w_031_299, w_031_300, w_031_301, w_031_302, w_031_303, w_031_304, w_031_305, w_031_306, w_031_307, w_031_308, w_031_309, w_031_310, w_031_311, w_031_312, w_031_313, w_031_314, w_031_315, w_031_316, w_031_317, w_031_318, w_031_319, w_031_320, w_031_321, w_031_322, w_031_323, w_031_324, w_031_325, w_031_326, w_031_327, w_031_328, w_031_329, w_031_330, w_031_331, w_031_332, w_031_333, w_031_334, w_031_335, w_031_336, w_031_337, w_031_338, w_031_339, w_031_340, w_031_341, w_031_342, w_031_343, w_031_344, w_031_345, w_031_346, w_031_347, w_031_348, w_031_349, w_031_350, w_031_351, w_031_352, w_031_353, w_031_354, w_031_355, w_031_356, w_031_357, w_031_358, w_031_359, w_031_360, w_031_361, w_031_362, w_031_363, w_031_364, w_031_365, w_031_366, w_031_367, w_031_368, w_031_369, w_031_370, w_031_371, w_031_372, w_031_373, w_031_374, w_031_375, w_031_376, w_031_377, w_031_378, w_031_379, w_031_380, w_031_381, w_031_382, w_031_383, w_031_384, w_031_385, w_031_386, w_031_387, w_031_388, w_031_389, w_031_390, w_031_391, w_031_392, w_031_393, w_031_394, w_031_395, w_031_396, w_031_397, w_031_398, w_031_399, w_031_400, w_031_401, w_031_402, w_031_403, w_031_404, w_031_405, w_031_407, w_031_408, w_031_409, w_031_410, w_031_411, w_031_412, w_031_413, w_031_414, w_031_415, w_031_416, w_031_417, w_031_418, w_031_419, w_031_420, w_031_421, w_031_422, w_031_423, w_031_424, w_031_425, w_031_426, w_031_427, w_031_429, w_031_430, w_031_431, w_031_432, w_031_433, w_031_434, w_031_435, w_031_436, w_031_437, w_031_438, w_031_439, w_031_440, w_031_441, w_031_442, w_031_443, w_031_444, w_031_445, w_031_446, w_031_447, w_031_448, w_031_449, w_031_450, w_031_451, w_031_452, w_031_454, w_031_455, w_031_456, w_031_457, w_031_458, w_031_459, w_031_460, w_031_461, w_031_462, w_031_463, w_031_464, w_031_465, w_031_466, w_031_467, w_031_468, w_031_469, w_031_470, w_031_471, w_031_472, w_031_473, w_031_474, w_031_475, w_031_476, w_031_477, w_031_478, w_031_479, w_031_480, w_031_481, w_031_482, w_031_483, w_031_484, w_031_485, w_031_486, w_031_487, w_031_488, w_031_490, w_031_491, w_031_492, w_031_493, w_031_494, w_031_495, w_031_496, w_031_497, w_031_498, w_031_499, w_031_500, w_031_501, w_031_502, w_031_503, w_031_504, w_031_505, w_031_506, w_031_507, w_031_508, w_031_509, w_031_510, w_031_511, w_031_512, w_031_513, w_031_514, w_031_515, w_031_516, w_031_517, w_031_518, w_031_519, w_031_520, w_031_521, w_031_522, w_031_523, w_031_524, w_031_525, w_031_526, w_031_527, w_031_528, w_031_529, w_031_530, w_031_531, w_031_532, w_031_533, w_031_534, w_031_535, w_031_536, w_031_537, w_031_538, w_031_539, w_031_540, w_031_541, w_031_542, w_031_543, w_031_544, w_031_545, w_031_546, w_031_547, w_031_548, w_031_549, w_031_550, w_031_551, w_031_552, w_031_553, w_031_554, w_031_555, w_031_556, w_031_557, w_031_558, w_031_559, w_031_560, w_031_561, w_031_562, w_031_563, w_031_564, w_031_565, w_031_566, w_031_567, w_031_568, w_031_569, w_031_570, w_031_571, w_031_572, w_031_573, w_031_574, w_031_575, w_031_576, w_031_577, w_031_578, w_031_579, w_031_580, w_031_581, w_031_582, w_031_583, w_031_584, w_031_585, w_031_587, w_031_588, w_031_589, w_031_590, w_031_591, w_031_592, w_031_593, w_031_594, w_031_595, w_031_596, w_031_597, w_031_598, w_031_599, w_031_600, w_031_601, w_031_602, w_031_603, w_031_604, w_031_605, w_031_606, w_031_607, w_031_608, w_031_609, w_031_610, w_031_611, w_031_612, w_031_613, w_031_614, w_031_615, w_031_616, w_031_617, w_031_618, w_031_619, w_031_620, w_031_621, w_031_622, w_031_623, w_031_624, w_031_625, w_031_626, w_031_627, w_031_628, w_031_629, w_031_630, w_031_631, w_031_632, w_031_633, w_031_634, w_031_635, w_031_636, w_031_637, w_031_638, w_031_639, w_031_640, w_031_641, w_031_642, w_031_643, w_031_644, w_031_645, w_031_646, w_031_647, w_031_648, w_031_649, w_031_650, w_031_651, w_031_652, w_031_653, w_031_654, w_031_655, w_031_656, w_031_657, w_031_658, w_031_659, w_031_660, w_031_661, w_031_662, w_031_663, w_031_664, w_031_665, w_031_666, w_031_667, w_031_668, w_031_670, w_031_671, w_031_672, w_031_673, w_031_674, w_031_675, w_031_676, w_031_677, w_031_678, w_031_679, w_031_680, w_031_681, w_031_682, w_031_683, w_031_685, w_031_686, w_031_688, w_031_689, w_031_690, w_031_691, w_031_692, w_031_693, w_031_694, w_031_695, w_031_696, w_031_697, w_031_698, w_031_699, w_031_700, w_031_701, w_031_702, w_031_703, w_031_704, w_031_705, w_031_706, w_031_707, w_031_709, w_031_710, w_031_711, w_031_712, w_031_713, w_031_714, w_031_715, w_031_716, w_031_717, w_031_718, w_031_719, w_031_720, w_031_721, w_031_722, w_031_723, w_031_724, w_031_725, w_031_726, w_031_727, w_031_728, w_031_729, w_031_730, w_031_731, w_031_732, w_031_733, w_031_734, w_031_735, w_031_736, w_031_737, w_031_738, w_031_739, w_031_740, w_031_741, w_031_742, w_031_743, w_031_744, w_031_745, w_031_746, w_031_747, w_031_748, w_031_749, w_031_750, w_031_751, w_031_752, w_031_753, w_031_754, w_031_755, w_031_756, w_031_757, w_031_758, w_031_759, w_031_760, w_031_761, w_031_762, w_031_763, w_031_764, w_031_765, w_031_766, w_031_767, w_031_768, w_031_769, w_031_770, w_031_771, w_031_772, w_031_773, w_031_774, w_031_775, w_031_776, w_031_777, w_031_778, w_031_779, w_031_780, w_031_781, w_031_782, w_031_783, w_031_784, w_031_785, w_031_786, w_031_787, w_031_788, w_031_789, w_031_790, w_031_791, w_031_792, w_031_793, w_031_794, w_031_795, w_031_796, w_031_797, w_031_798, w_031_799, w_031_800, w_031_801, w_031_802, w_031_803, w_031_804, w_031_805, w_031_807, w_031_808, w_031_809, w_031_810, w_031_811, w_031_812, w_031_813, w_031_814, w_031_815, w_031_816, w_031_817, w_031_818, w_031_819, w_031_820, w_031_821, w_031_822, w_031_823, w_031_824, w_031_825, w_031_826, w_031_827, w_031_828, w_031_829, w_031_830, w_031_831, w_031_832, w_031_833, w_031_834, w_031_835, w_031_836, w_031_837, w_031_838, w_031_839, w_031_840, w_031_841, w_031_842, w_031_843, w_031_844, w_031_845, w_031_846, w_031_847, w_031_848, w_031_849, w_031_850, w_031_851, w_031_852, w_031_853, w_031_854, w_031_855, w_031_856, w_031_857, w_031_858, w_031_859, w_031_860, w_031_861, w_031_862, w_031_863, w_031_864, w_031_865, w_031_866, w_031_867, w_031_868, w_031_869, w_031_870, w_031_871, w_031_872, w_031_873, w_031_874, w_031_875, w_031_877, w_031_878, w_031_879, w_031_880, w_031_881, w_031_882, w_031_883, w_031_884, w_031_885, w_031_886, w_031_887, w_031_888, w_031_889, w_031_890, w_031_891, w_031_892, w_031_893, w_031_895, w_031_896, w_031_897, w_031_898, w_031_899, w_031_900, w_031_901, w_031_902, w_031_903, w_031_904, w_031_905, w_031_906, w_031_907, w_031_908, w_031_909, w_031_912, w_031_913, w_031_914, w_031_915, w_031_916, w_031_917, w_031_918, w_031_919, w_031_920, w_031_921, w_031_922, w_031_923, w_031_924, w_031_925, w_031_926, w_031_927, w_031_928, w_031_929, w_031_930, w_031_931, w_031_932, w_031_933, w_031_934, w_031_935, w_031_936, w_031_937, w_031_938, w_031_939, w_031_940, w_031_941, w_031_942, w_031_943, w_031_944, w_031_945, w_031_946, w_031_947, w_031_948, w_031_949, w_031_950, w_031_951, w_031_952, w_031_953, w_031_954, w_031_955, w_031_956, w_031_957, w_031_958, w_031_959, w_031_960, w_031_961, w_031_962, w_031_963, w_031_964, w_031_965, w_031_966, w_031_967, w_031_968, w_031_969, w_031_970, w_031_971, w_031_972, w_031_973, w_031_974, w_031_975, w_031_976, w_031_977, w_031_978, w_031_980, w_031_981, w_031_982, w_031_983, w_031_984, w_031_985, w_031_986, w_031_987, w_031_988, w_031_989, w_031_990, w_031_991, w_031_992, w_031_993, w_031_994, w_031_995, w_031_996, w_031_997, w_031_998, w_031_999, w_031_1000, w_031_1001, w_031_1002, w_031_1003, w_031_1004, w_031_1005, w_031_1006, w_031_1007, w_031_1008, w_031_1009, w_031_1010, w_031_1011, w_031_1012, w_031_1013, w_031_1014, w_031_1015, w_031_1016, w_031_1017, w_031_1018, w_031_1019, w_031_1021, w_031_1022, w_031_1023, w_031_1024, w_031_1025, w_031_1026, w_031_1027, w_031_1028, w_031_1029, w_031_1031, w_031_1032, w_031_1033, w_031_1034, w_031_1035, w_031_1036, w_031_1037, w_031_1038, w_031_1039, w_031_1040, w_031_1041, w_031_1042, w_031_1043, w_031_1044, w_031_1045, w_031_1046, w_031_1047, w_031_1048, w_031_1049, w_031_1050, w_031_1051, w_031_1052, w_031_1053, w_031_1054, w_031_1055, w_031_1056, w_031_1057, w_031_1058, w_031_1059, w_031_1060, w_031_1061, w_031_1062, w_031_1063, w_031_1064, w_031_1065, w_031_1066, w_031_1067, w_031_1068, w_031_1069, w_031_1070, w_031_1071, w_031_1072, w_031_1073, w_031_1074, w_031_1075, w_031_1076, w_031_1077, w_031_1078, w_031_1079, w_031_1080, w_031_1081, w_031_1082, w_031_1083, w_031_1084, w_031_1085, w_031_1086, w_031_1087, w_031_1088, w_031_1089, w_031_1090, w_031_1091, w_031_1092, w_031_1093, w_031_1094, w_031_1095, w_031_1096, w_031_1097, w_031_1098, w_031_1099, w_031_1100, w_031_1101, w_031_1102, w_031_1103, w_031_1104, w_031_1105, w_031_1106, w_031_1107, w_031_1108, w_031_1109, w_031_1110, w_031_1111, w_031_1112, w_031_1113, w_031_1115, w_031_1116, w_031_1117, w_031_1118, w_031_1119, w_031_1120, w_031_1121, w_031_1122, w_031_1123, w_031_1124, w_031_1125, w_031_1126, w_031_1127, w_031_1128, w_031_1129, w_031_1130, w_031_1131, w_031_1132, w_031_1133, w_031_1134, w_031_1135, w_031_1136, w_031_1137, w_031_1138, w_031_1139, w_031_1140, w_031_1142, w_031_1144, w_031_1145, w_031_1146, w_031_1147, w_031_1148, w_031_1149, w_031_1150, w_031_1151, w_031_1152, w_031_1153, w_031_1154, w_031_1155, w_031_1156, w_031_1157, w_031_1158, w_031_1159, w_031_1160, w_031_1161, w_031_1162, w_031_1163, w_031_1164, w_031_1165, w_031_1166, w_031_1167, w_031_1168, w_031_1169, w_031_1170, w_031_1171, w_031_1172;
  wire w_032_000, w_032_001, w_032_002, w_032_003, w_032_004, w_032_005, w_032_006, w_032_007, w_032_008, w_032_009, w_032_010, w_032_011, w_032_012, w_032_013, w_032_014, w_032_015, w_032_016, w_032_017, w_032_018, w_032_019, w_032_020, w_032_021, w_032_022, w_032_023, w_032_024, w_032_025, w_032_026, w_032_027, w_032_028, w_032_029, w_032_030, w_032_031, w_032_032, w_032_033, w_032_034, w_032_035, w_032_036, w_032_037, w_032_038, w_032_039, w_032_040, w_032_041, w_032_042, w_032_043, w_032_044, w_032_045, w_032_046, w_032_047, w_032_048, w_032_049, w_032_050, w_032_051, w_032_052, w_032_053, w_032_054, w_032_055, w_032_056, w_032_057, w_032_058, w_032_059, w_032_060, w_032_062, w_032_063, w_032_064, w_032_065, w_032_066, w_032_067, w_032_068, w_032_069, w_032_070, w_032_071, w_032_072, w_032_073, w_032_074, w_032_075, w_032_076, w_032_077, w_032_078, w_032_079, w_032_080, w_032_081, w_032_082, w_032_083, w_032_084, w_032_085, w_032_086, w_032_087, w_032_088, w_032_089, w_032_090, w_032_091, w_032_092, w_032_093, w_032_094, w_032_095, w_032_096, w_032_097, w_032_098, w_032_099, w_032_100, w_032_101, w_032_102, w_032_103, w_032_104, w_032_105, w_032_106, w_032_107, w_032_108, w_032_109, w_032_110, w_032_111, w_032_112, w_032_113, w_032_114, w_032_115, w_032_116, w_032_117, w_032_118, w_032_119, w_032_120, w_032_121, w_032_122, w_032_123, w_032_124, w_032_125, w_032_126, w_032_127, w_032_128, w_032_129, w_032_130, w_032_131, w_032_132, w_032_133, w_032_134, w_032_135, w_032_136, w_032_137, w_032_138, w_032_139, w_032_141, w_032_142, w_032_143, w_032_144, w_032_145, w_032_146, w_032_147, w_032_148, w_032_149, w_032_150, w_032_151, w_032_152, w_032_153, w_032_154, w_032_155, w_032_156, w_032_157, w_032_158, w_032_159, w_032_160, w_032_161, w_032_162, w_032_163, w_032_164, w_032_165, w_032_166, w_032_167, w_032_168, w_032_169, w_032_170, w_032_171, w_032_172, w_032_173, w_032_174, w_032_175, w_032_176, w_032_177, w_032_178, w_032_179, w_032_180, w_032_181, w_032_182, w_032_183, w_032_184, w_032_185, w_032_186, w_032_187, w_032_188, w_032_189, w_032_190, w_032_191, w_032_192, w_032_193, w_032_194, w_032_195, w_032_196, w_032_197, w_032_198, w_032_199, w_032_200, w_032_201, w_032_202, w_032_203, w_032_204, w_032_205, w_032_206, w_032_207, w_032_208, w_032_209, w_032_210, w_032_211, w_032_212, w_032_213, w_032_214, w_032_215, w_032_216, w_032_217, w_032_218, w_032_219, w_032_221, w_032_222, w_032_223, w_032_224, w_032_225, w_032_226, w_032_227, w_032_228, w_032_229, w_032_230, w_032_231, w_032_232, w_032_233, w_032_234, w_032_235, w_032_236, w_032_237, w_032_238, w_032_239, w_032_240, w_032_241, w_032_242, w_032_243, w_032_244, w_032_245, w_032_246, w_032_247, w_032_248, w_032_249, w_032_250, w_032_251, w_032_252, w_032_253, w_032_254, w_032_255, w_032_256, w_032_257, w_032_258, w_032_259, w_032_260, w_032_261, w_032_262, w_032_263, w_032_264, w_032_265, w_032_266, w_032_267, w_032_268, w_032_269, w_032_270, w_032_271, w_032_272, w_032_273, w_032_274, w_032_275, w_032_276, w_032_277, w_032_278, w_032_279, w_032_280, w_032_281, w_032_282, w_032_283, w_032_284, w_032_285, w_032_286, w_032_287, w_032_288, w_032_289, w_032_290, w_032_291, w_032_292, w_032_293, w_032_294, w_032_295, w_032_296, w_032_297, w_032_298, w_032_299, w_032_300, w_032_301, w_032_302, w_032_303, w_032_304, w_032_305, w_032_306, w_032_307, w_032_308, w_032_309, w_032_310, w_032_312, w_032_313, w_032_314, w_032_315, w_032_316, w_032_317, w_032_318, w_032_319, w_032_320, w_032_321, w_032_322, w_032_323, w_032_324, w_032_325, w_032_326, w_032_327, w_032_328, w_032_329, w_032_330, w_032_331, w_032_332, w_032_333, w_032_334, w_032_335, w_032_336, w_032_337, w_032_338, w_032_339, w_032_340, w_032_341, w_032_342, w_032_343, w_032_344, w_032_345, w_032_346, w_032_347, w_032_348, w_032_349, w_032_350, w_032_351, w_032_352, w_032_353, w_032_354, w_032_355, w_032_356, w_032_357, w_032_358, w_032_359, w_032_360, w_032_361, w_032_362, w_032_363, w_032_364, w_032_365, w_032_366, w_032_367, w_032_368, w_032_369, w_032_370, w_032_371, w_032_372, w_032_373, w_032_374, w_032_375, w_032_376, w_032_377, w_032_378, w_032_379, w_032_380, w_032_381, w_032_382, w_032_383, w_032_384, w_032_385, w_032_386, w_032_387, w_032_388, w_032_389, w_032_390, w_032_391, w_032_392, w_032_393, w_032_394, w_032_395, w_032_396, w_032_397, w_032_398, w_032_399, w_032_400, w_032_401, w_032_402, w_032_403, w_032_404, w_032_405, w_032_406, w_032_407, w_032_408, w_032_409, w_032_410, w_032_411, w_032_412, w_032_413, w_032_414, w_032_415, w_032_416, w_032_417, w_032_419, w_032_420, w_032_421, w_032_422, w_032_423, w_032_424, w_032_425, w_032_426, w_032_427, w_032_428, w_032_429, w_032_430, w_032_431, w_032_432, w_032_433, w_032_434, w_032_435, w_032_436, w_032_437, w_032_438, w_032_439, w_032_440, w_032_441, w_032_442, w_032_443, w_032_444, w_032_445, w_032_446, w_032_447, w_032_448, w_032_449, w_032_450, w_032_451, w_032_452, w_032_453, w_032_454, w_032_455, w_032_456, w_032_457, w_032_458, w_032_459, w_032_460, w_032_461, w_032_462, w_032_463, w_032_464, w_032_465, w_032_466, w_032_467, w_032_468, w_032_469, w_032_471, w_032_472, w_032_473, w_032_474, w_032_475, w_032_476, w_032_477, w_032_478, w_032_479, w_032_480, w_032_481, w_032_482, w_032_483, w_032_484, w_032_485, w_032_486, w_032_487, w_032_488, w_032_489, w_032_490, w_032_491, w_032_492, w_032_493, w_032_494, w_032_495, w_032_496, w_032_497, w_032_498, w_032_499, w_032_500, w_032_501, w_032_502, w_032_503, w_032_504, w_032_505, w_032_506, w_032_507, w_032_508, w_032_509, w_032_510, w_032_511, w_032_512, w_032_513, w_032_514, w_032_515, w_032_516, w_032_517, w_032_518, w_032_519, w_032_520, w_032_521, w_032_522, w_032_523, w_032_525, w_032_526, w_032_527, w_032_528, w_032_530, w_032_531, w_032_532, w_032_533, w_032_534, w_032_535, w_032_536, w_032_537, w_032_538, w_032_539, w_032_540, w_032_541, w_032_542, w_032_543, w_032_544, w_032_545, w_032_546, w_032_547, w_032_548, w_032_549, w_032_550, w_032_551, w_032_552, w_032_553, w_032_554, w_032_555, w_032_556, w_032_557, w_032_558, w_032_559, w_032_560, w_032_561, w_032_562, w_032_563, w_032_564, w_032_565, w_032_566, w_032_567, w_032_568, w_032_569, w_032_570, w_032_571, w_032_572, w_032_573, w_032_574, w_032_575, w_032_576, w_032_577, w_032_578, w_032_579, w_032_580, w_032_581, w_032_582, w_032_583, w_032_584, w_032_585, w_032_586, w_032_587, w_032_588, w_032_589, w_032_590, w_032_591, w_032_592, w_032_593, w_032_594, w_032_595, w_032_596, w_032_597, w_032_598, w_032_599, w_032_600, w_032_601, w_032_602, w_032_603, w_032_604, w_032_605, w_032_606, w_032_607, w_032_608, w_032_609, w_032_610, w_032_611, w_032_612, w_032_613, w_032_614, w_032_615, w_032_616, w_032_617, w_032_618, w_032_619, w_032_620, w_032_621, w_032_622, w_032_623, w_032_624, w_032_625, w_032_626, w_032_627, w_032_628, w_032_629, w_032_630, w_032_631, w_032_632, w_032_633, w_032_634, w_032_635, w_032_636, w_032_637, w_032_638, w_032_639, w_032_640, w_032_641, w_032_642, w_032_643, w_032_644, w_032_645, w_032_646, w_032_647, w_032_648, w_032_649, w_032_650, w_032_651, w_032_652, w_032_653, w_032_654, w_032_655, w_032_656, w_032_657, w_032_658, w_032_659, w_032_660, w_032_661, w_032_662, w_032_663, w_032_664, w_032_665, w_032_666, w_032_667, w_032_668, w_032_669, w_032_670, w_032_671, w_032_672, w_032_673, w_032_674, w_032_675, w_032_676, w_032_677, w_032_678, w_032_679, w_032_680, w_032_681, w_032_682, w_032_683, w_032_684, w_032_685, w_032_686, w_032_687, w_032_688, w_032_689, w_032_690, w_032_691, w_032_692, w_032_693, w_032_694, w_032_695, w_032_696, w_032_697, w_032_698, w_032_699, w_032_700, w_032_701, w_032_702, w_032_703, w_032_704, w_032_705, w_032_706, w_032_707, w_032_708, w_032_709, w_032_710, w_032_711, w_032_712, w_032_713, w_032_714, w_032_715, w_032_716, w_032_717, w_032_718, w_032_719, w_032_720, w_032_721, w_032_722, w_032_724, w_032_725, w_032_726, w_032_727, w_032_728, w_032_729, w_032_730, w_032_731, w_032_732, w_032_733, w_032_734, w_032_735, w_032_736, w_032_737, w_032_738, w_032_739, w_032_740, w_032_741, w_032_742, w_032_743, w_032_744, w_032_745, w_032_747, w_032_748, w_032_749, w_032_750, w_032_751, w_032_752, w_032_753, w_032_754, w_032_755, w_032_756, w_032_757, w_032_758, w_032_759, w_032_760, w_032_761, w_032_762, w_032_763, w_032_764, w_032_765, w_032_766, w_032_767, w_032_768, w_032_769, w_032_771, w_032_772, w_032_773, w_032_774, w_032_775, w_032_776, w_032_777, w_032_778, w_032_779, w_032_780, w_032_781, w_032_782, w_032_783, w_032_784, w_032_785, w_032_786, w_032_787, w_032_788, w_032_789, w_032_790, w_032_791, w_032_792, w_032_793, w_032_794, w_032_795, w_032_796, w_032_797, w_032_798, w_032_799, w_032_800, w_032_801, w_032_802, w_032_803, w_032_804, w_032_805, w_032_806, w_032_807, w_032_808, w_032_809, w_032_810, w_032_811, w_032_812, w_032_813, w_032_814, w_032_815, w_032_816, w_032_817, w_032_818, w_032_819, w_032_820, w_032_821, w_032_822, w_032_823, w_032_824, w_032_825, w_032_826, w_032_827, w_032_828, w_032_829, w_032_830, w_032_831, w_032_832, w_032_833, w_032_834, w_032_835, w_032_836, w_032_837, w_032_838, w_032_839, w_032_840, w_032_841, w_032_842, w_032_843, w_032_844, w_032_845, w_032_846, w_032_847, w_032_848, w_032_849, w_032_850, w_032_851, w_032_852, w_032_853, w_032_854, w_032_855, w_032_856, w_032_857, w_032_858, w_032_859, w_032_860, w_032_861, w_032_862, w_032_863, w_032_864, w_032_865, w_032_866, w_032_867, w_032_868, w_032_869, w_032_870, w_032_871, w_032_872, w_032_873, w_032_874, w_032_875, w_032_876, w_032_877, w_032_878, w_032_879, w_032_880, w_032_881, w_032_882, w_032_883, w_032_884, w_032_885, w_032_886, w_032_887, w_032_888, w_032_889, w_032_890, w_032_891, w_032_892, w_032_893, w_032_894, w_032_896, w_032_897, w_032_899, w_032_900, w_032_901, w_032_902, w_032_903, w_032_904, w_032_905, w_032_906, w_032_907, w_032_908, w_032_909, w_032_910, w_032_911, w_032_912, w_032_913, w_032_914, w_032_915, w_032_916, w_032_917, w_032_918, w_032_919, w_032_920, w_032_921, w_032_922, w_032_923, w_032_924, w_032_925, w_032_926, w_032_927, w_032_928, w_032_929, w_032_930, w_032_931, w_032_932, w_032_933, w_032_934, w_032_936, w_032_937, w_032_938, w_032_939, w_032_940, w_032_941, w_032_942, w_032_943, w_032_944, w_032_945, w_032_946, w_032_947, w_032_948, w_032_949, w_032_950, w_032_951, w_032_952, w_032_953, w_032_954, w_032_955, w_032_956, w_032_957, w_032_958, w_032_959, w_032_960, w_032_961, w_032_962, w_032_963, w_032_964, w_032_965, w_032_966, w_032_967, w_032_968, w_032_969, w_032_970, w_032_971, w_032_972, w_032_973, w_032_974, w_032_975, w_032_976, w_032_977, w_032_978, w_032_979, w_032_980, w_032_981, w_032_982, w_032_983, w_032_984, w_032_985, w_032_986, w_032_987, w_032_988, w_032_989, w_032_990, w_032_991, w_032_992, w_032_993, w_032_994, w_032_995, w_032_996, w_032_997, w_032_998, w_032_999, w_032_1000, w_032_1001, w_032_1002, w_032_1003, w_032_1004, w_032_1005, w_032_1006, w_032_1007, w_032_1008, w_032_1009, w_032_1010, w_032_1011, w_032_1012, w_032_1013, w_032_1014, w_032_1015, w_032_1016, w_032_1017, w_032_1018, w_032_1019, w_032_1020, w_032_1021, w_032_1022, w_032_1023, w_032_1025, w_032_1026, w_032_1027, w_032_1028, w_032_1029, w_032_1030, w_032_1031, w_032_1032, w_032_1033, w_032_1034, w_032_1035, w_032_1036, w_032_1037, w_032_1038, w_032_1039, w_032_1040, w_032_1041, w_032_1042, w_032_1043, w_032_1044, w_032_1045, w_032_1046, w_032_1047, w_032_1048, w_032_1049, w_032_1050, w_032_1051, w_032_1052, w_032_1053, w_032_1054, w_032_1055, w_032_1056, w_032_1057, w_032_1058, w_032_1060, w_032_1061, w_032_1062, w_032_1063, w_032_1064, w_032_1065, w_032_1066, w_032_1067, w_032_1068, w_032_1069, w_032_1070, w_032_1071, w_032_1072, w_032_1073, w_032_1074, w_032_1075, w_032_1076, w_032_1077, w_032_1078, w_032_1079, w_032_1080, w_032_1081, w_032_1082, w_032_1083, w_032_1084, w_032_1085, w_032_1086, w_032_1087, w_032_1088, w_032_1089, w_032_1090, w_032_1091, w_032_1092, w_032_1093, w_032_1094, w_032_1095, w_032_1096, w_032_1097, w_032_1098, w_032_1099, w_032_1100, w_032_1101, w_032_1102, w_032_1103, w_032_1104, w_032_1105, w_032_1106, w_032_1107, w_032_1108, w_032_1109, w_032_1110, w_032_1111, w_032_1112, w_032_1113, w_032_1114, w_032_1115, w_032_1116, w_032_1117, w_032_1118, w_032_1119, w_032_1120, w_032_1121, w_032_1122, w_032_1123, w_032_1124, w_032_1125, w_032_1126, w_032_1127, w_032_1128, w_032_1129, w_032_1130, w_032_1131, w_032_1132, w_032_1133, w_032_1134, w_032_1135, w_032_1136, w_032_1137, w_032_1138, w_032_1139, w_032_1140, w_032_1141, w_032_1142, w_032_1143, w_032_1144, w_032_1145, w_032_1146, w_032_1147, w_032_1148, w_032_1149, w_032_1150, w_032_1151, w_032_1152, w_032_1153, w_032_1154, w_032_1155, w_032_1156, w_032_1157, w_032_1158, w_032_1159, w_032_1160, w_032_1161, w_032_1162, w_032_1163, w_032_1164, w_032_1165, w_032_1166, w_032_1167, w_032_1168, w_032_1169, w_032_1170;
  wire w_033_000, w_033_001, w_033_002, w_033_003, w_033_004, w_033_005, w_033_006, w_033_007, w_033_009, w_033_013, w_033_015, w_033_016, w_033_017, w_033_019, w_033_021, w_033_022, w_033_023, w_033_024, w_033_025, w_033_026, w_033_028, w_033_029, w_033_030, w_033_031, w_033_032, w_033_034, w_033_035, w_033_036, w_033_037, w_033_038, w_033_039, w_033_040, w_033_041, w_033_042, w_033_043, w_033_044, w_033_045, w_033_046, w_033_047, w_033_048, w_033_049, w_033_050, w_033_052, w_033_053, w_033_054, w_033_055, w_033_056, w_033_058, w_033_059, w_033_061, w_033_062, w_033_064, w_033_065, w_033_066, w_033_068, w_033_069, w_033_070, w_033_072, w_033_073, w_033_075, w_033_076, w_033_077, w_033_078, w_033_080, w_033_081, w_033_082, w_033_083, w_033_084, w_033_085, w_033_086, w_033_087, w_033_088, w_033_089, w_033_090, w_033_091, w_033_093, w_033_095, w_033_096, w_033_097, w_033_098, w_033_099, w_033_100, w_033_101, w_033_102, w_033_103, w_033_104, w_033_105, w_033_106, w_033_107, w_033_108, w_033_109, w_033_110, w_033_111, w_033_112, w_033_113, w_033_114, w_033_115, w_033_116, w_033_117, w_033_118, w_033_119, w_033_120, w_033_121, w_033_122, w_033_124, w_033_125, w_033_126, w_033_127, w_033_128, w_033_129, w_033_130, w_033_132, w_033_133, w_033_135, w_033_138, w_033_139, w_033_140, w_033_141, w_033_143, w_033_144, w_033_145, w_033_146, w_033_147, w_033_148, w_033_149, w_033_150, w_033_151, w_033_152, w_033_153, w_033_154, w_033_155, w_033_156, w_033_157, w_033_158, w_033_159, w_033_161, w_033_162, w_033_163, w_033_165, w_033_167, w_033_168, w_033_169, w_033_170, w_033_171, w_033_172, w_033_173, w_033_174, w_033_177, w_033_178, w_033_179, w_033_181, w_033_182, w_033_183, w_033_184, w_033_185, w_033_186, w_033_187, w_033_188, w_033_190, w_033_191, w_033_192, w_033_193, w_033_194, w_033_195, w_033_196, w_033_197, w_033_198, w_033_199, w_033_200, w_033_201, w_033_202, w_033_203, w_033_204, w_033_205, w_033_206, w_033_207, w_033_208, w_033_209, w_033_210, w_033_211, w_033_212, w_033_213, w_033_214, w_033_215, w_033_216, w_033_217, w_033_218, w_033_219, w_033_220, w_033_221, w_033_222, w_033_223, w_033_224, w_033_225, w_033_226, w_033_227, w_033_228, w_033_229, w_033_230, w_033_231, w_033_232, w_033_233, w_033_235, w_033_237, w_033_238, w_033_239, w_033_242, w_033_243, w_033_244, w_033_245, w_033_246, w_033_247, w_033_248, w_033_249, w_033_250, w_033_253, w_033_254, w_033_255, w_033_257, w_033_258, w_033_262, w_033_263, w_033_264, w_033_265, w_033_266, w_033_267, w_033_268, w_033_269, w_033_270, w_033_271, w_033_272, w_033_273, w_033_275, w_033_276, w_033_278, w_033_279, w_033_280, w_033_281, w_033_282, w_033_283, w_033_284, w_033_285, w_033_286, w_033_287, w_033_289, w_033_291, w_033_293, w_033_295, w_033_297, w_033_298, w_033_299, w_033_300, w_033_301, w_033_302, w_033_303, w_033_304, w_033_305, w_033_306, w_033_310, w_033_312, w_033_313, w_033_314, w_033_315, w_033_316, w_033_318, w_033_319, w_033_320, w_033_321, w_033_322, w_033_323, w_033_324, w_033_325, w_033_327, w_033_328, w_033_329, w_033_330, w_033_333, w_033_334, w_033_335, w_033_336, w_033_337, w_033_339, w_033_340, w_033_342, w_033_344, w_033_345, w_033_346, w_033_347, w_033_348, w_033_349, w_033_350, w_033_352, w_033_353, w_033_354, w_033_355, w_033_356, w_033_357, w_033_358, w_033_359, w_033_360, w_033_361, w_033_362, w_033_363, w_033_364, w_033_365, w_033_366, w_033_367, w_033_368, w_033_370, w_033_371, w_033_372, w_033_373, w_033_374, w_033_375, w_033_376, w_033_377, w_033_378, w_033_379, w_033_380, w_033_381, w_033_382, w_033_383, w_033_384, w_033_385, w_033_386, w_033_389, w_033_390, w_033_391, w_033_393, w_033_394, w_033_395, w_033_396, w_033_397, w_033_398, w_033_399, w_033_401, w_033_402, w_033_403, w_033_404, w_033_405, w_033_406, w_033_408, w_033_409, w_033_410, w_033_411, w_033_412, w_033_413, w_033_415, w_033_416, w_033_417, w_033_419, w_033_420, w_033_421, w_033_422, w_033_423, w_033_424, w_033_426, w_033_427, w_033_428, w_033_429, w_033_430, w_033_431, w_033_432, w_033_433, w_033_434, w_033_435, w_033_437, w_033_438, w_033_439, w_033_441, w_033_443, w_033_444, w_033_445, w_033_446, w_033_447, w_033_448, w_033_449, w_033_450, w_033_452, w_033_453, w_033_454, w_033_455, w_033_456, w_033_457, w_033_458, w_033_459, w_033_460, w_033_461, w_033_462, w_033_463, w_033_464, w_033_465, w_033_466, w_033_467, w_033_468, w_033_470, w_033_471, w_033_472, w_033_473, w_033_475, w_033_476, w_033_477, w_033_478, w_033_479, w_033_481, w_033_482, w_033_483, w_033_484, w_033_485, w_033_486, w_033_487, w_033_488, w_033_489, w_033_490, w_033_491, w_033_492, w_033_493, w_033_495, w_033_496, w_033_498, w_033_499, w_033_500, w_033_501, w_033_502, w_033_503, w_033_504, w_033_505, w_033_506, w_033_507, w_033_508, w_033_509, w_033_510, w_033_511, w_033_512, w_033_513, w_033_514, w_033_515, w_033_516, w_033_517, w_033_518, w_033_519, w_033_520, w_033_521, w_033_522, w_033_523, w_033_527, w_033_528, w_033_529, w_033_531, w_033_532, w_033_533, w_033_534, w_033_537, w_033_538, w_033_539, w_033_540, w_033_541, w_033_542, w_033_543, w_033_545, w_033_546, w_033_547, w_033_548, w_033_549, w_033_550, w_033_551, w_033_553, w_033_554, w_033_555, w_033_556, w_033_558, w_033_559, w_033_560, w_033_562, w_033_563, w_033_564, w_033_565, w_033_566, w_033_568, w_033_569, w_033_570, w_033_571, w_033_572, w_033_573, w_033_574, w_033_575, w_033_576, w_033_578, w_033_579, w_033_580, w_033_581, w_033_582, w_033_583, w_033_584, w_033_585, w_033_586, w_033_587, w_033_589, w_033_591, w_033_593, w_033_594, w_033_595, w_033_596, w_033_597, w_033_598, w_033_599, w_033_601, w_033_602, w_033_603, w_033_604, w_033_606, w_033_607, w_033_608, w_033_610, w_033_612, w_033_613, w_033_614, w_033_615, w_033_618, w_033_619, w_033_620, w_033_621, w_033_622, w_033_623, w_033_624, w_033_625, w_033_626, w_033_627, w_033_628, w_033_629, w_033_631, w_033_632, w_033_633, w_033_635, w_033_636, w_033_637, w_033_638, w_033_639, w_033_640, w_033_641, w_033_642, w_033_643, w_033_644, w_033_645, w_033_646, w_033_647, w_033_648, w_033_649, w_033_650, w_033_651, w_033_653, w_033_654, w_033_655, w_033_657, w_033_658, w_033_659, w_033_661, w_033_662, w_033_663, w_033_664, w_033_665, w_033_666, w_033_667, w_033_668, w_033_669, w_033_671, w_033_673, w_033_674, w_033_676, w_033_677, w_033_678, w_033_679, w_033_681, w_033_682, w_033_684, w_033_686, w_033_687, w_033_688, w_033_689, w_033_690, w_033_691, w_033_692, w_033_693, w_033_694, w_033_695, w_033_696, w_033_698, w_033_699, w_033_700, w_033_701, w_033_702, w_033_703, w_033_704, w_033_705, w_033_707, w_033_708, w_033_709, w_033_710, w_033_712, w_033_714, w_033_715, w_033_717, w_033_718, w_033_719, w_033_720, w_033_721, w_033_723, w_033_724, w_033_725, w_033_726, w_033_727, w_033_729, w_033_731, w_033_733, w_033_734, w_033_735, w_033_737, w_033_738, w_033_739, w_033_740, w_033_741, w_033_742, w_033_743, w_033_746, w_033_747, w_033_749, w_033_750, w_033_751, w_033_752, w_033_753, w_033_754, w_033_755, w_033_756, w_033_759, w_033_760, w_033_761, w_033_762, w_033_763, w_033_765, w_033_766, w_033_767, w_033_769, w_033_770, w_033_772, w_033_773, w_033_775, w_033_776, w_033_777, w_033_778, w_033_779, w_033_780, w_033_781, w_033_783, w_033_784, w_033_786, w_033_787, w_033_788, w_033_789, w_033_790, w_033_791, w_033_792, w_033_794, w_033_795, w_033_796, w_033_797, w_033_798, w_033_799, w_033_800, w_033_801, w_033_802, w_033_803, w_033_804, w_033_805, w_033_806, w_033_807, w_033_808, w_033_809, w_033_810, w_033_811, w_033_812, w_033_815, w_033_816, w_033_817, w_033_819, w_033_820, w_033_821, w_033_822, w_033_823, w_033_824, w_033_825, w_033_826, w_033_827, w_033_828, w_033_829, w_033_830, w_033_831, w_033_832, w_033_833, w_033_835, w_033_836, w_033_837, w_033_838, w_033_840, w_033_841, w_033_842, w_033_843, w_033_844, w_033_845, w_033_846, w_033_847, w_033_848, w_033_849, w_033_852, w_033_854, w_033_855, w_033_856, w_033_857, w_033_858, w_033_859, w_033_860, w_033_861, w_033_862, w_033_863, w_033_864, w_033_865, w_033_866, w_033_867, w_033_868, w_033_869, w_033_870, w_033_873, w_033_874, w_033_875, w_033_876, w_033_877, w_033_878, w_033_879, w_033_880, w_033_881, w_033_882, w_033_883, w_033_884, w_033_885, w_033_886, w_033_887, w_033_888, w_033_889, w_033_890, w_033_891, w_033_892, w_033_893, w_033_894, w_033_897, w_033_898, w_033_899, w_033_901, w_033_902, w_033_903, w_033_904, w_033_905, w_033_906, w_033_907, w_033_908, w_033_909, w_033_910, w_033_913, w_033_915, w_033_916, w_033_917, w_033_918, w_033_921, w_033_922, w_033_923, w_033_924, w_033_926, w_033_928, w_033_929, w_033_930, w_033_931, w_033_932, w_033_933, w_033_934, w_033_936, w_033_937, w_033_938, w_033_939, w_033_941, w_033_942, w_033_943, w_033_944, w_033_945, w_033_946, w_033_947, w_033_948, w_033_949, w_033_950, w_033_951, w_033_952, w_033_953, w_033_954, w_033_955, w_033_956, w_033_957, w_033_958, w_033_959, w_033_960, w_033_961, w_033_962, w_033_963, w_033_964, w_033_965, w_033_966, w_033_968, w_033_969, w_033_970, w_033_971, w_033_972, w_033_973, w_033_974, w_033_975, w_033_978, w_033_979, w_033_980, w_033_981, w_033_982, w_033_983, w_033_984, w_033_985, w_033_986, w_033_987, w_033_988, w_033_989, w_033_990, w_033_991, w_033_992, w_033_994, w_033_995, w_033_996, w_033_997, w_033_998, w_033_1000, w_033_1001, w_033_1002, w_033_1003, w_033_1004, w_033_1005, w_033_1007, w_033_1008, w_033_1009, w_033_1010, w_033_1011, w_033_1012, w_033_1013, w_033_1015, w_033_1016, w_033_1018, w_033_1020, w_033_1021, w_033_1023, w_033_1024, w_033_1025, w_033_1026, w_033_1027, w_033_1028, w_033_1029, w_033_1031, w_033_1032, w_033_1033, w_033_1034, w_033_1035, w_033_1036, w_033_1037, w_033_1038, w_033_1039, w_033_1040, w_033_1041, w_033_1042, w_033_1044, w_033_1045, w_033_1046, w_033_1047, w_033_1048, w_033_1049, w_033_1050, w_033_1051, w_033_1052, w_033_1054, w_033_1056, w_033_1057, w_033_1058, w_033_1059, w_033_1060, w_033_1061, w_033_1062, w_033_1063, w_033_1064, w_033_1065, w_033_1067, w_033_1068, w_033_1070, w_033_1071, w_033_1072, w_033_1073, w_033_1074, w_033_1075, w_033_1076, w_033_1077, w_033_1078, w_033_1079, w_033_1080, w_033_1081, w_033_1082, w_033_1083, w_033_1084, w_033_1086, w_033_1087, w_033_1088, w_033_1090, w_033_1091, w_033_1092, w_033_1093, w_033_1094, w_033_1095, w_033_1096, w_033_1097, w_033_1098, w_033_1099, w_033_1100, w_033_1101, w_033_1102, w_033_1103, w_033_1104, w_033_1105, w_033_1107, w_033_1108, w_033_1109, w_033_1110, w_033_1114, w_033_1115, w_033_1116, w_033_1117, w_033_1118, w_033_1119, w_033_1120, w_033_1122, w_033_1123, w_033_1124, w_033_1125, w_033_1127, w_033_1128, w_033_1129, w_033_1130, w_033_1131, w_033_1132, w_033_1133, w_033_1135, w_033_1138, w_033_1139, w_033_1142, w_033_1143, w_033_1144, w_033_1146, w_033_1148, w_033_1149, w_033_1152, w_033_1154, w_033_1155, w_033_1156, w_033_1158, w_033_1159, w_033_1160, w_033_1163, w_033_1164, w_033_1166, w_033_1167, w_033_1168, w_033_1171, w_033_1174, w_033_1175, w_033_1176, w_033_1177, w_033_1178, w_033_1182, w_033_1183, w_033_1185, w_033_1187, w_033_1189, w_033_1190, w_033_1191, w_033_1193, w_033_1194, w_033_1195, w_033_1196, w_033_1197, w_033_1199, w_033_1201, w_033_1202, w_033_1203, w_033_1205, w_033_1206, w_033_1207, w_033_1208, w_033_1211, w_033_1212, w_033_1215, w_033_1216, w_033_1217, w_033_1218, w_033_1219, w_033_1220, w_033_1221, w_033_1223, w_033_1224, w_033_1228, w_033_1229, w_033_1230, w_033_1231, w_033_1232, w_033_1233, w_033_1234, w_033_1235, w_033_1238, w_033_1239, w_033_1240, w_033_1243, w_033_1244, w_033_1245, w_033_1246, w_033_1248, w_033_1249, w_033_1251, w_033_1254, w_033_1258, w_033_1259, w_033_1260, w_033_1261, w_033_1262, w_033_1264, w_033_1265, w_033_1266, w_033_1268, w_033_1271, w_033_1272, w_033_1273, w_033_1274, w_033_1276, w_033_1277, w_033_1278, w_033_1279, w_033_1280, w_033_1281, w_033_1282, w_033_1284, w_033_1285, w_033_1290, w_033_1292, w_033_1293, w_033_1298, w_033_1299, w_033_1302, w_033_1305, w_033_1307, w_033_1308, w_033_1309, w_033_1310, w_033_1311, w_033_1313, w_033_1314, w_033_1317, w_033_1318, w_033_1319, w_033_1320, w_033_1322, w_033_1323, w_033_1324, w_033_1326, w_033_1328, w_033_1330, w_033_1335, w_033_1336, w_033_1337, w_033_1340, w_033_1341, w_033_1342, w_033_1345, w_033_1346, w_033_1347, w_033_1348, w_033_1350, w_033_1351, w_033_1352, w_033_1353, w_033_1354, w_033_1355, w_033_1356, w_033_1360, w_033_1361, w_033_1363, w_033_1366, w_033_1368, w_033_1369, w_033_1370, w_033_1371, w_033_1373, w_033_1374, w_033_1375, w_033_1376, w_033_1378, w_033_1379, w_033_1383, w_033_1384, w_033_1385, w_033_1387, w_033_1389, w_033_1390, w_033_1392, w_033_1394, w_033_1395, w_033_1397, w_033_1398, w_033_1400, w_033_1402, w_033_1403, w_033_1406, w_033_1408, w_033_1409, w_033_1410, w_033_1412, w_033_1413, w_033_1414, w_033_1415, w_033_1416, w_033_1420, w_033_1421, w_033_1424, w_033_1430, w_033_1431, w_033_1432, w_033_1437, w_033_1438, w_033_1439, w_033_1440, w_033_1442, w_033_1443, w_033_1444, w_033_1446, w_033_1447, w_033_1451, w_033_1452, w_033_1453, w_033_1454, w_033_1456, w_033_1458, w_033_1459, w_033_1460, w_033_1463, w_033_1464, w_033_1465, w_033_1466, w_033_1468, w_033_1471, w_033_1473, w_033_1475, w_033_1477, w_033_1479, w_033_1481, w_033_1482, w_033_1484, w_033_1485, w_033_1486, w_033_1488, w_033_1489, w_033_1490, w_033_1493, w_033_1495, w_033_1496, w_033_1499, w_033_1500, w_033_1501, w_033_1503, w_033_1505, w_033_1507, w_033_1508, w_033_1509, w_033_1513, w_033_1514, w_033_1516, w_033_1517, w_033_1518, w_033_1519, w_033_1521, w_033_1523, w_033_1525, w_033_1527, w_033_1529, w_033_1530, w_033_1533, w_033_1535, w_033_1539, w_033_1540, w_033_1541, w_033_1542, w_033_1543, w_033_1544, w_033_1545, w_033_1546, w_033_1548, w_033_1549, w_033_1550, w_033_1552, w_033_1553, w_033_1554, w_033_1556, w_033_1557, w_033_1558, w_033_1561, w_033_1562, w_033_1563, w_033_1564, w_033_1568, w_033_1569, w_033_1570, w_033_1572, w_033_1574, w_033_1575, w_033_1576, w_033_1580, w_033_1581, w_033_1582, w_033_1584, w_033_1585, w_033_1586, w_033_1590, w_033_1591, w_033_1592, w_033_1594, w_033_1595, w_033_1597, w_033_1600, w_033_1601, w_033_1602, w_033_1603, w_033_1604, w_033_1605, w_033_1606, w_033_1608, w_033_1611, w_033_1617, w_033_1618, w_033_1619, w_033_1620, w_033_1624, w_033_1626, w_033_1627, w_033_1628, w_033_1630, w_033_1631, w_033_1632, w_033_1633, w_033_1634, w_033_1636, w_033_1637, w_033_1641, w_033_1642, w_033_1644, w_033_1645, w_033_1647, w_033_1648, w_033_1649, w_033_1650, w_033_1651, w_033_1652, w_033_1654, w_033_1655, w_033_1657, w_033_1659, w_033_1660, w_033_1661, w_033_1662, w_033_1665, w_033_1671, w_033_1672, w_033_1673, w_033_1674, w_033_1675, w_033_1676, w_033_1677, w_033_1680, w_033_1682, w_033_1683, w_033_1685, w_033_1687, w_033_1689, w_033_1691, w_033_1694, w_033_1695, w_033_1700, w_033_1701, w_033_1702, w_033_1705, w_033_1707, w_033_1708, w_033_1709, w_033_1711, w_033_1713, w_033_1714, w_033_1717, w_033_1718, w_033_1720, w_033_1723, w_033_1724, w_033_1725, w_033_1726, w_033_1727, w_033_1728, w_033_1729, w_033_1733, w_033_1734, w_033_1735, w_033_1736, w_033_1737, w_033_1740, w_033_1743, w_033_1745, w_033_1747, w_033_1751, w_033_1753, w_033_1755, w_033_1758, w_033_1760, w_033_1761, w_033_1763, w_033_1764, w_033_1765, w_033_1766, w_033_1767, w_033_1771, w_033_1772, w_033_1775, w_033_1777, w_033_1779, w_033_1780, w_033_1781, w_033_1784, w_033_1787, w_033_1788, w_033_1790, w_033_1792, w_033_1793, w_033_1794, w_033_1797, w_033_1799, w_033_1801, w_033_1804, w_033_1805, w_033_1806, w_033_1807, w_033_1810, w_033_1811, w_033_1814, w_033_1815, w_033_1816, w_033_1819, w_033_1821, w_033_1822, w_033_1824, w_033_1825, w_033_1826, w_033_1828, w_033_1830, w_033_1831, w_033_1832, w_033_1833, w_033_1836, w_033_1837, w_033_1838, w_033_1839, w_033_1840, w_033_1841, w_033_1842, w_033_1843, w_033_1846, w_033_1847, w_033_1849, w_033_1852, w_033_1853, w_033_1855, w_033_1856, w_033_1857, w_033_1858, w_033_1859, w_033_1860, w_033_1861, w_033_1862, w_033_1866, w_033_1868, w_033_1869, w_033_1872, w_033_1873, w_033_1874, w_033_1875, w_033_1876, w_033_1878, w_033_1879, w_033_1880, w_033_1881, w_033_1882, w_033_1883, w_033_1885, w_033_1886, w_033_1888, w_033_1889, w_033_1890, w_033_1892, w_033_1893, w_033_1895, w_033_1896, w_033_1897, w_033_1898, w_033_1899, w_033_1901, w_033_1906, w_033_1907, w_033_1911, w_033_1912, w_033_1913, w_033_1914, w_033_1915, w_033_1916, w_033_1918, w_033_1919, w_033_1920, w_033_1921, w_033_1922, w_033_1925, w_033_1927, w_033_1931, w_033_1933, w_033_1935, w_033_1940, w_033_1941, w_033_1942, w_033_1944, w_033_1945, w_033_1948, w_033_1949, w_033_1950, w_033_1951, w_033_1954, w_033_1956, w_033_1957, w_033_1960, w_033_1962, w_033_1963, w_033_1965, w_033_1966, w_033_1967, w_033_1969, w_033_1970, w_033_1971, w_033_1974, w_033_1976, w_033_1978, w_033_1979, w_033_1981, w_033_1983, w_033_1984, w_033_1985, w_033_1986, w_033_1987, w_033_1988, w_033_1989, w_033_1990, w_033_1993, w_033_1997, w_033_1998, w_033_1999, w_033_2000, w_033_2001, w_033_2006, w_033_2007, w_033_2009, w_033_2011, w_033_2014, w_033_2016, w_033_2019, w_033_2022, w_033_2023, w_033_2026, w_033_2029, w_033_2031, w_033_2032, w_033_2035, w_033_2039, w_033_2041, w_033_2042, w_033_2046, w_033_2047, w_033_2049, w_033_2051, w_033_2052, w_033_2053, w_033_2054, w_033_2055, w_033_2058, w_033_2060, w_033_2061, w_033_2062, w_033_2063, w_033_2064, w_033_2065, w_033_2067, w_033_2068, w_033_2071, w_033_2073, w_033_2074, w_033_2075, w_033_2076, w_033_2077, w_033_2080, w_033_2081, w_033_2083, w_033_2084, w_033_2086, w_033_2087, w_033_2088, w_033_2091, w_033_2092, w_033_2093, w_033_2094, w_033_2095, w_033_2096, w_033_2098, w_033_2099, w_033_2100, w_033_2104, w_033_2107, w_033_2108, w_033_2109, w_033_2111, w_033_2112, w_033_2116, w_033_2117, w_033_2119, w_033_2120, w_033_2122, w_033_2124, w_033_2125, w_033_2126, w_033_2127, w_033_2128, w_033_2129, w_033_2130, w_033_2131, w_033_2134, w_033_2135, w_033_2137, w_033_2138, w_033_2139, w_033_2141, w_033_2142, w_033_2144, w_033_2147, w_033_2148, w_033_2150, w_033_2151, w_033_2153, w_033_2156, w_033_2158, w_033_2160, w_033_2161, w_033_2162, w_033_2163, w_033_2164, w_033_2165, w_033_2166, w_033_2167, w_033_2172, w_033_2173, w_033_2174, w_033_2176, w_033_2177, w_033_2178, w_033_2179, w_033_2180, w_033_2181, w_033_2182, w_033_2186, w_033_2188, w_033_2189, w_033_2191, w_033_2192, w_033_2197, w_033_2198, w_033_2201, w_033_2204, w_033_2209, w_033_2210, w_033_2212, w_033_2213, w_033_2214, w_033_2215, w_033_2216, w_033_2217, w_033_2220, w_033_2221, w_033_2223, w_033_2225, w_033_2226, w_033_2227, w_033_2228, w_033_2229, w_033_2230, w_033_2232, w_033_2233, w_033_2234, w_033_2237, w_033_2238, w_033_2239, w_033_2240, w_033_2241, w_033_2243, w_033_2244, w_033_2245, w_033_2246, w_033_2247, w_033_2250, w_033_2253, w_033_2254, w_033_2259, w_033_2260, w_033_2261, w_033_2263, w_033_2264, w_033_2266, w_033_2267, w_033_2268, w_033_2271, w_033_2272, w_033_2273, w_033_2274, w_033_2275, w_033_2277, w_033_2278, w_033_2280, w_033_2284, w_033_2285, w_033_2286, w_033_2289, w_033_2293, w_033_2294, w_033_2295, w_033_2296, w_033_2297, w_033_2299, w_033_2301, w_033_2302, w_033_2303, w_033_2304, w_033_2305, w_033_2306, w_033_2308, w_033_2309, w_033_2310, w_033_2312, w_033_2316, w_033_2319, w_033_2320, w_033_2321, w_033_2322, w_033_2323, w_033_2324, w_033_2325, w_033_2327, w_033_2328, w_033_2334, w_033_2336, w_033_2337, w_033_2338, w_033_2339, w_033_2340, w_033_2342, w_033_2346, w_033_2347, w_033_2348, w_033_2349, w_033_2350, w_033_2351, w_033_2352, w_033_2353, w_033_2355, w_033_2357, w_033_2358, w_033_2359, w_033_2361, w_033_2362, w_033_2364, w_033_2365, w_033_2366, w_033_2367, w_033_2368, w_033_2369, w_033_2372, w_033_2373, w_033_2379, w_033_2380, w_033_2381, w_033_2383, w_033_2384, w_033_2385, w_033_2387, w_033_2389, w_033_2390, w_033_2391, w_033_2392, w_033_2395, w_033_2396, w_033_2397, w_033_2399, w_033_2402, w_033_2404, w_033_2405, w_033_2406, w_033_2407, w_033_2410, w_033_2411, w_033_2412, w_033_2414, w_033_2415, w_033_2417, w_033_2418, w_033_2421, w_033_2423, w_033_2424, w_033_2425, w_033_2426, w_033_2427, w_033_2428, w_033_2429, w_033_2432, w_033_2433, w_033_2434, w_033_2437, w_033_2438, w_033_2439, w_033_2441, w_033_2443, w_033_2444, w_033_2447, w_033_2448, w_033_2450, w_033_2451, w_033_2452, w_033_2453, w_033_2456, w_033_2457, w_033_2458, w_033_2459, w_033_2460, w_033_2462, w_033_2463, w_033_2464, w_033_2465, w_033_2467, w_033_2468, w_033_2470, w_033_2471, w_033_2472, w_033_2473, w_033_2474, w_033_2475, w_033_2476, w_033_2477, w_033_2478, w_033_2480, w_033_2481, w_033_2483, w_033_2486, w_033_2487, w_033_2490, w_033_2491, w_033_2492, w_033_2493, w_033_2494, w_033_2496, w_033_2498, w_033_2500, w_033_2502, w_033_2503, w_033_2504, w_033_2505, w_033_2507, w_033_2508, w_033_2509, w_033_2510, w_033_2511, w_033_2513, w_033_2515, w_033_2517, w_033_2518, w_033_2519, w_033_2520, w_033_2521, w_033_2523, w_033_2524, w_033_2525, w_033_2527, w_033_2529, w_033_2530, w_033_2531, w_033_2533, w_033_2534, w_033_2535, w_033_2539, w_033_2540, w_033_2543, w_033_2546, w_033_2547, w_033_2549, w_033_2550, w_033_2551, w_033_2552, w_033_2554, w_033_2557, w_033_2558, w_033_2561, w_033_2562, w_033_2563, w_033_2566, w_033_2569, w_033_2570, w_033_2571, w_033_2573, w_033_2574, w_033_2576, w_033_2577, w_033_2578, w_033_2581, w_033_2585, w_033_2586, w_033_2587, w_033_2588, w_033_2591, w_033_2592, w_033_2593, w_033_2594, w_033_2596, w_033_2597, w_033_2600, w_033_2603, w_033_2604, w_033_2609, w_033_2612, w_033_2616, w_033_2617, w_033_2619, w_033_2620, w_033_2622, w_033_2623, w_033_2624, w_033_2625, w_033_2627, w_033_2628, w_033_2630, w_033_2631, w_033_2633, w_033_2635, w_033_2636, w_033_2637, w_033_2639, w_033_2640, w_033_2642, w_033_2643, w_033_2644, w_033_2645, w_033_2648, w_033_2649, w_033_2650, w_033_2651, w_033_2652, w_033_2654, w_033_2655, w_033_2659, w_033_2660, w_033_2661, w_033_2663, w_033_2666, w_033_2668, w_033_2669, w_033_2671, w_033_2672, w_033_2673, w_033_2674, w_033_2677, w_033_2679, w_033_2680, w_033_2681, w_033_2682, w_033_2683, w_033_2685, w_033_2686, w_033_2687, w_033_2688, w_033_2689, w_033_2690, w_033_2692, w_033_2693, w_033_2694, w_033_2695, w_033_2696, w_033_2701, w_033_2704, w_033_2706, w_033_2708, w_033_2710, w_033_2711, w_033_2713, w_033_2715, w_033_2716, w_033_2720, w_033_2721, w_033_2724, w_033_2725, w_033_2727, w_033_2728, w_033_2729, w_033_2731, w_033_2732, w_033_2738, w_033_2740, w_033_2741, w_033_2742, w_033_2743, w_033_2744, w_033_2745, w_033_2747, w_033_2750, w_033_2751, w_033_2752, w_033_2754, w_033_2758, w_033_2759, w_033_2762, w_033_2763, w_033_2764, w_033_2765, w_033_2769, w_033_2770, w_033_2771, w_033_2772, w_033_2773, w_033_2774, w_033_2775, w_033_2776, w_033_2777, w_033_2778, w_033_2779, w_033_2780, w_033_2782, w_033_2783, w_033_2784, w_033_2791, w_033_2792, w_033_2794, w_033_2795, w_033_2796, w_033_2797, w_033_2798, w_033_2799, w_033_2800, w_033_2801, w_033_2802, w_033_2803, w_033_2805, w_033_2807, w_033_2808, w_033_2810, w_033_2811, w_033_2812, w_033_2814, w_033_2816, w_033_2817, w_033_2818, w_033_2821, w_033_2823, w_033_2825, w_033_2826, w_033_2830, w_033_2834, w_033_2835, w_033_2837, w_033_2841, w_033_2842, w_033_2843, w_033_2845, w_033_2847, w_033_2849, w_033_2851, w_033_2852, w_033_2853, w_033_2854, w_033_2855, w_033_2856, w_033_2861, w_033_2862, w_033_2863, w_033_2866, w_033_2870, w_033_2871, w_033_2872, w_033_2873, w_033_2874, w_033_2875, w_033_2876, w_033_2878, w_033_2879, w_033_2880, w_033_2882, w_033_2884, w_033_2890, w_033_2892, w_033_2893, w_033_2894, w_033_2895, w_033_2896, w_033_2897, w_033_2899, w_033_2900, w_033_2901, w_033_2902, w_033_2903, w_033_2904, w_033_2905, w_033_2906, w_033_2907, w_033_2908, w_033_2910, w_033_2911, w_033_2913, w_033_2915, w_033_2920, w_033_2923, w_033_2924, w_033_2926, w_033_2928, w_033_2930, w_033_2932, w_033_2936, w_033_2937, w_033_2939, w_033_2941, w_033_2942, w_033_2943, w_033_2945, w_033_2947, w_033_2949, w_033_2950, w_033_2951, w_033_2953, w_033_2954, w_033_2955, w_033_2956, w_033_2957, w_033_2958, w_033_2961, w_033_2962, w_033_2967, w_033_2968, w_033_2971, w_033_2974, w_033_2975, w_033_2977, w_033_2978, w_033_2982, w_033_2983, w_033_2984, w_033_2985, w_033_2986, w_033_2987, w_033_2989, w_033_2990, w_033_2991, w_033_2992, w_033_2994, w_033_2997, w_033_3000, w_033_3002, w_033_3004, w_033_3005, w_033_3006, w_033_3008, w_033_3010, w_033_3011, w_033_3012, w_033_3013, w_033_3014, w_033_3015, w_033_3016, w_033_3021, w_033_3022, w_033_3024, w_033_3025, w_033_3026, w_033_3028, w_033_3029, w_033_3030, w_033_3031, w_033_3032, w_033_3037, w_033_3039, w_033_3040, w_033_3041, w_033_3042, w_033_3043, w_033_3045, w_033_3046, w_033_3047, w_033_3048, w_033_3050, w_033_3052, w_033_3053, w_033_3054, w_033_3055, w_033_3056, w_033_3057, w_033_3060, w_033_3061, w_033_3062, w_033_3063, w_033_3064, w_033_3067, w_033_3068, w_033_3071, w_033_3072, w_033_3073, w_033_3075, w_033_3077, w_033_3078, w_033_3079, w_033_3081, w_033_3083, w_033_3084, w_033_3086, w_033_3089, w_033_3092, w_033_3093, w_033_3094, w_033_3096, w_033_3097, w_033_3098, w_033_3099, w_033_3100, w_033_3101, w_033_3102, w_033_3103, w_033_3104, w_033_3107, w_033_3108, w_033_3110, w_033_3112, w_033_3114, w_033_3115, w_033_3116, w_033_3117, w_033_3118, w_033_3120, w_033_3122, w_033_3123, w_033_3124, w_033_3125, w_033_3127, w_033_3129, w_033_3131, w_033_3132, w_033_3134, w_033_3135, w_033_3137, w_033_3138, w_033_3139, w_033_3142, w_033_3150, w_033_3152, w_033_3153, w_033_3154, w_033_3155, w_033_3156, w_033_3157, w_033_3158, w_033_3159, w_033_3163, w_033_3164, w_033_3165, w_033_3166, w_033_3167, w_033_3169, w_033_3170, w_033_3171, w_033_3172, w_033_3174, w_033_3175, w_033_3178, w_033_3180, w_033_3181, w_033_3182, w_033_3183, w_033_3185, w_033_3186, w_033_3190, w_033_3191, w_033_3192, w_033_3193, w_033_3195, w_033_3196, w_033_3197, w_033_3200, w_033_3201, w_033_3206, w_033_3207, w_033_3208, w_033_3209, w_033_3210, w_033_3211, w_033_3213, w_033_3214, w_033_3216, w_033_3217, w_033_3219, w_033_3220, w_033_3223, w_033_3224, w_033_3227, w_033_3231, w_033_3232, w_033_3233, w_033_3234, w_033_3235, w_033_3236, w_033_3237, w_033_3238, w_033_3239, w_033_3242, w_033_3244, w_033_3246, w_033_3249, w_033_3252, w_033_3254, w_033_3255, w_033_3256, w_033_3258, w_033_3261, w_033_3263, w_033_3265, w_033_3268, w_033_3269, w_033_3271, w_033_3273, w_033_3274, w_033_3275, w_033_3277, w_033_3279, w_033_3280, w_033_3282, w_033_3284, w_033_3285, w_033_3288, w_033_3290, w_033_3291, w_033_3292, w_033_3293, w_033_3294, w_033_3296, w_033_3297, w_033_3298, w_033_3299, w_033_3300, w_033_3301, w_033_3302, w_033_3303, w_033_3304, w_033_3305, w_033_3307, w_033_3309, w_033_3312, w_033_3314, w_033_3315, w_033_3316, w_033_3319, w_033_3323, w_033_3325, w_033_3326, w_033_3328, w_033_3330, w_033_3332, w_033_3333, w_033_3335, w_033_3336, w_033_3337, w_033_3338, w_033_3339, w_033_3342, w_033_3344, w_033_3345, w_033_3346, w_033_3347, w_033_3351, w_033_3354, w_033_3355, w_033_3358, w_033_3359, w_033_3360, w_033_3361, w_033_3366, w_033_3367, w_033_3368, w_033_3370, w_033_3371, w_033_3372, w_033_3373, w_033_3374, w_033_3377, w_033_3378, w_033_3383, w_033_3384, w_033_3385, w_033_3388, w_033_3392, w_033_3394, w_033_3395, w_033_3396, w_033_3397, w_033_3398, w_033_3403, w_033_3404, w_033_3410, w_033_3411, w_033_3412, w_033_3413, w_033_3414, w_033_3415, w_033_3416, w_033_3417, w_033_3420, w_033_3421, w_033_3422, w_033_3423, w_033_3424, w_033_3426, w_033_3427, w_033_3430, w_033_3431, w_033_3434, w_033_3436, w_033_3437, w_033_3438, w_033_3439, w_033_3440, w_033_3441, w_033_3443, w_033_3445, w_033_3446, w_033_3447, w_033_3448, w_033_3450, w_033_3451, w_033_3452, w_033_3453, w_033_3454, w_033_3455, w_033_3457, w_033_3458, w_033_3459, w_033_3461, w_033_3462, w_033_3463, w_033_3464, w_033_3467, w_033_3468, w_033_3469, w_033_3471, w_033_3472, w_033_3473, w_033_3474, w_033_3475, w_033_3477, w_033_3479, w_033_3480, w_033_3481, w_033_3482, w_033_3484, w_033_3485, w_033_3486, w_033_3487, w_033_3489, w_033_3490, w_033_3494, w_033_3495, w_033_3498, w_033_3499, w_033_3500, w_033_3502, w_033_3503, w_033_3504, w_033_3505, w_033_3509, w_033_3510, w_033_3513, w_033_3514, w_033_3515, w_033_3516, w_033_3519, w_033_3522, w_033_3523, w_033_3524, w_033_3525, w_033_3526, w_033_3527, w_033_3528, w_033_3529, w_033_3531, w_033_3532, w_033_3533, w_033_3535, w_033_3536, w_033_3537, w_033_3539, w_033_3540, w_033_3542, w_033_3543, w_033_3545, w_033_3546, w_033_3547, w_033_3549, w_033_3551, w_033_3554, w_033_3556, w_033_3557, w_033_3558, w_033_3560, w_033_3561, w_033_3562, w_033_3564, w_033_3566, w_033_3567, w_033_3568, w_033_3569, w_033_3570, w_033_3572, w_033_3574, w_033_3575, w_033_3576, w_033_3577, w_033_3578, w_033_3579, w_033_3580, w_033_3581, w_033_3582, w_033_3585, w_033_3586, w_033_3590, w_033_3591, w_033_3592, w_033_3593, w_033_3595, w_033_3596, w_033_3597, w_033_3598, w_033_3600, w_033_3603, w_033_3604, w_033_3606, w_033_3607, w_033_3608, w_033_3609, w_033_3610, w_033_3611, w_033_3612, w_033_3615, w_033_3617, w_033_3621, w_033_3625, w_033_3626, w_033_3627, w_033_3628, w_033_3629, w_033_3630, w_033_3631, w_033_3634, w_033_3635, w_033_3637, w_033_3638, w_033_3640, w_033_3641, w_033_3643, w_033_3644, w_033_3645, w_033_3646, w_033_3648, w_033_3649, w_033_3650, w_033_3651, w_033_3653, w_033_3654, w_033_3655, w_033_3659, w_033_3661, w_033_3662, w_033_3663, w_033_3666, w_033_3667, w_033_3669, w_033_3670, w_033_3671, w_033_3673, w_033_3676, w_033_3677, w_033_3678, w_033_3680, w_033_3684, w_033_3685, w_033_3687, w_033_3688, w_033_3691, w_033_3692, w_033_3693, w_033_3694, w_033_3698, w_033_3699, w_033_3700, w_033_3702, w_033_3703, w_033_3704, w_033_3705, w_033_3706, w_033_3709, w_033_3713, w_033_3717, w_033_3718, w_033_3719, w_033_3720, w_033_3721, w_033_3722, w_033_3723, w_033_3725, w_033_3728, w_033_3729, w_033_3730, w_033_3731, w_033_3733, w_033_3734, w_033_3736, w_033_3739, w_033_3740, w_033_3741, w_033_3743, w_033_3746, w_033_3747, w_033_3749, w_033_3750, w_033_3751, w_033_3753, w_033_3755, w_033_3756, w_033_3757, w_033_3758, w_033_3759, w_033_3760, w_033_3761, w_033_3763, w_033_3765, w_033_3766, w_033_3767, w_033_3768, w_033_3770, w_033_3773, w_033_3775, w_033_3776, w_033_3777, w_033_3781, w_033_3784, w_033_3785, w_033_3786, w_033_3787, w_033_3788, w_033_3789, w_033_3791, w_033_3792, w_033_3793, w_033_3794, w_033_3797, w_033_3799, w_033_3800, w_033_3802, w_033_3803, w_033_3804, w_033_3808, w_033_3809, w_033_3810, w_033_3811, w_033_3812, w_033_3813, w_033_3814, w_033_3815, w_033_3817, w_033_3818, w_033_3819, w_033_3820, w_033_3821, w_033_3822, w_033_3823, w_033_3824, w_033_3825, w_033_3829, w_033_3830, w_033_3831, w_033_3832, w_033_3834, w_033_3835, w_033_3836, w_033_3837, w_033_3838, w_033_3841, w_033_3843, w_033_3844, w_033_3845, w_033_3847, w_033_3848, w_033_3849, w_033_3850, w_033_3851, w_033_3852, w_033_3853, w_033_3863, w_033_3864, w_033_3866, w_033_3868, w_033_3871;
  wire w_034_000, w_034_001, w_034_002, w_034_003, w_034_004, w_034_005, w_034_006, w_034_007, w_034_008, w_034_009, w_034_010, w_034_011, w_034_012, w_034_013, w_034_014, w_034_015, w_034_016, w_034_017, w_034_018, w_034_019, w_034_020, w_034_021, w_034_022, w_034_023, w_034_024, w_034_025, w_034_026, w_034_027, w_034_028, w_034_029, w_034_030, w_034_031, w_034_032, w_034_033, w_034_034, w_034_035, w_034_036, w_034_037, w_034_038, w_034_039, w_034_040, w_034_041, w_034_042, w_034_043, w_034_044, w_034_045, w_034_046, w_034_047, w_034_048, w_034_049, w_034_050, w_034_051, w_034_052, w_034_053, w_034_054, w_034_055, w_034_056, w_034_057, w_034_058, w_034_059, w_034_060, w_034_061, w_034_062, w_034_063, w_034_064, w_034_065, w_034_066, w_034_067, w_034_068, w_034_069, w_034_070, w_034_071, w_034_072, w_034_073, w_034_074, w_034_075, w_034_076, w_034_077, w_034_078, w_034_079, w_034_080, w_034_081, w_034_082, w_034_083, w_034_084, w_034_085, w_034_086, w_034_087, w_034_088, w_034_089, w_034_090, w_034_091, w_034_092, w_034_093, w_034_094, w_034_095, w_034_096, w_034_097, w_034_098, w_034_099, w_034_100, w_034_101, w_034_102, w_034_103, w_034_104, w_034_105, w_034_106, w_034_107, w_034_108, w_034_109, w_034_110, w_034_111, w_034_112, w_034_113, w_034_114, w_034_116, w_034_117, w_034_118, w_034_119, w_034_120, w_034_121, w_034_122, w_034_123, w_034_124, w_034_125, w_034_126, w_034_127, w_034_128, w_034_129, w_034_130, w_034_131, w_034_132, w_034_133, w_034_134, w_034_135, w_034_136, w_034_137, w_034_138, w_034_139, w_034_140, w_034_141, w_034_142, w_034_143, w_034_144, w_034_145, w_034_146, w_034_147, w_034_148, w_034_149, w_034_150, w_034_151, w_034_152, w_034_153, w_034_154, w_034_155, w_034_156, w_034_157, w_034_158, w_034_159, w_034_160, w_034_161, w_034_162, w_034_163, w_034_164, w_034_165, w_034_166, w_034_167, w_034_168, w_034_169, w_034_170, w_034_171, w_034_172, w_034_173, w_034_174, w_034_175, w_034_176, w_034_177, w_034_178, w_034_180, w_034_181, w_034_182, w_034_183, w_034_184, w_034_185, w_034_186, w_034_187, w_034_188, w_034_189, w_034_190, w_034_191, w_034_192, w_034_193, w_034_194, w_034_195, w_034_196, w_034_197, w_034_198, w_034_199, w_034_200, w_034_201, w_034_202, w_034_203, w_034_204, w_034_205, w_034_206, w_034_207, w_034_208, w_034_209, w_034_210, w_034_211, w_034_212, w_034_213, w_034_214, w_034_215, w_034_216, w_034_217, w_034_218, w_034_219, w_034_220, w_034_221, w_034_222, w_034_223, w_034_224, w_034_225, w_034_226, w_034_227, w_034_228, w_034_229, w_034_230, w_034_231, w_034_232, w_034_233, w_034_234, w_034_235, w_034_236, w_034_237, w_034_238, w_034_239, w_034_240, w_034_241, w_034_242, w_034_243, w_034_244, w_034_245, w_034_247, w_034_248, w_034_249, w_034_250, w_034_251, w_034_252, w_034_253, w_034_254, w_034_255, w_034_256, w_034_257, w_034_258, w_034_259, w_034_260, w_034_261, w_034_262, w_034_263, w_034_264, w_034_265, w_034_266, w_034_267, w_034_268, w_034_269, w_034_270, w_034_271, w_034_272, w_034_273, w_034_274, w_034_275, w_034_276, w_034_277, w_034_278, w_034_279, w_034_280, w_034_281, w_034_282, w_034_283, w_034_284, w_034_285, w_034_286, w_034_287, w_034_288, w_034_289, w_034_290, w_034_291, w_034_292, w_034_293, w_034_294, w_034_295, w_034_296, w_034_297, w_034_298, w_034_299, w_034_300, w_034_301, w_034_302, w_034_303, w_034_304, w_034_305, w_034_306, w_034_307, w_034_308, w_034_309, w_034_310, w_034_311, w_034_312, w_034_313, w_034_314, w_034_315, w_034_316, w_034_317, w_034_318, w_034_319, w_034_320, w_034_321, w_034_322, w_034_323, w_034_324, w_034_325, w_034_326, w_034_327, w_034_328, w_034_329, w_034_330, w_034_331, w_034_332, w_034_333, w_034_334, w_034_335, w_034_336, w_034_338, w_034_339, w_034_341, w_034_342, w_034_343, w_034_344, w_034_345, w_034_346, w_034_347, w_034_348, w_034_349, w_034_350, w_034_351, w_034_352, w_034_353, w_034_354, w_034_355, w_034_356, w_034_357, w_034_358, w_034_359, w_034_360, w_034_361, w_034_362, w_034_363, w_034_364, w_034_365, w_034_366, w_034_368, w_034_369, w_034_370, w_034_371, w_034_373, w_034_374, w_034_375, w_034_376, w_034_377, w_034_378, w_034_379, w_034_380, w_034_381, w_034_382, w_034_383, w_034_384, w_034_385, w_034_386, w_034_387, w_034_388, w_034_389, w_034_390, w_034_391, w_034_392, w_034_393, w_034_394, w_034_395, w_034_396, w_034_397, w_034_398, w_034_399, w_034_400, w_034_401, w_034_402, w_034_403, w_034_404, w_034_405, w_034_406, w_034_407, w_034_408, w_034_409, w_034_410, w_034_411, w_034_412, w_034_413, w_034_414, w_034_415, w_034_416, w_034_417, w_034_418, w_034_419, w_034_420, w_034_421, w_034_422, w_034_423, w_034_424, w_034_425, w_034_426, w_034_427, w_034_428, w_034_429, w_034_430, w_034_431, w_034_432, w_034_433, w_034_434, w_034_435, w_034_436, w_034_437, w_034_438, w_034_439, w_034_440, w_034_441, w_034_442, w_034_443, w_034_444, w_034_446, w_034_447, w_034_448, w_034_449, w_034_450, w_034_451, w_034_452, w_034_453, w_034_455, w_034_456, w_034_457, w_034_458, w_034_459, w_034_460, w_034_461, w_034_462, w_034_463, w_034_464, w_034_465, w_034_466, w_034_467, w_034_468, w_034_469, w_034_470, w_034_471, w_034_472, w_034_473, w_034_474, w_034_475, w_034_476, w_034_477, w_034_478, w_034_479, w_034_480, w_034_481, w_034_482, w_034_483, w_034_484, w_034_485, w_034_486, w_034_487, w_034_488, w_034_489, w_034_490, w_034_491, w_034_492, w_034_493, w_034_494, w_034_495, w_034_496, w_034_497, w_034_498, w_034_499, w_034_500, w_034_501, w_034_502, w_034_503, w_034_504, w_034_505, w_034_506, w_034_507, w_034_508, w_034_509, w_034_510, w_034_511, w_034_512, w_034_513, w_034_514, w_034_515, w_034_516, w_034_517, w_034_518, w_034_519, w_034_520, w_034_521, w_034_522, w_034_523, w_034_524, w_034_525, w_034_526, w_034_527, w_034_528, w_034_529, w_034_530, w_034_531, w_034_532, w_034_533, w_034_534, w_034_535, w_034_536, w_034_537, w_034_538, w_034_539, w_034_540, w_034_541, w_034_542, w_034_544, w_034_545, w_034_546, w_034_548, w_034_549, w_034_550, w_034_551, w_034_552, w_034_553, w_034_554, w_034_555, w_034_556, w_034_557, w_034_558, w_034_559, w_034_560, w_034_561, w_034_562, w_034_563, w_034_564, w_034_565, w_034_566, w_034_567, w_034_568, w_034_569, w_034_570, w_034_571, w_034_572, w_034_573, w_034_574, w_034_575, w_034_576, w_034_577, w_034_578, w_034_579, w_034_580, w_034_581, w_034_582, w_034_583, w_034_584, w_034_585, w_034_586, w_034_587, w_034_588, w_034_589, w_034_590, w_034_591, w_034_592, w_034_593, w_034_594, w_034_595, w_034_596, w_034_597, w_034_598, w_034_599, w_034_600, w_034_602, w_034_603, w_034_604, w_034_605, w_034_606, w_034_607, w_034_608, w_034_609, w_034_611, w_034_612, w_034_613, w_034_614, w_034_616, w_034_617, w_034_618, w_034_619, w_034_620, w_034_621, w_034_622, w_034_623, w_034_624, w_034_625, w_034_626, w_034_627, w_034_628, w_034_629, w_034_630, w_034_631, w_034_632, w_034_633, w_034_634, w_034_635, w_034_636, w_034_637, w_034_638, w_034_639, w_034_640, w_034_641, w_034_642, w_034_643, w_034_644, w_034_645, w_034_646, w_034_647, w_034_648, w_034_649, w_034_650, w_034_651, w_034_652, w_034_653, w_034_654, w_034_655, w_034_656, w_034_657, w_034_658, w_034_659, w_034_661, w_034_662, w_034_663, w_034_664, w_034_665, w_034_666, w_034_667, w_034_668, w_034_669, w_034_670, w_034_671, w_034_672, w_034_673, w_034_674, w_034_675, w_034_676, w_034_677, w_034_678, w_034_679, w_034_680, w_034_681, w_034_682, w_034_683, w_034_684, w_034_685, w_034_686, w_034_687, w_034_688, w_034_689, w_034_690, w_034_691, w_034_692, w_034_693, w_034_694, w_034_696, w_034_697, w_034_698, w_034_699, w_034_700, w_034_701, w_034_702, w_034_703, w_034_705, w_034_706, w_034_707, w_034_709, w_034_710, w_034_711, w_034_712, w_034_713, w_034_714, w_034_715, w_034_716, w_034_717, w_034_718, w_034_719, w_034_720, w_034_721, w_034_722, w_034_723, w_034_724, w_034_725, w_034_726, w_034_727, w_034_728, w_034_729, w_034_730, w_034_731, w_034_733, w_034_734, w_034_735, w_034_736, w_034_737, w_034_739, w_034_740, w_034_741, w_034_742, w_034_743, w_034_744, w_034_745, w_034_746, w_034_747, w_034_748, w_034_750, w_034_752, w_034_753, w_034_755, w_034_756, w_034_757, w_034_758, w_034_760, w_034_762, w_034_764, w_034_765, w_034_766, w_034_767, w_034_768, w_034_769, w_034_770, w_034_771, w_034_773, w_034_774, w_034_775, w_034_777, w_034_778, w_034_779, w_034_781, w_034_782, w_034_783, w_034_784, w_034_785, w_034_787, w_034_788, w_034_789, w_034_790, w_034_791, w_034_792, w_034_793, w_034_794, w_034_795, w_034_796, w_034_797, w_034_798, w_034_799, w_034_800, w_034_801, w_034_802, w_034_803, w_034_804, w_034_805, w_034_806, w_034_807, w_034_808, w_034_809, w_034_810, w_034_811, w_034_812, w_034_813, w_034_814, w_034_815, w_034_816, w_034_817, w_034_818, w_034_819, w_034_820, w_034_821, w_034_822, w_034_823, w_034_824, w_034_825, w_034_826, w_034_827, w_034_828, w_034_829, w_034_830, w_034_831, w_034_832, w_034_833, w_034_834, w_034_835, w_034_836, w_034_837, w_034_838, w_034_839, w_034_840, w_034_842, w_034_843, w_034_844, w_034_845, w_034_846, w_034_847, w_034_848, w_034_849, w_034_850, w_034_851, w_034_852, w_034_853, w_034_854, w_034_855, w_034_856, w_034_857, w_034_858, w_034_860, w_034_861, w_034_862, w_034_863, w_034_864, w_034_865, w_034_866, w_034_867, w_034_868, w_034_869, w_034_870, w_034_871, w_034_872, w_034_873, w_034_875, w_034_876, w_034_877, w_034_878, w_034_879, w_034_880, w_034_881, w_034_882, w_034_883, w_034_884, w_034_885, w_034_886, w_034_887, w_034_888, w_034_889, w_034_890, w_034_891, w_034_892, w_034_893, w_034_894, w_034_895, w_034_896, w_034_897, w_034_898, w_034_899, w_034_900, w_034_901, w_034_902, w_034_903, w_034_905, w_034_906, w_034_907, w_034_908, w_034_909, w_034_910, w_034_911, w_034_912, w_034_913, w_034_914, w_034_915, w_034_916, w_034_917, w_034_918, w_034_919, w_034_921, w_034_922, w_034_923, w_034_924, w_034_925, w_034_926, w_034_927, w_034_928, w_034_929, w_034_931, w_034_932, w_034_933, w_034_934, w_034_935, w_034_936, w_034_937, w_034_938, w_034_939, w_034_940, w_034_941, w_034_942, w_034_943, w_034_944, w_034_945, w_034_946, w_034_947, w_034_948, w_034_949, w_034_950, w_034_951, w_034_952, w_034_953, w_034_954, w_034_955, w_034_956, w_034_957, w_034_958, w_034_959, w_034_960, w_034_961, w_034_962, w_034_963, w_034_964, w_034_965, w_034_966, w_034_967, w_034_968, w_034_969, w_034_970, w_034_971, w_034_972, w_034_973, w_034_974, w_034_977, w_034_978, w_034_979, w_034_980, w_034_981, w_034_982, w_034_983, w_034_984, w_034_985, w_034_986, w_034_987, w_034_988, w_034_989, w_034_990, w_034_991, w_034_992, w_034_993, w_034_994, w_034_996, w_034_998, w_034_999, w_034_1000, w_034_1001, w_034_1002, w_034_1003, w_034_1004, w_034_1005, w_034_1006, w_034_1008, w_034_1009, w_034_1010, w_034_1011, w_034_1012, w_034_1013, w_034_1014, w_034_1015, w_034_1016, w_034_1017, w_034_1018, w_034_1019, w_034_1020, w_034_1021, w_034_1023, w_034_1024, w_034_1025, w_034_1026, w_034_1027, w_034_1028, w_034_1029, w_034_1030, w_034_1031, w_034_1032, w_034_1033, w_034_1034, w_034_1035, w_034_1036, w_034_1037, w_034_1038, w_034_1039, w_034_1040, w_034_1041, w_034_1042, w_034_1043, w_034_1044, w_034_1045, w_034_1046, w_034_1047, w_034_1048, w_034_1049, w_034_1050, w_034_1051, w_034_1052, w_034_1053, w_034_1054, w_034_1055, w_034_1056, w_034_1057, w_034_1058, w_034_1059, w_034_1060, w_034_1063, w_034_1064, w_034_1065, w_034_1066, w_034_1067, w_034_1068, w_034_1069, w_034_1070, w_034_1071, w_034_1072, w_034_1073, w_034_1074, w_034_1075, w_034_1076, w_034_1077, w_034_1078, w_034_1079, w_034_1080, w_034_1081, w_034_1082, w_034_1083, w_034_1084, w_034_1085, w_034_1086, w_034_1087, w_034_1088, w_034_1089, w_034_1090, w_034_1091, w_034_1092, w_034_1093, w_034_1094, w_034_1095, w_034_1096, w_034_1097, w_034_1098, w_034_1099, w_034_1100, w_034_1101, w_034_1102, w_034_1104, w_034_1105, w_034_1106, w_034_1107, w_034_1108, w_034_1109, w_034_1110, w_034_1111, w_034_1112, w_034_1113, w_034_1114, w_034_1115, w_034_1116, w_034_1117, w_034_1118, w_034_1119, w_034_1120, w_034_1121, w_034_1122, w_034_1123, w_034_1124, w_034_1125, w_034_1126, w_034_1127, w_034_1128, w_034_1129, w_034_1130, w_034_1131, w_034_1132, w_034_1133, w_034_1134, w_034_1135, w_034_1137, w_034_1138, w_034_1139, w_034_1140, w_034_1141, w_034_1142, w_034_1143, w_034_1144, w_034_1145, w_034_1146, w_034_1147, w_034_1148, w_034_1149, w_034_1150, w_034_1151, w_034_1152, w_034_1153, w_034_1154, w_034_1155, w_034_1156, w_034_1157, w_034_1158, w_034_1159, w_034_1160, w_034_1161, w_034_1162, w_034_1163, w_034_1164, w_034_1165, w_034_1166, w_034_1167, w_034_1168, w_034_1169, w_034_1170, w_034_1171, w_034_1172, w_034_1173, w_034_1174, w_034_1175, w_034_1176, w_034_1177, w_034_1178, w_034_1179, w_034_1180, w_034_1181, w_034_1182, w_034_1183, w_034_1184, w_034_1185, w_034_1186, w_034_1187, w_034_1188, w_034_1189, w_034_1190, w_034_1191, w_034_1192, w_034_1193, w_034_1194, w_034_1195, w_034_1198, w_034_1199, w_034_1200, w_034_1202, w_034_1203, w_034_1204, w_034_1205, w_034_1207, w_034_1208, w_034_1211, w_034_1212, w_034_1213, w_034_1214, w_034_1215, w_034_1216, w_034_1217, w_034_1218, w_034_1219, w_034_1220, w_034_1221, w_034_1222, w_034_1223, w_034_1224, w_034_1225, w_034_1226, w_034_1227, w_034_1228, w_034_1229, w_034_1230, w_034_1231, w_034_1232, w_034_1233, w_034_1234, w_034_1235, w_034_1236, w_034_1237, w_034_1238, w_034_1239, w_034_1240, w_034_1241, w_034_1242, w_034_1243, w_034_1244, w_034_1245, w_034_1247, w_034_1249, w_034_1250, w_034_1251, w_034_1252, w_034_1253, w_034_1254, w_034_1255, w_034_1257, w_034_1258, w_034_1259, w_034_1260, w_034_1261, w_034_1262, w_034_1263, w_034_1264, w_034_1265, w_034_1266, w_034_1267, w_034_1268, w_034_1269, w_034_1270, w_034_1271, w_034_1272, w_034_1273, w_034_1274, w_034_1275, w_034_1276, w_034_1277, w_034_1278, w_034_1279, w_034_1280, w_034_1281, w_034_1282, w_034_1283, w_034_1284, w_034_1285, w_034_1286, w_034_1287, w_034_1288, w_034_1289, w_034_1290, w_034_1291, w_034_1292, w_034_1293, w_034_1294, w_034_1295, w_034_1296, w_034_1297, w_034_1298, w_034_1299, w_034_1300, w_034_1301, w_034_1302, w_034_1304, w_034_1305, w_034_1306, w_034_1307, w_034_1308, w_034_1309, w_034_1310, w_034_1311, w_034_1312, w_034_1314, w_034_1315, w_034_1316, w_034_1317, w_034_1318, w_034_1319, w_034_1320, w_034_1321, w_034_1322, w_034_1323, w_034_1324, w_034_1325, w_034_1326, w_034_1327, w_034_1328, w_034_1329, w_034_1330, w_034_1331, w_034_1332, w_034_1333, w_034_1334, w_034_1335, w_034_1336, w_034_1338, w_034_1339, w_034_1340, w_034_1341, w_034_1342, w_034_1343, w_034_1344, w_034_1345, w_034_1346, w_034_1347, w_034_1348, w_034_1349, w_034_1350, w_034_1351, w_034_1352, w_034_1353, w_034_1354, w_034_1355, w_034_1356, w_034_1357, w_034_1359, w_034_1360, w_034_1361, w_034_1362, w_034_1363, w_034_1364, w_034_1366, w_034_1368, w_034_1369, w_034_1370, w_034_1371, w_034_1372, w_034_1373, w_034_1374, w_034_1376, w_034_1377, w_034_1378, w_034_1379, w_034_1380, w_034_1381, w_034_1382, w_034_1383, w_034_1384, w_034_1386, w_034_1387, w_034_1388, w_034_1389, w_034_1390, w_034_1391, w_034_1394, w_034_1395, w_034_1396, w_034_1397, w_034_1398, w_034_1400, w_034_1402, w_034_1403, w_034_1404, w_034_1405, w_034_1407, w_034_1408, w_034_1409, w_034_1410, w_034_1411, w_034_1412, w_034_1413, w_034_1414, w_034_1415, w_034_1416, w_034_1417, w_034_1418, w_034_1419, w_034_1420, w_034_1421, w_034_1422, w_034_1423, w_034_1424, w_034_1425, w_034_1426, w_034_1427, w_034_1428, w_034_1429, w_034_1430, w_034_1432, w_034_1433, w_034_1434, w_034_1435, w_034_1436, w_034_1437, w_034_1438, w_034_1439, w_034_1441, w_034_1442, w_034_1443, w_034_1444, w_034_1445, w_034_1446;
  wire w_035_000, w_035_002, w_035_003, w_035_004, w_035_005, w_035_006, w_035_007, w_035_008, w_035_009, w_035_010, w_035_011, w_035_012, w_035_014, w_035_015, w_035_016, w_035_017, w_035_018, w_035_020, w_035_021, w_035_023, w_035_024, w_035_025, w_035_026, w_035_027, w_035_028, w_035_029, w_035_030, w_035_031, w_035_032, w_035_033, w_035_034, w_035_035, w_035_038, w_035_039, w_035_040, w_035_041, w_035_043, w_035_044, w_035_045, w_035_046, w_035_047, w_035_048, w_035_049, w_035_051, w_035_052, w_035_054, w_035_055, w_035_056, w_035_058, w_035_059, w_035_060, w_035_061, w_035_062, w_035_063, w_035_064, w_035_066, w_035_067, w_035_068, w_035_069, w_035_070, w_035_072, w_035_073, w_035_075, w_035_076, w_035_077, w_035_078, w_035_079, w_035_080, w_035_081, w_035_082, w_035_084, w_035_085, w_035_086, w_035_087, w_035_088, w_035_090, w_035_091, w_035_092, w_035_093, w_035_094, w_035_095, w_035_096, w_035_097, w_035_098, w_035_099, w_035_100, w_035_101, w_035_103, w_035_104, w_035_105, w_035_106, w_035_107, w_035_109, w_035_111, w_035_112, w_035_113, w_035_114, w_035_115, w_035_116, w_035_117, w_035_118, w_035_119, w_035_120, w_035_121, w_035_122, w_035_123, w_035_124, w_035_125, w_035_126, w_035_128, w_035_130, w_035_131, w_035_132, w_035_133, w_035_134, w_035_135, w_035_136, w_035_137, w_035_138, w_035_139, w_035_141, w_035_143, w_035_144, w_035_146, w_035_147, w_035_148, w_035_150, w_035_151, w_035_152, w_035_153, w_035_154, w_035_155, w_035_156, w_035_157, w_035_158, w_035_159, w_035_160, w_035_162, w_035_163, w_035_164, w_035_166, w_035_167, w_035_168, w_035_169, w_035_170, w_035_171, w_035_172, w_035_174, w_035_175, w_035_176, w_035_177, w_035_178, w_035_179, w_035_180, w_035_181, w_035_182, w_035_184, w_035_185, w_035_186, w_035_187, w_035_189, w_035_191, w_035_193, w_035_194, w_035_195, w_035_196, w_035_197, w_035_198, w_035_199, w_035_200, w_035_201, w_035_204, w_035_205, w_035_206, w_035_208, w_035_209, w_035_210, w_035_212, w_035_213, w_035_216, w_035_217, w_035_218, w_035_219, w_035_220, w_035_221, w_035_222, w_035_224, w_035_225, w_035_226, w_035_227, w_035_228, w_035_229, w_035_230, w_035_231, w_035_232, w_035_235, w_035_236, w_035_238, w_035_239, w_035_240, w_035_241, w_035_242, w_035_243, w_035_244, w_035_245, w_035_246, w_035_249, w_035_250, w_035_251, w_035_252, w_035_253, w_035_254, w_035_255, w_035_256, w_035_257, w_035_258, w_035_259, w_035_260, w_035_261, w_035_262, w_035_263, w_035_264, w_035_265, w_035_266, w_035_267, w_035_268, w_035_269, w_035_270, w_035_271, w_035_272, w_035_273, w_035_274, w_035_275, w_035_276, w_035_277, w_035_278, w_035_279, w_035_281, w_035_282, w_035_283, w_035_284, w_035_286, w_035_287, w_035_289, w_035_291, w_035_292, w_035_293, w_035_294, w_035_295, w_035_296, w_035_297, w_035_298, w_035_299, w_035_300, w_035_301, w_035_302, w_035_303, w_035_304, w_035_305, w_035_306, w_035_307, w_035_308, w_035_309, w_035_310, w_035_311, w_035_312, w_035_313, w_035_314, w_035_315, w_035_316, w_035_319, w_035_320, w_035_321, w_035_322, w_035_324, w_035_325, w_035_326, w_035_327, w_035_328, w_035_329, w_035_330, w_035_331, w_035_332, w_035_333, w_035_334, w_035_335, w_035_336, w_035_337, w_035_338, w_035_339, w_035_340, w_035_341, w_035_342, w_035_343, w_035_344, w_035_345, w_035_346, w_035_347, w_035_348, w_035_349, w_035_350, w_035_351, w_035_352, w_035_354, w_035_355, w_035_356, w_035_357, w_035_358, w_035_360, w_035_361, w_035_362, w_035_363, w_035_364, w_035_366, w_035_367, w_035_369, w_035_371, w_035_372, w_035_373, w_035_374, w_035_375, w_035_376, w_035_377, w_035_378, w_035_379, w_035_380, w_035_381, w_035_383, w_035_384, w_035_385, w_035_386, w_035_387, w_035_388, w_035_389, w_035_391, w_035_392, w_035_393, w_035_394, w_035_395, w_035_396, w_035_397, w_035_398, w_035_399, w_035_400, w_035_401, w_035_402, w_035_403, w_035_404, w_035_405, w_035_406, w_035_407, w_035_408, w_035_410, w_035_412, w_035_414, w_035_415, w_035_416, w_035_417, w_035_418, w_035_419, w_035_420, w_035_421, w_035_422, w_035_424, w_035_425, w_035_426, w_035_427, w_035_428, w_035_429, w_035_430, w_035_431, w_035_432, w_035_433, w_035_434, w_035_435, w_035_437, w_035_438, w_035_439, w_035_441, w_035_442, w_035_444, w_035_445, w_035_446, w_035_448, w_035_450, w_035_451, w_035_452, w_035_454, w_035_455, w_035_457, w_035_458, w_035_459, w_035_460, w_035_461, w_035_462, w_035_463, w_035_464, w_035_465, w_035_466, w_035_467, w_035_468, w_035_469, w_035_470, w_035_471, w_035_473, w_035_474, w_035_476, w_035_477, w_035_479, w_035_480, w_035_481, w_035_482, w_035_483, w_035_484, w_035_485, w_035_486, w_035_488, w_035_489, w_035_490, w_035_491, w_035_492, w_035_493, w_035_494, w_035_495, w_035_496, w_035_498, w_035_499, w_035_500, w_035_502, w_035_503, w_035_504, w_035_507, w_035_508, w_035_509, w_035_510, w_035_511, w_035_512, w_035_514, w_035_515, w_035_516, w_035_517, w_035_518, w_035_520, w_035_521, w_035_522, w_035_523, w_035_524, w_035_525, w_035_527, w_035_528, w_035_529, w_035_530, w_035_531, w_035_533, w_035_534, w_035_536, w_035_538, w_035_539, w_035_540, w_035_542, w_035_543, w_035_544, w_035_545, w_035_546, w_035_547, w_035_548, w_035_549, w_035_550, w_035_551, w_035_552, w_035_553, w_035_554, w_035_556, w_035_557, w_035_558, w_035_559, w_035_560, w_035_561, w_035_562, w_035_563, w_035_564, w_035_565, w_035_566, w_035_567, w_035_568, w_035_569, w_035_570, w_035_571, w_035_572, w_035_573, w_035_574, w_035_575, w_035_576, w_035_577, w_035_578, w_035_579, w_035_580, w_035_581, w_035_582, w_035_583, w_035_584, w_035_585, w_035_586, w_035_587, w_035_589, w_035_590, w_035_591, w_035_592, w_035_593, w_035_594, w_035_595, w_035_596, w_035_597, w_035_598, w_035_599, w_035_600, w_035_601, w_035_602, w_035_603, w_035_604, w_035_605, w_035_607, w_035_608, w_035_609, w_035_610, w_035_611, w_035_612, w_035_613, w_035_614, w_035_615, w_035_616, w_035_617, w_035_618, w_035_619, w_035_620, w_035_621, w_035_622, w_035_623, w_035_624, w_035_625, w_035_626, w_035_627, w_035_628, w_035_629, w_035_630, w_035_631, w_035_632, w_035_633, w_035_634, w_035_635, w_035_636, w_035_637, w_035_638, w_035_639, w_035_641, w_035_642, w_035_643, w_035_644, w_035_645, w_035_646, w_035_648, w_035_650, w_035_651, w_035_653, w_035_654, w_035_655, w_035_657, w_035_661, w_035_662, w_035_663, w_035_664, w_035_665, w_035_666, w_035_667, w_035_668, w_035_669, w_035_670, w_035_673, w_035_674, w_035_675, w_035_676, w_035_677, w_035_680, w_035_681, w_035_682, w_035_684, w_035_687, w_035_688, w_035_689, w_035_690, w_035_692, w_035_693, w_035_694, w_035_695, w_035_696, w_035_697, w_035_698, w_035_699, w_035_700, w_035_701, w_035_702, w_035_703, w_035_704, w_035_705, w_035_706, w_035_708, w_035_709, w_035_710, w_035_711, w_035_712, w_035_713, w_035_714, w_035_715, w_035_716, w_035_717, w_035_718, w_035_719, w_035_720, w_035_721, w_035_722, w_035_723, w_035_724, w_035_727, w_035_728, w_035_729, w_035_731, w_035_733, w_035_734, w_035_737, w_035_738, w_035_739, w_035_740, w_035_741, w_035_742, w_035_743, w_035_744, w_035_745, w_035_746, w_035_747, w_035_748, w_035_752, w_035_753, w_035_754, w_035_755, w_035_756, w_035_757, w_035_758, w_035_759, w_035_760, w_035_761, w_035_763, w_035_765, w_035_766, w_035_767, w_035_768, w_035_769, w_035_770, w_035_772, w_035_773, w_035_774, w_035_775, w_035_776, w_035_778, w_035_779, w_035_780, w_035_781, w_035_782, w_035_783, w_035_784, w_035_786, w_035_787, w_035_788, w_035_789, w_035_790, w_035_791, w_035_792, w_035_794, w_035_795, w_035_796, w_035_799, w_035_801, w_035_803, w_035_805, w_035_806, w_035_808, w_035_809, w_035_810, w_035_811, w_035_813, w_035_814, w_035_815, w_035_816, w_035_817, w_035_818, w_035_820, w_035_821, w_035_822, w_035_823, w_035_824, w_035_825, w_035_826, w_035_827, w_035_829, w_035_832, w_035_833, w_035_834, w_035_835, w_035_836, w_035_838, w_035_839, w_035_840, w_035_841, w_035_842, w_035_844, w_035_845, w_035_846, w_035_847, w_035_848, w_035_849, w_035_850, w_035_851, w_035_852, w_035_853, w_035_854, w_035_855, w_035_856, w_035_857, w_035_858, w_035_859, w_035_860, w_035_861, w_035_862, w_035_863, w_035_864, w_035_866, w_035_867, w_035_868, w_035_869, w_035_870, w_035_871, w_035_872, w_035_873, w_035_874, w_035_875, w_035_876, w_035_878, w_035_879, w_035_880, w_035_882, w_035_883, w_035_884, w_035_885, w_035_886, w_035_887, w_035_888, w_035_889, w_035_890, w_035_891, w_035_892, w_035_893, w_035_894, w_035_895, w_035_896, w_035_898, w_035_899, w_035_901, w_035_902, w_035_903, w_035_904, w_035_906, w_035_907, w_035_908, w_035_909, w_035_910, w_035_911, w_035_912, w_035_914, w_035_915, w_035_916, w_035_918, w_035_919, w_035_920, w_035_921, w_035_922, w_035_923, w_035_924, w_035_925, w_035_926, w_035_927, w_035_928, w_035_929, w_035_930, w_035_931, w_035_932, w_035_933, w_035_934, w_035_940, w_035_941, w_035_942, w_035_944, w_035_945, w_035_946, w_035_947, w_035_948, w_035_950, w_035_952, w_035_953, w_035_954, w_035_955, w_035_956, w_035_957, w_035_958, w_035_960, w_035_961, w_035_962, w_035_963, w_035_964, w_035_965, w_035_967, w_035_968, w_035_969, w_035_970, w_035_974, w_035_975, w_035_976, w_035_984, w_035_985, w_035_986, w_035_987, w_035_989, w_035_990, w_035_991, w_035_993, w_035_994, w_035_996, w_035_997, w_035_998, w_035_1000, w_035_1001, w_035_1003, w_035_1006, w_035_1007, w_035_1008, w_035_1010, w_035_1014, w_035_1016, w_035_1018, w_035_1019, w_035_1020, w_035_1021, w_035_1022, w_035_1023, w_035_1027, w_035_1028, w_035_1030, w_035_1031, w_035_1034, w_035_1038, w_035_1040, w_035_1044, w_035_1045, w_035_1046, w_035_1047, w_035_1048, w_035_1049, w_035_1051, w_035_1053, w_035_1054, w_035_1055, w_035_1056, w_035_1057, w_035_1058, w_035_1059, w_035_1061, w_035_1062, w_035_1063, w_035_1065, w_035_1068, w_035_1069, w_035_1071, w_035_1072, w_035_1073, w_035_1075, w_035_1076, w_035_1077, w_035_1079, w_035_1081, w_035_1084, w_035_1086, w_035_1090, w_035_1094, w_035_1095, w_035_1096, w_035_1097, w_035_1098, w_035_1099, w_035_1100, w_035_1101, w_035_1102, w_035_1103, w_035_1104, w_035_1105, w_035_1106, w_035_1110, w_035_1111, w_035_1114, w_035_1115, w_035_1116, w_035_1117, w_035_1118, w_035_1119, w_035_1120, w_035_1121, w_035_1122, w_035_1124, w_035_1127, w_035_1129, w_035_1130, w_035_1131, w_035_1133, w_035_1134, w_035_1135, w_035_1139, w_035_1140, w_035_1141, w_035_1142, w_035_1143, w_035_1144, w_035_1146, w_035_1147, w_035_1149, w_035_1150, w_035_1151, w_035_1152, w_035_1153, w_035_1157, w_035_1158, w_035_1160, w_035_1161, w_035_1163, w_035_1166, w_035_1167, w_035_1168, w_035_1173, w_035_1174, w_035_1177, w_035_1181, w_035_1184, w_035_1185, w_035_1186, w_035_1189, w_035_1192, w_035_1195, w_035_1196, w_035_1197, w_035_1199, w_035_1200, w_035_1201, w_035_1202, w_035_1203, w_035_1205, w_035_1207, w_035_1211, w_035_1212, w_035_1215, w_035_1216, w_035_1218, w_035_1219, w_035_1222, w_035_1224, w_035_1226, w_035_1227, w_035_1228, w_035_1229, w_035_1230, w_035_1231, w_035_1234, w_035_1237, w_035_1241, w_035_1242, w_035_1243, w_035_1244, w_035_1245, w_035_1246, w_035_1248, w_035_1249, w_035_1250, w_035_1251, w_035_1252, w_035_1253, w_035_1254, w_035_1255, w_035_1256, w_035_1257, w_035_1260, w_035_1262, w_035_1263, w_035_1264, w_035_1265, w_035_1266, w_035_1267, w_035_1270, w_035_1271, w_035_1272, w_035_1273, w_035_1275, w_035_1276, w_035_1277, w_035_1278, w_035_1279, w_035_1280, w_035_1281, w_035_1283, w_035_1286, w_035_1287, w_035_1289, w_035_1292, w_035_1293, w_035_1295, w_035_1298, w_035_1302, w_035_1303, w_035_1304, w_035_1306, w_035_1308, w_035_1309, w_035_1314, w_035_1316, w_035_1317, w_035_1318, w_035_1319, w_035_1320, w_035_1321, w_035_1324, w_035_1326, w_035_1327, w_035_1329, w_035_1330, w_035_1333, w_035_1334, w_035_1337, w_035_1338, w_035_1340, w_035_1341, w_035_1342, w_035_1343, w_035_1344, w_035_1346, w_035_1347, w_035_1349, w_035_1350, w_035_1352, w_035_1353, w_035_1359, w_035_1360, w_035_1363, w_035_1364, w_035_1367, w_035_1369, w_035_1370, w_035_1371, w_035_1373, w_035_1375, w_035_1376, w_035_1378, w_035_1379, w_035_1380, w_035_1382, w_035_1383, w_035_1385, w_035_1386, w_035_1388, w_035_1389, w_035_1390, w_035_1391, w_035_1392, w_035_1393, w_035_1394, w_035_1395, w_035_1396, w_035_1400, w_035_1401, w_035_1402, w_035_1404, w_035_1405, w_035_1406, w_035_1407, w_035_1409, w_035_1410, w_035_1412, w_035_1413, w_035_1414, w_035_1416, w_035_1418, w_035_1420, w_035_1421, w_035_1422, w_035_1424, w_035_1425, w_035_1427, w_035_1428, w_035_1432, w_035_1433, w_035_1435, w_035_1436, w_035_1437, w_035_1438, w_035_1440, w_035_1443, w_035_1444, w_035_1445, w_035_1446, w_035_1447, w_035_1448, w_035_1449, w_035_1450, w_035_1451, w_035_1452, w_035_1454, w_035_1455, w_035_1457, w_035_1458, w_035_1459, w_035_1460, w_035_1461, w_035_1462, w_035_1464, w_035_1465, w_035_1466, w_035_1467, w_035_1469, w_035_1470, w_035_1471, w_035_1472, w_035_1474, w_035_1478, w_035_1480, w_035_1481, w_035_1482, w_035_1483, w_035_1484, w_035_1486, w_035_1489, w_035_1490, w_035_1491, w_035_1492, w_035_1493, w_035_1496, w_035_1498, w_035_1499, w_035_1500, w_035_1501, w_035_1502, w_035_1503, w_035_1504, w_035_1507, w_035_1508, w_035_1509, w_035_1511, w_035_1512, w_035_1514, w_035_1515, w_035_1516, w_035_1519, w_035_1520, w_035_1524, w_035_1526, w_035_1527, w_035_1528, w_035_1529, w_035_1530, w_035_1531, w_035_1532, w_035_1533, w_035_1534, w_035_1535, w_035_1536, w_035_1537, w_035_1538, w_035_1540, w_035_1542, w_035_1543, w_035_1545, w_035_1546, w_035_1547, w_035_1548, w_035_1549, w_035_1550, w_035_1551, w_035_1552, w_035_1554, w_035_1556, w_035_1557, w_035_1558, w_035_1559, w_035_1560, w_035_1561, w_035_1564, w_035_1566, w_035_1567, w_035_1569, w_035_1570, w_035_1572, w_035_1574, w_035_1575, w_035_1576, w_035_1580, w_035_1581, w_035_1582, w_035_1584, w_035_1585, w_035_1586, w_035_1587, w_035_1588, w_035_1589, w_035_1591, w_035_1592, w_035_1597, w_035_1598, w_035_1599, w_035_1600, w_035_1601, w_035_1602, w_035_1603, w_035_1607, w_035_1608, w_035_1609, w_035_1610, w_035_1613, w_035_1614, w_035_1618, w_035_1620, w_035_1621, w_035_1622, w_035_1623, w_035_1625, w_035_1626, w_035_1627, w_035_1629, w_035_1630, w_035_1631, w_035_1632, w_035_1635, w_035_1639, w_035_1641, w_035_1643, w_035_1644, w_035_1645, w_035_1646, w_035_1647, w_035_1648, w_035_1649, w_035_1650, w_035_1651, w_035_1653, w_035_1655, w_035_1657, w_035_1658, w_035_1659, w_035_1660, w_035_1661, w_035_1662, w_035_1663, w_035_1664, w_035_1666, w_035_1667, w_035_1668, w_035_1671, w_035_1672, w_035_1675, w_035_1676, w_035_1677, w_035_1680, w_035_1681, w_035_1682, w_035_1685, w_035_1686, w_035_1688, w_035_1689, w_035_1690, w_035_1692, w_035_1693, w_035_1694, w_035_1695, w_035_1696, w_035_1700, w_035_1701, w_035_1703, w_035_1706, w_035_1707, w_035_1708, w_035_1710, w_035_1713, w_035_1714, w_035_1716, w_035_1719, w_035_1720, w_035_1722, w_035_1728, w_035_1729, w_035_1730, w_035_1732, w_035_1733, w_035_1735, w_035_1740, w_035_1741, w_035_1742, w_035_1749, w_035_1750, w_035_1751, w_035_1752, w_035_1753, w_035_1754, w_035_1758, w_035_1759, w_035_1760, w_035_1761, w_035_1762, w_035_1763, w_035_1764, w_035_1765, w_035_1766, w_035_1767, w_035_1768, w_035_1769, w_035_1771, w_035_1772, w_035_1774, w_035_1775, w_035_1777, w_035_1778, w_035_1779, w_035_1781, w_035_1782, w_035_1785, w_035_1787, w_035_1789, w_035_1791, w_035_1792, w_035_1794, w_035_1795, w_035_1797, w_035_1798, w_035_1800, w_035_1801, w_035_1802, w_035_1803, w_035_1804, w_035_1805, w_035_1806, w_035_1807, w_035_1809, w_035_1810, w_035_1811, w_035_1813, w_035_1814, w_035_1816, w_035_1824, w_035_1825, w_035_1827, w_035_1828, w_035_1831, w_035_1833, w_035_1835, w_035_1836, w_035_1838, w_035_1840, w_035_1842, w_035_1843, w_035_1844, w_035_1846, w_035_1849, w_035_1850, w_035_1852, w_035_1853, w_035_1854, w_035_1855, w_035_1856, w_035_1857, w_035_1858, w_035_1859, w_035_1860, w_035_1862, w_035_1863, w_035_1867, w_035_1868, w_035_1874, w_035_1875, w_035_1879, w_035_1880, w_035_1883, w_035_1884, w_035_1885, w_035_1887, w_035_1890, w_035_1891, w_035_1892, w_035_1895, w_035_1896, w_035_1900, w_035_1901, w_035_1902, w_035_1903, w_035_1904, w_035_1906, w_035_1907, w_035_1908, w_035_1909, w_035_1910, w_035_1912, w_035_1917, w_035_1922, w_035_1926, w_035_1929, w_035_1930, w_035_1931, w_035_1933, w_035_1934, w_035_1935, w_035_1936, w_035_1937, w_035_1939, w_035_1940, w_035_1941, w_035_1942, w_035_1943, w_035_1946, w_035_1947, w_035_1948, w_035_1949, w_035_1950, w_035_1951, w_035_1952, w_035_1954, w_035_1958, w_035_1959, w_035_1961, w_035_1966, w_035_1968, w_035_1969, w_035_1970, w_035_1976, w_035_1977, w_035_1978, w_035_1979, w_035_1981, w_035_1982, w_035_1984, w_035_1988, w_035_1989, w_035_1991, w_035_1993, w_035_1999, w_035_2000, w_035_2002, w_035_2003, w_035_2005, w_035_2006, w_035_2008, w_035_2009, w_035_2010, w_035_2011, w_035_2012, w_035_2013, w_035_2015, w_035_2016, w_035_2017, w_035_2018, w_035_2021, w_035_2024, w_035_2025, w_035_2029, w_035_2031, w_035_2032, w_035_2033, w_035_2034, w_035_2036, w_035_2039, w_035_2045, w_035_2046, w_035_2047, w_035_2048, w_035_2053, w_035_2054, w_035_2055, w_035_2056, w_035_2059, w_035_2062, w_035_2064, w_035_2066, w_035_2068, w_035_2070, w_035_2071, w_035_2072, w_035_2073, w_035_2074, w_035_2075, w_035_2076, w_035_2080, w_035_2082, w_035_2083, w_035_2085, w_035_2087, w_035_2088, w_035_2090, w_035_2092, w_035_2093, w_035_2095, w_035_2096, w_035_2097, w_035_2098, w_035_2099, w_035_2100, w_035_2101, w_035_2102, w_035_2103, w_035_2104, w_035_2106, w_035_2107, w_035_2110, w_035_2113, w_035_2114, w_035_2115, w_035_2116, w_035_2117, w_035_2118, w_035_2120, w_035_2122, w_035_2123, w_035_2125, w_035_2127, w_035_2130, w_035_2131, w_035_2134, w_035_2136, w_035_2139, w_035_2140, w_035_2142, w_035_2145, w_035_2146, w_035_2147, w_035_2148, w_035_2149, w_035_2150, w_035_2151, w_035_2152, w_035_2154, w_035_2155, w_035_2156, w_035_2159, w_035_2160, w_035_2161, w_035_2163, w_035_2164, w_035_2167, w_035_2169, w_035_2170, w_035_2172, w_035_2173, w_035_2175, w_035_2176, w_035_2177, w_035_2180, w_035_2181, w_035_2182, w_035_2183, w_035_2184, w_035_2186, w_035_2187, w_035_2188, w_035_2191, w_035_2192, w_035_2195, w_035_2199, w_035_2200, w_035_2201, w_035_2202, w_035_2205, w_035_2206, w_035_2208, w_035_2214, w_035_2216, w_035_2217, w_035_2218, w_035_2219, w_035_2221, w_035_2224, w_035_2227, w_035_2228, w_035_2229, w_035_2230, w_035_2231, w_035_2233, w_035_2234, w_035_2236, w_035_2242, w_035_2245, w_035_2248, w_035_2249, w_035_2250, w_035_2251, w_035_2252, w_035_2253, w_035_2254, w_035_2255, w_035_2256, w_035_2257, w_035_2258, w_035_2260, w_035_2264, w_035_2265, w_035_2266, w_035_2267, w_035_2268, w_035_2269, w_035_2270, w_035_2272, w_035_2273, w_035_2275, w_035_2276, w_035_2277, w_035_2278, w_035_2281, w_035_2283, w_035_2284, w_035_2286, w_035_2287, w_035_2290, w_035_2295, w_035_2297, w_035_2298, w_035_2300, w_035_2301, w_035_2302, w_035_2303, w_035_2304, w_035_2306, w_035_2307, w_035_2308, w_035_2309, w_035_2310, w_035_2312, w_035_2313, w_035_2314, w_035_2315, w_035_2316, w_035_2318, w_035_2319, w_035_2320, w_035_2324, w_035_2326, w_035_2328, w_035_2329, w_035_2330, w_035_2331, w_035_2332, w_035_2334, w_035_2335, w_035_2336, w_035_2339, w_035_2342, w_035_2344, w_035_2346, w_035_2347, w_035_2349, w_035_2351, w_035_2352, w_035_2356, w_035_2358, w_035_2359, w_035_2360, w_035_2361, w_035_2362, w_035_2363, w_035_2364, w_035_2366, w_035_2368, w_035_2369, w_035_2370, w_035_2371, w_035_2372, w_035_2373, w_035_2375, w_035_2376, w_035_2379, w_035_2381, w_035_2382, w_035_2384, w_035_2385, w_035_2386, w_035_2388, w_035_2389, w_035_2390, w_035_2391, w_035_2393, w_035_2394, w_035_2395, w_035_2402, w_035_2404, w_035_2405, w_035_2406, w_035_2407, w_035_2414, w_035_2415, w_035_2416, w_035_2417, w_035_2418, w_035_2419, w_035_2420, w_035_2425, w_035_2426, w_035_2427, w_035_2431, w_035_2433, w_035_2434, w_035_2436, w_035_2437, w_035_2438, w_035_2439, w_035_2441, w_035_2444, w_035_2447, w_035_2448, w_035_2449, w_035_2450, w_035_2451, w_035_2452, w_035_2453, w_035_2454, w_035_2455, w_035_2456, w_035_2459, w_035_2460, w_035_2462, w_035_2463, w_035_2464, w_035_2465, w_035_2471, w_035_2475, w_035_2476, w_035_2478, w_035_2479, w_035_2481, w_035_2482, w_035_2483, w_035_2485, w_035_2486, w_035_2488, w_035_2490, w_035_2491, w_035_2494, w_035_2495, w_035_2497, w_035_2498, w_035_2499, w_035_2500, w_035_2501, w_035_2504, w_035_2505, w_035_2507, w_035_2511, w_035_2513, w_035_2516, w_035_2518, w_035_2519, w_035_2520, w_035_2521, w_035_2522, w_035_2524, w_035_2526, w_035_2532, w_035_2536, w_035_2539, w_035_2541, w_035_2542, w_035_2543, w_035_2545, w_035_2546, w_035_2547, w_035_2548, w_035_2549, w_035_2550, w_035_2553, w_035_2555, w_035_2557, w_035_2559, w_035_2562, w_035_2564, w_035_2565, w_035_2566, w_035_2567, w_035_2569, w_035_2571, w_035_2572, w_035_2574, w_035_2576, w_035_2577, w_035_2578, w_035_2579, w_035_2580, w_035_2581, w_035_2582, w_035_2583, w_035_2585, w_035_2587, w_035_2589, w_035_2590, w_035_2591, w_035_2592, w_035_2593, w_035_2596, w_035_2599, w_035_2600, w_035_2602, w_035_2604, w_035_2606, w_035_2607, w_035_2609, w_035_2610, w_035_2612, w_035_2613, w_035_2614, w_035_2617, w_035_2618, w_035_2620, w_035_2621, w_035_2622, w_035_2624, w_035_2625, w_035_2627, w_035_2628, w_035_2629, w_035_2630, w_035_2633, w_035_2635, w_035_2637, w_035_2638, w_035_2639, w_035_2640, w_035_2641, w_035_2643, w_035_2644, w_035_2645, w_035_2646, w_035_2647, w_035_2648, w_035_2649, w_035_2651, w_035_2653, w_035_2654, w_035_2655, w_035_2659, w_035_2660, w_035_2661, w_035_2663, w_035_2664, w_035_2666, w_035_2667, w_035_2669, w_035_2672, w_035_2674, w_035_2677, w_035_2680, w_035_2681, w_035_2683, w_035_2686, w_035_2688, w_035_2689, w_035_2690, w_035_2696, w_035_2697, w_035_2698, w_035_2700, w_035_2703, w_035_2705, w_035_2706, w_035_2707, w_035_2709, w_035_2710, w_035_2712, w_035_2713, w_035_2714, w_035_2716, w_035_2717, w_035_2720, w_035_2721, w_035_2722, w_035_2724, w_035_2725, w_035_2726, w_035_2727, w_035_2732, w_035_2733, w_035_2735, w_035_2737, w_035_2738, w_035_2740, w_035_2741, w_035_2742, w_035_2744, w_035_2745, w_035_2747, w_035_2751, w_035_2752, w_035_2753, w_035_2754, w_035_2755, w_035_2757, w_035_2758, w_035_2759, w_035_2763, w_035_2765, w_035_2768, w_035_2770, w_035_2776, w_035_2777, w_035_2779, w_035_2780, w_035_2782, w_035_2784, w_035_2786, w_035_2787, w_035_2789, w_035_2790, w_035_2791, w_035_2792, w_035_2794, w_035_2795, w_035_2796, w_035_2797, w_035_2799, w_035_2801, w_035_2803, w_035_2804, w_035_2805, w_035_2806, w_035_2808, w_035_2809, w_035_2814, w_035_2815, w_035_2816, w_035_2817, w_035_2820, w_035_2821, w_035_2822, w_035_2823, w_035_2824, w_035_2825, w_035_2826, w_035_2828, w_035_2829, w_035_2830, w_035_2831, w_035_2833, w_035_2834, w_035_2835, w_035_2836, w_035_2837, w_035_2839, w_035_2840, w_035_2843, w_035_2844, w_035_2846, w_035_2847, w_035_2848, w_035_2849, w_035_2857, w_035_2859, w_035_2860, w_035_2862, w_035_2864, w_035_2866, w_035_2868, w_035_2870, w_035_2871, w_035_2872, w_035_2873, w_035_2875, w_035_2876, w_035_2877, w_035_2883, w_035_2884, w_035_2888, w_035_2889, w_035_2894, w_035_2895, w_035_2897, w_035_2898, w_035_2899, w_035_2902, w_035_2905, w_035_2906, w_035_2909, w_035_2912, w_035_2913, w_035_2914, w_035_2915, w_035_2916, w_035_2917, w_035_2919, w_035_2920, w_035_2921, w_035_2922, w_035_2923, w_035_2924, w_035_2925, w_035_2926, w_035_2928, w_035_2929, w_035_2930, w_035_2931, w_035_2932, w_035_2933, w_035_2934, w_035_2935, w_035_2937, w_035_2938, w_035_2939, w_035_2940, w_035_2941, w_035_2943, w_035_2944, w_035_2945, w_035_2946, w_035_2947, w_035_2948, w_035_2953, w_035_2956, w_035_2957, w_035_2958, w_035_2959, w_035_2960, w_035_2961, w_035_2963, w_035_2965, w_035_2966, w_035_2967, w_035_2968, w_035_2970, w_035_2972, w_035_2974, w_035_2975, w_035_2976, w_035_2979, w_035_2980, w_035_2981, w_035_2982, w_035_2983, w_035_2986, w_035_2993, w_035_2997, w_035_2998, w_035_2999, w_035_3001, w_035_3005, w_035_3007, w_035_3009, w_035_3011, w_035_3015, w_035_3016, w_035_3017, w_035_3018, w_035_3019, w_035_3020, w_035_3023, w_035_3025, w_035_3027, w_035_3031, w_035_3032, w_035_3033, w_035_3034, w_035_3035, w_035_3036, w_035_3037, w_035_3038, w_035_3039, w_035_3040, w_035_3041, w_035_3042, w_035_3044, w_035_3045, w_035_3047, w_035_3048, w_035_3049, w_035_3051, w_035_3053, w_035_3057, w_035_3058, w_035_3059, w_035_3061, w_035_3063, w_035_3065, w_035_3066, w_035_3069, w_035_3070, w_035_3071, w_035_3072, w_035_3073, w_035_3075, w_035_3076, w_035_3079, w_035_3081, w_035_3083, w_035_3084, w_035_3085, w_035_3086, w_035_3087, w_035_3088, w_035_3089, w_035_3093, w_035_3094, w_035_3095, w_035_3096, w_035_3097, w_035_3098, w_035_3099, w_035_3100, w_035_3101, w_035_3103, w_035_3105, w_035_3106, w_035_3107, w_035_3108, w_035_3113, w_035_3115, w_035_3117, w_035_3119, w_035_3120, w_035_3122, w_035_3123, w_035_3124, w_035_3125, w_035_3126, w_035_3127, w_035_3131, w_035_3133, w_035_3134, w_035_3135, w_035_3136, w_035_3138, w_035_3140, w_035_3141, w_035_3142, w_035_3143, w_035_3146, w_035_3149, w_035_3150, w_035_3151, w_035_3153, w_035_3156, w_035_3157, w_035_3158, w_035_3162, w_035_3164, w_035_3165, w_035_3167, w_035_3169, w_035_3170, w_035_3172, w_035_3173, w_035_3178, w_035_3179, w_035_3181, w_035_3182, w_035_3183, w_035_3184, w_035_3185, w_035_3187, w_035_3188, w_035_3189, w_035_3190, w_035_3191, w_035_3192, w_035_3193, w_035_3194, w_035_3199, w_035_3200, w_035_3203, w_035_3205, w_035_3207, w_035_3211, w_035_3214, w_035_3215, w_035_3216, w_035_3219, w_035_3221, w_035_3222, w_035_3224, w_035_3225, w_035_3227, w_035_3228, w_035_3229, w_035_3231, w_035_3232, w_035_3235, w_035_3236, w_035_3237, w_035_3238, w_035_3243, w_035_3244, w_035_3246, w_035_3247, w_035_3248, w_035_3250, w_035_3253, w_035_3254, w_035_3255, w_035_3256, w_035_3258, w_035_3259, w_035_3262, w_035_3263, w_035_3264, w_035_3268, w_035_3270, w_035_3271, w_035_3276, w_035_3277, w_035_3278, w_035_3279, w_035_3280, w_035_3281, w_035_3284, w_035_3285, w_035_3287, w_035_3288, w_035_3289, w_035_3291, w_035_3292, w_035_3293, w_035_3294, w_035_3295, w_035_3299, w_035_3300, w_035_3302, w_035_3303, w_035_3304, w_035_3305, w_035_3306, w_035_3307, w_035_3308, w_035_3309, w_035_3310, w_035_3311, w_035_3312, w_035_3313, w_035_3314, w_035_3315, w_035_3316, w_035_3318, w_035_3319, w_035_3323, w_035_3326, w_035_3329, w_035_3331, w_035_3332, w_035_3333, w_035_3336, w_035_3337, w_035_3338, w_035_3339, w_035_3340, w_035_3344, w_035_3348, w_035_3349, w_035_3350, w_035_3351, w_035_3352, w_035_3355, w_035_3356, w_035_3357, w_035_3358, w_035_3359, w_035_3360, w_035_3362, w_035_3366, w_035_3371, w_035_3374, w_035_3375, w_035_3376, w_035_3377, w_035_3380, w_035_3381, w_035_3382, w_035_3384, w_035_3385, w_035_3389, w_035_3391, w_035_3392, w_035_3393, w_035_3394, w_035_3395, w_035_3396, w_035_3399, w_035_3404, w_035_3405, w_035_3406, w_035_3407, w_035_3409, w_035_3412, w_035_3413, w_035_3414, w_035_3415, w_035_3416, w_035_3417, w_035_3418, w_035_3421, w_035_3422, w_035_3424, w_035_3427, w_035_3428, w_035_3429, w_035_3430, w_035_3431, w_035_3434, w_035_3436, w_035_3437, w_035_3438, w_035_3439, w_035_3441, w_035_3443, w_035_3444, w_035_3445, w_035_3447, w_035_3452, w_035_3454, w_035_3457, w_035_3460, w_035_3462, w_035_3463, w_035_3466, w_035_3467, w_035_3469, w_035_3470, w_035_3472, w_035_3474, w_035_3475, w_035_3477, w_035_3478, w_035_3479, w_035_3481, w_035_3483, w_035_3484, w_035_3486, w_035_3488, w_035_3489, w_035_3491, w_035_3493, w_035_3494, w_035_3495, w_035_3497, w_035_3499, w_035_3502, w_035_3504, w_035_3506, w_035_3507, w_035_3510, w_035_3512, w_035_3513, w_035_3514, w_035_3517, w_035_3519, w_035_3520, w_035_3521, w_035_3524, w_035_3527, w_035_3528, w_035_3529, w_035_3532, w_035_3533, w_035_3534, w_035_3539, w_035_3540, w_035_3541, w_035_3542, w_035_3543, w_035_3545, w_035_3546, w_035_3547, w_035_3548, w_035_3549, w_035_3551, w_035_3552, w_035_3553, w_035_3555, w_035_3556, w_035_3559, w_035_3561, w_035_3563, w_035_3564, w_035_3566, w_035_3568, w_035_3570, w_035_3572, w_035_3573, w_035_3576, w_035_3578, w_035_3579, w_035_3581, w_035_3582, w_035_3584, w_035_3585, w_035_3586, w_035_3589, w_035_3590, w_035_3593, w_035_3594, w_035_3596, w_035_3597, w_035_3598, w_035_3599, w_035_3600, w_035_3601, w_035_3607, w_035_3608, w_035_3613, w_035_3615, w_035_3616, w_035_3617, w_035_3618, w_035_3619, w_035_3620, w_035_3621, w_035_3623, w_035_3624, w_035_3625, w_035_3626, w_035_3627, w_035_3629, w_035_3630, w_035_3631, w_035_3632, w_035_3635, w_035_3636, w_035_3637, w_035_3638, w_035_3641, w_035_3643, w_035_3644, w_035_3645, w_035_3646, w_035_3648, w_035_3649, w_035_3650, w_035_3651, w_035_3653, w_035_3654, w_035_3655, w_035_3657, w_035_3658, w_035_3660, w_035_3664, w_035_3666, w_035_3668, w_035_3669, w_035_3670, w_035_3671, w_035_3672, w_035_3674, w_035_3675, w_035_3676, w_035_3677, w_035_3679, w_035_3686, w_035_3690, w_035_3692, w_035_3693, w_035_3694, w_035_3696, w_035_3697, w_035_3698, w_035_3699, w_035_3700, w_035_3701, w_035_3705, w_035_3706, w_035_3707, w_035_3708, w_035_3709, w_035_3712, w_035_3713, w_035_3714, w_035_3715, w_035_3717, w_035_3719, w_035_3721, w_035_3722, w_035_3725, w_035_3727, w_035_3728, w_035_3729, w_035_3730, w_035_3731, w_035_3734, w_035_3735, w_035_3736, w_035_3737, w_035_3738, w_035_3740, w_035_3742, w_035_3743, w_035_3745, w_035_3746, w_035_3749, w_035_3753, w_035_3755, w_035_3757, w_035_3759, w_035_3760, w_035_3761, w_035_3763, w_035_3764, w_035_3765, w_035_3766, w_035_3767, w_035_3769, w_035_3770, w_035_3771, w_035_3772, w_035_3773, w_035_3774, w_035_3776, w_035_3777, w_035_3778, w_035_3779, w_035_3780, w_035_3781, w_035_3782, w_035_3785, w_035_3791, w_035_3793, w_035_3796, w_035_3797, w_035_3798, w_035_3800, w_035_3801, w_035_3805, w_035_3806, w_035_3808, w_035_3810, w_035_3812, w_035_3814, w_035_3815, w_035_3817, w_035_3818, w_035_3819, w_035_3820, w_035_3821, w_035_3822, w_035_3823, w_035_3824, w_035_3826, w_035_3827, w_035_3829, w_035_3830, w_035_3831, w_035_3834, w_035_3835, w_035_3836, w_035_3838, w_035_3839, w_035_3840, w_035_3842, w_035_3843, w_035_3844, w_035_3847, w_035_3848, w_035_3849, w_035_3850, w_035_3852, w_035_3853, w_035_3854, w_035_3857, w_035_3858, w_035_3860, w_035_3861, w_035_3863, w_035_3866, w_035_3868, w_035_3869, w_035_3871, w_035_3872, w_035_3873, w_035_3874, w_035_3875, w_035_3876, w_035_3877, w_035_3879, w_035_3880, w_035_3881, w_035_3883, w_035_3885, w_035_3886, w_035_3889, w_035_3892, w_035_3894, w_035_3895, w_035_3896, w_035_3897, w_035_3898, w_035_3899, w_035_3901, w_035_3902, w_035_3903, w_035_3905, w_035_3906, w_035_3907, w_035_3908, w_035_3909, w_035_3912, w_035_3914, w_035_3915, w_035_3917, w_035_3918, w_035_3920, w_035_3921, w_035_3922, w_035_3923, w_035_3924, w_035_3927, w_035_3928, w_035_3931, w_035_3932, w_035_3936, w_035_3939, w_035_3940, w_035_3941, w_035_3943, w_035_3944, w_035_3945, w_035_3947, w_035_3950, w_035_3956, w_035_3957, w_035_3961, w_035_3963, w_035_3964, w_035_3965, w_035_3967, w_035_3968, w_035_3970, w_035_3971, w_035_3972, w_035_3974, w_035_3975, w_035_3976, w_035_3977, w_035_3979, w_035_3981, w_035_3982, w_035_3985, w_035_3986, w_035_3987, w_035_3988, w_035_3989, w_035_3990, w_035_3992, w_035_3993, w_035_3995, w_035_3996, w_035_3997, w_035_3999, w_035_4000, w_035_4001, w_035_4002, w_035_4004, w_035_4005, w_035_4006, w_035_4007, w_035_4008, w_035_4009, w_035_4010, w_035_4012, w_035_4013, w_035_4014, w_035_4015, w_035_4016, w_035_4017, w_035_4019, w_035_4020, w_035_4021, w_035_4023, w_035_4027, w_035_4028, w_035_4029, w_035_4033, w_035_4034, w_035_4035, w_035_4037, w_035_4039, w_035_4040, w_035_4041, w_035_4042, w_035_4044, w_035_4045, w_035_4046, w_035_4047, w_035_4048, w_035_4050, w_035_4051, w_035_4054, w_035_4055, w_035_4058, w_035_4060, w_035_4062, w_035_4063, w_035_4064, w_035_4065, w_035_4067;
  wire w_036_000, w_036_001, w_036_002, w_036_003, w_036_004, w_036_005, w_036_006, w_036_008, w_036_009, w_036_010, w_036_011, w_036_013, w_036_015, w_036_016, w_036_017, w_036_018, w_036_020, w_036_021, w_036_022, w_036_023, w_036_024, w_036_025, w_036_026, w_036_027, w_036_028, w_036_030, w_036_031, w_036_033, w_036_034, w_036_036, w_036_037, w_036_039, w_036_040, w_036_041, w_036_043, w_036_044, w_036_045, w_036_046, w_036_047, w_036_048, w_036_049, w_036_050, w_036_051, w_036_052, w_036_053, w_036_054, w_036_056, w_036_057, w_036_058, w_036_059, w_036_060, w_036_061, w_036_062, w_036_063, w_036_064, w_036_065, w_036_066, w_036_067, w_036_069, w_036_070, w_036_071, w_036_074, w_036_075, w_036_076, w_036_078, w_036_079, w_036_080, w_036_082, w_036_083, w_036_084, w_036_085, w_036_086, w_036_087, w_036_088, w_036_089, w_036_090, w_036_091, w_036_092, w_036_093, w_036_094, w_036_095, w_036_096, w_036_097, w_036_098, w_036_099, w_036_102, w_036_103, w_036_104, w_036_105, w_036_106, w_036_107, w_036_109, w_036_110, w_036_111, w_036_112, w_036_113, w_036_114, w_036_115, w_036_117, w_036_118, w_036_119, w_036_120, w_036_121, w_036_123, w_036_124, w_036_125, w_036_126, w_036_127, w_036_128, w_036_129, w_036_130, w_036_131, w_036_134, w_036_136, w_036_137, w_036_138, w_036_139, w_036_140, w_036_141, w_036_142, w_036_143, w_036_144, w_036_145, w_036_146, w_036_147, w_036_149, w_036_151, w_036_152, w_036_153, w_036_154, w_036_155, w_036_156, w_036_157, w_036_158, w_036_159, w_036_160, w_036_161, w_036_162, w_036_163, w_036_164, w_036_165, w_036_166, w_036_167, w_036_168, w_036_169, w_036_170, w_036_171, w_036_172, w_036_173, w_036_175, w_036_176, w_036_177, w_036_179, w_036_180, w_036_181, w_036_182, w_036_183, w_036_184, w_036_187, w_036_188, w_036_189, w_036_191, w_036_192, w_036_193, w_036_194, w_036_195, w_036_196, w_036_197, w_036_198, w_036_199, w_036_200, w_036_201, w_036_202, w_036_203, w_036_204, w_036_205, w_036_206, w_036_207, w_036_208, w_036_210, w_036_211, w_036_212, w_036_215, w_036_216, w_036_217, w_036_218, w_036_219, w_036_220, w_036_221, w_036_222, w_036_223, w_036_225, w_036_226, w_036_227, w_036_228, w_036_229, w_036_230, w_036_231, w_036_232, w_036_233, w_036_234, w_036_236, w_036_237, w_036_239, w_036_240, w_036_241, w_036_242, w_036_243, w_036_244, w_036_245, w_036_247, w_036_248, w_036_249, w_036_250, w_036_251, w_036_252, w_036_253, w_036_254, w_036_255, w_036_256, w_036_257, w_036_258, w_036_259, w_036_260, w_036_261, w_036_263, w_036_264, w_036_265, w_036_266, w_036_267, w_036_268, w_036_269, w_036_270, w_036_272, w_036_273, w_036_275, w_036_276, w_036_277, w_036_278, w_036_279, w_036_280, w_036_282, w_036_283, w_036_284, w_036_285, w_036_286, w_036_287, w_036_288, w_036_289, w_036_290, w_036_292, w_036_293, w_036_295, w_036_296, w_036_297, w_036_298, w_036_299, w_036_300, w_036_301, w_036_302, w_036_303, w_036_304, w_036_305, w_036_306, w_036_307, w_036_308, w_036_309, w_036_310, w_036_311, w_036_312, w_036_313, w_036_314, w_036_315, w_036_316, w_036_317, w_036_318, w_036_319, w_036_320, w_036_321, w_036_322, w_036_324, w_036_325, w_036_326, w_036_327, w_036_328, w_036_329, w_036_331, w_036_332, w_036_333, w_036_334, w_036_335, w_036_336, w_036_337, w_036_338, w_036_339, w_036_340, w_036_341, w_036_342, w_036_343, w_036_344, w_036_345, w_036_346, w_036_347, w_036_348, w_036_349, w_036_351, w_036_352, w_036_353, w_036_354, w_036_355, w_036_356, w_036_357, w_036_358, w_036_359, w_036_361, w_036_362, w_036_363, w_036_364, w_036_365, w_036_366, w_036_367, w_036_368, w_036_370, w_036_371, w_036_373, w_036_374, w_036_375, w_036_376, w_036_377, w_036_379, w_036_380, w_036_381, w_036_382, w_036_384, w_036_385, w_036_386, w_036_387, w_036_388, w_036_391, w_036_392, w_036_393, w_036_394, w_036_395, w_036_396, w_036_398, w_036_399, w_036_400, w_036_401, w_036_402, w_036_403, w_036_404, w_036_405, w_036_406, w_036_407, w_036_408, w_036_409, w_036_410, w_036_411, w_036_412, w_036_413, w_036_414, w_036_415, w_036_416, w_036_417, w_036_418, w_036_419, w_036_420, w_036_421, w_036_422, w_036_423, w_036_424, w_036_425, w_036_426, w_036_428, w_036_430, w_036_432, w_036_435, w_036_436, w_036_437, w_036_438, w_036_439, w_036_440, w_036_442, w_036_443, w_036_445, w_036_447, w_036_448, w_036_449, w_036_450, w_036_451, w_036_453, w_036_455, w_036_456, w_036_457, w_036_458, w_036_459, w_036_460, w_036_461, w_036_462, w_036_463, w_036_465, w_036_466, w_036_467, w_036_468, w_036_469, w_036_470, w_036_472, w_036_473, w_036_474, w_036_475, w_036_476, w_036_477, w_036_478, w_036_481, w_036_482, w_036_484, w_036_485, w_036_487, w_036_488, w_036_489, w_036_490, w_036_491, w_036_492, w_036_493, w_036_494, w_036_495, w_036_496, w_036_499, w_036_500, w_036_501, w_036_502, w_036_503, w_036_504, w_036_505, w_036_506, w_036_507, w_036_508, w_036_509, w_036_510, w_036_511, w_036_512, w_036_513, w_036_514, w_036_515, w_036_516, w_036_517, w_036_518, w_036_520, w_036_521, w_036_522, w_036_523, w_036_524, w_036_525, w_036_526, w_036_527, w_036_529, w_036_530, w_036_531, w_036_532, w_036_533, w_036_534, w_036_536, w_036_537, w_036_539, w_036_540, w_036_542, w_036_543, w_036_544, w_036_545, w_036_546, w_036_548, w_036_549, w_036_550, w_036_551, w_036_552, w_036_553, w_036_554, w_036_556, w_036_557, w_036_558, w_036_559, w_036_560, w_036_561, w_036_562, w_036_564, w_036_565, w_036_566, w_036_568, w_036_569, w_036_570, w_036_571, w_036_572, w_036_573, w_036_575, w_036_576, w_036_577, w_036_578, w_036_579, w_036_581, w_036_582, w_036_584, w_036_585, w_036_586, w_036_587, w_036_590, w_036_591, w_036_592, w_036_593, w_036_594, w_036_595, w_036_596, w_036_597, w_036_598, w_036_599, w_036_600, w_036_601, w_036_602, w_036_603, w_036_604, w_036_605, w_036_606, w_036_607, w_036_608, w_036_610, w_036_611, w_036_612, w_036_613, w_036_614, w_036_615, w_036_617, w_036_618, w_036_619, w_036_620, w_036_621, w_036_624, w_036_625, w_036_626, w_036_627, w_036_628, w_036_629, w_036_630, w_036_631, w_036_632, w_036_633, w_036_635, w_036_636, w_036_637, w_036_638, w_036_639, w_036_640, w_036_641, w_036_643, w_036_644, w_036_646, w_036_647, w_036_648, w_036_649, w_036_650, w_036_652, w_036_654, w_036_655, w_036_656, w_036_657, w_036_659, w_036_660, w_036_661, w_036_662, w_036_663, w_036_664, w_036_665, w_036_666, w_036_667, w_036_668, w_036_669, w_036_670, w_036_671, w_036_672, w_036_674, w_036_675, w_036_677, w_036_678, w_036_679, w_036_680, w_036_681, w_036_682, w_036_683, w_036_685, w_036_687, w_036_688, w_036_689, w_036_690, w_036_691, w_036_693, w_036_694, w_036_695, w_036_696, w_036_698, w_036_699, w_036_700, w_036_701, w_036_703, w_036_704, w_036_705, w_036_707, w_036_708, w_036_709, w_036_710, w_036_712, w_036_713, w_036_714, w_036_716, w_036_717, w_036_720, w_036_721, w_036_723, w_036_724, w_036_725, w_036_726, w_036_727, w_036_728, w_036_729, w_036_732, w_036_733, w_036_734, w_036_735, w_036_736, w_036_737, w_036_738, w_036_739, w_036_740, w_036_742, w_036_744, w_036_746, w_036_748, w_036_750, w_036_751, w_036_752, w_036_754, w_036_755, w_036_756, w_036_758, w_036_759, w_036_760, w_036_761, w_036_764, w_036_765, w_036_766, w_036_767, w_036_768, w_036_769, w_036_770, w_036_771, w_036_772, w_036_773, w_036_774, w_036_775, w_036_776, w_036_777, w_036_779, w_036_780, w_036_781, w_036_782, w_036_783, w_036_785, w_036_787, w_036_788, w_036_789, w_036_790, w_036_791, w_036_792, w_036_793, w_036_794, w_036_795, w_036_796, w_036_797, w_036_799, w_036_800, w_036_801, w_036_802, w_036_803, w_036_804, w_036_805, w_036_806, w_036_807, w_036_808, w_036_809, w_036_810, w_036_811, w_036_812, w_036_813, w_036_815, w_036_816, w_036_817, w_036_818, w_036_819, w_036_820, w_036_821, w_036_823, w_036_824, w_036_825, w_036_826, w_036_827, w_036_828, w_036_829, w_036_830, w_036_831, w_036_832, w_036_833, w_036_834, w_036_835, w_036_836, w_036_837, w_036_838, w_036_839, w_036_840, w_036_841, w_036_842, w_036_843, w_036_844, w_036_845, w_036_846, w_036_847, w_036_848, w_036_850, w_036_851, w_036_852, w_036_853, w_036_854, w_036_855, w_036_856, w_036_857, w_036_858, w_036_859, w_036_860, w_036_861, w_036_862, w_036_863, w_036_864, w_036_865, w_036_866, w_036_867, w_036_868, w_036_871, w_036_872, w_036_875, w_036_876, w_036_877, w_036_878, w_036_879, w_036_881, w_036_882, w_036_884, w_036_885, w_036_886, w_036_887, w_036_889, w_036_890, w_036_891, w_036_893, w_036_894, w_036_895, w_036_896, w_036_897, w_036_898, w_036_899, w_036_900, w_036_901, w_036_902, w_036_903, w_036_904, w_036_905, w_036_906, w_036_907, w_036_908, w_036_909, w_036_910, w_036_911, w_036_912, w_036_914, w_036_915, w_036_916, w_036_917, w_036_918, w_036_919, w_036_920, w_036_922, w_036_923, w_036_924, w_036_925, w_036_926, w_036_927, w_036_928, w_036_930, w_036_931, w_036_932, w_036_933, w_036_934, w_036_935, w_036_936, w_036_937, w_036_938, w_036_939, w_036_940, w_036_943, w_036_945, w_036_946, w_036_948, w_036_949, w_036_950, w_036_951, w_036_952, w_036_953, w_036_954, w_036_955, w_036_956, w_036_957, w_036_958, w_036_959, w_036_960, w_036_961, w_036_962, w_036_963, w_036_964, w_036_965, w_036_966, w_036_967, w_036_968, w_036_969, w_036_970, w_036_971, w_036_973, w_036_974, w_036_976, w_036_977, w_036_978, w_036_979, w_036_980, w_036_981, w_036_982, w_036_983, w_036_984, w_036_985, w_036_986, w_036_988, w_036_989, w_036_990, w_036_991, w_036_992, w_036_993, w_036_994, w_036_995, w_036_997, w_036_998, w_036_1000, w_036_1001, w_036_1002, w_036_1003, w_036_1004, w_036_1005, w_036_1006, w_036_1007, w_036_1008, w_036_1009, w_036_1010, w_036_1011, w_036_1012, w_036_1013, w_036_1014, w_036_1015, w_036_1016, w_036_1017, w_036_1018, w_036_1019, w_036_1020, w_036_1021, w_036_1022, w_036_1024, w_036_1025, w_036_1026, w_036_1027, w_036_1028, w_036_1031, w_036_1033, w_036_1034, w_036_1035, w_036_1036, w_036_1037, w_036_1038, w_036_1040, w_036_1041, w_036_1042, w_036_1043, w_036_1044, w_036_1045, w_036_1046, w_036_1047, w_036_1048, w_036_1049, w_036_1050, w_036_1051, w_036_1052, w_036_1053, w_036_1054, w_036_1055, w_036_1056, w_036_1057, w_036_1058, w_036_1059, w_036_1060, w_036_1061, w_036_1062, w_036_1063, w_036_1064, w_036_1065, w_036_1066, w_036_1067, w_036_1068, w_036_1069, w_036_1070, w_036_1071, w_036_1072, w_036_1073, w_036_1074, w_036_1075, w_036_1077, w_036_1078, w_036_1079, w_036_1080, w_036_1081, w_036_1082, w_036_1083, w_036_1084, w_036_1085, w_036_1087, w_036_1088, w_036_1089, w_036_1090, w_036_1091, w_036_1093, w_036_1094, w_036_1095, w_036_1096, w_036_1097, w_036_1098, w_036_1099, w_036_1100, w_036_1101, w_036_1103, w_036_1104, w_036_1105, w_036_1106, w_036_1108, w_036_1110, w_036_1112, w_036_1113, w_036_1114, w_036_1115, w_036_1116, w_036_1117, w_036_1118, w_036_1119, w_036_1120, w_036_1121, w_036_1123, w_036_1125, w_036_1126, w_036_1129, w_036_1130, w_036_1131, w_036_1132, w_036_1133, w_036_1134, w_036_1135, w_036_1136, w_036_1137, w_036_1138, w_036_1139, w_036_1142, w_036_1143, w_036_1144, w_036_1145, w_036_1146, w_036_1147, w_036_1148, w_036_1149, w_036_1150, w_036_1151, w_036_1153, w_036_1154, w_036_1155, w_036_1156, w_036_1157, w_036_1158, w_036_1159, w_036_1160, w_036_1162, w_036_1164, w_036_1165, w_036_1166, w_036_1167, w_036_1168, w_036_1169, w_036_1170, w_036_1171, w_036_1172, w_036_1173, w_036_1174, w_036_1175, w_036_1176, w_036_1177, w_036_1178, w_036_1179, w_036_1180, w_036_1181, w_036_1182, w_036_1183, w_036_1184, w_036_1185, w_036_1186, w_036_1187, w_036_1188, w_036_1189, w_036_1190, w_036_1191, w_036_1192, w_036_1193, w_036_1194, w_036_1196, w_036_1197, w_036_1198, w_036_1199, w_036_1200, w_036_1201, w_036_1202, w_036_1203, w_036_1206, w_036_1207, w_036_1208, w_036_1209, w_036_1211, w_036_1212, w_036_1214, w_036_1215, w_036_1216, w_036_1217, w_036_1218, w_036_1219, w_036_1221, w_036_1223, w_036_1224, w_036_1225, w_036_1226, w_036_1227, w_036_1228, w_036_1230, w_036_1232, w_036_1233, w_036_1234, w_036_1235, w_036_1237, w_036_1238, w_036_1239, w_036_1240, w_036_1241, w_036_1242, w_036_1243, w_036_1244, w_036_1245, w_036_1246, w_036_1247, w_036_1249, w_036_1250, w_036_1252, w_036_1253, w_036_1254, w_036_1255, w_036_1256, w_036_1257, w_036_1258, w_036_1259, w_036_1261, w_036_1262, w_036_1263, w_036_1264, w_036_1265, w_036_1266, w_036_1268, w_036_1269, w_036_1270, w_036_1271, w_036_1272, w_036_1273, w_036_1275, w_036_1276, w_036_1277, w_036_1278, w_036_1279, w_036_1280, w_036_1281, w_036_1282, w_036_1284, w_036_1285, w_036_1286, w_036_1287, w_036_1288, w_036_1289, w_036_1290, w_036_1291, w_036_1292, w_036_1293, w_036_1294, w_036_1296, w_036_1297, w_036_1298, w_036_1299, w_036_1300, w_036_1301, w_036_1302, w_036_1303, w_036_1304, w_036_1305, w_036_1306, w_036_1309, w_036_1310, w_036_1312, w_036_1313, w_036_1314, w_036_1315, w_036_1316, w_036_1317, w_036_1318, w_036_1319, w_036_1320, w_036_1321, w_036_1322, w_036_1323, w_036_1325, w_036_1326, w_036_1327, w_036_1328, w_036_1331, w_036_1332, w_036_1335, w_036_1336, w_036_1337, w_036_1338, w_036_1339, w_036_1340, w_036_1341, w_036_1342, w_036_1343, w_036_1345, w_036_1346, w_036_1347, w_036_1348, w_036_1349, w_036_1350, w_036_1351, w_036_1352, w_036_1353, w_036_1354, w_036_1355, w_036_1356, w_036_1357, w_036_1358, w_036_1359, w_036_1361, w_036_1362, w_036_1363, w_036_1364, w_036_1365, w_036_1366, w_036_1368, w_036_1369, w_036_1370, w_036_1371, w_036_1372, w_036_1374, w_036_1375, w_036_1376, w_036_1377, w_036_1378, w_036_1379, w_036_1380, w_036_1381, w_036_1382, w_036_1383, w_036_1384, w_036_1385, w_036_1386, w_036_1388, w_036_1389, w_036_1390, w_036_1391, w_036_1392, w_036_1393, w_036_1394, w_036_1396, w_036_1397, w_036_1398, w_036_1400, w_036_1403, w_036_1404, w_036_1405, w_036_1406, w_036_1407, w_036_1408, w_036_1409, w_036_1410, w_036_1411, w_036_1412, w_036_1413, w_036_1414, w_036_1415, w_036_1416, w_036_1417, w_036_1418, w_036_1419, w_036_1420, w_036_1421, w_036_1422, w_036_1424, w_036_1425, w_036_1426, w_036_1427, w_036_1429, w_036_1430, w_036_1431, w_036_1432, w_036_1433, w_036_1434, w_036_1435, w_036_1437, w_036_1438, w_036_1439, w_036_1440, w_036_1441, w_036_1442, w_036_1444, w_036_1445, w_036_1446, w_036_1448, w_036_1450, w_036_1451, w_036_1452, w_036_1455, w_036_1456, w_036_1457, w_036_1458, w_036_1460, w_036_1461, w_036_1462, w_036_1464, w_036_1465, w_036_1467, w_036_1468, w_036_1469, w_036_1470, w_036_1472, w_036_1473, w_036_1474, w_036_1475, w_036_1476, w_036_1478, w_036_1479, w_036_1480, w_036_1481, w_036_1482, w_036_1483, w_036_1484, w_036_1486, w_036_1487, w_036_1488, w_036_1489, w_036_1490, w_036_1492, w_036_1495, w_036_1496, w_036_1497, w_036_1499, w_036_1501, w_036_1502, w_036_1503, w_036_1504, w_036_1506, w_036_1507, w_036_1508, w_036_1510, w_036_1511, w_036_1512, w_036_1513, w_036_1514, w_036_1516, w_036_1517, w_036_1518, w_036_1519, w_036_1520, w_036_1522, w_036_1523, w_036_1525, w_036_1526, w_036_1527, w_036_1528, w_036_1530, w_036_1531, w_036_1532, w_036_1533, w_036_1534, w_036_1535, w_036_1536, w_036_1537, w_036_1538, w_036_1539, w_036_1543, w_036_1545, w_036_1546, w_036_1547, w_036_1549, w_036_1550, w_036_1551, w_036_1552, w_036_1553, w_036_1554, w_036_1555, w_036_1556, w_036_1557, w_036_1558, w_036_1559, w_036_1560, w_036_1561, w_036_1562, w_036_1563, w_036_1564, w_036_1566, w_036_1567, w_036_1568, w_036_1569, w_036_1570, w_036_1571, w_036_1572, w_036_1573, w_036_1575, w_036_1576, w_036_1577, w_036_1578, w_036_1579, w_036_1580, w_036_1581, w_036_1582, w_036_1583, w_036_1584, w_036_1585, w_036_1586, w_036_1587, w_036_1588, w_036_1590, w_036_1591, w_036_1592, w_036_1593, w_036_1594, w_036_1595, w_036_1596, w_036_1597, w_036_1598, w_036_1599, w_036_1602, w_036_1603, w_036_1604, w_036_1605, w_036_1606, w_036_1607, w_036_1608, w_036_1609, w_036_1610, w_036_1611, w_036_1612, w_036_1613, w_036_1615, w_036_1616, w_036_1617, w_036_1618, w_036_1619, w_036_1620, w_036_1621, w_036_1622, w_036_1623, w_036_1624, w_036_1625, w_036_1626, w_036_1627, w_036_1628, w_036_1629, w_036_1630, w_036_1631, w_036_1633, w_036_1634, w_036_1635, w_036_1636, w_036_1637, w_036_1638, w_036_1639, w_036_1640, w_036_1641, w_036_1643, w_036_1644, w_036_1645, w_036_1646, w_036_1647, w_036_1648, w_036_1650, w_036_1651, w_036_1652, w_036_1653, w_036_1654, w_036_1655, w_036_1656, w_036_1657, w_036_1658, w_036_1659, w_036_1660, w_036_1661, w_036_1662, w_036_1663, w_036_1665, w_036_1666, w_036_1668, w_036_1669, w_036_1670, w_036_1671, w_036_1672, w_036_1673, w_036_1674, w_036_1675, w_036_1677, w_036_1678, w_036_1680, w_036_1681, w_036_1682, w_036_1683, w_036_1684, w_036_1685, w_036_1686, w_036_1687, w_036_1688, w_036_1689, w_036_1690, w_036_1693, w_036_1694, w_036_1696, w_036_1697, w_036_1698, w_036_1699, w_036_1700, w_036_1701, w_036_1702, w_036_1703, w_036_1704, w_036_1705, w_036_1706, w_036_1707, w_036_1708, w_036_1709, w_036_1710, w_036_1711, w_036_1712, w_036_1713, w_036_1715, w_036_1716, w_036_1717, w_036_1719, w_036_1721, w_036_1722, w_036_1725, w_036_1726, w_036_1727, w_036_1728, w_036_1729, w_036_1730, w_036_1731, w_036_1732, w_036_1733, w_036_1734, w_036_1735, w_036_1736, w_036_1737, w_036_1738, w_036_1740, w_036_1741, w_036_1742, w_036_1743, w_036_1744, w_036_1745, w_036_1746, w_036_1747, w_036_1748, w_036_1749, w_036_1750, w_036_1751, w_036_1752, w_036_1753, w_036_1756, w_036_1757, w_036_1758, w_036_1759, w_036_1760, w_036_1762, w_036_1765, w_036_1766, w_036_1769, w_036_1770, w_036_1771, w_036_1772, w_036_1774, w_036_1775, w_036_1777, w_036_1778, w_036_1779, w_036_1781, w_036_1782, w_036_1783, w_036_1784, w_036_1785, w_036_1786, w_036_1788, w_036_1789, w_036_1790, w_036_1791, w_036_1793, w_036_1794, w_036_1795, w_036_1797, w_036_1798, w_036_1799, w_036_1800, w_036_1801, w_036_1802, w_036_1803, w_036_1805, w_036_1807, w_036_1808, w_036_1809, w_036_1810, w_036_1811, w_036_1812, w_036_1813, w_036_1814, w_036_1815, w_036_1816, w_036_1817, w_036_1819, w_036_1820, w_036_1821, w_036_1822, w_036_1823, w_036_1824, w_036_1825, w_036_1827, w_036_1828, w_036_1829, w_036_1830, w_036_1831, w_036_1832, w_036_1833, w_036_1834, w_036_1835, w_036_1836, w_036_1837, w_036_1838, w_036_1839, w_036_1841, w_036_1843, w_036_1844, w_036_1845, w_036_1846, w_036_1847, w_036_1849, w_036_1850, w_036_1851, w_036_1853, w_036_1854, w_036_1855, w_036_1856, w_036_1857, w_036_1858, w_036_1859, w_036_1860, w_036_1861, w_036_1862, w_036_1863, w_036_1864, w_036_1865, w_036_1866, w_036_1867, w_036_1868, w_036_1869, w_036_1870, w_036_1871, w_036_1872, w_036_1874, w_036_1875, w_036_1876, w_036_1878, w_036_1879, w_036_1880, w_036_1881, w_036_1882, w_036_1883, w_036_1884, w_036_1886, w_036_1887, w_036_1888, w_036_1889, w_036_1890, w_036_1891, w_036_1892, w_036_1893, w_036_1894, w_036_1895, w_036_1896, w_036_1898, w_036_1899, w_036_1900, w_036_1902, w_036_1903, w_036_1905, w_036_1906, w_036_1907, w_036_1908, w_036_1909, w_036_1910, w_036_1911, w_036_1912, w_036_1913, w_036_1914, w_036_1915, w_036_1917, w_036_1918, w_036_1919, w_036_1920, w_036_1921, w_036_1922, w_036_1923, w_036_1924, w_036_1925, w_036_1928, w_036_1930, w_036_1931, w_036_1932, w_036_1933, w_036_1934, w_036_1935, w_036_1936, w_036_1937, w_036_1938, w_036_1939, w_036_1940, w_036_1941, w_036_1942, w_036_1944, w_036_1945, w_036_1946, w_036_1947, w_036_1948, w_036_1949, w_036_1950, w_036_1952, w_036_1953, w_036_1955, w_036_1956, w_036_1957, w_036_1959, w_036_1960, w_036_1961, w_036_1962, w_036_1963, w_036_1964, w_036_1965, w_036_1966, w_036_1968, w_036_1969, w_036_1970, w_036_1971, w_036_1972, w_036_1973, w_036_1974, w_036_1978, w_036_1979, w_036_1981, w_036_1983, w_036_1984, w_036_1985, w_036_1986, w_036_1988, w_036_1989, w_036_1990, w_036_1991, w_036_1992, w_036_1994, w_036_1995, w_036_1996, w_036_1997, w_036_1998, w_036_1999, w_036_2000, w_036_2001, w_036_2002, w_036_2003, w_036_2004, w_036_2005, w_036_2006, w_036_2007, w_036_2008, w_036_2009, w_036_2011, w_036_2013, w_036_2016, w_036_2017, w_036_2018, w_036_2019, w_036_2020, w_036_2021, w_036_2022, w_036_2023, w_036_2024, w_036_2025, w_036_2026, w_036_2027, w_036_2028, w_036_2029, w_036_2030, w_036_2031, w_036_2032, w_036_2033, w_036_2036, w_036_2037, w_036_2040, w_036_2041, w_036_2044, w_036_2046, w_036_2047, w_036_2048, w_036_2049, w_036_2051, w_036_2052, w_036_2054, w_036_2060, w_036_2061, w_036_2067, w_036_2070, w_036_2071, w_036_2074, w_036_2076, w_036_2077, w_036_2078, w_036_2080, w_036_2081, w_036_2083, w_036_2084, w_036_2085, w_036_2088, w_036_2091, w_036_2095, w_036_2097, w_036_2098, w_036_2099, w_036_2101, w_036_2105, w_036_2107, w_036_2108, w_036_2114, w_036_2115, w_036_2116, w_036_2117, w_036_2118, w_036_2122, w_036_2123, w_036_2124, w_036_2126, w_036_2130, w_036_2131, w_036_2132, w_036_2133, w_036_2134, w_036_2135, w_036_2136, w_036_2137, w_036_2139, w_036_2141, w_036_2144, w_036_2145, w_036_2146, w_036_2148, w_036_2149, w_036_2152, w_036_2159, w_036_2161, w_036_2162, w_036_2163, w_036_2164, w_036_2166, w_036_2168, w_036_2171, w_036_2172, w_036_2174, w_036_2175, w_036_2176, w_036_2179, w_036_2180, w_036_2183, w_036_2185, w_036_2186, w_036_2188, w_036_2191, w_036_2192, w_036_2194, w_036_2195, w_036_2197, w_036_2198, w_036_2199, w_036_2201, w_036_2202, w_036_2205, w_036_2210, w_036_2211, w_036_2213, w_036_2214, w_036_2215, w_036_2217, w_036_2218, w_036_2219, w_036_2221, w_036_2222, w_036_2223, w_036_2224, w_036_2225, w_036_2226, w_036_2228, w_036_2229, w_036_2230, w_036_2231, w_036_2232, w_036_2235, w_036_2236, w_036_2237, w_036_2238, w_036_2239, w_036_2241, w_036_2242, w_036_2243, w_036_2245, w_036_2247, w_036_2248, w_036_2251, w_036_2253, w_036_2254, w_036_2257, w_036_2258, w_036_2262, w_036_2265, w_036_2266, w_036_2268, w_036_2269, w_036_2270, w_036_2271, w_036_2272, w_036_2275, w_036_2277, w_036_2278, w_036_2280, w_036_2281, w_036_2284, w_036_2286, w_036_2287, w_036_2288, w_036_2289, w_036_2291, w_036_2292, w_036_2293, w_036_2294, w_036_2297, w_036_2298, w_036_2300, w_036_2301, w_036_2303, w_036_2304, w_036_2305, w_036_2306, w_036_2307, w_036_2308, w_036_2310, w_036_2311, w_036_2312, w_036_2315, w_036_2317, w_036_2318, w_036_2319, w_036_2321, w_036_2322, w_036_2323, w_036_2325, w_036_2326, w_036_2327, w_036_2328, w_036_2329, w_036_2330, w_036_2331, w_036_2334, w_036_2335, w_036_2337, w_036_2341, w_036_2344, w_036_2345, w_036_2347, w_036_2349, w_036_2350, w_036_2351, w_036_2352, w_036_2353, w_036_2354, w_036_2355, w_036_2356, w_036_2357, w_036_2358, w_036_2359, w_036_2360, w_036_2361, w_036_2364, w_036_2365, w_036_2366, w_036_2367, w_036_2371, w_036_2373, w_036_2374, w_036_2375, w_036_2376, w_036_2377, w_036_2378, w_036_2380, w_036_2381, w_036_2385, w_036_2386, w_036_2388, w_036_2389, w_036_2390, w_036_2392, w_036_2396, w_036_2397, w_036_2399, w_036_2402, w_036_2403, w_036_2405, w_036_2406, w_036_2408, w_036_2410, w_036_2413, w_036_2414, w_036_2416, w_036_2418, w_036_2419, w_036_2425, w_036_2426, w_036_2427, w_036_2428, w_036_2433, w_036_2434, w_036_2436, w_036_2437, w_036_2438, w_036_2439, w_036_2440, w_036_2441, w_036_2446, w_036_2447, w_036_2448, w_036_2449, w_036_2450, w_036_2451, w_036_2452, w_036_2453, w_036_2454, w_036_2455, w_036_2457, w_036_2458, w_036_2459, w_036_2460, w_036_2461, w_036_2462, w_036_2463, w_036_2464, w_036_2466, w_036_2468, w_036_2469, w_036_2470, w_036_2472, w_036_2475, w_036_2477, w_036_2478, w_036_2479, w_036_2482, w_036_2483, w_036_2485, w_036_2488, w_036_2489, w_036_2490, w_036_2493, w_036_2494, w_036_2496, w_036_2498, w_036_2499, w_036_2500, w_036_2501, w_036_2502, w_036_2508, w_036_2509, w_036_2510, w_036_2512, w_036_2515, w_036_2516, w_036_2517, w_036_2519, w_036_2522, w_036_2523, w_036_2524, w_036_2527, w_036_2528, w_036_2529, w_036_2530, w_036_2531, w_036_2533, w_036_2534, w_036_2537, w_036_2538, w_036_2539, w_036_2541, w_036_2543, w_036_2544, w_036_2547, w_036_2549, w_036_2550, w_036_2551, w_036_2552, w_036_2553, w_036_2558, w_036_2560, w_036_2564, w_036_2565, w_036_2567, w_036_2573, w_036_2574, w_036_2575, w_036_2577, w_036_2578, w_036_2579, w_036_2580, w_036_2584, w_036_2585, w_036_2586, w_036_2587, w_036_2590, w_036_2591, w_036_2592, w_036_2593, w_036_2598, w_036_2601, w_036_2602, w_036_2604, w_036_2605, w_036_2606, w_036_2607, w_036_2608, w_036_2610, w_036_2612, w_036_2613, w_036_2615, w_036_2618, w_036_2620, w_036_2621, w_036_2622, w_036_2625, w_036_2626, w_036_2627, w_036_2628, w_036_2629, w_036_2630, w_036_2631, w_036_2634, w_036_2635, w_036_2636, w_036_2642, w_036_2643, w_036_2644, w_036_2645, w_036_2647, w_036_2648, w_036_2649, w_036_2651, w_036_2652, w_036_2653, w_036_2654, w_036_2656, w_036_2657, w_036_2659, w_036_2662, w_036_2663, w_036_2664, w_036_2666, w_036_2667, w_036_2668, w_036_2669, w_036_2671, w_036_2672, w_036_2673, w_036_2674, w_036_2675, w_036_2676, w_036_2677, w_036_2679, w_036_2681, w_036_2682, w_036_2683, w_036_2686, w_036_2687, w_036_2688, w_036_2689, w_036_2690, w_036_2691, w_036_2692, w_036_2693, w_036_2696, w_036_2699, w_036_2700, w_036_2702, w_036_2703, w_036_2705, w_036_2707, w_036_2712, w_036_2715, w_036_2717, w_036_2720, w_036_2721, w_036_2722, w_036_2723, w_036_2724, w_036_2726, w_036_2727, w_036_2729, w_036_2730, w_036_2732, w_036_2734, w_036_2737, w_036_2739, w_036_2740, w_036_2741, w_036_2742, w_036_2743, w_036_2746, w_036_2747, w_036_2748, w_036_2749, w_036_2753, w_036_2756, w_036_2757, w_036_2758, w_036_2759, w_036_2762, w_036_2763, w_036_2765, w_036_2766, w_036_2767, w_036_2768, w_036_2769, w_036_2771, w_036_2772, w_036_2773, w_036_2774, w_036_2775, w_036_2776, w_036_2778, w_036_2779, w_036_2780, w_036_2782, w_036_2783, w_036_2785, w_036_2786, w_036_2787, w_036_2789, w_036_2791, w_036_2793, w_036_2794, w_036_2795, w_036_2797, w_036_2798, w_036_2799, w_036_2800, w_036_2801, w_036_2805, w_036_2806, w_036_2807, w_036_2809, w_036_2810, w_036_2812, w_036_2813, w_036_2814, w_036_2817, w_036_2818, w_036_2819, w_036_2820, w_036_2821, w_036_2822, w_036_2823, w_036_2824, w_036_2825, w_036_2829, w_036_2830, w_036_2831, w_036_2833, w_036_2834, w_036_2836, w_036_2837, w_036_2838, w_036_2839, w_036_2840, w_036_2841, w_036_2843, w_036_2846, w_036_2848, w_036_2850, w_036_2851, w_036_2852, w_036_2853, w_036_2854, w_036_2855, w_036_2856, w_036_2857, w_036_2858, w_036_2859, w_036_2861, w_036_2863, w_036_2866, w_036_2867, w_036_2869, w_036_2872, w_036_2873, w_036_2874, w_036_2876, w_036_2877, w_036_2878, w_036_2879, w_036_2880, w_036_2882, w_036_2884, w_036_2885, w_036_2887, w_036_2888, w_036_2891, w_036_2892, w_036_2893, w_036_2894, w_036_2896, w_036_2899, w_036_2900, w_036_2901, w_036_2902, w_036_2903, w_036_2905, w_036_2907, w_036_2908, w_036_2909, w_036_2910, w_036_2912, w_036_2913, w_036_2916, w_036_2918, w_036_2920, w_036_2921, w_036_2922, w_036_2924, w_036_2925, w_036_2927, w_036_2933, w_036_2934, w_036_2938, w_036_2939, w_036_2941, w_036_2943, w_036_2945, w_036_2947, w_036_2949, w_036_2950, w_036_2951, w_036_2952, w_036_2954, w_036_2958, w_036_2959, w_036_2960, w_036_2961;
  wire w_037_000, w_037_001, w_037_002, w_037_003, w_037_004, w_037_005, w_037_006, w_037_007, w_037_008, w_037_009, w_037_010, w_037_011, w_037_013, w_037_014, w_037_015, w_037_016, w_037_017, w_037_018, w_037_019, w_037_022, w_037_023, w_037_024, w_037_025, w_037_026, w_037_028, w_037_029, w_037_031, w_037_032, w_037_033, w_037_035, w_037_036, w_037_037, w_037_038, w_037_039, w_037_041, w_037_042, w_037_043, w_037_044, w_037_045, w_037_046, w_037_047, w_037_048, w_037_049, w_037_051, w_037_052, w_037_053, w_037_057, w_037_059, w_037_060, w_037_061, w_037_062, w_037_063, w_037_064, w_037_065, w_037_066, w_037_067, w_037_068, w_037_069, w_037_070, w_037_071, w_037_073, w_037_074, w_037_075, w_037_076, w_037_078, w_037_080, w_037_081, w_037_082, w_037_083, w_037_084, w_037_085, w_037_087, w_037_088, w_037_089, w_037_090, w_037_091, w_037_093, w_037_095, w_037_097, w_037_098, w_037_099, w_037_101, w_037_102, w_037_103, w_037_104, w_037_105, w_037_107, w_037_108, w_037_109, w_037_110, w_037_112, w_037_113, w_037_114, w_037_116, w_037_117, w_037_119, w_037_120, w_037_121, w_037_122, w_037_123, w_037_125, w_037_126, w_037_127, w_037_130, w_037_131, w_037_132, w_037_133, w_037_134, w_037_135, w_037_136, w_037_137, w_037_138, w_037_139, w_037_140, w_037_141, w_037_142, w_037_143, w_037_144, w_037_145, w_037_148, w_037_150, w_037_151, w_037_152, w_037_153, w_037_154, w_037_156, w_037_157, w_037_158, w_037_159, w_037_161, w_037_162, w_037_163, w_037_164, w_037_165, w_037_166, w_037_168, w_037_169, w_037_170, w_037_171, w_037_172, w_037_173, w_037_174, w_037_175, w_037_176, w_037_177, w_037_179, w_037_180, w_037_181, w_037_182, w_037_183, w_037_184, w_037_185, w_037_186, w_037_187, w_037_188, w_037_189, w_037_190, w_037_191, w_037_193, w_037_195, w_037_196, w_037_198, w_037_199, w_037_200, w_037_201, w_037_202, w_037_203, w_037_204, w_037_205, w_037_206, w_037_207, w_037_209, w_037_211, w_037_212, w_037_214, w_037_215, w_037_216, w_037_217, w_037_218, w_037_220, w_037_221, w_037_223, w_037_224, w_037_225, w_037_226, w_037_227, w_037_228, w_037_229, w_037_230, w_037_232, w_037_233, w_037_234, w_037_236, w_037_237, w_037_238, w_037_239, w_037_240, w_037_242, w_037_243, w_037_244, w_037_245, w_037_246, w_037_247, w_037_248, w_037_249, w_037_251, w_037_252, w_037_253, w_037_254, w_037_256, w_037_258, w_037_259, w_037_260, w_037_261, w_037_262, w_037_265, w_037_266, w_037_267, w_037_268, w_037_269, w_037_270, w_037_272, w_037_273, w_037_275, w_037_276, w_037_278, w_037_280, w_037_281, w_037_282, w_037_283, w_037_284, w_037_285, w_037_286, w_037_287, w_037_288, w_037_289, w_037_290, w_037_291, w_037_292, w_037_294, w_037_295, w_037_297, w_037_298, w_037_299, w_037_300, w_037_301, w_037_303, w_037_305, w_037_306, w_037_307, w_037_308, w_037_309, w_037_310, w_037_311, w_037_312, w_037_313, w_037_314, w_037_315, w_037_316, w_037_318, w_037_319, w_037_320, w_037_321, w_037_322, w_037_325, w_037_327, w_037_328, w_037_329, w_037_331, w_037_332, w_037_334, w_037_335, w_037_336, w_037_337, w_037_338, w_037_339, w_037_342, w_037_343, w_037_344, w_037_345, w_037_346, w_037_347, w_037_348, w_037_349, w_037_350, w_037_352, w_037_353, w_037_354, w_037_355, w_037_357, w_037_358, w_037_359, w_037_360, w_037_361, w_037_362, w_037_365, w_037_366, w_037_368, w_037_369, w_037_371, w_037_372, w_037_373, w_037_374, w_037_375, w_037_376, w_037_378, w_037_379, w_037_380, w_037_381, w_037_382, w_037_384, w_037_385, w_037_386, w_037_387, w_037_390, w_037_392, w_037_393, w_037_394, w_037_395, w_037_396, w_037_398, w_037_399, w_037_400, w_037_401, w_037_402, w_037_403, w_037_405, w_037_406, w_037_407, w_037_409, w_037_410, w_037_411, w_037_412, w_037_413, w_037_414, w_037_415, w_037_418, w_037_419, w_037_421, w_037_422, w_037_423, w_037_424, w_037_425, w_037_427, w_037_430, w_037_431, w_037_432, w_037_433, w_037_435, w_037_437, w_037_438, w_037_439, w_037_440, w_037_441, w_037_443, w_037_444, w_037_445, w_037_446, w_037_447, w_037_448, w_037_449, w_037_450, w_037_451, w_037_453, w_037_456, w_037_457, w_037_458, w_037_460, w_037_461, w_037_462, w_037_463, w_037_464, w_037_465, w_037_466, w_037_467, w_037_468, w_037_469, w_037_470, w_037_473, w_037_474, w_037_476, w_037_477, w_037_478, w_037_479, w_037_480, w_037_481, w_037_482, w_037_483, w_037_484, w_037_486, w_037_487, w_037_488, w_037_490, w_037_491, w_037_493, w_037_494, w_037_495, w_037_497, w_037_498, w_037_499, w_037_500, w_037_501, w_037_504, w_037_505, w_037_506, w_037_508, w_037_509, w_037_510, w_037_511, w_037_512, w_037_513, w_037_514, w_037_515, w_037_516, w_037_517, w_037_518, w_037_519, w_037_521, w_037_522, w_037_523, w_037_525, w_037_527, w_037_528, w_037_531, w_037_532, w_037_533, w_037_534, w_037_536, w_037_537, w_037_538, w_037_540, w_037_541, w_037_542, w_037_543, w_037_544, w_037_545, w_037_547, w_037_548, w_037_549, w_037_550, w_037_551, w_037_552, w_037_554, w_037_555, w_037_556, w_037_557, w_037_558, w_037_559, w_037_560, w_037_561, w_037_562, w_037_563, w_037_566, w_037_567, w_037_568, w_037_569, w_037_572, w_037_573, w_037_574, w_037_576, w_037_577, w_037_579, w_037_580, w_037_582, w_037_583, w_037_584, w_037_585, w_037_586, w_037_587, w_037_588, w_037_589, w_037_590, w_037_592, w_037_593, w_037_594, w_037_595, w_037_596, w_037_597, w_037_598, w_037_600, w_037_602, w_037_603, w_037_604, w_037_605, w_037_607, w_037_609, w_037_610, w_037_611, w_037_613, w_037_615, w_037_616, w_037_617, w_037_619, w_037_620, w_037_621, w_037_623, w_037_625, w_037_626, w_037_627, w_037_628, w_037_629, w_037_630, w_037_631, w_037_632, w_037_633, w_037_634, w_037_635, w_037_636, w_037_637, w_037_638, w_037_641, w_037_642, w_037_643, w_037_644, w_037_645, w_037_646, w_037_647, w_037_648, w_037_649, w_037_650, w_037_651, w_037_652, w_037_653, w_037_654, w_037_656, w_037_657, w_037_658, w_037_659, w_037_661, w_037_662, w_037_663, w_037_664, w_037_665, w_037_666, w_037_667, w_037_668, w_037_669, w_037_670, w_037_671, w_037_672, w_037_673, w_037_674, w_037_676, w_037_677, w_037_678, w_037_679, w_037_682, w_037_683, w_037_685, w_037_686, w_037_687, w_037_688, w_037_689, w_037_690, w_037_691, w_037_692, w_037_693, w_037_695, w_037_696, w_037_697, w_037_699, w_037_701, w_037_703, w_037_707, w_037_708, w_037_709, w_037_710, w_037_711, w_037_713, w_037_715, w_037_717, w_037_718, w_037_719, w_037_721, w_037_722, w_037_723, w_037_725, w_037_728, w_037_729, w_037_730, w_037_731, w_037_733, w_037_734, w_037_736, w_037_737, w_037_738, w_037_740, w_037_741, w_037_743, w_037_744, w_037_745, w_037_746, w_037_748, w_037_749, w_037_750, w_037_752, w_037_753, w_037_754, w_037_755, w_037_756, w_037_757, w_037_758, w_037_759, w_037_760, w_037_761, w_037_762, w_037_763, w_037_764, w_037_765, w_037_766, w_037_767, w_037_768, w_037_769, w_037_770, w_037_771, w_037_773, w_037_775, w_037_776, w_037_778, w_037_779, w_037_780, w_037_781, w_037_782, w_037_783, w_037_784, w_037_785, w_037_786, w_037_787, w_037_788, w_037_790, w_037_791, w_037_792, w_037_793, w_037_797, w_037_798, w_037_801, w_037_802, w_037_803, w_037_805, w_037_806, w_037_807, w_037_808, w_037_809, w_037_810, w_037_811, w_037_813, w_037_814, w_037_815, w_037_817, w_037_818, w_037_819, w_037_820, w_037_821, w_037_822, w_037_824, w_037_825, w_037_826, w_037_828, w_037_829, w_037_830, w_037_831, w_037_832, w_037_833, w_037_836, w_037_837, w_037_838, w_037_839, w_037_840, w_037_841, w_037_843, w_037_844, w_037_845, w_037_846, w_037_847, w_037_848, w_037_849, w_037_850, w_037_851, w_037_852, w_037_853, w_037_854, w_037_855, w_037_856, w_037_857, w_037_858, w_037_859, w_037_861, w_037_863, w_037_865, w_037_866, w_037_867, w_037_868, w_037_869, w_037_870, w_037_871, w_037_872, w_037_873, w_037_875, w_037_876, w_037_877, w_037_878, w_037_879, w_037_881, w_037_883, w_037_886, w_037_887, w_037_888, w_037_889, w_037_890, w_037_891, w_037_892, w_037_893, w_037_895, w_037_896, w_037_897, w_037_898, w_037_899, w_037_900, w_037_901, w_037_902, w_037_903, w_037_904, w_037_905, w_037_906, w_037_907, w_037_908, w_037_909, w_037_910, w_037_911, w_037_912, w_037_914, w_037_915, w_037_916, w_037_918, w_037_919, w_037_920, w_037_921, w_037_922, w_037_924, w_037_925, w_037_926, w_037_927, w_037_928, w_037_930, w_037_932, w_037_933, w_037_934, w_037_935, w_037_937, w_037_938, w_037_939, w_037_940, w_037_941, w_037_942, w_037_943, w_037_944, w_037_945, w_037_946, w_037_947, w_037_948, w_037_949, w_037_950, w_037_951, w_037_952, w_037_953, w_037_955, w_037_956, w_037_957, w_037_958, w_037_959, w_037_960, w_037_961, w_037_962, w_037_963, w_037_965, w_037_966, w_037_967, w_037_968, w_037_969, w_037_970, w_037_971, w_037_972, w_037_973, w_037_974, w_037_975, w_037_977, w_037_978, w_037_979, w_037_980, w_037_981, w_037_983, w_037_984, w_037_985, w_037_986, w_037_987, w_037_988, w_037_989, w_037_990, w_037_991, w_037_992, w_037_993, w_037_994, w_037_995, w_037_996, w_037_997, w_037_998, w_037_1000, w_037_1001, w_037_1002, w_037_1004, w_037_1005, w_037_1006, w_037_1009, w_037_1010, w_037_1011, w_037_1012, w_037_1013, w_037_1014, w_037_1015, w_037_1016, w_037_1017, w_037_1018, w_037_1019, w_037_1020, w_037_1021, w_037_1022, w_037_1023, w_037_1024, w_037_1025, w_037_1026, w_037_1027, w_037_1028, w_037_1029, w_037_1030, w_037_1031, w_037_1032, w_037_1033, w_037_1034, w_037_1035, w_037_1036, w_037_1037, w_037_1038, w_037_1039, w_037_1041, w_037_1042, w_037_1043, w_037_1044, w_037_1045, w_037_1046, w_037_1047, w_037_1048, w_037_1049, w_037_1050, w_037_1051, w_037_1052, w_037_1053, w_037_1054, w_037_1055, w_037_1056, w_037_1057, w_037_1058, w_037_1059, w_037_1060, w_037_1061, w_037_1063, w_037_1064, w_037_1065, w_037_1067, w_037_1069, w_037_1070, w_037_1071, w_037_1072, w_037_1073, w_037_1075, w_037_1076, w_037_1079, w_037_1080, w_037_1082, w_037_1084, w_037_1085, w_037_1086, w_037_1087, w_037_1088, w_037_1090, w_037_1091, w_037_1093, w_037_1094, w_037_1095, w_037_1096, w_037_1097, w_037_1098, w_037_1099, w_037_1100, w_037_1101, w_037_1102, w_037_1103, w_037_1105, w_037_1106, w_037_1107, w_037_1108, w_037_1109, w_037_1110, w_037_1111, w_037_1112, w_037_1113, w_037_1114, w_037_1115, w_037_1116, w_037_1117, w_037_1118, w_037_1119, w_037_1120, w_037_1121, w_037_1122, w_037_1123, w_037_1124, w_037_1125, w_037_1126, w_037_1127, w_037_1128, w_037_1129, w_037_1131, w_037_1132, w_037_1133, w_037_1134, w_037_1135, w_037_1136, w_037_1138, w_037_1139, w_037_1140, w_037_1141, w_037_1142, w_037_1143, w_037_1146, w_037_1147, w_037_1148, w_037_1149, w_037_1150, w_037_1151, w_037_1152, w_037_1153, w_037_1154, w_037_1155, w_037_1156, w_037_1157, w_037_1158, w_037_1159, w_037_1161, w_037_1163, w_037_1164, w_037_1165, w_037_1167, w_037_1168, w_037_1169, w_037_1170, w_037_1171, w_037_1172, w_037_1173, w_037_1175, w_037_1176, w_037_1177, w_037_1178, w_037_1179, w_037_1180, w_037_1182, w_037_1183, w_037_1184, w_037_1185, w_037_1186, w_037_1187, w_037_1188, w_037_1189, w_037_1190, w_037_1191, w_037_1192, w_037_1193, w_037_1196, w_037_1197, w_037_1198, w_037_1199, w_037_1200, w_037_1202, w_037_1203, w_037_1204, w_037_1206, w_037_1207, w_037_1208, w_037_1209, w_037_1210, w_037_1212, w_037_1213, w_037_1214, w_037_1216, w_037_1217, w_037_1218, w_037_1219, w_037_1220, w_037_1221, w_037_1222, w_037_1223, w_037_1224, w_037_1225, w_037_1226, w_037_1228, w_037_1229, w_037_1230, w_037_1231, w_037_1232, w_037_1233, w_037_1234, w_037_1235, w_037_1236, w_037_1237, w_037_1238, w_037_1239, w_037_1240, w_037_1242, w_037_1243, w_037_1244, w_037_1246, w_037_1247, w_037_1248, w_037_1249, w_037_1250, w_037_1252, w_037_1253, w_037_1256, w_037_1257, w_037_1258, w_037_1259, w_037_1260, w_037_1261, w_037_1262, w_037_1263, w_037_1264, w_037_1265, w_037_1266, w_037_1269, w_037_1270, w_037_1271, w_037_1272, w_037_1273, w_037_1274, w_037_1275, w_037_1276, w_037_1277, w_037_1278, w_037_1279, w_037_1280, w_037_1281, w_037_1282, w_037_1283, w_037_1284, w_037_1285, w_037_1286, w_037_1287, w_037_1288, w_037_1290, w_037_1292, w_037_1293, w_037_1294, w_037_1295, w_037_1296, w_037_1297, w_037_1298, w_037_1300, w_037_1301, w_037_1302, w_037_1303, w_037_1304, w_037_1305, w_037_1307, w_037_1308, w_037_1309, w_037_1310, w_037_1311, w_037_1312, w_037_1313, w_037_1314, w_037_1316, w_037_1317, w_037_1318, w_037_1320, w_037_1321, w_037_1322, w_037_1324, w_037_1325, w_037_1326, w_037_1327, w_037_1328, w_037_1330, w_037_1331, w_037_1332, w_037_1333, w_037_1334, w_037_1335, w_037_1336, w_037_1337, w_037_1338, w_037_1340, w_037_1341, w_037_1342, w_037_1343, w_037_1344, w_037_1345, w_037_1349, w_037_1350, w_037_1351, w_037_1352, w_037_1353, w_037_1354, w_037_1356, w_037_1358, w_037_1359, w_037_1360, w_037_1361, w_037_1362, w_037_1363, w_037_1364, w_037_1365, w_037_1366, w_037_1367, w_037_1368, w_037_1369, w_037_1370, w_037_1371, w_037_1372, w_037_1374, w_037_1375, w_037_1376, w_037_1377, w_037_1378, w_037_1380, w_037_1381, w_037_1382, w_037_1383, w_037_1386, w_037_1387, w_037_1388, w_037_1389, w_037_1391, w_037_1392, w_037_1393, w_037_1395, w_037_1397, w_037_1398, w_037_1399, w_037_1401, w_037_1403, w_037_1404, w_037_1406, w_037_1407, w_037_1408, w_037_1410, w_037_1412, w_037_1413, w_037_1414, w_037_1415, w_037_1416, w_037_1417, w_037_1418, w_037_1419, w_037_1420, w_037_1422, w_037_1423, w_037_1425, w_037_1426, w_037_1427, w_037_1428, w_037_1429, w_037_1431, w_037_1432, w_037_1435, w_037_1436, w_037_1437, w_037_1438, w_037_1439, w_037_1440, w_037_1441, w_037_1442, w_037_1443, w_037_1444, w_037_1445, w_037_1446, w_037_1447, w_037_1449, w_037_1450, w_037_1451, w_037_1453, w_037_1454, w_037_1455, w_037_1456, w_037_1457, w_037_1458, w_037_1459, w_037_1460, w_037_1461, w_037_1462, w_037_1463, w_037_1464, w_037_1465, w_037_1466, w_037_1467, w_037_1468, w_037_1469, w_037_1470, w_037_1471, w_037_1472, w_037_1473, w_037_1474, w_037_1475, w_037_1476, w_037_1477, w_037_1479, w_037_1480, w_037_1483, w_037_1484, w_037_1485, w_037_1486, w_037_1487, w_037_1488, w_037_1489, w_037_1491, w_037_1492, w_037_1493, w_037_1494, w_037_1495, w_037_1496, w_037_1498, w_037_1500, w_037_1501, w_037_1502, w_037_1503, w_037_1504, w_037_1505, w_037_1506, w_037_1507, w_037_1508, w_037_1509, w_037_1510, w_037_1511, w_037_1512, w_037_1513, w_037_1514, w_037_1515, w_037_1516, w_037_1517, w_037_1518, w_037_1519, w_037_1520, w_037_1523, w_037_1524, w_037_1525, w_037_1526, w_037_1527, w_037_1528, w_037_1529, w_037_1530, w_037_1532, w_037_1533, w_037_1534, w_037_1536, w_037_1537, w_037_1538, w_037_1539, w_037_1540, w_037_1541, w_037_1542, w_037_1547, w_037_1548, w_037_1550, w_037_1551, w_037_1552, w_037_1553, w_037_1554, w_037_1555, w_037_1556, w_037_1557, w_037_1558, w_037_1560, w_037_1561, w_037_1562, w_037_1563, w_037_1564, w_037_1565, w_037_1567, w_037_1568, w_037_1569, w_037_1570, w_037_1572, w_037_1573, w_037_1574, w_037_1575, w_037_1576, w_037_1577, w_037_1578, w_037_1579, w_037_1580, w_037_1581, w_037_1583, w_037_1584, w_037_1585, w_037_1586, w_037_1587, w_037_1588, w_037_1589, w_037_1592, w_037_1593, w_037_1594, w_037_1595, w_037_1596, w_037_1597, w_037_1598, w_037_1599, w_037_1600, w_037_1603, w_037_1605, w_037_1606, w_037_1607, w_037_1608, w_037_1609, w_037_1610, w_037_1611, w_037_1612, w_037_1614, w_037_1615, w_037_1616, w_037_1618, w_037_1619, w_037_1621, w_037_1624, w_037_1625, w_037_1626, w_037_1628, w_037_1631, w_037_1632, w_037_1633, w_037_1634, w_037_1635, w_037_1636, w_037_1637, w_037_1638, w_037_1639, w_037_1640, w_037_1641, w_037_1643, w_037_1645, w_037_1646, w_037_1647, w_037_1648, w_037_1649, w_037_1651, w_037_1652, w_037_1653, w_037_1654, w_037_1655, w_037_1656, w_037_1657, w_037_1658, w_037_1660, w_037_1661, w_037_1662, w_037_1663, w_037_1665, w_037_1666, w_037_1667, w_037_1669, w_037_1670, w_037_1671, w_037_1673, w_037_1675, w_037_1676, w_037_1677, w_037_1678, w_037_1679, w_037_1680, w_037_1681, w_037_1683, w_037_1685, w_037_1686, w_037_1688, w_037_1689, w_037_1690, w_037_1691, w_037_1693, w_037_1694, w_037_1695, w_037_1696, w_037_1697, w_037_1698, w_037_1699, w_037_1701, w_037_1702, w_037_1703, w_037_1704, w_037_1706, w_037_1707, w_037_1708, w_037_1709, w_037_1710, w_037_1711, w_037_1713, w_037_1714, w_037_1715, w_037_1716, w_037_1717, w_037_1718, w_037_1719, w_037_1720, w_037_1721, w_037_1722, w_037_1724, w_037_1725, w_037_1726, w_037_1727, w_037_1729, w_037_1730, w_037_1731, w_037_1732, w_037_1733, w_037_1734, w_037_1735, w_037_1737, w_037_1738, w_037_1739, w_037_1741, w_037_1742, w_037_1743, w_037_1744, w_037_1745, w_037_1746, w_037_1748, w_037_1749, w_037_1750, w_037_1751, w_037_1752, w_037_1753, w_037_1754, w_037_1756, w_037_1757, w_037_1759, w_037_1760, w_037_1761, w_037_1762, w_037_1763, w_037_1764, w_037_1767, w_037_1768, w_037_1770, w_037_1772, w_037_1773, w_037_1775, w_037_1776, w_037_1777, w_037_1778, w_037_1779, w_037_1780, w_037_1781, w_037_1783, w_037_1784, w_037_1785, w_037_1787, w_037_1790, w_037_1791, w_037_1792, w_037_1794, w_037_1795, w_037_1796, w_037_1798, w_037_1799, w_037_1800, w_037_1801, w_037_1802, w_037_1803, w_037_1804, w_037_1806, w_037_1807, w_037_1808, w_037_1809, w_037_1811, w_037_1812, w_037_1813, w_037_1814, w_037_1816, w_037_1817, w_037_1818, w_037_1819, w_037_1820, w_037_1821, w_037_1824, w_037_1825, w_037_1826, w_037_1827, w_037_1829, w_037_1830, w_037_1831, w_037_1832, w_037_1833, w_037_1834, w_037_1836, w_037_1837, w_037_1838, w_037_1840, w_037_1841, w_037_1842, w_037_1844, w_037_1846, w_037_1847, w_037_1848, w_037_1850, w_037_1851, w_037_1852, w_037_1853, w_037_1854, w_037_1855, w_037_1856, w_037_1857, w_037_1858, w_037_1860, w_037_1863, w_037_1864, w_037_1865, w_037_1866, w_037_1867, w_037_1868, w_037_1871, w_037_1872, w_037_1874, w_037_1875, w_037_1876, w_037_1877, w_037_1878, w_037_1879, w_037_1880, w_037_1881, w_037_1883, w_037_1884, w_037_1885, w_037_1886, w_037_1887, w_037_1888, w_037_1889, w_037_1890, w_037_1891, w_037_1893, w_037_1894, w_037_1895, w_037_1896, w_037_1897, w_037_1898, w_037_1899, w_037_1900, w_037_1901, w_037_1903, w_037_1904, w_037_1905, w_037_1906, w_037_1909, w_037_1910, w_037_1911, w_037_1912, w_037_1913, w_037_1915, w_037_1916, w_037_1917, w_037_1918, w_037_1919, w_037_1921, w_037_1922, w_037_1923, w_037_1924, w_037_1926, w_037_1927, w_037_1928, w_037_1930, w_037_1931, w_037_1932, w_037_1933, w_037_1934, w_037_1935, w_037_1936, w_037_1937, w_037_1938, w_037_1939, w_037_1941, w_037_1942, w_037_1943, w_037_1944, w_037_1946, w_037_1947, w_037_1948, w_037_1949, w_037_1951, w_037_1952, w_037_1953, w_037_1954, w_037_1955, w_037_1956, w_037_1958, w_037_1959, w_037_1961, w_037_1962, w_037_1963, w_037_1964, w_037_1965, w_037_1966, w_037_1967, w_037_1968, w_037_1969, w_037_1972, w_037_1975, w_037_1976, w_037_1978, w_037_1979, w_037_1980, w_037_1982, w_037_1983, w_037_1984, w_037_1985, w_037_1986, w_037_1988, w_037_1989, w_037_1990, w_037_1991, w_037_1992, w_037_1995, w_037_1996, w_037_1997, w_037_1998, w_037_1999, w_037_2000, w_037_2001, w_037_2002, w_037_2006, w_037_2007, w_037_2008, w_037_2009, w_037_2010, w_037_2011, w_037_2013, w_037_2015, w_037_2016, w_037_2017, w_037_2018, w_037_2019, w_037_2020, w_037_2022, w_037_2023, w_037_2024, w_037_2025, w_037_2026, w_037_2029, w_037_2030, w_037_2032, w_037_2033, w_037_2034, w_037_2035, w_037_2036, w_037_2037, w_037_2038, w_037_2039, w_037_2040, w_037_2041, w_037_2042, w_037_2043, w_037_2044, w_037_2045, w_037_2046, w_037_2048, w_037_2049, w_037_2050, w_037_2051, w_037_2053, w_037_2056, w_037_2057, w_037_2058, w_037_2059, w_037_2060, w_037_2062, w_037_2064, w_037_2065, w_037_2066, w_037_2067, w_037_2069, w_037_2070, w_037_2072, w_037_2073, w_037_2074, w_037_2075, w_037_2078, w_037_2079, w_037_2080, w_037_2081, w_037_2082, w_037_2083, w_037_2084, w_037_2085, w_037_2086, w_037_2087, w_037_2089, w_037_2090, w_037_2092, w_037_2093, w_037_2094, w_037_2095, w_037_2096, w_037_2097, w_037_2098, w_037_2099, w_037_2100, w_037_2101, w_037_2103, w_037_2104, w_037_2106, w_037_2107, w_037_2110, w_037_2111, w_037_2113, w_037_2115, w_037_2117, w_037_2118, w_037_2119, w_037_2120, w_037_2121, w_037_2122, w_037_2123, w_037_2124, w_037_2125, w_037_2126, w_037_2127, w_037_2128, w_037_2129, w_037_2130, w_037_2131, w_037_2132, w_037_2133, w_037_2135, w_037_2136, w_037_2137, w_037_2139, w_037_2140, w_037_2141, w_037_2142, w_037_2143, w_037_2144, w_037_2146, w_037_2147, w_037_2148, w_037_2149, w_037_2152, w_037_2153, w_037_2154, w_037_2156, w_037_2157, w_037_2158, w_037_2159, w_037_2160, w_037_2163, w_037_2164, w_037_2165, w_037_2166, w_037_2167, w_037_2168, w_037_2169, w_037_2171, w_037_2173, w_037_2175, w_037_2176, w_037_2177, w_037_2178, w_037_2179, w_037_2180, w_037_2181, w_037_2182, w_037_2183, w_037_2184, w_037_2185, w_037_2187, w_037_2188, w_037_2189, w_037_2190, w_037_2191, w_037_2192, w_037_2193, w_037_2194, w_037_2195, w_037_2196, w_037_2197, w_037_2198, w_037_2199, w_037_2200, w_037_2201, w_037_2202, w_037_2203, w_037_2204, w_037_2205, w_037_2206, w_037_2207, w_037_2208, w_037_2209, w_037_2210, w_037_2211, w_037_2212, w_037_2213, w_037_2214, w_037_2215, w_037_2216, w_037_2217, w_037_2219, w_037_2220, w_037_2221, w_037_2222, w_037_2223, w_037_2224, w_037_2226, w_037_2227, w_037_2228, w_037_2229, w_037_2232, w_037_2233, w_037_2235, w_037_2236, w_037_2237, w_037_2238, w_037_2240, w_037_2241, w_037_2242, w_037_2243, w_037_2244, w_037_2245, w_037_2246, w_037_2247, w_037_2248, w_037_2250, w_037_2251, w_037_2252, w_037_2253, w_037_2254, w_037_2255, w_037_2256, w_037_2257, w_037_2258, w_037_2259, w_037_2260, w_037_2262, w_037_2264, w_037_2265, w_037_2266, w_037_2267, w_037_2271, w_037_2272, w_037_2273, w_037_2274, w_037_2276, w_037_2277, w_037_2279, w_037_2280, w_037_2282, w_037_2283, w_037_2286, w_037_2287, w_037_2288, w_037_2289, w_037_2290, w_037_2291, w_037_2293, w_037_2294, w_037_2295, w_037_2296, w_037_2297, w_037_2298, w_037_2299, w_037_2300, w_037_2301, w_037_2302, w_037_2303, w_037_2304, w_037_2305, w_037_2306, w_037_2307, w_037_2309, w_037_2310, w_037_2311, w_037_2312, w_037_2313, w_037_2314, w_037_2315, w_037_2316, w_037_2317, w_037_2318, w_037_2319, w_037_2320, w_037_2321, w_037_2322, w_037_2323, w_037_2324, w_037_2325, w_037_2326, w_037_2327, w_037_2328, w_037_2329, w_037_2331, w_037_2332, w_037_2333, w_037_2334, w_037_2337, w_037_2338, w_037_2339, w_037_2340, w_037_2341, w_037_2342, w_037_2343, w_037_2344, w_037_2346, w_037_2347, w_037_2348, w_037_2349, w_037_2350, w_037_2351, w_037_2352, w_037_2353, w_037_2354, w_037_2355, w_037_2356, w_037_2357, w_037_2358, w_037_2359, w_037_2360, w_037_2361, w_037_2362, w_037_2363, w_037_2364, w_037_2365, w_037_2366, w_037_2369, w_037_2370, w_037_2373, w_037_2374, w_037_2376, w_037_2379, w_037_2380, w_037_2382, w_037_2383, w_037_2384, w_037_2386, w_037_2387, w_037_2390, w_037_2391, w_037_2392, w_037_2393, w_037_2395, w_037_2397, w_037_2398, w_037_2399, w_037_2401, w_037_2402, w_037_2403, w_037_2405, w_037_2406, w_037_2407, w_037_2408, w_037_2410, w_037_2413, w_037_2415, w_037_2416, w_037_2417, w_037_2418, w_037_2419, w_037_2420, w_037_2421, w_037_2422, w_037_2425, w_037_2427, w_037_2428, w_037_2429, w_037_2434, w_037_2436, w_037_2437, w_037_2439, w_037_2441, w_037_2442, w_037_2444, w_037_2445, w_037_2446, w_037_2447, w_037_2448, w_037_2452, w_037_2455, w_037_2457, w_037_2458, w_037_2462, w_037_2463, w_037_2464, w_037_2466, w_037_2468, w_037_2470, w_037_2471, w_037_2472, w_037_2478, w_037_2479, w_037_2481, w_037_2482, w_037_2483, w_037_2488, w_037_2491, w_037_2492, w_037_2493, w_037_2495, w_037_2497, w_037_2498, w_037_2500, w_037_2502, w_037_2503, w_037_2504, w_037_2505, w_037_2506, w_037_2507, w_037_2508, w_037_2511, w_037_2512, w_037_2513, w_037_2514, w_037_2516, w_037_2519, w_037_2520, w_037_2521, w_037_2522, w_037_2523, w_037_2524, w_037_2526, w_037_2528, w_037_2530, w_037_2531, w_037_2537, w_037_2538, w_037_2540, w_037_2542, w_037_2544, w_037_2546, w_037_2547, w_037_2548, w_037_2554, w_037_2555, w_037_2557, w_037_2558, w_037_2559, w_037_2560, w_037_2563, w_037_2565, w_037_2566, w_037_2567, w_037_2568, w_037_2570, w_037_2571, w_037_2572, w_037_2573, w_037_2577, w_037_2580, w_037_2581, w_037_2584, w_037_2585, w_037_2586, w_037_2587, w_037_2588, w_037_2589, w_037_2593, w_037_2594, w_037_2595, w_037_2596, w_037_2598, w_037_2599, w_037_2601, w_037_2605, w_037_2606, w_037_2607, w_037_2608, w_037_2610, w_037_2611, w_037_2613, w_037_2616, w_037_2619, w_037_2621, w_037_2624, w_037_2629, w_037_2630, w_037_2632;
  wire w_038_000, w_038_001, w_038_002, w_038_003, w_038_004, w_038_005, w_038_006, w_038_007, w_038_008, w_038_009, w_038_010, w_038_011, w_038_012, w_038_013, w_038_014, w_038_015, w_038_016, w_038_017, w_038_018, w_038_019, w_038_020, w_038_021, w_038_022, w_038_023, w_038_024, w_038_025, w_038_026, w_038_027, w_038_028, w_038_029, w_038_030, w_038_031, w_038_032, w_038_033, w_038_034, w_038_035, w_038_036, w_038_037, w_038_038, w_038_039, w_038_040, w_038_041, w_038_042, w_038_043, w_038_044, w_038_045, w_038_046, w_038_047, w_038_048, w_038_049, w_038_050, w_038_051, w_038_052, w_038_053, w_038_054, w_038_055, w_038_057, w_038_058, w_038_059, w_038_060, w_038_062, w_038_063, w_038_064, w_038_065, w_038_066, w_038_067, w_038_068, w_038_069, w_038_070, w_038_073, w_038_074, w_038_075, w_038_076, w_038_077, w_038_078, w_038_079, w_038_080, w_038_081, w_038_082, w_038_083, w_038_084, w_038_085, w_038_086, w_038_088, w_038_089, w_038_090, w_038_092, w_038_094, w_038_095, w_038_096, w_038_098, w_038_099, w_038_100, w_038_101, w_038_102, w_038_103, w_038_104, w_038_105, w_038_106, w_038_107, w_038_108, w_038_109, w_038_110, w_038_111, w_038_112, w_038_113, w_038_114, w_038_115, w_038_116, w_038_117, w_038_118, w_038_119, w_038_120, w_038_121, w_038_122, w_038_123, w_038_124, w_038_125, w_038_126, w_038_127, w_038_128, w_038_129, w_038_130, w_038_131, w_038_132, w_038_133, w_038_134, w_038_135, w_038_136, w_038_137, w_038_138, w_038_139, w_038_140, w_038_141, w_038_142, w_038_143, w_038_144, w_038_145, w_038_146, w_038_147, w_038_148, w_038_149, w_038_150, w_038_151, w_038_152, w_038_153, w_038_154, w_038_155, w_038_156, w_038_157, w_038_158, w_038_159, w_038_160, w_038_161, w_038_162, w_038_163, w_038_164, w_038_165, w_038_166, w_038_167, w_038_168, w_038_169, w_038_170, w_038_171, w_038_172, w_038_173, w_038_174, w_038_175, w_038_176, w_038_177, w_038_178, w_038_179, w_038_181, w_038_182, w_038_183, w_038_184, w_038_186, w_038_187, w_038_188, w_038_189, w_038_190, w_038_191, w_038_192, w_038_193, w_038_194, w_038_196, w_038_197, w_038_198, w_038_199, w_038_200, w_038_201, w_038_202, w_038_203, w_038_204, w_038_205, w_038_206, w_038_207, w_038_208, w_038_209, w_038_210, w_038_211, w_038_212, w_038_213, w_038_214, w_038_215, w_038_216, w_038_217, w_038_218, w_038_219, w_038_221, w_038_222, w_038_223, w_038_224, w_038_225, w_038_226, w_038_227, w_038_229, w_038_230, w_038_231, w_038_232, w_038_233, w_038_234, w_038_235, w_038_236, w_038_237, w_038_238, w_038_240, w_038_241, w_038_242, w_038_243, w_038_244, w_038_245, w_038_246, w_038_248, w_038_249, w_038_250, w_038_251, w_038_253, w_038_254, w_038_255, w_038_256, w_038_257, w_038_258, w_038_259, w_038_260, w_038_261, w_038_262, w_038_263, w_038_264, w_038_265, w_038_266, w_038_267, w_038_268, w_038_269, w_038_270, w_038_271, w_038_272, w_038_273, w_038_274, w_038_275, w_038_276, w_038_277, w_038_278, w_038_279, w_038_280, w_038_281, w_038_283, w_038_284, w_038_285, w_038_286, w_038_287, w_038_288, w_038_289, w_038_290, w_038_291, w_038_292, w_038_293, w_038_294, w_038_295, w_038_296, w_038_297, w_038_298, w_038_299, w_038_300, w_038_302, w_038_303, w_038_304, w_038_305, w_038_306, w_038_307, w_038_308, w_038_309, w_038_310, w_038_311, w_038_312, w_038_313, w_038_314, w_038_315, w_038_316, w_038_317, w_038_318, w_038_319, w_038_320, w_038_321, w_038_322, w_038_323, w_038_324, w_038_326, w_038_327, w_038_328, w_038_330, w_038_331, w_038_332, w_038_333, w_038_335, w_038_336, w_038_337, w_038_338, w_038_339, w_038_340, w_038_341, w_038_342, w_038_343, w_038_344, w_038_345, w_038_346, w_038_348, w_038_349, w_038_350, w_038_351, w_038_352, w_038_354, w_038_355, w_038_356, w_038_357, w_038_358, w_038_359, w_038_360, w_038_361, w_038_362, w_038_363, w_038_364, w_038_365, w_038_366, w_038_367, w_038_368, w_038_369, w_038_370, w_038_371, w_038_372, w_038_373, w_038_374, w_038_375, w_038_376, w_038_377, w_038_378, w_038_379, w_038_380, w_038_381, w_038_382, w_038_383, w_038_384, w_038_385, w_038_386, w_038_387, w_038_388, w_038_389, w_038_390, w_038_391, w_038_392, w_038_393, w_038_394, w_038_395, w_038_396, w_038_397, w_038_398, w_038_399, w_038_400, w_038_401, w_038_402, w_038_403, w_038_404, w_038_405, w_038_406, w_038_407, w_038_408, w_038_409, w_038_410, w_038_411, w_038_412, w_038_413, w_038_414, w_038_415, w_038_416, w_038_417, w_038_418, w_038_419, w_038_420, w_038_421, w_038_422, w_038_423, w_038_424, w_038_425, w_038_426, w_038_427, w_038_428, w_038_429, w_038_430, w_038_431, w_038_432, w_038_433, w_038_434, w_038_435, w_038_436, w_038_437, w_038_438, w_038_439, w_038_440, w_038_441, w_038_442, w_038_443, w_038_444, w_038_445, w_038_447, w_038_448, w_038_449, w_038_451, w_038_452, w_038_453, w_038_454, w_038_455, w_038_456, w_038_457, w_038_458, w_038_459, w_038_460, w_038_461, w_038_462, w_038_463, w_038_464, w_038_465, w_038_466, w_038_467, w_038_468, w_038_469, w_038_470, w_038_471, w_038_473, w_038_474, w_038_475, w_038_476, w_038_477, w_038_478, w_038_479, w_038_480, w_038_481, w_038_482, w_038_483, w_038_484, w_038_485, w_038_486, w_038_487, w_038_488, w_038_489, w_038_490, w_038_491, w_038_492, w_038_493, w_038_494, w_038_495, w_038_496, w_038_497, w_038_498, w_038_499, w_038_500, w_038_501, w_038_502, w_038_503, w_038_504, w_038_505, w_038_506, w_038_507, w_038_508, w_038_509, w_038_510, w_038_511, w_038_513, w_038_515, w_038_516, w_038_517, w_038_518, w_038_519, w_038_520, w_038_521, w_038_522, w_038_523, w_038_524, w_038_525, w_038_526, w_038_527, w_038_528, w_038_529, w_038_530, w_038_531, w_038_532, w_038_533, w_038_534, w_038_535, w_038_537, w_038_538, w_038_539, w_038_540, w_038_541, w_038_542, w_038_543, w_038_544, w_038_545, w_038_546, w_038_547, w_038_548, w_038_549, w_038_550, w_038_551, w_038_552, w_038_554, w_038_555, w_038_556, w_038_557, w_038_558, w_038_559, w_038_560, w_038_561, w_038_562, w_038_563, w_038_564, w_038_565, w_038_566, w_038_567, w_038_568, w_038_569, w_038_570, w_038_571, w_038_572, w_038_573, w_038_574, w_038_575, w_038_576, w_038_577, w_038_578, w_038_579, w_038_580, w_038_581, w_038_582, w_038_585, w_038_586, w_038_587, w_038_588, w_038_589, w_038_590, w_038_592, w_038_597, w_038_598, w_038_599, w_038_600, w_038_601, w_038_602, w_038_603, w_038_605, w_038_606, w_038_607, w_038_608, w_038_609, w_038_610, w_038_611, w_038_612, w_038_613, w_038_614, w_038_615, w_038_616, w_038_617, w_038_618, w_038_619, w_038_620, w_038_621, w_038_622, w_038_623, w_038_624, w_038_625, w_038_626, w_038_627, w_038_628, w_038_629, w_038_630, w_038_631, w_038_632, w_038_633, w_038_634, w_038_636, w_038_637, w_038_638, w_038_639, w_038_640, w_038_641, w_038_642, w_038_643, w_038_644, w_038_645, w_038_646, w_038_647, w_038_648, w_038_649, w_038_650, w_038_651, w_038_652, w_038_653, w_038_654, w_038_655, w_038_657, w_038_658, w_038_659, w_038_660, w_038_661, w_038_662, w_038_663, w_038_664, w_038_665, w_038_666, w_038_667, w_038_668, w_038_669, w_038_670, w_038_671, w_038_672, w_038_673, w_038_675, w_038_676, w_038_677, w_038_678, w_038_679, w_038_680, w_038_681, w_038_683, w_038_684, w_038_685, w_038_686, w_038_687, w_038_688, w_038_689, w_038_690, w_038_691, w_038_693, w_038_694, w_038_695, w_038_696, w_038_697, w_038_698, w_038_699, w_038_700, w_038_701, w_038_702, w_038_703, w_038_704, w_038_705, w_038_706, w_038_707, w_038_708, w_038_709, w_038_710, w_038_712, w_038_713, w_038_714, w_038_715, w_038_717, w_038_718, w_038_719, w_038_720, w_038_721, w_038_722, w_038_723, w_038_724, w_038_727, w_038_728, w_038_729, w_038_730, w_038_731, w_038_732, w_038_733, w_038_734, w_038_735, w_038_736, w_038_737, w_038_738, w_038_739, w_038_740, w_038_741, w_038_742, w_038_743, w_038_744, w_038_745, w_038_746, w_038_747, w_038_748, w_038_749, w_038_750, w_038_751, w_038_752, w_038_753, w_038_754, w_038_755, w_038_756, w_038_757, w_038_758, w_038_760, w_038_761, w_038_762, w_038_764, w_038_766, w_038_767, w_038_768, w_038_769, w_038_770, w_038_771, w_038_772, w_038_773, w_038_774, w_038_775, w_038_777, w_038_778, w_038_779, w_038_781, w_038_782, w_038_783, w_038_784, w_038_785, w_038_786, w_038_787, w_038_788, w_038_789, w_038_790, w_038_791, w_038_792, w_038_794, w_038_795, w_038_796, w_038_797, w_038_798, w_038_799, w_038_800, w_038_801, w_038_802, w_038_803, w_038_804, w_038_805, w_038_807, w_038_808, w_038_809, w_038_810, w_038_811, w_038_812, w_038_813, w_038_814, w_038_815, w_038_816, w_038_817, w_038_818, w_038_819, w_038_820, w_038_821, w_038_822, w_038_823, w_038_824, w_038_825, w_038_826, w_038_827, w_038_828, w_038_829, w_038_830, w_038_831, w_038_832, w_038_833, w_038_834, w_038_835, w_038_836, w_038_837, w_038_838, w_038_839, w_038_840, w_038_842, w_038_843, w_038_844, w_038_845, w_038_846, w_038_847, w_038_848, w_038_849, w_038_850, w_038_851, w_038_852, w_038_853, w_038_854, w_038_855, w_038_856, w_038_857, w_038_858, w_038_859, w_038_860, w_038_861, w_038_862, w_038_863, w_038_864, w_038_865, w_038_866, w_038_867, w_038_868, w_038_869, w_038_870, w_038_871, w_038_872, w_038_873, w_038_874, w_038_875, w_038_876, w_038_878, w_038_879, w_038_880, w_038_881, w_038_882, w_038_883, w_038_884, w_038_885, w_038_886, w_038_887, w_038_888, w_038_889, w_038_890, w_038_891, w_038_892, w_038_893, w_038_894, w_038_895, w_038_896, w_038_897, w_038_898, w_038_899, w_038_900, w_038_901, w_038_902, w_038_904, w_038_905, w_038_906, w_038_908, w_038_909, w_038_910, w_038_911, w_038_912, w_038_914, w_038_915, w_038_916, w_038_918, w_038_919, w_038_920, w_038_921, w_038_922, w_038_923, w_038_924, w_038_925, w_038_926, w_038_927, w_038_928, w_038_929, w_038_930, w_038_931, w_038_932, w_038_933, w_038_935, w_038_936, w_038_937, w_038_938, w_038_939, w_038_940, w_038_941, w_038_942, w_038_943, w_038_945, w_038_946, w_038_947, w_038_948, w_038_949, w_038_950, w_038_951, w_038_952, w_038_954, w_038_955, w_038_956, w_038_959, w_038_960, w_038_961, w_038_962, w_038_963, w_038_965, w_038_966, w_038_967, w_038_968, w_038_969, w_038_970, w_038_971, w_038_972, w_038_973, w_038_974, w_038_975, w_038_976, w_038_977, w_038_978, w_038_979, w_038_980, w_038_981, w_038_982, w_038_983, w_038_984, w_038_985, w_038_987, w_038_988, w_038_989, w_038_990, w_038_991, w_038_992, w_038_993, w_038_995, w_038_996, w_038_997, w_038_998, w_038_999, w_038_1000, w_038_1001, w_038_1002, w_038_1004, w_038_1005, w_038_1006, w_038_1007, w_038_1008, w_038_1009, w_038_1010, w_038_1011, w_038_1012, w_038_1013, w_038_1014, w_038_1015, w_038_1016, w_038_1017, w_038_1018, w_038_1019, w_038_1020, w_038_1021, w_038_1022, w_038_1023, w_038_1024, w_038_1025, w_038_1026, w_038_1027, w_038_1028, w_038_1029, w_038_1030, w_038_1031, w_038_1032, w_038_1033, w_038_1034, w_038_1035, w_038_1036, w_038_1037, w_038_1038, w_038_1039, w_038_1040, w_038_1041, w_038_1043, w_038_1044, w_038_1045, w_038_1046, w_038_1047, w_038_1048, w_038_1049, w_038_1050, w_038_1051, w_038_1052, w_038_1053, w_038_1054, w_038_1055, w_038_1056, w_038_1057, w_038_1058, w_038_1059, w_038_1060, w_038_1061, w_038_1062, w_038_1063, w_038_1064, w_038_1065, w_038_1066, w_038_1067, w_038_1068, w_038_1069, w_038_1070, w_038_1071, w_038_1072, w_038_1073, w_038_1074, w_038_1075, w_038_1076, w_038_1077, w_038_1078, w_038_1079, w_038_1080, w_038_1081, w_038_1083, w_038_1084, w_038_1085, w_038_1086, w_038_1087, w_038_1088, w_038_1089, w_038_1090, w_038_1091, w_038_1092, w_038_1093, w_038_1094, w_038_1095, w_038_1096, w_038_1097, w_038_1098, w_038_1099, w_038_1100, w_038_1101, w_038_1104, w_038_1105, w_038_1106, w_038_1107, w_038_1108, w_038_1109, w_038_1110, w_038_1111, w_038_1112, w_038_1114, w_038_1115, w_038_1116, w_038_1117, w_038_1119, w_038_1120, w_038_1121, w_038_1122, w_038_1123, w_038_1124, w_038_1126, w_038_1127, w_038_1128, w_038_1129, w_038_1130, w_038_1131, w_038_1133, w_038_1134, w_038_1135, w_038_1136, w_038_1137, w_038_1138, w_038_1139, w_038_1140, w_038_1141, w_038_1142, w_038_1143, w_038_1144, w_038_1146, w_038_1148, w_038_1149, w_038_1150, w_038_1151, w_038_1152, w_038_1153, w_038_1155, w_038_1156, w_038_1157, w_038_1159, w_038_1160, w_038_1161, w_038_1162, w_038_1163, w_038_1164, w_038_1165, w_038_1166, w_038_1167, w_038_1168, w_038_1169, w_038_1171, w_038_1172, w_038_1173, w_038_1174, w_038_1175, w_038_1176, w_038_1177, w_038_1178, w_038_1179, w_038_1180, w_038_1182, w_038_1183, w_038_1184, w_038_1185, w_038_1186, w_038_1187, w_038_1188, w_038_1189, w_038_1190, w_038_1191, w_038_1192, w_038_1193, w_038_1194, w_038_1195, w_038_1197, w_038_1198, w_038_1199, w_038_1200, w_038_1201, w_038_1202, w_038_1203, w_038_1204, w_038_1205, w_038_1206, w_038_1207, w_038_1208, w_038_1209, w_038_1210, w_038_1211, w_038_1212, w_038_1213, w_038_1214, w_038_1215, w_038_1216, w_038_1217, w_038_1218, w_038_1219, w_038_1220, w_038_1221, w_038_1222, w_038_1223, w_038_1224, w_038_1225, w_038_1226, w_038_1228, w_038_1229, w_038_1230, w_038_1231, w_038_1232, w_038_1233, w_038_1234, w_038_1235, w_038_1236, w_038_1237, w_038_1238, w_038_1239, w_038_1240, w_038_1241, w_038_1242, w_038_1243, w_038_1244, w_038_1245, w_038_1246, w_038_1247, w_038_1248, w_038_1249, w_038_1250, w_038_1251, w_038_1252, w_038_1253, w_038_1254, w_038_1255, w_038_1257, w_038_1258, w_038_1260, w_038_1261, w_038_1262, w_038_1263, w_038_1264, w_038_1265, w_038_1266, w_038_1268, w_038_1269, w_038_1270, w_038_1271, w_038_1272, w_038_1273, w_038_1274, w_038_1275, w_038_1276, w_038_1278, w_038_1279, w_038_1280, w_038_1281, w_038_1282, w_038_1283, w_038_1284, w_038_1285, w_038_1286, w_038_1287, w_038_1291, w_038_1292, w_038_1293, w_038_1294, w_038_1295, w_038_1296, w_038_1297, w_038_1298, w_038_1299, w_038_1301, w_038_1303, w_038_1304, w_038_1306, w_038_1307, w_038_1308, w_038_1309, w_038_1310, w_038_1311, w_038_1312, w_038_1313, w_038_1314, w_038_1315, w_038_1316, w_038_1317, w_038_1318, w_038_1319, w_038_1320, w_038_1321, w_038_1322, w_038_1323, w_038_1324, w_038_1325, w_038_1326, w_038_1327, w_038_1328, w_038_1329, w_038_1330, w_038_1331, w_038_1332, w_038_1333, w_038_1335, w_038_1336, w_038_1337, w_038_1338, w_038_1339, w_038_1340, w_038_1341, w_038_1342, w_038_1343, w_038_1344, w_038_1345, w_038_1346, w_038_1347, w_038_1348, w_038_1349, w_038_1350, w_038_1351, w_038_1352, w_038_1353, w_038_1354, w_038_1355, w_038_1356, w_038_1358, w_038_1359, w_038_1360, w_038_1361, w_038_1362, w_038_1363, w_038_1364, w_038_1366, w_038_1367, w_038_1368, w_038_1369, w_038_1370, w_038_1371, w_038_1372, w_038_1373, w_038_1374, w_038_1375, w_038_1376, w_038_1377, w_038_1378, w_038_1379, w_038_1380, w_038_1381, w_038_1382, w_038_1383, w_038_1384, w_038_1385, w_038_1387, w_038_1388, w_038_1389, w_038_1390, w_038_1391, w_038_1392, w_038_1393, w_038_1394, w_038_1395, w_038_1396, w_038_1397, w_038_1398, w_038_1399, w_038_1400, w_038_1401, w_038_1402, w_038_1403, w_038_1404, w_038_1405, w_038_1406, w_038_1407, w_038_1408, w_038_1410, w_038_1411, w_038_1412, w_038_1413, w_038_1414, w_038_1415, w_038_1416, w_038_1417, w_038_1418, w_038_1419, w_038_1420, w_038_1421, w_038_1422, w_038_1423, w_038_1424, w_038_1425, w_038_1426, w_038_1428, w_038_1429, w_038_1430, w_038_1431, w_038_1432, w_038_1433, w_038_1434, w_038_1435, w_038_1437, w_038_1438, w_038_1439, w_038_1440, w_038_1441, w_038_1442, w_038_1443, w_038_1444, w_038_1445, w_038_1446, w_038_1447, w_038_1448, w_038_1449, w_038_1450, w_038_1451, w_038_1452, w_038_1454, w_038_1455, w_038_1456, w_038_1457, w_038_1458, w_038_1459, w_038_1460, w_038_1461, w_038_1462, w_038_1463, w_038_1464, w_038_1465, w_038_1466, w_038_1467, w_038_1468, w_038_1469, w_038_1470, w_038_1471, w_038_1472, w_038_1473, w_038_1474, w_038_1475, w_038_1476, w_038_1477, w_038_1478, w_038_1479, w_038_1480, w_038_1483, w_038_1484, w_038_1485, w_038_1486, w_038_1487, w_038_1488, w_038_1489, w_038_1490, w_038_1491, w_038_1492, w_038_1493, w_038_1494, w_038_1495, w_038_1496, w_038_1497, w_038_1498, w_038_1500, w_038_1501, w_038_1502, w_038_1503, w_038_1505, w_038_1506, w_038_1507, w_038_1508, w_038_1509, w_038_1511, w_038_1512, w_038_1514, w_038_1515, w_038_1516, w_038_1517, w_038_1518, w_038_1519, w_038_1520, w_038_1521, w_038_1522, w_038_1523, w_038_1524, w_038_1526, w_038_1527, w_038_1528, w_038_1531, w_038_1533, w_038_1534, w_038_1535, w_038_1536, w_038_1537, w_038_1538, w_038_1539, w_038_1540, w_038_1541, w_038_1542, w_038_1543, w_038_1544, w_038_1546, w_038_1547, w_038_1548, w_038_1549, w_038_1550, w_038_1551, w_038_1552, w_038_1553, w_038_1554, w_038_1555, w_038_1556, w_038_1558, w_038_1559, w_038_1561, w_038_1562, w_038_1563, w_038_1564, w_038_1565, w_038_1568, w_038_1569, w_038_1571, w_038_1572, w_038_1574, w_038_1575, w_038_1576, w_038_1577, w_038_1578, w_038_1579, w_038_1580, w_038_1581, w_038_1582, w_038_1584, w_038_1585, w_038_1586, w_038_1587, w_038_1588, w_038_1589, w_038_1590, w_038_1591, w_038_1592, w_038_1593, w_038_1594, w_038_1596, w_038_1597, w_038_1599, w_038_1600, w_038_1601, w_038_1602, w_038_1603, w_038_1604, w_038_1605, w_038_1606, w_038_1607, w_038_1608, w_038_1609, w_038_1610, w_038_1611, w_038_1612, w_038_1613, w_038_1614, w_038_1615, w_038_1616, w_038_1617, w_038_1619, w_038_1621, w_038_1622, w_038_1623, w_038_1625, w_038_1626, w_038_1627, w_038_1628, w_038_1629, w_038_1630, w_038_1631, w_038_1634, w_038_1635, w_038_1636, w_038_1637, w_038_1638, w_038_1639, w_038_1640, w_038_1641, w_038_1644, w_038_1645, w_038_1646, w_038_1647, w_038_1648, w_038_1649, w_038_1650, w_038_1651, w_038_1653, w_038_1657, w_038_1658, w_038_1659, w_038_1660, w_038_1661, w_038_1663, w_038_1665, w_038_1666, w_038_1667, w_038_1668, w_038_1669, w_038_1670, w_038_1671, w_038_1672, w_038_1673, w_038_1674, w_038_1675, w_038_1676, w_038_1677, w_038_1678, w_038_1679, w_038_1681, w_038_1682, w_038_1683, w_038_1684, w_038_1685, w_038_1686, w_038_1688, w_038_1690, w_038_1691, w_038_1692, w_038_1693, w_038_1695, w_038_1696, w_038_1697, w_038_1698, w_038_1699, w_038_1701, w_038_1702, w_038_1703, w_038_1704, w_038_1705, w_038_1706, w_038_1707, w_038_1708, w_038_1709, w_038_1710, w_038_1711, w_038_1712, w_038_1713, w_038_1714, w_038_1715, w_038_1716, w_038_1718, w_038_1719, w_038_1720, w_038_1722, w_038_1723, w_038_1724, w_038_1726, w_038_1727, w_038_1728, w_038_1729, w_038_1730, w_038_1732, w_038_1733, w_038_1735, w_038_1736, w_038_1737, w_038_1738, w_038_1741, w_038_1742, w_038_1743, w_038_1744, w_038_1745, w_038_1746, w_038_1747, w_038_1748, w_038_1749, w_038_1751, w_038_1753, w_038_1754, w_038_1755, w_038_1756, w_038_1757, w_038_1758, w_038_1759, w_038_1760, w_038_1761, w_038_1762, w_038_1763, w_038_1765;
  wire w_039_003, w_039_004, w_039_005, w_039_006, w_039_008, w_039_009, w_039_010, w_039_011, w_039_014, w_039_015, w_039_016, w_039_017, w_039_018, w_039_019, w_039_020, w_039_021, w_039_022, w_039_023, w_039_024, w_039_025, w_039_026, w_039_027, w_039_029, w_039_030, w_039_031, w_039_033, w_039_034, w_039_035, w_039_036, w_039_037, w_039_038, w_039_042, w_039_044, w_039_045, w_039_046, w_039_047, w_039_048, w_039_049, w_039_050, w_039_051, w_039_052, w_039_053, w_039_054, w_039_055, w_039_056, w_039_058, w_039_059, w_039_061, w_039_062, w_039_063, w_039_064, w_039_065, w_039_066, w_039_067, w_039_068, w_039_069, w_039_070, w_039_071, w_039_073, w_039_074, w_039_076, w_039_077, w_039_078, w_039_079, w_039_081, w_039_082, w_039_083, w_039_084, w_039_085, w_039_086, w_039_088, w_039_091, w_039_092, w_039_095, w_039_096, w_039_097, w_039_098, w_039_100, w_039_101, w_039_102, w_039_103, w_039_105, w_039_106, w_039_107, w_039_109, w_039_110, w_039_111, w_039_112, w_039_113, w_039_114, w_039_115, w_039_116, w_039_118, w_039_119, w_039_120, w_039_121, w_039_122, w_039_123, w_039_126, w_039_128, w_039_129, w_039_130, w_039_131, w_039_132, w_039_133, w_039_134, w_039_136, w_039_137, w_039_138, w_039_139, w_039_140, w_039_141, w_039_142, w_039_143, w_039_144, w_039_145, w_039_146, w_039_148, w_039_149, w_039_152, w_039_153, w_039_154, w_039_155, w_039_158, w_039_159, w_039_160, w_039_161, w_039_162, w_039_163, w_039_164, w_039_165, w_039_166, w_039_167, w_039_168, w_039_169, w_039_170, w_039_171, w_039_172, w_039_174, w_039_176, w_039_177, w_039_178, w_039_179, w_039_180, w_039_181, w_039_182, w_039_183, w_039_186, w_039_187, w_039_188, w_039_189, w_039_191, w_039_192, w_039_193, w_039_194, w_039_195, w_039_196, w_039_197, w_039_198, w_039_199, w_039_200, w_039_201, w_039_202, w_039_203, w_039_205, w_039_206, w_039_207, w_039_208, w_039_209, w_039_210, w_039_211, w_039_214, w_039_216, w_039_218, w_039_219, w_039_221, w_039_222, w_039_223, w_039_224, w_039_229, w_039_231, w_039_234, w_039_235, w_039_236, w_039_237, w_039_238, w_039_239, w_039_241, w_039_242, w_039_243, w_039_245, w_039_246, w_039_247, w_039_248, w_039_249, w_039_251, w_039_253, w_039_254, w_039_255, w_039_257, w_039_258, w_039_261, w_039_262, w_039_263, w_039_265, w_039_266, w_039_267, w_039_268, w_039_270, w_039_271, w_039_273, w_039_274, w_039_275, w_039_276, w_039_277, w_039_278, w_039_279, w_039_280, w_039_281, w_039_282, w_039_283, w_039_285, w_039_286, w_039_287, w_039_288, w_039_289, w_039_290, w_039_291, w_039_293, w_039_294, w_039_295, w_039_296, w_039_298, w_039_299, w_039_301, w_039_302, w_039_303, w_039_304, w_039_305, w_039_306, w_039_307, w_039_308, w_039_310, w_039_311, w_039_312, w_039_313, w_039_314, w_039_315, w_039_316, w_039_317, w_039_318, w_039_319, w_039_320, w_039_321, w_039_323, w_039_326, w_039_327, w_039_329, w_039_330, w_039_331, w_039_332, w_039_333, w_039_334, w_039_336, w_039_337, w_039_338, w_039_339, w_039_341, w_039_342, w_039_343, w_039_345, w_039_346, w_039_347, w_039_348, w_039_349, w_039_350, w_039_351, w_039_352, w_039_354, w_039_355, w_039_356, w_039_357, w_039_358, w_039_359, w_039_360, w_039_361, w_039_362, w_039_363, w_039_364, w_039_365, w_039_366, w_039_367, w_039_368, w_039_370, w_039_371, w_039_372, w_039_373, w_039_374, w_039_375, w_039_376, w_039_377, w_039_378, w_039_379, w_039_380, w_039_381, w_039_382, w_039_383, w_039_384, w_039_385, w_039_386, w_039_387, w_039_388, w_039_389, w_039_392, w_039_393, w_039_395, w_039_396, w_039_397, w_039_398, w_039_399, w_039_400, w_039_402, w_039_404, w_039_405, w_039_406, w_039_408, w_039_409, w_039_410, w_039_411, w_039_414, w_039_416, w_039_417, w_039_418, w_039_419, w_039_420, w_039_422, w_039_423, w_039_425, w_039_426, w_039_427, w_039_428, w_039_429, w_039_431, w_039_432, w_039_433, w_039_434, w_039_435, w_039_437, w_039_438, w_039_439, w_039_440, w_039_442, w_039_443, w_039_444, w_039_445, w_039_446, w_039_449, w_039_450, w_039_451, w_039_452, w_039_453, w_039_454, w_039_455, w_039_456, w_039_457, w_039_458, w_039_459, w_039_460, w_039_461, w_039_462, w_039_464, w_039_465, w_039_466, w_039_467, w_039_468, w_039_470, w_039_474, w_039_475, w_039_476, w_039_477, w_039_479, w_039_480, w_039_482, w_039_483, w_039_484, w_039_487, w_039_489, w_039_490, w_039_492, w_039_493, w_039_495, w_039_497, w_039_498, w_039_501, w_039_503, w_039_504, w_039_505, w_039_507, w_039_508, w_039_509, w_039_511, w_039_513, w_039_514, w_039_515, w_039_516, w_039_517, w_039_518, w_039_519, w_039_520, w_039_521, w_039_522, w_039_523, w_039_524, w_039_525, w_039_526, w_039_527, w_039_528, w_039_529, w_039_530, w_039_531, w_039_534, w_039_535, w_039_536, w_039_537, w_039_538, w_039_539, w_039_540, w_039_542, w_039_543, w_039_545, w_039_546, w_039_547, w_039_548, w_039_549, w_039_550, w_039_552, w_039_553, w_039_554, w_039_555, w_039_556, w_039_558, w_039_559, w_039_560, w_039_561, w_039_562, w_039_563, w_039_564, w_039_566, w_039_567, w_039_568, w_039_570, w_039_571, w_039_572, w_039_574, w_039_575, w_039_576, w_039_578, w_039_579, w_039_580, w_039_582, w_039_583, w_039_584, w_039_586, w_039_587, w_039_588, w_039_589, w_039_590, w_039_591, w_039_592, w_039_594, w_039_597, w_039_599, w_039_600, w_039_601, w_039_602, w_039_603, w_039_604, w_039_605, w_039_606, w_039_607, w_039_608, w_039_609, w_039_610, w_039_611, w_039_612, w_039_614, w_039_615, w_039_617, w_039_618, w_039_619, w_039_620, w_039_621, w_039_622, w_039_623, w_039_626, w_039_628, w_039_629, w_039_630, w_039_631, w_039_634, w_039_635, w_039_636, w_039_637, w_039_638, w_039_639, w_039_640, w_039_642, w_039_643, w_039_644, w_039_646, w_039_647, w_039_648, w_039_649, w_039_650, w_039_652, w_039_655, w_039_657, w_039_658, w_039_660, w_039_661, w_039_662, w_039_663, w_039_664, w_039_665, w_039_666, w_039_667, w_039_668, w_039_670, w_039_672, w_039_673, w_039_674, w_039_675, w_039_677, w_039_678, w_039_679, w_039_681, w_039_682, w_039_683, w_039_684, w_039_685, w_039_687, w_039_688, w_039_689, w_039_690, w_039_691, w_039_692, w_039_693, w_039_694, w_039_695, w_039_697, w_039_699, w_039_700, w_039_701, w_039_702, w_039_703, w_039_704, w_039_705, w_039_706, w_039_708, w_039_709, w_039_710, w_039_711, w_039_712, w_039_713, w_039_714, w_039_716, w_039_717, w_039_718, w_039_719, w_039_720, w_039_721, w_039_722, w_039_723, w_039_724, w_039_726, w_039_727, w_039_728, w_039_730, w_039_731, w_039_732, w_039_733, w_039_734, w_039_735, w_039_736, w_039_738, w_039_739, w_039_740, w_039_741, w_039_742, w_039_743, w_039_744, w_039_746, w_039_747, w_039_748, w_039_749, w_039_750, w_039_753, w_039_754, w_039_756, w_039_758, w_039_760, w_039_761, w_039_765, w_039_766, w_039_767, w_039_768, w_039_769, w_039_770, w_039_771, w_039_772, w_039_773, w_039_774, w_039_775, w_039_776, w_039_777, w_039_778, w_039_779, w_039_780, w_039_781, w_039_782, w_039_783, w_039_784, w_039_785, w_039_786, w_039_787, w_039_789, w_039_790, w_039_791, w_039_793, w_039_794, w_039_795, w_039_798, w_039_799, w_039_800, w_039_801, w_039_802, w_039_803, w_039_804, w_039_805, w_039_808, w_039_809, w_039_811, w_039_813, w_039_814, w_039_815, w_039_816, w_039_817, w_039_818, w_039_820, w_039_821, w_039_822, w_039_823, w_039_824, w_039_827, w_039_829, w_039_830, w_039_831, w_039_832, w_039_834, w_039_835, w_039_836, w_039_838, w_039_841, w_039_842, w_039_843, w_039_844, w_039_845, w_039_847, w_039_849, w_039_851, w_039_853, w_039_854, w_039_855, w_039_856, w_039_857, w_039_858, w_039_859, w_039_860, w_039_861, w_039_862, w_039_864, w_039_865, w_039_866, w_039_867, w_039_868, w_039_869, w_039_870, w_039_871, w_039_872, w_039_873, w_039_874, w_039_875, w_039_876, w_039_877, w_039_878, w_039_880, w_039_881, w_039_882, w_039_884, w_039_885, w_039_886, w_039_887, w_039_889, w_039_891, w_039_892, w_039_893, w_039_895, w_039_897, w_039_898, w_039_899, w_039_900, w_039_901, w_039_903, w_039_904, w_039_906, w_039_907, w_039_909, w_039_911, w_039_912, w_039_913, w_039_914, w_039_915, w_039_916, w_039_917, w_039_918, w_039_919, w_039_921, w_039_922, w_039_923, w_039_924, w_039_925, w_039_926, w_039_927, w_039_928, w_039_929, w_039_930, w_039_931, w_039_932, w_039_934, w_039_935, w_039_936, w_039_937, w_039_938, w_039_940, w_039_941, w_039_942, w_039_943, w_039_945, w_039_946, w_039_947, w_039_948, w_039_949, w_039_950, w_039_951, w_039_953, w_039_954, w_039_955, w_039_956, w_039_957, w_039_958, w_039_959, w_039_961, w_039_962, w_039_963, w_039_964, w_039_965, w_039_968, w_039_969, w_039_970, w_039_971, w_039_972, w_039_973, w_039_974, w_039_975, w_039_977, w_039_980, w_039_981, w_039_982, w_039_983, w_039_984, w_039_986, w_039_987, w_039_988, w_039_992, w_039_993, w_039_994, w_039_995, w_039_996, w_039_997, w_039_998, w_039_999, w_039_1000, w_039_1001, w_039_1003, w_039_1004, w_039_1005, w_039_1007, w_039_1009, w_039_1010, w_039_1013, w_039_1014, w_039_1015, w_039_1017, w_039_1018, w_039_1019, w_039_1020, w_039_1021, w_039_1022, w_039_1023, w_039_1024, w_039_1025, w_039_1026, w_039_1028, w_039_1029, w_039_1030, w_039_1031, w_039_1032, w_039_1033, w_039_1034, w_039_1035, w_039_1037, w_039_1038, w_039_1039, w_039_1040, w_039_1041, w_039_1042, w_039_1043, w_039_1044, w_039_1045, w_039_1046, w_039_1047, w_039_1048, w_039_1049, w_039_1050, w_039_1051, w_039_1052, w_039_1054, w_039_1055, w_039_1056, w_039_1058, w_039_1059, w_039_1061, w_039_1062, w_039_1063, w_039_1064, w_039_1065, w_039_1066, w_039_1067, w_039_1068, w_039_1069, w_039_1071, w_039_1072, w_039_1073, w_039_1074, w_039_1075, w_039_1076, w_039_1077, w_039_1078, w_039_1079, w_039_1081, w_039_1082, w_039_1084, w_039_1085, w_039_1087, w_039_1088, w_039_1089, w_039_1090, w_039_1091, w_039_1092, w_039_1093, w_039_1094, w_039_1096, w_039_1097, w_039_1098, w_039_1099, w_039_1100, w_039_1101, w_039_1102, w_039_1103, w_039_1104, w_039_1105, w_039_1106, w_039_1107, w_039_1108, w_039_1109, w_039_1110, w_039_1111, w_039_1112, w_039_1113, w_039_1114, w_039_1115, w_039_1116, w_039_1117, w_039_1118, w_039_1119, w_039_1120, w_039_1121, w_039_1122, w_039_1123, w_039_1124, w_039_1126, w_039_1127, w_039_1128, w_039_1129, w_039_1130, w_039_1131, w_039_1132, w_039_1133, w_039_1135, w_039_1136, w_039_1137, w_039_1138, w_039_1139, w_039_1140, w_039_1141, w_039_1142, w_039_1143, w_039_1144, w_039_1145, w_039_1146, w_039_1148, w_039_1149, w_039_1151, w_039_1152, w_039_1153, w_039_1154, w_039_1155, w_039_1157, w_039_1158, w_039_1159, w_039_1160, w_039_1161, w_039_1162, w_039_1163, w_039_1164, w_039_1165, w_039_1166, w_039_1167, w_039_1168, w_039_1169, w_039_1170, w_039_1171, w_039_1175, w_039_1176, w_039_1177, w_039_1178, w_039_1179, w_039_1180, w_039_1182, w_039_1185, w_039_1186, w_039_1187, w_039_1188, w_039_1189, w_039_1190, w_039_1192, w_039_1193, w_039_1194, w_039_1195, w_039_1196, w_039_1197, w_039_1198, w_039_1200, w_039_1201, w_039_1202, w_039_1203, w_039_1204, w_039_1205, w_039_1206, w_039_1207, w_039_1209, w_039_1211, w_039_1213, w_039_1214, w_039_1215, w_039_1216, w_039_1217, w_039_1219, w_039_1220, w_039_1221, w_039_1222, w_039_1223, w_039_1224, w_039_1225, w_039_1226, w_039_1227, w_039_1228, w_039_1229, w_039_1230, w_039_1231, w_039_1232, w_039_1233, w_039_1234, w_039_1235, w_039_1236, w_039_1237, w_039_1238, w_039_1239, w_039_1240, w_039_1241, w_039_1244, w_039_1246, w_039_1247, w_039_1248, w_039_1249, w_039_1250, w_039_1251, w_039_1253, w_039_1254, w_039_1255, w_039_1256, w_039_1257, w_039_1258, w_039_1259, w_039_1260, w_039_1261, w_039_1262, w_039_1263, w_039_1265, w_039_1266, w_039_1267, w_039_1268, w_039_1271, w_039_1272, w_039_1273, w_039_1274, w_039_1276, w_039_1277, w_039_1278, w_039_1279, w_039_1280, w_039_1283, w_039_1285, w_039_1286, w_039_1287, w_039_1288, w_039_1290, w_039_1291, w_039_1292, w_039_1293, w_039_1295, w_039_1297, w_039_1298, w_039_1299, w_039_1300, w_039_1301, w_039_1302, w_039_1303, w_039_1304, w_039_1305, w_039_1306, w_039_1307, w_039_1308, w_039_1309, w_039_1310, w_039_1311, w_039_1312, w_039_1313, w_039_1314, w_039_1315, w_039_1316, w_039_1317, w_039_1318, w_039_1319, w_039_1320, w_039_1321, w_039_1322, w_039_1323, w_039_1324, w_039_1325, w_039_1326, w_039_1328, w_039_1329, w_039_1330, w_039_1331, w_039_1332, w_039_1334, w_039_1338, w_039_1339, w_039_1340, w_039_1341, w_039_1342, w_039_1343, w_039_1344, w_039_1345, w_039_1346, w_039_1347, w_039_1348, w_039_1349, w_039_1350, w_039_1352, w_039_1354, w_039_1355, w_039_1357, w_039_1358, w_039_1359, w_039_1360, w_039_1361, w_039_1364, w_039_1365, w_039_1371, w_039_1374, w_039_1377, w_039_1379, w_039_1380, w_039_1381, w_039_1383, w_039_1385, w_039_1386, w_039_1388, w_039_1390, w_039_1393, w_039_1395, w_039_1396, w_039_1397, w_039_1398, w_039_1399, w_039_1401, w_039_1402, w_039_1403, w_039_1406, w_039_1410, w_039_1413, w_039_1414, w_039_1416, w_039_1418, w_039_1419, w_039_1422, w_039_1423, w_039_1426, w_039_1427, w_039_1431, w_039_1432, w_039_1433, w_039_1436, w_039_1437, w_039_1438, w_039_1439, w_039_1441, w_039_1442, w_039_1443, w_039_1444, w_039_1445, w_039_1448, w_039_1451, w_039_1452, w_039_1453, w_039_1454, w_039_1456, w_039_1457, w_039_1458, w_039_1460, w_039_1461, w_039_1462, w_039_1464, w_039_1465, w_039_1467, w_039_1468, w_039_1471, w_039_1473, w_039_1474, w_039_1476, w_039_1477, w_039_1481, w_039_1482, w_039_1483, w_039_1484, w_039_1486, w_039_1491, w_039_1492, w_039_1494, w_039_1495, w_039_1496, w_039_1497, w_039_1498, w_039_1501, w_039_1504, w_039_1508, w_039_1512, w_039_1513, w_039_1514, w_039_1515, w_039_1517, w_039_1518, w_039_1519, w_039_1521, w_039_1522, w_039_1523, w_039_1524, w_039_1525, w_039_1526, w_039_1530, w_039_1532, w_039_1534, w_039_1536, w_039_1539, w_039_1541, w_039_1542, w_039_1543, w_039_1545, w_039_1549, w_039_1550, w_039_1553, w_039_1554, w_039_1555, w_039_1556, w_039_1557, w_039_1558, w_039_1559, w_039_1565, w_039_1567, w_039_1569, w_039_1570, w_039_1573, w_039_1574, w_039_1575, w_039_1576, w_039_1577, w_039_1578, w_039_1579, w_039_1581, w_039_1586, w_039_1587, w_039_1588, w_039_1589, w_039_1596, w_039_1598, w_039_1599, w_039_1601, w_039_1602, w_039_1605, w_039_1610, w_039_1611, w_039_1612, w_039_1613, w_039_1616, w_039_1617, w_039_1618, w_039_1619, w_039_1620, w_039_1625, w_039_1627, w_039_1629, w_039_1630, w_039_1631, w_039_1632, w_039_1634, w_039_1635, w_039_1636, w_039_1637, w_039_1639, w_039_1640, w_039_1641, w_039_1642, w_039_1643, w_039_1644, w_039_1645, w_039_1646, w_039_1649, w_039_1650, w_039_1651, w_039_1652, w_039_1653, w_039_1654, w_039_1656, w_039_1659, w_039_1660, w_039_1661, w_039_1664, w_039_1667, w_039_1668, w_039_1676, w_039_1678, w_039_1681, w_039_1682, w_039_1684, w_039_1685, w_039_1686, w_039_1688, w_039_1691, w_039_1692, w_039_1696, w_039_1698, w_039_1702, w_039_1703, w_039_1705, w_039_1707, w_039_1708, w_039_1710, w_039_1711, w_039_1714, w_039_1715, w_039_1716, w_039_1726, w_039_1727, w_039_1729, w_039_1732, w_039_1733, w_039_1736, w_039_1737, w_039_1739, w_039_1740, w_039_1743, w_039_1744, w_039_1747, w_039_1749, w_039_1752, w_039_1753, w_039_1757, w_039_1758, w_039_1761, w_039_1764, w_039_1765, w_039_1766, w_039_1768, w_039_1770, w_039_1771, w_039_1772, w_039_1775, w_039_1779, w_039_1780, w_039_1781, w_039_1783, w_039_1784, w_039_1785, w_039_1786, w_039_1787, w_039_1788, w_039_1789, w_039_1790, w_039_1791, w_039_1792, w_039_1794, w_039_1795, w_039_1797, w_039_1798, w_039_1799, w_039_1800, w_039_1801, w_039_1802, w_039_1803, w_039_1804, w_039_1805, w_039_1806, w_039_1807, w_039_1810, w_039_1812, w_039_1813, w_039_1815, w_039_1816, w_039_1818, w_039_1822, w_039_1823, w_039_1824, w_039_1827, w_039_1830, w_039_1832, w_039_1836, w_039_1838, w_039_1839, w_039_1840, w_039_1841, w_039_1842, w_039_1843, w_039_1845, w_039_1846, w_039_1847, w_039_1848, w_039_1850, w_039_1855, w_039_1857, w_039_1858, w_039_1859, w_039_1864, w_039_1867, w_039_1872, w_039_1874, w_039_1878, w_039_1880, w_039_1881, w_039_1882, w_039_1884, w_039_1885, w_039_1887, w_039_1889, w_039_1890, w_039_1891, w_039_1892, w_039_1895, w_039_1897, w_039_1899, w_039_1900, w_039_1901, w_039_1902, w_039_1903, w_039_1904, w_039_1906, w_039_1907, w_039_1909, w_039_1910, w_039_1913, w_039_1914, w_039_1915, w_039_1916, w_039_1917, w_039_1918, w_039_1919, w_039_1921, w_039_1926, w_039_1928, w_039_1931, w_039_1932, w_039_1933, w_039_1934, w_039_1936, w_039_1938, w_039_1940, w_039_1942, w_039_1943, w_039_1944, w_039_1945, w_039_1947, w_039_1948, w_039_1949, w_039_1953, w_039_1956, w_039_1959, w_039_1961, w_039_1962, w_039_1963, w_039_1964, w_039_1965, w_039_1966, w_039_1971, w_039_1972, w_039_1973, w_039_1974, w_039_1976, w_039_1978, w_039_1979, w_039_1981, w_039_1982, w_039_1984, w_039_1985, w_039_1986, w_039_1988, w_039_1989, w_039_1991, w_039_1993, w_039_1995, w_039_1996, w_039_1998, w_039_2000, w_039_2003, w_039_2006, w_039_2010, w_039_2011, w_039_2012, w_039_2013, w_039_2015, w_039_2017, w_039_2019, w_039_2020, w_039_2023, w_039_2027, w_039_2029, w_039_2030, w_039_2031, w_039_2032, w_039_2034, w_039_2036, w_039_2038, w_039_2039, w_039_2040, w_039_2042, w_039_2045, w_039_2046, w_039_2047, w_039_2048, w_039_2050, w_039_2053, w_039_2054, w_039_2055, w_039_2056, w_039_2057, w_039_2058, w_039_2060, w_039_2064, w_039_2067, w_039_2068, w_039_2072, w_039_2073, w_039_2074, w_039_2076, w_039_2077, w_039_2079, w_039_2083, w_039_2084, w_039_2085, w_039_2087, w_039_2088, w_039_2089, w_039_2090, w_039_2091, w_039_2093, w_039_2095, w_039_2096, w_039_2098, w_039_2103, w_039_2104, w_039_2105, w_039_2107, w_039_2108, w_039_2111, w_039_2112, w_039_2114, w_039_2115, w_039_2116, w_039_2117, w_039_2118, w_039_2121, w_039_2122, w_039_2123, w_039_2124, w_039_2125, w_039_2126, w_039_2131, w_039_2133, w_039_2135, w_039_2136, w_039_2137, w_039_2140, w_039_2141, w_039_2142, w_039_2144, w_039_2145, w_039_2146, w_039_2148, w_039_2149, w_039_2150, w_039_2154, w_039_2157, w_039_2159, w_039_2160, w_039_2161, w_039_2162, w_039_2164, w_039_2165, w_039_2166, w_039_2167, w_039_2168, w_039_2169, w_039_2170, w_039_2171, w_039_2173, w_039_2174, w_039_2176, w_039_2178, w_039_2179, w_039_2180, w_039_2185, w_039_2187, w_039_2188, w_039_2189, w_039_2190, w_039_2192, w_039_2193, w_039_2195, w_039_2196, w_039_2197, w_039_2198, w_039_2199, w_039_2200, w_039_2201, w_039_2202, w_039_2205, w_039_2206, w_039_2207, w_039_2208, w_039_2209, w_039_2211, w_039_2215, w_039_2219, w_039_2223, w_039_2225, w_039_2228, w_039_2235, w_039_2236, w_039_2237, w_039_2238, w_039_2240, w_039_2241, w_039_2242, w_039_2246, w_039_2247, w_039_2249, w_039_2250, w_039_2253, w_039_2254, w_039_2256, w_039_2258, w_039_2259, w_039_2260, w_039_2261, w_039_2262, w_039_2264, w_039_2268, w_039_2270, w_039_2271, w_039_2273, w_039_2274, w_039_2275, w_039_2278, w_039_2279, w_039_2280, w_039_2281, w_039_2282, w_039_2288, w_039_2292, w_039_2293, w_039_2295, w_039_2297, w_039_2298, w_039_2299, w_039_2300, w_039_2305, w_039_2306, w_039_2307, w_039_2310, w_039_2311, w_039_2313, w_039_2314, w_039_2315, w_039_2316, w_039_2317, w_039_2320, w_039_2321, w_039_2322, w_039_2323, w_039_2325, w_039_2327, w_039_2329, w_039_2330, w_039_2332, w_039_2333, w_039_2337, w_039_2339, w_039_2340, w_039_2346, w_039_2348, w_039_2349, w_039_2350, w_039_2351, w_039_2352, w_039_2354, w_039_2355, w_039_2356, w_039_2357, w_039_2359, w_039_2360, w_039_2361, w_039_2362, w_039_2363, w_039_2364, w_039_2367, w_039_2368, w_039_2369, w_039_2370, w_039_2371, w_039_2372, w_039_2373, w_039_2374, w_039_2375, w_039_2376, w_039_2377, w_039_2378, w_039_2382, w_039_2383, w_039_2384, w_039_2385, w_039_2386, w_039_2387, w_039_2388, w_039_2389, w_039_2390, w_039_2391, w_039_2392, w_039_2393, w_039_2395, w_039_2397, w_039_2398, w_039_2399, w_039_2401, w_039_2402, w_039_2404, w_039_2408, w_039_2409, w_039_2410, w_039_2412, w_039_2413, w_039_2415, w_039_2416, w_039_2419, w_039_2420, w_039_2422, w_039_2423, w_039_2424, w_039_2425, w_039_2428, w_039_2429, w_039_2431, w_039_2432, w_039_2434, w_039_2435, w_039_2437, w_039_2439, w_039_2440, w_039_2441, w_039_2444, w_039_2445, w_039_2451, w_039_2453, w_039_2454, w_039_2457, w_039_2458, w_039_2460, w_039_2467, w_039_2472, w_039_2473, w_039_2474, w_039_2480, w_039_2481, w_039_2483, w_039_2485, w_039_2487, w_039_2488, w_039_2489, w_039_2491, w_039_2498, w_039_2501, w_039_2502, w_039_2503, w_039_2504, w_039_2505, w_039_2506, w_039_2507, w_039_2509, w_039_2510, w_039_2511, w_039_2512, w_039_2513, w_039_2514, w_039_2517, w_039_2518, w_039_2519, w_039_2521, w_039_2522, w_039_2523, w_039_2524, w_039_2525, w_039_2526, w_039_2528, w_039_2529, w_039_2530, w_039_2532, w_039_2534, w_039_2536, w_039_2538, w_039_2539, w_039_2540, w_039_2541, w_039_2542, w_039_2544, w_039_2545, w_039_2546, w_039_2547, w_039_2548, w_039_2549, w_039_2553, w_039_2555, w_039_2558, w_039_2559, w_039_2560, w_039_2562, w_039_2563, w_039_2570, w_039_2571, w_039_2572, w_039_2575, w_039_2576, w_039_2578, w_039_2581, w_039_2582, w_039_2584, w_039_2592, w_039_2593, w_039_2595, w_039_2597, w_039_2600, w_039_2601, w_039_2602, w_039_2605, w_039_2606, w_039_2610, w_039_2612, w_039_2616, w_039_2618, w_039_2621, w_039_2622, w_039_2623, w_039_2625, w_039_2626, w_039_2627, w_039_2628, w_039_2629, w_039_2630, w_039_2631, w_039_2633, w_039_2634, w_039_2637, w_039_2638, w_039_2639, w_039_2640, w_039_2641, w_039_2642, w_039_2643, w_039_2644, w_039_2646, w_039_2648, w_039_2650, w_039_2651, w_039_2652, w_039_2653, w_039_2655, w_039_2656, w_039_2657, w_039_2658, w_039_2659, w_039_2661, w_039_2663, w_039_2664, w_039_2665, w_039_2667, w_039_2673, w_039_2675, w_039_2676, w_039_2677, w_039_2678, w_039_2679, w_039_2681, w_039_2683, w_039_2684, w_039_2685, w_039_2686, w_039_2687, w_039_2688, w_039_2689, w_039_2691, w_039_2692, w_039_2693, w_039_2695, w_039_2699, w_039_2701, w_039_2703, w_039_2707, w_039_2708, w_039_2710, w_039_2713, w_039_2714, w_039_2717, w_039_2718, w_039_2719, w_039_2721, w_039_2723, w_039_2724, w_039_2726, w_039_2730, w_039_2735, w_039_2736, w_039_2739, w_039_2743, w_039_2744, w_039_2745, w_039_2747, w_039_2748, w_039_2750, w_039_2751, w_039_2752, w_039_2753, w_039_2754, w_039_2755, w_039_2757, w_039_2758, w_039_2759, w_039_2761, w_039_2762, w_039_2763, w_039_2764, w_039_2769, w_039_2770, w_039_2771, w_039_2773, w_039_2774, w_039_2775, w_039_2781, w_039_2786, w_039_2790, w_039_2792, w_039_2793, w_039_2794, w_039_2798, w_039_2800, w_039_2801, w_039_2802, w_039_2806, w_039_2809, w_039_2813, w_039_2814, w_039_2815, w_039_2816, w_039_2818, w_039_2819, w_039_2822, w_039_2826, w_039_2827, w_039_2829, w_039_2830, w_039_2832, w_039_2834, w_039_2836, w_039_2840, w_039_2842, w_039_2845, w_039_2846, w_039_2847, w_039_2848, w_039_2849, w_039_2851, w_039_2854, w_039_2857, w_039_2859, w_039_2861, w_039_2862, w_039_2863, w_039_2866, w_039_2867, w_039_2868, w_039_2869, w_039_2874, w_039_2875, w_039_2877, w_039_2878, w_039_2879, w_039_2880, w_039_2881, w_039_2883, w_039_2884, w_039_2888, w_039_2890, w_039_2896, w_039_2898, w_039_2901, w_039_2902, w_039_2903, w_039_2904, w_039_2907, w_039_2908, w_039_2909, w_039_2911, w_039_2912, w_039_2913, w_039_2914, w_039_2915, w_039_2916, w_039_2918, w_039_2921, w_039_2922, w_039_2924, w_039_2925, w_039_2926, w_039_2927, w_039_2928, w_039_2930, w_039_2932, w_039_2933, w_039_2935, w_039_2937, w_039_2938, w_039_2940, w_039_2941, w_039_2942, w_039_2948, w_039_2950, w_039_2951, w_039_2952, w_039_2953, w_039_2955, w_039_2961, w_039_2963, w_039_2964, w_039_2966, w_039_2969, w_039_2971, w_039_2972, w_039_2973, w_039_2975, w_039_2977, w_039_2978, w_039_2979, w_039_2980, w_039_2981, w_039_2982, w_039_2983, w_039_2985, w_039_2986, w_039_2987, w_039_2989, w_039_2992, w_039_2993, w_039_2996, w_039_2998, w_039_2999, w_039_3000, w_039_3001, w_039_3002, w_039_3007, w_039_3009, w_039_3017, w_039_3018, w_039_3019, w_039_3023, w_039_3024, w_039_3025, w_039_3026, w_039_3027, w_039_3028, w_039_3029, w_039_3030, w_039_3031, w_039_3032, w_039_3035, w_039_3037, w_039_3038, w_039_3039, w_039_3040, w_039_3044, w_039_3045, w_039_3046, w_039_3047, w_039_3050, w_039_3051, w_039_3052, w_039_3053, w_039_3054, w_039_3058, w_039_3059, w_039_3060, w_039_3061, w_039_3063, w_039_3064, w_039_3065, w_039_3066, w_039_3067, w_039_3070, w_039_3071, w_039_3072, w_039_3073, w_039_3076, w_039_3077, w_039_3079, w_039_3080, w_039_3082, w_039_3083, w_039_3084, w_039_3087, w_039_3088, w_039_3089, w_039_3090, w_039_3092, w_039_3094, w_039_3098, w_039_3099, w_039_3100, w_039_3101, w_039_3102, w_039_3104, w_039_3105, w_039_3107, w_039_3109, w_039_3112, w_039_3113, w_039_3115, w_039_3117, w_039_3118, w_039_3120, w_039_3122, w_039_3125, w_039_3126, w_039_3128, w_039_3129, w_039_3130, w_039_3132, w_039_3134, w_039_3135, w_039_3137, w_039_3139, w_039_3140, w_039_3142, w_039_3143, w_039_3144, w_039_3145, w_039_3147, w_039_3148, w_039_3149, w_039_3150, w_039_3151, w_039_3154, w_039_3155, w_039_3157, w_039_3159, w_039_3161, w_039_3162, w_039_3165, w_039_3167, w_039_3168, w_039_3169, w_039_3170, w_039_3171, w_039_3172, w_039_3175, w_039_3177, w_039_3178, w_039_3180, w_039_3181, w_039_3183, w_039_3185, w_039_3187, w_039_3188, w_039_3189, w_039_3190, w_039_3192, w_039_3193, w_039_3194, w_039_3195, w_039_3197, w_039_3198, w_039_3199, w_039_3202, w_039_3203, w_039_3207, w_039_3208, w_039_3215, w_039_3218, w_039_3220, w_039_3222, w_039_3223, w_039_3224, w_039_3226, w_039_3227, w_039_3228, w_039_3229, w_039_3230, w_039_3231, w_039_3232, w_039_3234, w_039_3235, w_039_3237, w_039_3238, w_039_3239, w_039_3240, w_039_3241, w_039_3243, w_039_3246, w_039_3247, w_039_3248, w_039_3249, w_039_3251, w_039_3253, w_039_3255, w_039_3256, w_039_3260, w_039_3261, w_039_3262, w_039_3263, w_039_3266, w_039_3267, w_039_3269, w_039_3270, w_039_3272, w_039_3273, w_039_3274, w_039_3275, w_039_3276, w_039_3278, w_039_3280, w_039_3283, w_039_3284, w_039_3285, w_039_3287, w_039_3289, w_039_3290, w_039_3291, w_039_3293, w_039_3294, w_039_3295, w_039_3296, w_039_3298, w_039_3299, w_039_3300, w_039_3301, w_039_3302, w_039_3303, w_039_3304, w_039_3305, w_039_3307, w_039_3308, w_039_3312, w_039_3314, w_039_3318, w_039_3320, w_039_3321, w_039_3322, w_039_3323, w_039_3325, w_039_3327, w_039_3328, w_039_3329, w_039_3331, w_039_3332, w_039_3333, w_039_3334, w_039_3336, w_039_3337, w_039_3339, w_039_3340, w_039_3341, w_039_3342, w_039_3343, w_039_3345, w_039_3347, w_039_3348, w_039_3349, w_039_3350, w_039_3352, w_039_3354, w_039_3357, w_039_3358, w_039_3359, w_039_3360, w_039_3361, w_039_3362, w_039_3365, w_039_3366, w_039_3369, w_039_3371, w_039_3372, w_039_3375, w_039_3376, w_039_3379, w_039_3381, w_039_3382, w_039_3384, w_039_3386, w_039_3387, w_039_3390, w_039_3392, w_039_3393, w_039_3396, w_039_3397, w_039_3400, w_039_3401, w_039_3402, w_039_3405, w_039_3406, w_039_3407, w_039_3409, w_039_3410, w_039_3414, w_039_3415, w_039_3416, w_039_3418, w_039_3419, w_039_3423, w_039_3424, w_039_3427, w_039_3428, w_039_3431, w_039_3436, w_039_3437, w_039_3438, w_039_3439, w_039_3441, w_039_3443, w_039_3444, w_039_3446, w_039_3447, w_039_3450, w_039_3451, w_039_3453, w_039_3454, w_039_3458, w_039_3459, w_039_3460, w_039_3461, w_039_3462, w_039_3465, w_039_3466, w_039_3467, w_039_3468, w_039_3469, w_039_3470, w_039_3474, w_039_3475, w_039_3476, w_039_3477, w_039_3479, w_039_3480, w_039_3482, w_039_3483, w_039_3484, w_039_3485, w_039_3489, w_039_3490, w_039_3492, w_039_3493, w_039_3494, w_039_3499, w_039_3503, w_039_3505, w_039_3506, w_039_3507, w_039_3508, w_039_3509, w_039_3512, w_039_3513, w_039_3514, w_039_3515, w_039_3518, w_039_3519, w_039_3521, w_039_3522, w_039_3523, w_039_3524, w_039_3525, w_039_3528, w_039_3530, w_039_3531, w_039_3532, w_039_3533, w_039_3534, w_039_3535, w_039_3536, w_039_3539, w_039_3540, w_039_3541, w_039_3544, w_039_3547, w_039_3549, w_039_3550, w_039_3551, w_039_3558, w_039_3559, w_039_3560, w_039_3562, w_039_3563, w_039_3566, w_039_3569, w_039_3572, w_039_3573, w_039_3574, w_039_3576, w_039_3577, w_039_3583, w_039_3584, w_039_3585, w_039_3586, w_039_3587, w_039_3589, w_039_3592, w_039_3594, w_039_3597, w_039_3598, w_039_3601, w_039_3602, w_039_3603, w_039_3605, w_039_3606, w_039_3609, w_039_3610, w_039_3611, w_039_3612, w_039_3613, w_039_3614, w_039_3615, w_039_3616, w_039_3617, w_039_3618, w_039_3620, w_039_3622, w_039_3623, w_039_3626, w_039_3627, w_039_3628, w_039_3629, w_039_3631, w_039_3633;
  wire w_040_000, w_040_001, w_040_002, w_040_003, w_040_004, w_040_005, w_040_006, w_040_007, w_040_008, w_040_009, w_040_010, w_040_011, w_040_012, w_040_013, w_040_014, w_040_016, w_040_017, w_040_018, w_040_019, w_040_020, w_040_021, w_040_022, w_040_023, w_040_025, w_040_027, w_040_029, w_040_030, w_040_031, w_040_032, w_040_033, w_040_034, w_040_035, w_040_036, w_040_037, w_040_038, w_040_039, w_040_040, w_040_042, w_040_043, w_040_045, w_040_046, w_040_047, w_040_048, w_040_049, w_040_050, w_040_051, w_040_052, w_040_054, w_040_055, w_040_056, w_040_057, w_040_059, w_040_060, w_040_061, w_040_062, w_040_063, w_040_064, w_040_065, w_040_066, w_040_067, w_040_068, w_040_069, w_040_070, w_040_072, w_040_074, w_040_075, w_040_076, w_040_077, w_040_078, w_040_080, w_040_081, w_040_082, w_040_083, w_040_084, w_040_085, w_040_086, w_040_088, w_040_089, w_040_090, w_040_091, w_040_092, w_040_093, w_040_094, w_040_095, w_040_097, w_040_101, w_040_102, w_040_104, w_040_105, w_040_106, w_040_107, w_040_108, w_040_109, w_040_110, w_040_112, w_040_113, w_040_114, w_040_115, w_040_116, w_040_117, w_040_118, w_040_119, w_040_120, w_040_121, w_040_122, w_040_124, w_040_125, w_040_126, w_040_127, w_040_128, w_040_129, w_040_130, w_040_131, w_040_132, w_040_133, w_040_134, w_040_135, w_040_136, w_040_137, w_040_139, w_040_140, w_040_141, w_040_143, w_040_144, w_040_145, w_040_146, w_040_147, w_040_148, w_040_150, w_040_151, w_040_153, w_040_154, w_040_155, w_040_157, w_040_158, w_040_160, w_040_162, w_040_165, w_040_166, w_040_167, w_040_168, w_040_169, w_040_170, w_040_172, w_040_174, w_040_175, w_040_176, w_040_177, w_040_178, w_040_179, w_040_180, w_040_181, w_040_182, w_040_183, w_040_184, w_040_185, w_040_186, w_040_187, w_040_188, w_040_189, w_040_190, w_040_191, w_040_192, w_040_193, w_040_195, w_040_196, w_040_198, w_040_199, w_040_200, w_040_201, w_040_202, w_040_203, w_040_204, w_040_205, w_040_206, w_040_207, w_040_209, w_040_211, w_040_212, w_040_213, w_040_216, w_040_217, w_040_218, w_040_220, w_040_221, w_040_222, w_040_224, w_040_225, w_040_227, w_040_230, w_040_231, w_040_233, w_040_234, w_040_235, w_040_236, w_040_238, w_040_240, w_040_241, w_040_243, w_040_244, w_040_245, w_040_247, w_040_248, w_040_251, w_040_252, w_040_253, w_040_254, w_040_255, w_040_256, w_040_257, w_040_258, w_040_259, w_040_260, w_040_261, w_040_262, w_040_263, w_040_264, w_040_266, w_040_267, w_040_269, w_040_270, w_040_271, w_040_272, w_040_274, w_040_275, w_040_276, w_040_277, w_040_279, w_040_280, w_040_281, w_040_285, w_040_286, w_040_288, w_040_290, w_040_291, w_040_293, w_040_294, w_040_295, w_040_296, w_040_297, w_040_298, w_040_300, w_040_301, w_040_302, w_040_303, w_040_304, w_040_305, w_040_306, w_040_307, w_040_309, w_040_310, w_040_312, w_040_313, w_040_314, w_040_315, w_040_316, w_040_317, w_040_318, w_040_319, w_040_321, w_040_324, w_040_325, w_040_326, w_040_327, w_040_328, w_040_330, w_040_331, w_040_332, w_040_333, w_040_334, w_040_335, w_040_336, w_040_337, w_040_338, w_040_339, w_040_340, w_040_342, w_040_343, w_040_344, w_040_345, w_040_346, w_040_347, w_040_349, w_040_350, w_040_351, w_040_352, w_040_353, w_040_354, w_040_355, w_040_356, w_040_357, w_040_359, w_040_360, w_040_361, w_040_362, w_040_363, w_040_364, w_040_365, w_040_366, w_040_368, w_040_371, w_040_373, w_040_374, w_040_375, w_040_377, w_040_378, w_040_380, w_040_381, w_040_382, w_040_383, w_040_385, w_040_386, w_040_387, w_040_389, w_040_390, w_040_391, w_040_392, w_040_393, w_040_394, w_040_395, w_040_397, w_040_398, w_040_399, w_040_400, w_040_401, w_040_403, w_040_406, w_040_407, w_040_408, w_040_409, w_040_410, w_040_413, w_040_414, w_040_415, w_040_416, w_040_417, w_040_419, w_040_420, w_040_422, w_040_423, w_040_424, w_040_426, w_040_427, w_040_428, w_040_429, w_040_432, w_040_433, w_040_434, w_040_436, w_040_438, w_040_441, w_040_442, w_040_443, w_040_444, w_040_445, w_040_446, w_040_447, w_040_448, w_040_449, w_040_450, w_040_451, w_040_454, w_040_456, w_040_457, w_040_458, w_040_459, w_040_460, w_040_462, w_040_463, w_040_464, w_040_465, w_040_466, w_040_467, w_040_468, w_040_469, w_040_470, w_040_471, w_040_472, w_040_473, w_040_474, w_040_475, w_040_476, w_040_477, w_040_478, w_040_479, w_040_480, w_040_483, w_040_484, w_040_485, w_040_486, w_040_487, w_040_489, w_040_490, w_040_491, w_040_492, w_040_493, w_040_494, w_040_496, w_040_497, w_040_500, w_040_501, w_040_502, w_040_503, w_040_504, w_040_505, w_040_506, w_040_508, w_040_509, w_040_510, w_040_511, w_040_512, w_040_513, w_040_515, w_040_518, w_040_519, w_040_520, w_040_521, w_040_523, w_040_524, w_040_525, w_040_526, w_040_528, w_040_529, w_040_530, w_040_531, w_040_532, w_040_533, w_040_535, w_040_536, w_040_537, w_040_538, w_040_539, w_040_540, w_040_542, w_040_543, w_040_544, w_040_545, w_040_546, w_040_547, w_040_548, w_040_549, w_040_550, w_040_552, w_040_553, w_040_554, w_040_555, w_040_559, w_040_560, w_040_561, w_040_562, w_040_563, w_040_564, w_040_565, w_040_566, w_040_567, w_040_568, w_040_570, w_040_571, w_040_572, w_040_574, w_040_575, w_040_576, w_040_577, w_040_578, w_040_579, w_040_580, w_040_581, w_040_582, w_040_584, w_040_587, w_040_590, w_040_591, w_040_592, w_040_593, w_040_594, w_040_595, w_040_597, w_040_598, w_040_599, w_040_600, w_040_601, w_040_602, w_040_603, w_040_604, w_040_605, w_040_606, w_040_607, w_040_609, w_040_610, w_040_614, w_040_615, w_040_616, w_040_617, w_040_618, w_040_620, w_040_621, w_040_622, w_040_623, w_040_624, w_040_626, w_040_629, w_040_631, w_040_633, w_040_634, w_040_635, w_040_636, w_040_637, w_040_638, w_040_639, w_040_640, w_040_641, w_040_643, w_040_645, w_040_646, w_040_647, w_040_649, w_040_651, w_040_652, w_040_653, w_040_654, w_040_657, w_040_658, w_040_659, w_040_660, w_040_663, w_040_664, w_040_665, w_040_666, w_040_667, w_040_668, w_040_669, w_040_670, w_040_671, w_040_673, w_040_674, w_040_676, w_040_677, w_040_678, w_040_679, w_040_680, w_040_681, w_040_682, w_040_683, w_040_684, w_040_685, w_040_686, w_040_687, w_040_688, w_040_690, w_040_691, w_040_692, w_040_693, w_040_694, w_040_695, w_040_696, w_040_697, w_040_698, w_040_700, w_040_701, w_040_702, w_040_703, w_040_704, w_040_705, w_040_706, w_040_708, w_040_709, w_040_710, w_040_712, w_040_715, w_040_716, w_040_717, w_040_719, w_040_720, w_040_721, w_040_722, w_040_723, w_040_725, w_040_726, w_040_728, w_040_729, w_040_730, w_040_731, w_040_732, w_040_733, w_040_735, w_040_736, w_040_737, w_040_738, w_040_739, w_040_740, w_040_741, w_040_743, w_040_744, w_040_745, w_040_747, w_040_749, w_040_750, w_040_752, w_040_753, w_040_754, w_040_755, w_040_756, w_040_758, w_040_759, w_040_760, w_040_761, w_040_762, w_040_763, w_040_764, w_040_766, w_040_767, w_040_768, w_040_769, w_040_770, w_040_771, w_040_773, w_040_774, w_040_775, w_040_776, w_040_777, w_040_778, w_040_779, w_040_780, w_040_781, w_040_782, w_040_783, w_040_784, w_040_786, w_040_787, w_040_788, w_040_789, w_040_790, w_040_791, w_040_792, w_040_793, w_040_795, w_040_796, w_040_797, w_040_798, w_040_799, w_040_800, w_040_801, w_040_802, w_040_805, w_040_806, w_040_809, w_040_810, w_040_811, w_040_812, w_040_813, w_040_814, w_040_817, w_040_818, w_040_819, w_040_820, w_040_822, w_040_825, w_040_826, w_040_827, w_040_828, w_040_830, w_040_831, w_040_832, w_040_833, w_040_835, w_040_836, w_040_837, w_040_838, w_040_839, w_040_840, w_040_841, w_040_842, w_040_843, w_040_844, w_040_845, w_040_846, w_040_848, w_040_850, w_040_852, w_040_853, w_040_854, w_040_855, w_040_856, w_040_857, w_040_858, w_040_860, w_040_861, w_040_862, w_040_863, w_040_864, w_040_865, w_040_866, w_040_867, w_040_868, w_040_869, w_040_870, w_040_871, w_040_872, w_040_873, w_040_875, w_040_876, w_040_877, w_040_878, w_040_880, w_040_882, w_040_884, w_040_885, w_040_886, w_040_887, w_040_888, w_040_889, w_040_890, w_040_891, w_040_892, w_040_893, w_040_895, w_040_896, w_040_897, w_040_898, w_040_899, w_040_900, w_040_901, w_040_902, w_040_903, w_040_904, w_040_905, w_040_907, w_040_908, w_040_909, w_040_911, w_040_912, w_040_913, w_040_914, w_040_915, w_040_916, w_040_917, w_040_918, w_040_919, w_040_920, w_040_921, w_040_922, w_040_923, w_040_924, w_040_925, w_040_928, w_040_929, w_040_930, w_040_931, w_040_933, w_040_934, w_040_935, w_040_936, w_040_937, w_040_938, w_040_939, w_040_940, w_040_941, w_040_942, w_040_944, w_040_945, w_040_946, w_040_948, w_040_949, w_040_951, w_040_952, w_040_953, w_040_954, w_040_955, w_040_956, w_040_959, w_040_960, w_040_961, w_040_962, w_040_964, w_040_965, w_040_966, w_040_967, w_040_970, w_040_971, w_040_972, w_040_973, w_040_974, w_040_975, w_040_976, w_040_977, w_040_980, w_040_981, w_040_982, w_040_983, w_040_984, w_040_985, w_040_986, w_040_988, w_040_989, w_040_990, w_040_991, w_040_992, w_040_993, w_040_994, w_040_995, w_040_997, w_040_998, w_040_999, w_040_1000, w_040_1001, w_040_1002, w_040_1003, w_040_1004, w_040_1005, w_040_1006, w_040_1007, w_040_1008, w_040_1009, w_040_1010, w_040_1013, w_040_1016, w_040_1017, w_040_1018, w_040_1019, w_040_1020, w_040_1021, w_040_1022, w_040_1023, w_040_1024, w_040_1025, w_040_1026, w_040_1027, w_040_1028, w_040_1029, w_040_1030, w_040_1033, w_040_1034, w_040_1035, w_040_1036, w_040_1037, w_040_1038, w_040_1039, w_040_1041, w_040_1042, w_040_1043, w_040_1044, w_040_1045, w_040_1046, w_040_1048, w_040_1049, w_040_1050, w_040_1051, w_040_1052, w_040_1054, w_040_1055, w_040_1056, w_040_1057, w_040_1058, w_040_1059, w_040_1060, w_040_1061, w_040_1062, w_040_1063, w_040_1065, w_040_1066, w_040_1067, w_040_1068, w_040_1069, w_040_1072, w_040_1073, w_040_1074, w_040_1075, w_040_1076, w_040_1077, w_040_1079, w_040_1080, w_040_1081, w_040_1082, w_040_1084, w_040_1085, w_040_1086, w_040_1087, w_040_1088, w_040_1089, w_040_1090, w_040_1091, w_040_1092, w_040_1093, w_040_1094, w_040_1095, w_040_1097, w_040_1098, w_040_1099, w_040_1100, w_040_1101, w_040_1103, w_040_1105, w_040_1106, w_040_1107, w_040_1108, w_040_1109, w_040_1112, w_040_1113, w_040_1114, w_040_1115, w_040_1116, w_040_1117, w_040_1118, w_040_1119, w_040_1120, w_040_1122, w_040_1123, w_040_1124, w_040_1125, w_040_1126, w_040_1127, w_040_1128, w_040_1129, w_040_1130, w_040_1131, w_040_1132, w_040_1133, w_040_1134, w_040_1135, w_040_1136, w_040_1137, w_040_1138, w_040_1140, w_040_1141, w_040_1142, w_040_1143, w_040_1144, w_040_1146, w_040_1148, w_040_1149, w_040_1150, w_040_1151, w_040_1152, w_040_1153, w_040_1154, w_040_1157, w_040_1158, w_040_1159, w_040_1160, w_040_1161, w_040_1162, w_040_1163, w_040_1164, w_040_1166, w_040_1168, w_040_1169, w_040_1171, w_040_1173, w_040_1174, w_040_1175, w_040_1176, w_040_1177, w_040_1178, w_040_1179, w_040_1180, w_040_1181, w_040_1182, w_040_1184, w_040_1185, w_040_1188, w_040_1190, w_040_1191, w_040_1192, w_040_1193, w_040_1194, w_040_1195, w_040_1196, w_040_1197, w_040_1198, w_040_1199, w_040_1200, w_040_1201, w_040_1202, w_040_1203, w_040_1204, w_040_1206, w_040_1207, w_040_1208, w_040_1210, w_040_1211, w_040_1212, w_040_1213, w_040_1214, w_040_1215, w_040_1216, w_040_1217, w_040_1218, w_040_1221, w_040_1222, w_040_1223, w_040_1224, w_040_1225, w_040_1227, w_040_1228, w_040_1229, w_040_1231, w_040_1232, w_040_1234, w_040_1235, w_040_1236, w_040_1237, w_040_1238, w_040_1239, w_040_1240, w_040_1241, w_040_1244, w_040_1245, w_040_1246, w_040_1247, w_040_1248, w_040_1249, w_040_1250, w_040_1253, w_040_1254, w_040_1255, w_040_1256, w_040_1259, w_040_1260, w_040_1261, w_040_1264, w_040_1266, w_040_1267, w_040_1269, w_040_1270, w_040_1272, w_040_1273, w_040_1274, w_040_1275, w_040_1277, w_040_1279, w_040_1280, w_040_1281, w_040_1282, w_040_1283, w_040_1284, w_040_1286, w_040_1287, w_040_1288, w_040_1289, w_040_1290, w_040_1292, w_040_1294, w_040_1295, w_040_1296, w_040_1297, w_040_1299, w_040_1300, w_040_1301, w_040_1302, w_040_1303, w_040_1305, w_040_1306, w_040_1307, w_040_1309, w_040_1310, w_040_1311, w_040_1312, w_040_1313, w_040_1314, w_040_1315, w_040_1316, w_040_1317, w_040_1318, w_040_1319, w_040_1320, w_040_1321, w_040_1322, w_040_1323, w_040_1324, w_040_1325, w_040_1326, w_040_1327, w_040_1329, w_040_1330, w_040_1331, w_040_1332, w_040_1333, w_040_1334, w_040_1335, w_040_1336, w_040_1338, w_040_1339, w_040_1341, w_040_1342, w_040_1343, w_040_1345, w_040_1348, w_040_1349, w_040_1350, w_040_1351, w_040_1352, w_040_1353, w_040_1354, w_040_1356, w_040_1358, w_040_1359, w_040_1360, w_040_1362, w_040_1363, w_040_1364, w_040_1365, w_040_1366, w_040_1367, w_040_1368, w_040_1369, w_040_1371, w_040_1372, w_040_1375, w_040_1376, w_040_1377, w_040_1378, w_040_1379, w_040_1380, w_040_1381, w_040_1382, w_040_1383, w_040_1384, w_040_1385, w_040_1386, w_040_1387, w_040_1388, w_040_1389, w_040_1390, w_040_1391, w_040_1392, w_040_1393, w_040_1396, w_040_1397, w_040_1399, w_040_1400, w_040_1401, w_040_1402, w_040_1403, w_040_1404, w_040_1405, w_040_1406, w_040_1408, w_040_1409, w_040_1411, w_040_1414, w_040_1417, w_040_1418, w_040_1419, w_040_1420, w_040_1422, w_040_1423, w_040_1424, w_040_1425, w_040_1426, w_040_1428, w_040_1429, w_040_1430, w_040_1431, w_040_1432, w_040_1433, w_040_1435, w_040_1436, w_040_1437, w_040_1439, w_040_1440, w_040_1441, w_040_1442, w_040_1443, w_040_1444, w_040_1445, w_040_1447, w_040_1448, w_040_1449, w_040_1450, w_040_1451, w_040_1452, w_040_1453, w_040_1454, w_040_1455, w_040_1456, w_040_1457, w_040_1458, w_040_1459, w_040_1460, w_040_1464, w_040_1465, w_040_1466, w_040_1468, w_040_1469, w_040_1470, w_040_1471, w_040_1472, w_040_1473, w_040_1474, w_040_1475, w_040_1476, w_040_1477, w_040_1478, w_040_1479, w_040_1480, w_040_1481, w_040_1482, w_040_1484, w_040_1485, w_040_1486, w_040_1487, w_040_1488, w_040_1490, w_040_1491, w_040_1492, w_040_1493, w_040_1494, w_040_1495, w_040_1496, w_040_1497, w_040_1498, w_040_1499, w_040_1501, w_040_1502, w_040_1503, w_040_1504, w_040_1505, w_040_1506, w_040_1507, w_040_1509, w_040_1510, w_040_1511, w_040_1512, w_040_1513, w_040_1514, w_040_1515, w_040_1516, w_040_1517, w_040_1518, w_040_1519, w_040_1520, w_040_1522, w_040_1524, w_040_1525, w_040_1526, w_040_1527, w_040_1528, w_040_1530, w_040_1531, w_040_1532, w_040_1533, w_040_1534, w_040_1536, w_040_1537, w_040_1538, w_040_1539, w_040_1540, w_040_1542, w_040_1544, w_040_1545, w_040_1547, w_040_1548, w_040_1549, w_040_1550, w_040_1551, w_040_1552, w_040_1554, w_040_1556, w_040_1557, w_040_1558, w_040_1559, w_040_1560, w_040_1561, w_040_1562, w_040_1563, w_040_1564, w_040_1567, w_040_1568, w_040_1570, w_040_1571, w_040_1572, w_040_1573, w_040_1575, w_040_1576, w_040_1577, w_040_1578, w_040_1579, w_040_1580, w_040_1581, w_040_1582, w_040_1583, w_040_1584, w_040_1585, w_040_1586, w_040_1587, w_040_1588, w_040_1589, w_040_1590, w_040_1591, w_040_1593, w_040_1594, w_040_1596, w_040_1598, w_040_1600, w_040_1601, w_040_1603, w_040_1605, w_040_1606, w_040_1607, w_040_1609, w_040_1611, w_040_1612, w_040_1613, w_040_1614, w_040_1615, w_040_1616, w_040_1617, w_040_1618, w_040_1619, w_040_1621, w_040_1623, w_040_1625, w_040_1627, w_040_1628, w_040_1630, w_040_1631, w_040_1632, w_040_1633, w_040_1634, w_040_1635, w_040_1636, w_040_1637, w_040_1638, w_040_1639, w_040_1640, w_040_1642, w_040_1643, w_040_1644, w_040_1648, w_040_1652, w_040_1654, w_040_1655, w_040_1656, w_040_1657, w_040_1658, w_040_1659, w_040_1660, w_040_1661, w_040_1662, w_040_1663, w_040_1664, w_040_1665, w_040_1666, w_040_1668, w_040_1671, w_040_1672, w_040_1673, w_040_1674, w_040_1675, w_040_1676, w_040_1677, w_040_1678, w_040_1681, w_040_1682, w_040_1683, w_040_1684, w_040_1685, w_040_1687, w_040_1688, w_040_1689, w_040_1690, w_040_1691, w_040_1694, w_040_1695, w_040_1696, w_040_1697, w_040_1698, w_040_1699, w_040_1700, w_040_1701, w_040_1702, w_040_1703, w_040_1704, w_040_1705, w_040_1706, w_040_1707, w_040_1709, w_040_1710, w_040_1711, w_040_1712, w_040_1713, w_040_1714, w_040_1715, w_040_1716, w_040_1717, w_040_1718, w_040_1719, w_040_1720, w_040_1722, w_040_1723, w_040_1725, w_040_1726, w_040_1727, w_040_1729, w_040_1730, w_040_1731, w_040_1732, w_040_1733, w_040_1734, w_040_1735, w_040_1736, w_040_1737, w_040_1738, w_040_1739, w_040_1740, w_040_1743, w_040_1744, w_040_1745, w_040_1746, w_040_1747, w_040_1749, w_040_1752, w_040_1753, w_040_1754, w_040_1755, w_040_1756, w_040_1758, w_040_1759, w_040_1761, w_040_1763, w_040_1764, w_040_1765, w_040_1766, w_040_1767, w_040_1768, w_040_1771, w_040_1772, w_040_1773, w_040_1774, w_040_1775, w_040_1776, w_040_1777, w_040_1778, w_040_1779, w_040_1780, w_040_1781, w_040_1782, w_040_1783, w_040_1784, w_040_1785, w_040_1786, w_040_1787, w_040_1788, w_040_1789, w_040_1790, w_040_1791, w_040_1792, w_040_1793, w_040_1794, w_040_1795, w_040_1796, w_040_1797, w_040_1798, w_040_1799, w_040_1800, w_040_1802, w_040_1803, w_040_1805, w_040_1806, w_040_1808, w_040_1809, w_040_1810, w_040_1812, w_040_1813, w_040_1814, w_040_1815, w_040_1816, w_040_1817, w_040_1818, w_040_1819, w_040_1820, w_040_1821, w_040_1822, w_040_1823, w_040_1824, w_040_1825, w_040_1826, w_040_1828, w_040_1829, w_040_1831, w_040_1833, w_040_1834, w_040_1835, w_040_1836, w_040_1837, w_040_1839, w_040_1840, w_040_1842, w_040_1843, w_040_1844, w_040_1846, w_040_1847, w_040_1849, w_040_1850, w_040_1851, w_040_1852, w_040_1853, w_040_1855, w_040_1856, w_040_1857, w_040_1858, w_040_1859, w_040_1860, w_040_1861, w_040_1862, w_040_1864, w_040_1865, w_040_1866, w_040_1867, w_040_1868, w_040_1869, w_040_1870, w_040_1871, w_040_1872, w_040_1873, w_040_1874, w_040_1875, w_040_1876, w_040_1878, w_040_1879, w_040_1881, w_040_1882, w_040_1883, w_040_1884, w_040_1887, w_040_1888, w_040_1889, w_040_1890, w_040_1891, w_040_1892, w_040_1893, w_040_1894, w_040_1895, w_040_1897, w_040_1898, w_040_1900, w_040_1901, w_040_1903, w_040_1904, w_040_1905, w_040_1906, w_040_1907, w_040_1908, w_040_1909, w_040_1910, w_040_1911, w_040_1913, w_040_1914, w_040_1915, w_040_1916, w_040_1919, w_040_1920, w_040_1921, w_040_1923, w_040_1924, w_040_1925, w_040_1926, w_040_1927, w_040_1928, w_040_1930, w_040_1931, w_040_1932, w_040_1933, w_040_1934, w_040_1937, w_040_1938, w_040_1939, w_040_1940, w_040_1941, w_040_1943, w_040_1945, w_040_1946, w_040_1947, w_040_1950, w_040_1951, w_040_1954, w_040_1955, w_040_1958, w_040_1959, w_040_1960, w_040_1962, w_040_1963, w_040_1964, w_040_1965, w_040_1966, w_040_1967, w_040_1968, w_040_1969, w_040_1970, w_040_1971, w_040_1972, w_040_1973, w_040_1974, w_040_1975, w_040_1976, w_040_1977, w_040_1979, w_040_1981, w_040_1982, w_040_1984, w_040_1985, w_040_1986, w_040_1987, w_040_1989, w_040_1990, w_040_1991, w_040_1992, w_040_1993, w_040_1995, w_040_1996, w_040_1997, w_040_1998, w_040_2000, w_040_2001, w_040_2003, w_040_2004, w_040_2005, w_040_2006, w_040_2008, w_040_2009, w_040_2010, w_040_2011, w_040_2012, w_040_2014, w_040_2016, w_040_2017, w_040_2018, w_040_2019, w_040_2020, w_040_2021, w_040_2022, w_040_2023, w_040_2024, w_040_2025, w_040_2027, w_040_2028, w_040_2029, w_040_2031, w_040_2032, w_040_2033, w_040_2034, w_040_2035, w_040_2038, w_040_2039, w_040_2040, w_040_2041, w_040_2042, w_040_2043, w_040_2044, w_040_2045, w_040_2046, w_040_2047, w_040_2049, w_040_2050, w_040_2051, w_040_2053, w_040_2054, w_040_2055, w_040_2056, w_040_2057, w_040_2058, w_040_2059, w_040_2062, w_040_2063, w_040_2064, w_040_2065, w_040_2066, w_040_2067, w_040_2068, w_040_2069, w_040_2071, w_040_2072, w_040_2073, w_040_2074, w_040_2075, w_040_2076, w_040_2078, w_040_2080, w_040_2081, w_040_2083, w_040_2084, w_040_2085, w_040_2086, w_040_2087, w_040_2088, w_040_2089, w_040_2090, w_040_2091, w_040_2093, w_040_2094, w_040_2095, w_040_2096, w_040_2097, w_040_2098, w_040_2100, w_040_2101, w_040_2102, w_040_2103, w_040_2104, w_040_2106, w_040_2107, w_040_2108, w_040_2109, w_040_2110, w_040_2111, w_040_2112, w_040_2113, w_040_2114, w_040_2116, w_040_2118, w_040_2119, w_040_2121, w_040_2123, w_040_2124, w_040_2129, w_040_2131, w_040_2132, w_040_2133, w_040_2135, w_040_2136, w_040_2137, w_040_2139, w_040_2142, w_040_2144, w_040_2145, w_040_2147, w_040_2149, w_040_2150, w_040_2151, w_040_2153, w_040_2155, w_040_2156, w_040_2158, w_040_2160, w_040_2161, w_040_2162, w_040_2163, w_040_2165, w_040_2166, w_040_2169, w_040_2170, w_040_2172, w_040_2175, w_040_2177, w_040_2178, w_040_2181, w_040_2182, w_040_2185, w_040_2186, w_040_2188, w_040_2189, w_040_2190, w_040_2191, w_040_2192, w_040_2193, w_040_2197, w_040_2199, w_040_2203, w_040_2205, w_040_2207, w_040_2208, w_040_2209, w_040_2210, w_040_2212, w_040_2213, w_040_2214, w_040_2215, w_040_2216, w_040_2220, w_040_2222, w_040_2226, w_040_2227, w_040_2228, w_040_2229, w_040_2230, w_040_2231, w_040_2232, w_040_2233, w_040_2236, w_040_2237, w_040_2238, w_040_2239, w_040_2241, w_040_2246, w_040_2247, w_040_2248, w_040_2252, w_040_2253, w_040_2254, w_040_2255, w_040_2256, w_040_2257, w_040_2259, w_040_2261, w_040_2262, w_040_2263, w_040_2266, w_040_2268, w_040_2270, w_040_2271, w_040_2272, w_040_2273, w_040_2276, w_040_2277, w_040_2278, w_040_2279, w_040_2280, w_040_2283, w_040_2284, w_040_2285, w_040_2286, w_040_2287, w_040_2288, w_040_2290, w_040_2291, w_040_2295, w_040_2299, w_040_2300, w_040_2302, w_040_2304, w_040_2305, w_040_2309, w_040_2310, w_040_2313, w_040_2315, w_040_2317, w_040_2318, w_040_2321, w_040_2323, w_040_2325, w_040_2326, w_040_2327, w_040_2328, w_040_2330, w_040_2332, w_040_2334, w_040_2335, w_040_2337, w_040_2339, w_040_2340, w_040_2341, w_040_2342, w_040_2343, w_040_2345, w_040_2347, w_040_2350, w_040_2352, w_040_2353, w_040_2354, w_040_2355, w_040_2356, w_040_2357, w_040_2359, w_040_2361, w_040_2365, w_040_2367, w_040_2368, w_040_2369, w_040_2370, w_040_2375, w_040_2376, w_040_2377, w_040_2382, w_040_2386, w_040_2387, w_040_2388, w_040_2389, w_040_2390, w_040_2391, w_040_2392, w_040_2395, w_040_2396, w_040_2397, w_040_2400, w_040_2401, w_040_2404, w_040_2405, w_040_2408, w_040_2409, w_040_2410, w_040_2411, w_040_2412, w_040_2413, w_040_2414, w_040_2415, w_040_2416, w_040_2418, w_040_2420, w_040_2424, w_040_2426, w_040_2429, w_040_2430, w_040_2433, w_040_2435, w_040_2436, w_040_2438, w_040_2440, w_040_2442, w_040_2445, w_040_2448, w_040_2453, w_040_2455, w_040_2457, w_040_2458, w_040_2459, w_040_2460, w_040_2461, w_040_2463, w_040_2465, w_040_2466, w_040_2468, w_040_2472, w_040_2473, w_040_2474, w_040_2476, w_040_2477, w_040_2478, w_040_2480, w_040_2483, w_040_2484, w_040_2487, w_040_2491, w_040_2492, w_040_2493, w_040_2495, w_040_2497, w_040_2501, w_040_2502, w_040_2503, w_040_2506, w_040_2510, w_040_2511, w_040_2512, w_040_2513, w_040_2514, w_040_2515, w_040_2516, w_040_2517, w_040_2518, w_040_2519, w_040_2522, w_040_2523, w_040_2526, w_040_2527, w_040_2530, w_040_2531, w_040_2533, w_040_2534, w_040_2535, w_040_2536, w_040_2539, w_040_2540, w_040_2545, w_040_2550, w_040_2551, w_040_2554, w_040_2555, w_040_2556, w_040_2557, w_040_2558, w_040_2560, w_040_2561, w_040_2563, w_040_2566, w_040_2568, w_040_2569, w_040_2570, w_040_2574, w_040_2575, w_040_2577, w_040_2578, w_040_2579, w_040_2580, w_040_2581, w_040_2584, w_040_2585, w_040_2589, w_040_2590, w_040_2591, w_040_2596, w_040_2597, w_040_2598, w_040_2599, w_040_2600, w_040_2601, w_040_2608, w_040_2609, w_040_2613, w_040_2615, w_040_2618, w_040_2619, w_040_2620, w_040_2621, w_040_2622, w_040_2624, w_040_2626, w_040_2627, w_040_2628, w_040_2629, w_040_2632, w_040_2633, w_040_2634, w_040_2635, w_040_2636, w_040_2637, w_040_2639, w_040_2642, w_040_2643, w_040_2645, w_040_2646, w_040_2648, w_040_2649, w_040_2650, w_040_2651, w_040_2655, w_040_2657, w_040_2659, w_040_2663, w_040_2665, w_040_2667, w_040_2668, w_040_2669, w_040_2671, w_040_2673, w_040_2674, w_040_2677, w_040_2678, w_040_2679, w_040_2681, w_040_2682, w_040_2686, w_040_2687, w_040_2688, w_040_2691, w_040_2692, w_040_2693, w_040_2694, w_040_2696, w_040_2699, w_040_2703, w_040_2704, w_040_2705, w_040_2707, w_040_2708, w_040_2709, w_040_2710, w_040_2711, w_040_2712, w_040_2713, w_040_2715, w_040_2716, w_040_2717, w_040_2721, w_040_2722, w_040_2723, w_040_2727, w_040_2729, w_040_2731, w_040_2732, w_040_2737, w_040_2739, w_040_2741, w_040_2743, w_040_2745, w_040_2748, w_040_2749, w_040_2753, w_040_2754, w_040_2756, w_040_2759, w_040_2761, w_040_2763, w_040_2765, w_040_2771, w_040_2773, w_040_2777, w_040_2778, w_040_2780, w_040_2782, w_040_2783, w_040_2785, w_040_2786, w_040_2787, w_040_2789, w_040_2790, w_040_2792, w_040_2793, w_040_2795, w_040_2796, w_040_2797, w_040_2798, w_040_2801, w_040_2802, w_040_2803, w_040_2804, w_040_2805, w_040_2806, w_040_2809, w_040_2811, w_040_2813, w_040_2814, w_040_2815, w_040_2817, w_040_2818, w_040_2819, w_040_2820, w_040_2821, w_040_2822, w_040_2823, w_040_2824, w_040_2825, w_040_2827, w_040_2828, w_040_2830, w_040_2831, w_040_2832, w_040_2833, w_040_2834, w_040_2835, w_040_2841, w_040_2842, w_040_2843, w_040_2845, w_040_2846, w_040_2848, w_040_2852, w_040_2853, w_040_2855, w_040_2856, w_040_2857, w_040_2858, w_040_2859, w_040_2860, w_040_2861, w_040_2862, w_040_2864, w_040_2865, w_040_2866, w_040_2867, w_040_2868, w_040_2869, w_040_2871, w_040_2872, w_040_2876, w_040_2878, w_040_2880, w_040_2881, w_040_2882, w_040_2883, w_040_2884, w_040_2885, w_040_2886, w_040_2889, w_040_2890, w_040_2891, w_040_2893, w_040_2895, w_040_2896, w_040_2897, w_040_2898, w_040_2899, w_040_2900, w_040_2901, w_040_2902, w_040_2903, w_040_2904, w_040_2905, w_040_2906, w_040_2908;
  wire w_041_000, w_041_001, w_041_002, w_041_003, w_041_004, w_041_005, w_041_006, w_041_007, w_041_008, w_041_009, w_041_010, w_041_011, w_041_012, w_041_013, w_041_015, w_041_016, w_041_017, w_041_019, w_041_020, w_041_021, w_041_022, w_041_023, w_041_024, w_041_025, w_041_026, w_041_027, w_041_028, w_041_029, w_041_030, w_041_031, w_041_032, w_041_033, w_041_035, w_041_036, w_041_037, w_041_038, w_041_039, w_041_040, w_041_041, w_041_043, w_041_044, w_041_047, w_041_049, w_041_050, w_041_051, w_041_053, w_041_056, w_041_058, w_041_059, w_041_060, w_041_061, w_041_062, w_041_063, w_041_064, w_041_065, w_041_066, w_041_067, w_041_069, w_041_070, w_041_071, w_041_073, w_041_074, w_041_075, w_041_076, w_041_077, w_041_080, w_041_081, w_041_082, w_041_083, w_041_084, w_041_085, w_041_086, w_041_087, w_041_088, w_041_089, w_041_090, w_041_091, w_041_092, w_041_095, w_041_097, w_041_098, w_041_099, w_041_100, w_041_101, w_041_103, w_041_104, w_041_105, w_041_106, w_041_107, w_041_109, w_041_110, w_041_112, w_041_113, w_041_114, w_041_116, w_041_117, w_041_118, w_041_119, w_041_120, w_041_121, w_041_122, w_041_123, w_041_124, w_041_126, w_041_128, w_041_129, w_041_130, w_041_131, w_041_134, w_041_135, w_041_136, w_041_138, w_041_140, w_041_141, w_041_142, w_041_143, w_041_144, w_041_145, w_041_146, w_041_148, w_041_149, w_041_153, w_041_154, w_041_156, w_041_157, w_041_158, w_041_159, w_041_160, w_041_161, w_041_163, w_041_166, w_041_167, w_041_168, w_041_169, w_041_171, w_041_172, w_041_173, w_041_176, w_041_179, w_041_180, w_041_181, w_041_183, w_041_184, w_041_185, w_041_186, w_041_187, w_041_188, w_041_189, w_041_190, w_041_191, w_041_192, w_041_194, w_041_195, w_041_196, w_041_197, w_041_198, w_041_199, w_041_200, w_041_201, w_041_202, w_041_203, w_041_204, w_041_205, w_041_207, w_041_208, w_041_209, w_041_211, w_041_212, w_041_213, w_041_214, w_041_216, w_041_217, w_041_218, w_041_219, w_041_220, w_041_221, w_041_222, w_041_223, w_041_224, w_041_225, w_041_227, w_041_228, w_041_230, w_041_231, w_041_232, w_041_233, w_041_234, w_041_235, w_041_236, w_041_238, w_041_239, w_041_240, w_041_241, w_041_242, w_041_243, w_041_244, w_041_245, w_041_246, w_041_247, w_041_248, w_041_250, w_041_251, w_041_252, w_041_253, w_041_254, w_041_257, w_041_258, w_041_259, w_041_260, w_041_262, w_041_263, w_041_264, w_041_265, w_041_266, w_041_267, w_041_268, w_041_269, w_041_270, w_041_271, w_041_273, w_041_274, w_041_275, w_041_276, w_041_277, w_041_278, w_041_279, w_041_280, w_041_281, w_041_282, w_041_283, w_041_284, w_041_285, w_041_287, w_041_289, w_041_291, w_041_292, w_041_294, w_041_295, w_041_297, w_041_299, w_041_300, w_041_301, w_041_302, w_041_304, w_041_305, w_041_306, w_041_307, w_041_308, w_041_309, w_041_310, w_041_311, w_041_312, w_041_313, w_041_315, w_041_316, w_041_317, w_041_318, w_041_319, w_041_320, w_041_321, w_041_322, w_041_324, w_041_325, w_041_326, w_041_328, w_041_329, w_041_331, w_041_332, w_041_333, w_041_335, w_041_336, w_041_337, w_041_338, w_041_339, w_041_340, w_041_342, w_041_343, w_041_344, w_041_345, w_041_346, w_041_347, w_041_348, w_041_349, w_041_350, w_041_351, w_041_352, w_041_353, w_041_354, w_041_355, w_041_356, w_041_358, w_041_359, w_041_360, w_041_361, w_041_362, w_041_363, w_041_364, w_041_366, w_041_367, w_041_368, w_041_369, w_041_371, w_041_373, w_041_374, w_041_375, w_041_377, w_041_380, w_041_381, w_041_382, w_041_383, w_041_384, w_041_385, w_041_386, w_041_387, w_041_388, w_041_389, w_041_390, w_041_392, w_041_393, w_041_394, w_041_396, w_041_397, w_041_399, w_041_400, w_041_401, w_041_402, w_041_404, w_041_405, w_041_406, w_041_407, w_041_408, w_041_409, w_041_410, w_041_411, w_041_412, w_041_413, w_041_414, w_041_416, w_041_417, w_041_418, w_041_419, w_041_420, w_041_421, w_041_422, w_041_423, w_041_424, w_041_426, w_041_427, w_041_428, w_041_430, w_041_431, w_041_432, w_041_433, w_041_434, w_041_435, w_041_438, w_041_439, w_041_440, w_041_441, w_041_442, w_041_444, w_041_445, w_041_447, w_041_448, w_041_449, w_041_450, w_041_451, w_041_453, w_041_455, w_041_456, w_041_458, w_041_459, w_041_460, w_041_461, w_041_463, w_041_464, w_041_465, w_041_466, w_041_467, w_041_469, w_041_470, w_041_472, w_041_473, w_041_474, w_041_475, w_041_476, w_041_477, w_041_478, w_041_479, w_041_481, w_041_482, w_041_483, w_041_484, w_041_485, w_041_487, w_041_488, w_041_490, w_041_491, w_041_492, w_041_493, w_041_494, w_041_495, w_041_496, w_041_497, w_041_500, w_041_501, w_041_502, w_041_503, w_041_504, w_041_505, w_041_507, w_041_508, w_041_509, w_041_510, w_041_513, w_041_514, w_041_516, w_041_517, w_041_518, w_041_519, w_041_520, w_041_521, w_041_522, w_041_523, w_041_524, w_041_525, w_041_526, w_041_527, w_041_528, w_041_529, w_041_530, w_041_531, w_041_532, w_041_533, w_041_535, w_041_536, w_041_537, w_041_538, w_041_539, w_041_540, w_041_542, w_041_543, w_041_544, w_041_547, w_041_548, w_041_549, w_041_550, w_041_551, w_041_552, w_041_553, w_041_554, w_041_555, w_041_556, w_041_557, w_041_559, w_041_560, w_041_561, w_041_562, w_041_563, w_041_564, w_041_565, w_041_569, w_041_570, w_041_571, w_041_572, w_041_574, w_041_575, w_041_576, w_041_577, w_041_578, w_041_580, w_041_583, w_041_585, w_041_586, w_041_587, w_041_588, w_041_589, w_041_590, w_041_591, w_041_592, w_041_594, w_041_595, w_041_596, w_041_597, w_041_598, w_041_599, w_041_601, w_041_602, w_041_603, w_041_604, w_041_605, w_041_606, w_041_607, w_041_608, w_041_609, w_041_610, w_041_611, w_041_612, w_041_614, w_041_615, w_041_616, w_041_617, w_041_618, w_041_619, w_041_620, w_041_621, w_041_622, w_041_623, w_041_624, w_041_625, w_041_626, w_041_630, w_041_631, w_041_632, w_041_633, w_041_634, w_041_635, w_041_636, w_041_637, w_041_639, w_041_640, w_041_641, w_041_643, w_041_644, w_041_645, w_041_646, w_041_647, w_041_648, w_041_649, w_041_650, w_041_651, w_041_652, w_041_654, w_041_655, w_041_656, w_041_657, w_041_658, w_041_659, w_041_660, w_041_661, w_041_662, w_041_663, w_041_664, w_041_665, w_041_670, w_041_671, w_041_672, w_041_673, w_041_675, w_041_676, w_041_677, w_041_678, w_041_679, w_041_680, w_041_683, w_041_684, w_041_685, w_041_686, w_041_687, w_041_688, w_041_689, w_041_690, w_041_692, w_041_693, w_041_694, w_041_697, w_041_698, w_041_699, w_041_700, w_041_701, w_041_702, w_041_703, w_041_704, w_041_705, w_041_706, w_041_707, w_041_708, w_041_709, w_041_710, w_041_711, w_041_712, w_041_713, w_041_715, w_041_716, w_041_720, w_041_721, w_041_722, w_041_723, w_041_724, w_041_725, w_041_726, w_041_727, w_041_728, w_041_729, w_041_730, w_041_731, w_041_732, w_041_733, w_041_734, w_041_735, w_041_736, w_041_737, w_041_738, w_041_740, w_041_741, w_041_742, w_041_743, w_041_744, w_041_745, w_041_746, w_041_747, w_041_748, w_041_749, w_041_750, w_041_751, w_041_752, w_041_753, w_041_754, w_041_755, w_041_756, w_041_757, w_041_758, w_041_759, w_041_760, w_041_761, w_041_762, w_041_763, w_041_766, w_041_767, w_041_769, w_041_771, w_041_772, w_041_773, w_041_774, w_041_775, w_041_776, w_041_777, w_041_778, w_041_779, w_041_780, w_041_781, w_041_782, w_041_784, w_041_785, w_041_786, w_041_787, w_041_789, w_041_791, w_041_792, w_041_793, w_041_794, w_041_795, w_041_796, w_041_797, w_041_799, w_041_800, w_041_801, w_041_802, w_041_803, w_041_804, w_041_805, w_041_807, w_041_808, w_041_809, w_041_810, w_041_811, w_041_813, w_041_815, w_041_816, w_041_817, w_041_818, w_041_819, w_041_820, w_041_821, w_041_822, w_041_823, w_041_824, w_041_825, w_041_826, w_041_827, w_041_829, w_041_830, w_041_831, w_041_833, w_041_835, w_041_836, w_041_837, w_041_840, w_041_841, w_041_842, w_041_844, w_041_845, w_041_847, w_041_850, w_041_851, w_041_852, w_041_853, w_041_855, w_041_857, w_041_858, w_041_859, w_041_861, w_041_862, w_041_863, w_041_866, w_041_867, w_041_869, w_041_870, w_041_872, w_041_873, w_041_874, w_041_875, w_041_876, w_041_877, w_041_878, w_041_879, w_041_880, w_041_882, w_041_884, w_041_885, w_041_886, w_041_887, w_041_888, w_041_892, w_041_893, w_041_894, w_041_895, w_041_896, w_041_897, w_041_898, w_041_900, w_041_901, w_041_902, w_041_903, w_041_904, w_041_905, w_041_906, w_041_907, w_041_908, w_041_909, w_041_910, w_041_911, w_041_913, w_041_914, w_041_915, w_041_917, w_041_918, w_041_919, w_041_920, w_041_921, w_041_922, w_041_923, w_041_924, w_041_925, w_041_926, w_041_927, w_041_928, w_041_929, w_041_930, w_041_931, w_041_933, w_041_934, w_041_935, w_041_936, w_041_938, w_041_940, w_041_941, w_041_942, w_041_943, w_041_944, w_041_945, w_041_946, w_041_947, w_041_948, w_041_949, w_041_950, w_041_952, w_041_954, w_041_955, w_041_956, w_041_957, w_041_958, w_041_959, w_041_960, w_041_962, w_041_963, w_041_964, w_041_965, w_041_966, w_041_967, w_041_968, w_041_970, w_041_971, w_041_973, w_041_974, w_041_975, w_041_976, w_041_977, w_041_978, w_041_979, w_041_980, w_041_981, w_041_982, w_041_984, w_041_986, w_041_987, w_041_989, w_041_990, w_041_991, w_041_993, w_041_994, w_041_995, w_041_997, w_041_998, w_041_999, w_041_1000, w_041_1001, w_041_1003, w_041_1004, w_041_1005, w_041_1006, w_041_1009, w_041_1010, w_041_1012, w_041_1013, w_041_1015, w_041_1017, w_041_1018, w_041_1019, w_041_1020, w_041_1023, w_041_1024, w_041_1025, w_041_1026, w_041_1029, w_041_1030, w_041_1031, w_041_1032, w_041_1033, w_041_1034, w_041_1036, w_041_1037, w_041_1040, w_041_1041, w_041_1043, w_041_1044, w_041_1046, w_041_1047, w_041_1048, w_041_1050, w_041_1051, w_041_1052, w_041_1053, w_041_1054, w_041_1056, w_041_1058, w_041_1059, w_041_1060, w_041_1061, w_041_1062, w_041_1063, w_041_1066, w_041_1067, w_041_1068, w_041_1069, w_041_1070, w_041_1071, w_041_1072, w_041_1073, w_041_1074, w_041_1075, w_041_1078, w_041_1079, w_041_1080, w_041_1081, w_041_1082, w_041_1084, w_041_1085, w_041_1086, w_041_1087, w_041_1088, w_041_1089, w_041_1090, w_041_1091, w_041_1092, w_041_1093, w_041_1094, w_041_1095, w_041_1096, w_041_1097, w_041_1098, w_041_1099, w_041_1100, w_041_1102, w_041_1103, w_041_1104, w_041_1106, w_041_1107, w_041_1108, w_041_1109, w_041_1110, w_041_1112, w_041_1113, w_041_1114, w_041_1115, w_041_1116, w_041_1117, w_041_1118, w_041_1121, w_041_1122, w_041_1123, w_041_1124, w_041_1125, w_041_1128, w_041_1129, w_041_1130, w_041_1131, w_041_1132, w_041_1133, w_041_1134, w_041_1136, w_041_1137, w_041_1139, w_041_1140, w_041_1141, w_041_1142, w_041_1143, w_041_1144, w_041_1145, w_041_1149, w_041_1150, w_041_1151, w_041_1152, w_041_1153, w_041_1154, w_041_1155, w_041_1158, w_041_1159, w_041_1161, w_041_1162, w_041_1163, w_041_1164, w_041_1166, w_041_1167, w_041_1168, w_041_1169, w_041_1170, w_041_1171, w_041_1172, w_041_1173, w_041_1174, w_041_1175, w_041_1176, w_041_1178, w_041_1179, w_041_1180, w_041_1181, w_041_1182, w_041_1184, w_041_1185, w_041_1186, w_041_1188, w_041_1189, w_041_1190, w_041_1192, w_041_1193, w_041_1194, w_041_1195, w_041_1196, w_041_1197, w_041_1198, w_041_1200, w_041_1201, w_041_1202, w_041_1203, w_041_1204, w_041_1205, w_041_1206, w_041_1207, w_041_1208, w_041_1209, w_041_1210, w_041_1211, w_041_1212, w_041_1214, w_041_1215, w_041_1216, w_041_1217, w_041_1219, w_041_1220, w_041_1221, w_041_1222, w_041_1223, w_041_1225, w_041_1227, w_041_1228, w_041_1229, w_041_1230, w_041_1231, w_041_1232, w_041_1233, w_041_1235, w_041_1236, w_041_1238, w_041_1239, w_041_1241, w_041_1242, w_041_1243, w_041_1244, w_041_1246, w_041_1247, w_041_1249, w_041_1250, w_041_1251, w_041_1252, w_041_1253, w_041_1254, w_041_1255, w_041_1257, w_041_1258, w_041_1260, w_041_1262, w_041_1263, w_041_1265, w_041_1266, w_041_1267, w_041_1268, w_041_1270, w_041_1271, w_041_1272, w_041_1273, w_041_1274, w_041_1276, w_041_1279, w_041_1281, w_041_1284, w_041_1285, w_041_1286, w_041_1287, w_041_1289, w_041_1290, w_041_1291, w_041_1292, w_041_1293, w_041_1294, w_041_1295, w_041_1297, w_041_1298, w_041_1299, w_041_1300, w_041_1303, w_041_1304, w_041_1305, w_041_1306, w_041_1307, w_041_1308, w_041_1309, w_041_1310, w_041_1311, w_041_1313, w_041_1314, w_041_1315, w_041_1316, w_041_1317, w_041_1318, w_041_1319, w_041_1320, w_041_1321, w_041_1322, w_041_1324, w_041_1325, w_041_1326, w_041_1328, w_041_1330, w_041_1331, w_041_1332, w_041_1333, w_041_1336, w_041_1337, w_041_1338, w_041_1339, w_041_1341, w_041_1342, w_041_1346, w_041_1347, w_041_1348, w_041_1349, w_041_1350, w_041_1351, w_041_1352, w_041_1354, w_041_1355, w_041_1356, w_041_1357, w_041_1358, w_041_1359, w_041_1361, w_041_1362, w_041_1363, w_041_1364, w_041_1365, w_041_1366, w_041_1367, w_041_1368, w_041_1369, w_041_1370, w_041_1372, w_041_1374, w_041_1375, w_041_1376, w_041_1377, w_041_1378, w_041_1379, w_041_1381, w_041_1382, w_041_1383, w_041_1384, w_041_1386, w_041_1387, w_041_1388, w_041_1389, w_041_1391, w_041_1392, w_041_1393, w_041_1395, w_041_1396, w_041_1398, w_041_1399, w_041_1400, w_041_1402, w_041_1403, w_041_1404, w_041_1405, w_041_1406, w_041_1407, w_041_1408, w_041_1409, w_041_1410, w_041_1411, w_041_1412, w_041_1413, w_041_1414, w_041_1415, w_041_1416, w_041_1417, w_041_1419, w_041_1420, w_041_1421, w_041_1422, w_041_1423, w_041_1424, w_041_1425, w_041_1426, w_041_1427, w_041_1428, w_041_1429, w_041_1430, w_041_1431, w_041_1432, w_041_1435, w_041_1439, w_041_1440, w_041_1442, w_041_1443, w_041_1444, w_041_1445, w_041_1446, w_041_1448, w_041_1450, w_041_1452, w_041_1453, w_041_1454, w_041_1455, w_041_1457, w_041_1458, w_041_1459, w_041_1461, w_041_1462, w_041_1463, w_041_1466, w_041_1467, w_041_1468, w_041_1470, w_041_1471, w_041_1474, w_041_1475, w_041_1476, w_041_1478, w_041_1479, w_041_1480, w_041_1482, w_041_1483, w_041_1484, w_041_1485, w_041_1486, w_041_1487, w_041_1488, w_041_1489, w_041_1490, w_041_1491, w_041_1492, w_041_1494, w_041_1495, w_041_1497, w_041_1498, w_041_1499, w_041_1501, w_041_1502, w_041_1503, w_041_1504, w_041_1506, w_041_1508, w_041_1509, w_041_1510, w_041_1512, w_041_1513, w_041_1514, w_041_1515, w_041_1516, w_041_1519, w_041_1520, w_041_1521, w_041_1523, w_041_1525, w_041_1527, w_041_1528, w_041_1529, w_041_1530, w_041_1531, w_041_1533, w_041_1534, w_041_1535, w_041_1536, w_041_1537, w_041_1538, w_041_1539, w_041_1540, w_041_1541, w_041_1542, w_041_1543, w_041_1544, w_041_1545, w_041_1546, w_041_1547, w_041_1548, w_041_1549, w_041_1550, w_041_1551, w_041_1552, w_041_1553, w_041_1554, w_041_1555, w_041_1556, w_041_1557, w_041_1558, w_041_1559, w_041_1560, w_041_1562, w_041_1563, w_041_1564, w_041_1566, w_041_1568, w_041_1569, w_041_1570, w_041_1571, w_041_1572, w_041_1573, w_041_1574, w_041_1575, w_041_1576, w_041_1577, w_041_1578, w_041_1579, w_041_1580, w_041_1581, w_041_1582, w_041_1584, w_041_1586, w_041_1588, w_041_1589, w_041_1590, w_041_1591, w_041_1592, w_041_1593, w_041_1594, w_041_1595, w_041_1596, w_041_1598, w_041_1599, w_041_1600, w_041_1601, w_041_1602, w_041_1603, w_041_1604, w_041_1606, w_041_1607, w_041_1608, w_041_1611, w_041_1612, w_041_1613, w_041_1615, w_041_1617, w_041_1618, w_041_1619, w_041_1620, w_041_1623, w_041_1624, w_041_1625, w_041_1627, w_041_1628, w_041_1630, w_041_1631, w_041_1632, w_041_1634, w_041_1635, w_041_1636, w_041_1637, w_041_1638, w_041_1639, w_041_1640, w_041_1641, w_041_1642, w_041_1643, w_041_1644, w_041_1645, w_041_1646, w_041_1647, w_041_1648, w_041_1649, w_041_1650, w_041_1652, w_041_1653, w_041_1654, w_041_1655, w_041_1656, w_041_1657, w_041_1659, w_041_1661, w_041_1662, w_041_1663, w_041_1664, w_041_1665, w_041_1666, w_041_1667, w_041_1668, w_041_1669, w_041_1670, w_041_1671, w_041_1672, w_041_1673, w_041_1674, w_041_1675, w_041_1677, w_041_1678, w_041_1679, w_041_1680, w_041_1681, w_041_1682, w_041_1683, w_041_1684, w_041_1685, w_041_1687, w_041_1689, w_041_1690, w_041_1692, w_041_1694, w_041_1695, w_041_1696, w_041_1697, w_041_1698, w_041_1699, w_041_1700, w_041_1701, w_041_1703, w_041_1705, w_041_1707, w_041_1708, w_041_1709, w_041_1711, w_041_1712, w_041_1714, w_041_1715, w_041_1717, w_041_1718, w_041_1719, w_041_1720, w_041_1721, w_041_1722, w_041_1723, w_041_1724, w_041_1725, w_041_1726, w_041_1727, w_041_1728, w_041_1729, w_041_1730, w_041_1733, w_041_1734, w_041_1735, w_041_1739, w_041_1740, w_041_1741, w_041_1742, w_041_1743, w_041_1745, w_041_1746, w_041_1747, w_041_1748, w_041_1749, w_041_1751, w_041_1752, w_041_1753, w_041_1754, w_041_1755, w_041_1757, w_041_1758, w_041_1760, w_041_1761, w_041_1762, w_041_1763, w_041_1764, w_041_1765, w_041_1766, w_041_1767, w_041_1768, w_041_1769, w_041_1770, w_041_1771, w_041_1772, w_041_1774, w_041_1775, w_041_1776, w_041_1777, w_041_1778, w_041_1779, w_041_1780, w_041_1781, w_041_1782, w_041_1783, w_041_1784, w_041_1785, w_041_1787, w_041_1788, w_041_1789, w_041_1791, w_041_1793, w_041_1797, w_041_1798, w_041_1799, w_041_1800, w_041_1801, w_041_1802, w_041_1803, w_041_1804, w_041_1805, w_041_1806, w_041_1807, w_041_1808, w_041_1810, w_041_1812, w_041_1813, w_041_1814, w_041_1817, w_041_1818, w_041_1820, w_041_1821, w_041_1822, w_041_1823, w_041_1828, w_041_1829, w_041_1830, w_041_1832, w_041_1833, w_041_1834, w_041_1835, w_041_1836, w_041_1837, w_041_1838, w_041_1839, w_041_1840, w_041_1841, w_041_1842, w_041_1844, w_041_1847, w_041_1848, w_041_1849, w_041_1851, w_041_1852, w_041_1853, w_041_1854, w_041_1855, w_041_1857, w_041_1858, w_041_1860, w_041_1861, w_041_1862, w_041_1863, w_041_1864, w_041_1866, w_041_1867, w_041_1868, w_041_1869, w_041_1870, w_041_1872, w_041_1873, w_041_1874, w_041_1875, w_041_1876, w_041_1877, w_041_1878, w_041_1879, w_041_1880, w_041_1881, w_041_1882, w_041_1883, w_041_1885, w_041_1888, w_041_1889, w_041_1890, w_041_1891, w_041_1893, w_041_1894, w_041_1898, w_041_1899, w_041_1901, w_041_1903, w_041_1904, w_041_1905, w_041_1907, w_041_1909, w_041_1913, w_041_1915, w_041_1916, w_041_1917, w_041_1919, w_041_1920, w_041_1921, w_041_1923, w_041_1925, w_041_1927, w_041_1928, w_041_1930, w_041_1933, w_041_1935, w_041_1936, w_041_1938, w_041_1940, w_041_1941, w_041_1944, w_041_1945, w_041_1946, w_041_1947, w_041_1949, w_041_1951, w_041_1952, w_041_1953, w_041_1955, w_041_1957, w_041_1959, w_041_1963, w_041_1966, w_041_1967, w_041_1968, w_041_1969, w_041_1970, w_041_1972, w_041_1973, w_041_1975, w_041_1976, w_041_1978, w_041_1979, w_041_1980, w_041_1984, w_041_1987, w_041_1992, w_041_1993, w_041_1994, w_041_1995, w_041_1999, w_041_2002, w_041_2003, w_041_2004, w_041_2006, w_041_2011, w_041_2014, w_041_2015, w_041_2016, w_041_2019, w_041_2022, w_041_2025, w_041_2030, w_041_2033, w_041_2034, w_041_2035, w_041_2040, w_041_2041, w_041_2044, w_041_2046, w_041_2047, w_041_2048, w_041_2052, w_041_2053, w_041_2055, w_041_2056, w_041_2058, w_041_2059, w_041_2060, w_041_2064, w_041_2066, w_041_2067, w_041_2068, w_041_2070, w_041_2072, w_041_2074, w_041_2075, w_041_2076, w_041_2079, w_041_2080, w_041_2081, w_041_2082, w_041_2083, w_041_2084, w_041_2086, w_041_2088, w_041_2090, w_041_2093, w_041_2094, w_041_2095, w_041_2096, w_041_2100, w_041_2101, w_041_2102, w_041_2104, w_041_2106, w_041_2109, w_041_2110, w_041_2111, w_041_2112, w_041_2113, w_041_2114, w_041_2115, w_041_2116, w_041_2120, w_041_2121, w_041_2122, w_041_2126, w_041_2127, w_041_2129, w_041_2130, w_041_2134, w_041_2135, w_041_2137, w_041_2139, w_041_2140, w_041_2142, w_041_2144, w_041_2147, w_041_2148, w_041_2149, w_041_2150, w_041_2151, w_041_2153, w_041_2154, w_041_2160, w_041_2161, w_041_2162, w_041_2164, w_041_2165, w_041_2166, w_041_2170, w_041_2172, w_041_2173, w_041_2174, w_041_2177, w_041_2182, w_041_2183, w_041_2185, w_041_2187, w_041_2188, w_041_2191, w_041_2192, w_041_2193, w_041_2195, w_041_2197, w_041_2200, w_041_2202, w_041_2204, w_041_2207, w_041_2208, w_041_2209, w_041_2211, w_041_2212, w_041_2214, w_041_2217, w_041_2218, w_041_2219, w_041_2222, w_041_2223, w_041_2224, w_041_2225, w_041_2229, w_041_2230, w_041_2231, w_041_2233, w_041_2234, w_041_2238, w_041_2239, w_041_2241, w_041_2242, w_041_2248, w_041_2249, w_041_2252, w_041_2256, w_041_2260, w_041_2265, w_041_2266, w_041_2268, w_041_2269, w_041_2271, w_041_2272, w_041_2274, w_041_2275, w_041_2278, w_041_2281, w_041_2282, w_041_2283, w_041_2284, w_041_2290, w_041_2292, w_041_2293, w_041_2294, w_041_2295, w_041_2298, w_041_2301, w_041_2303, w_041_2305, w_041_2306, w_041_2307, w_041_2308, w_041_2314, w_041_2315, w_041_2316, w_041_2318, w_041_2319, w_041_2321, w_041_2324, w_041_2325, w_041_2327, w_041_2328, w_041_2329, w_041_2332, w_041_2334, w_041_2335, w_041_2337, w_041_2340, w_041_2342, w_041_2344, w_041_2346, w_041_2347, w_041_2349, w_041_2350, w_041_2352, w_041_2354, w_041_2355, w_041_2356, w_041_2359, w_041_2362, w_041_2365, w_041_2370, w_041_2375, w_041_2376, w_041_2377, w_041_2381, w_041_2385, w_041_2386, w_041_2389, w_041_2390, w_041_2391, w_041_2392, w_041_2393, w_041_2395, w_041_2398, w_041_2399, w_041_2401, w_041_2402, w_041_2404, w_041_2405, w_041_2409, w_041_2410, w_041_2411, w_041_2412, w_041_2417, w_041_2418, w_041_2421, w_041_2423, w_041_2424, w_041_2425, w_041_2427, w_041_2428, w_041_2430, w_041_2432, w_041_2434, w_041_2435, w_041_2437, w_041_2439, w_041_2441, w_041_2442, w_041_2444, w_041_2445, w_041_2447, w_041_2450, w_041_2451, w_041_2453, w_041_2454, w_041_2456, w_041_2457, w_041_2459, w_041_2460, w_041_2463, w_041_2464, w_041_2465, w_041_2466, w_041_2467, w_041_2468, w_041_2469, w_041_2470, w_041_2472, w_041_2473, w_041_2474, w_041_2475, w_041_2479, w_041_2480, w_041_2481, w_041_2483, w_041_2484, w_041_2488, w_041_2489, w_041_2490, w_041_2493, w_041_2495, w_041_2496, w_041_2498, w_041_2501, w_041_2504, w_041_2506, w_041_2507, w_041_2509, w_041_2510, w_041_2511, w_041_2512, w_041_2513, w_041_2514, w_041_2517, w_041_2522, w_041_2523, w_041_2526, w_041_2528, w_041_2530, w_041_2532, w_041_2536, w_041_2537, w_041_2539, w_041_2542, w_041_2544, w_041_2547, w_041_2549, w_041_2550, w_041_2552, w_041_2553, w_041_2554, w_041_2556, w_041_2557, w_041_2558, w_041_2560, w_041_2562, w_041_2570, w_041_2571, w_041_2572, w_041_2574, w_041_2575, w_041_2576, w_041_2577, w_041_2578, w_041_2580, w_041_2581, w_041_2583, w_041_2584, w_041_2586, w_041_2587, w_041_2588, w_041_2591, w_041_2595, w_041_2596, w_041_2597, w_041_2599, w_041_2600, w_041_2603, w_041_2604, w_041_2605, w_041_2606, w_041_2608, w_041_2609, w_041_2610, w_041_2612, w_041_2614, w_041_2618, w_041_2620, w_041_2622, w_041_2625, w_041_2626, w_041_2627, w_041_2628, w_041_2629, w_041_2631, w_041_2632, w_041_2634, w_041_2635, w_041_2636, w_041_2637, w_041_2638, w_041_2639, w_041_2640, w_041_2641, w_041_2643, w_041_2644, w_041_2646, w_041_2648, w_041_2651, w_041_2652, w_041_2655, w_041_2658, w_041_2659, w_041_2660, w_041_2662, w_041_2663, w_041_2666, w_041_2667, w_041_2668, w_041_2669, w_041_2670, w_041_2671, w_041_2672, w_041_2673, w_041_2677, w_041_2680, w_041_2681, w_041_2683, w_041_2684, w_041_2685, w_041_2686, w_041_2687, w_041_2688, w_041_2690, w_041_2693, w_041_2694, w_041_2695, w_041_2698, w_041_2699, w_041_2700, w_041_2701, w_041_2702, w_041_2703, w_041_2704, w_041_2705, w_041_2709, w_041_2710, w_041_2712, w_041_2715, w_041_2717, w_041_2718, w_041_2719, w_041_2720, w_041_2721, w_041_2722, w_041_2723, w_041_2724, w_041_2726, w_041_2728, w_041_2729, w_041_2730, w_041_2732, w_041_2736, w_041_2737, w_041_2739, w_041_2740, w_041_2741, w_041_2745, w_041_2746, w_041_2747, w_041_2749, w_041_2750, w_041_2751, w_041_2752, w_041_2753, w_041_2754, w_041_2756, w_041_2757, w_041_2759, w_041_2761, w_041_2764, w_041_2765, w_041_2767, w_041_2768, w_041_2769, w_041_2770, w_041_2771, w_041_2773, w_041_2774, w_041_2776, w_041_2777, w_041_2779, w_041_2780, w_041_2781, w_041_2784, w_041_2788, w_041_2789, w_041_2792, w_041_2797, w_041_2798, w_041_2801, w_041_2804, w_041_2806, w_041_2808, w_041_2810, w_041_2811, w_041_2813, w_041_2815, w_041_2816, w_041_2817, w_041_2818, w_041_2819, w_041_2821, w_041_2825, w_041_2826, w_041_2827, w_041_2828, w_041_2829, w_041_2830, w_041_2833, w_041_2835, w_041_2836, w_041_2837, w_041_2838, w_041_2839, w_041_2840, w_041_2841, w_041_2844, w_041_2847, w_041_2849, w_041_2850, w_041_2851, w_041_2855, w_041_2859, w_041_2860, w_041_2861, w_041_2862, w_041_2864, w_041_2865, w_041_2866, w_041_2867, w_041_2868, w_041_2870, w_041_2871, w_041_2872, w_041_2873, w_041_2876, w_041_2877, w_041_2878, w_041_2879, w_041_2880, w_041_2881, w_041_2883, w_041_2887, w_041_2889, w_041_2891, w_041_2892, w_041_2894, w_041_2895, w_041_2896, w_041_2899, w_041_2900, w_041_2902, w_041_2903, w_041_2910, w_041_2911, w_041_2912, w_041_2913, w_041_2914, w_041_2915, w_041_2917, w_041_2918, w_041_2923, w_041_2924, w_041_2925, w_041_2928, w_041_2933, w_041_2934, w_041_2939, w_041_2941, w_041_2942, w_041_2943, w_041_2946, w_041_2947, w_041_2949, w_041_2950, w_041_2951, w_041_2952, w_041_2953, w_041_2955, w_041_2957, w_041_2958, w_041_2960, w_041_2962, w_041_2963, w_041_2964, w_041_2966, w_041_2967, w_041_2968, w_041_2969, w_041_2970, w_041_2971, w_041_2973, w_041_2974, w_041_2975, w_041_2976, w_041_2977, w_041_2978, w_041_2979, w_041_2980, w_041_2982, w_041_2983, w_041_2984, w_041_2988, w_041_2990, w_041_2992, w_041_2993, w_041_2994, w_041_2995, w_041_3005, w_041_3006, w_041_3007, w_041_3008, w_041_3009, w_041_3010, w_041_3014, w_041_3015, w_041_3017, w_041_3021, w_041_3022, w_041_3024, w_041_3025, w_041_3026, w_041_3028, w_041_3029, w_041_3033, w_041_3034, w_041_3035, w_041_3037, w_041_3038, w_041_3040, w_041_3043, w_041_3044, w_041_3045, w_041_3046, w_041_3047, w_041_3049, w_041_3052, w_041_3053, w_041_3055, w_041_3056, w_041_3057, w_041_3059, w_041_3062, w_041_3064, w_041_3065, w_041_3066, w_041_3067, w_041_3068, w_041_3074, w_041_3075, w_041_3076, w_041_3078, w_041_3079, w_041_3080, w_041_3081, w_041_3082, w_041_3083, w_041_3085, w_041_3087, w_041_3088, w_041_3090, w_041_3092, w_041_3095, w_041_3096, w_041_3099, w_041_3102, w_041_3110, w_041_3111, w_041_3112, w_041_3113, w_041_3114, w_041_3115, w_041_3116, w_041_3117, w_041_3118, w_041_3119, w_041_3120, w_041_3121, w_041_3125, w_041_3126, w_041_3127, w_041_3128, w_041_3129, w_041_3131, w_041_3133, w_041_3134, w_041_3135, w_041_3136, w_041_3137, w_041_3138, w_041_3139, w_041_3141;
  wire w_042_000, w_042_001, w_042_002, w_042_003, w_042_005, w_042_006, w_042_007, w_042_008, w_042_009, w_042_011, w_042_012, w_042_013, w_042_014, w_042_019, w_042_020, w_042_021, w_042_022, w_042_023, w_042_024, w_042_026, w_042_027, w_042_028, w_042_029, w_042_030, w_042_031, w_042_033, w_042_034, w_042_035, w_042_036, w_042_037, w_042_038, w_042_039, w_042_040, w_042_041, w_042_042, w_042_044, w_042_046, w_042_049, w_042_051, w_042_052, w_042_053, w_042_054, w_042_055, w_042_058, w_042_059, w_042_060, w_042_062, w_042_063, w_042_064, w_042_065, w_042_066, w_042_067, w_042_068, w_042_069, w_042_070, w_042_071, w_042_072, w_042_073, w_042_074, w_042_076, w_042_077, w_042_078, w_042_080, w_042_081, w_042_082, w_042_083, w_042_084, w_042_085, w_042_087, w_042_088, w_042_089, w_042_090, w_042_091, w_042_092, w_042_093, w_042_095, w_042_096, w_042_097, w_042_098, w_042_099, w_042_101, w_042_102, w_042_103, w_042_104, w_042_105, w_042_106, w_042_107, w_042_108, w_042_109, w_042_110, w_042_112, w_042_113, w_042_116, w_042_119, w_042_120, w_042_121, w_042_123, w_042_124, w_042_125, w_042_126, w_042_128, w_042_129, w_042_131, w_042_132, w_042_133, w_042_134, w_042_135, w_042_136, w_042_137, w_042_138, w_042_139, w_042_140, w_042_141, w_042_143, w_042_144, w_042_145, w_042_146, w_042_147, w_042_148, w_042_149, w_042_150, w_042_152, w_042_153, w_042_155, w_042_156, w_042_157, w_042_159, w_042_160, w_042_162, w_042_163, w_042_165, w_042_167, w_042_168, w_042_170, w_042_171, w_042_175, w_042_176, w_042_177, w_042_178, w_042_179, w_042_180, w_042_181, w_042_182, w_042_183, w_042_186, w_042_188, w_042_190, w_042_193, w_042_194, w_042_195, w_042_196, w_042_197, w_042_198, w_042_199, w_042_200, w_042_201, w_042_202, w_042_203, w_042_204, w_042_205, w_042_206, w_042_207, w_042_208, w_042_210, w_042_211, w_042_212, w_042_213, w_042_214, w_042_216, w_042_217, w_042_218, w_042_219, w_042_220, w_042_221, w_042_223, w_042_226, w_042_227, w_042_228, w_042_229, w_042_230, w_042_231, w_042_233, w_042_234, w_042_235, w_042_236, w_042_237, w_042_240, w_042_242, w_042_243, w_042_244, w_042_245, w_042_247, w_042_249, w_042_252, w_042_253, w_042_254, w_042_255, w_042_257, w_042_258, w_042_259, w_042_260, w_042_261, w_042_262, w_042_263, w_042_264, w_042_265, w_042_267, w_042_268, w_042_269, w_042_270, w_042_271, w_042_272, w_042_274, w_042_275, w_042_277, w_042_279, w_042_280, w_042_282, w_042_283, w_042_286, w_042_287, w_042_288, w_042_290, w_042_291, w_042_292, w_042_294, w_042_295, w_042_296, w_042_298, w_042_301, w_042_303, w_042_304, w_042_305, w_042_307, w_042_308, w_042_309, w_042_310, w_042_311, w_042_312, w_042_313, w_042_314, w_042_315, w_042_317, w_042_318, w_042_319, w_042_320, w_042_321, w_042_322, w_042_323, w_042_324, w_042_326, w_042_330, w_042_332, w_042_334, w_042_335, w_042_336, w_042_337, w_042_339, w_042_343, w_042_344, w_042_346, w_042_347, w_042_349, w_042_352, w_042_355, w_042_356, w_042_358, w_042_360, w_042_362, w_042_364, w_042_365, w_042_374, w_042_376, w_042_378, w_042_380, w_042_383, w_042_384, w_042_386, w_042_387, w_042_389, w_042_390, w_042_392, w_042_394, w_042_395, w_042_396, w_042_398, w_042_399, w_042_402, w_042_403, w_042_405, w_042_409, w_042_410, w_042_413, w_042_414, w_042_415, w_042_418, w_042_421, w_042_422, w_042_423, w_042_424, w_042_425, w_042_426, w_042_427, w_042_428, w_042_431, w_042_435, w_042_436, w_042_438, w_042_441, w_042_442, w_042_446, w_042_447, w_042_449, w_042_450, w_042_451, w_042_452, w_042_454, w_042_455, w_042_456, w_042_460, w_042_461, w_042_463, w_042_464, w_042_465, w_042_467, w_042_470, w_042_476, w_042_477, w_042_479, w_042_481, w_042_483, w_042_484, w_042_485, w_042_486, w_042_487, w_042_490, w_042_491, w_042_497, w_042_500, w_042_502, w_042_503, w_042_504, w_042_505, w_042_507, w_042_508, w_042_509, w_042_511, w_042_512, w_042_514, w_042_515, w_042_518, w_042_520, w_042_521, w_042_524, w_042_528, w_042_530, w_042_531, w_042_538, w_042_539, w_042_540, w_042_541, w_042_542, w_042_543, w_042_544, w_042_545, w_042_546, w_042_547, w_042_549, w_042_553, w_042_554, w_042_555, w_042_556, w_042_557, w_042_558, w_042_560, w_042_564, w_042_565, w_042_566, w_042_567, w_042_570, w_042_571, w_042_575, w_042_578, w_042_580, w_042_581, w_042_583, w_042_585, w_042_586, w_042_588, w_042_591, w_042_592, w_042_593, w_042_594, w_042_595, w_042_597, w_042_598, w_042_599, w_042_601, w_042_602, w_042_606, w_042_607, w_042_608, w_042_609, w_042_612, w_042_613, w_042_614, w_042_616, w_042_617, w_042_620, w_042_621, w_042_623, w_042_624, w_042_628, w_042_629, w_042_631, w_042_632, w_042_633, w_042_634, w_042_637, w_042_640, w_042_642, w_042_643, w_042_645, w_042_646, w_042_647, w_042_651, w_042_652, w_042_653, w_042_654, w_042_657, w_042_658, w_042_659, w_042_660, w_042_661, w_042_662, w_042_664, w_042_665, w_042_667, w_042_671, w_042_675, w_042_677, w_042_682, w_042_683, w_042_689, w_042_692, w_042_695, w_042_699, w_042_702, w_042_704, w_042_705, w_042_707, w_042_708, w_042_711, w_042_712, w_042_714, w_042_716, w_042_717, w_042_719, w_042_720, w_042_722, w_042_723, w_042_724, w_042_725, w_042_729, w_042_730, w_042_731, w_042_732, w_042_733, w_042_734, w_042_735, w_042_737, w_042_738, w_042_740, w_042_741, w_042_742, w_042_743, w_042_745, w_042_746, w_042_749, w_042_750, w_042_752, w_042_755, w_042_759, w_042_761, w_042_762, w_042_764, w_042_766, w_042_768, w_042_769, w_042_770, w_042_771, w_042_772, w_042_773, w_042_775, w_042_776, w_042_778, w_042_779, w_042_780, w_042_781, w_042_782, w_042_784, w_042_785, w_042_786, w_042_788, w_042_791, w_042_793, w_042_795, w_042_800, w_042_801, w_042_802, w_042_804, w_042_810, w_042_811, w_042_813, w_042_816, w_042_819, w_042_821, w_042_822, w_042_824, w_042_828, w_042_829, w_042_832, w_042_833, w_042_834, w_042_835, w_042_838, w_042_839, w_042_840, w_042_841, w_042_842, w_042_844, w_042_845, w_042_846, w_042_847, w_042_848, w_042_850, w_042_854, w_042_856, w_042_857, w_042_859, w_042_860, w_042_861, w_042_864, w_042_866, w_042_869, w_042_872, w_042_873, w_042_874, w_042_876, w_042_878, w_042_879, w_042_881, w_042_882, w_042_883, w_042_884, w_042_885, w_042_886, w_042_888, w_042_890, w_042_896, w_042_897, w_042_898, w_042_899, w_042_900, w_042_902, w_042_903, w_042_906, w_042_907, w_042_910, w_042_913, w_042_914, w_042_916, w_042_917, w_042_918, w_042_919, w_042_924, w_042_929, w_042_930, w_042_931, w_042_934, w_042_936, w_042_938, w_042_939, w_042_940, w_042_941, w_042_947, w_042_950, w_042_951, w_042_952, w_042_953, w_042_954, w_042_958, w_042_959, w_042_961, w_042_963, w_042_965, w_042_966, w_042_968, w_042_969, w_042_970, w_042_971, w_042_972, w_042_973, w_042_979, w_042_980, w_042_983, w_042_984, w_042_990, w_042_992, w_042_993, w_042_994, w_042_995, w_042_996, w_042_998, w_042_999, w_042_1004, w_042_1005, w_042_1006, w_042_1007, w_042_1009, w_042_1010, w_042_1013, w_042_1017, w_042_1019, w_042_1022, w_042_1023, w_042_1025, w_042_1026, w_042_1029, w_042_1030, w_042_1034, w_042_1036, w_042_1041, w_042_1042, w_042_1043, w_042_1044, w_042_1045, w_042_1046, w_042_1049, w_042_1053, w_042_1056, w_042_1057, w_042_1058, w_042_1059, w_042_1063, w_042_1064, w_042_1066, w_042_1067, w_042_1068, w_042_1070, w_042_1071, w_042_1074, w_042_1076, w_042_1077, w_042_1078, w_042_1079, w_042_1081, w_042_1085, w_042_1087, w_042_1088, w_042_1089, w_042_1091, w_042_1092, w_042_1095, w_042_1096, w_042_1097, w_042_1101, w_042_1102, w_042_1103, w_042_1105, w_042_1106, w_042_1107, w_042_1108, w_042_1110, w_042_1114, w_042_1115, w_042_1117, w_042_1121, w_042_1122, w_042_1124, w_042_1126, w_042_1127, w_042_1128, w_042_1129, w_042_1131, w_042_1133, w_042_1134, w_042_1135, w_042_1137, w_042_1139, w_042_1140, w_042_1142, w_042_1143, w_042_1145, w_042_1146, w_042_1148, w_042_1152, w_042_1154, w_042_1155, w_042_1156, w_042_1158, w_042_1160, w_042_1162, w_042_1165, w_042_1166, w_042_1168, w_042_1169, w_042_1170, w_042_1171, w_042_1172, w_042_1173, w_042_1174, w_042_1176, w_042_1177, w_042_1179, w_042_1181, w_042_1182, w_042_1183, w_042_1184, w_042_1186, w_042_1187, w_042_1189, w_042_1191, w_042_1195, w_042_1196, w_042_1197, w_042_1198, w_042_1199, w_042_1200, w_042_1207, w_042_1208, w_042_1209, w_042_1212, w_042_1213, w_042_1214, w_042_1215, w_042_1216, w_042_1218, w_042_1219, w_042_1220, w_042_1222, w_042_1224, w_042_1225, w_042_1227, w_042_1229, w_042_1231, w_042_1232, w_042_1233, w_042_1234, w_042_1236, w_042_1238, w_042_1239, w_042_1243, w_042_1244, w_042_1246, w_042_1252, w_042_1256, w_042_1259, w_042_1261, w_042_1263, w_042_1264, w_042_1265, w_042_1266, w_042_1267, w_042_1270, w_042_1273, w_042_1276, w_042_1277, w_042_1278, w_042_1279, w_042_1282, w_042_1284, w_042_1285, w_042_1286, w_042_1287, w_042_1290, w_042_1292, w_042_1294, w_042_1297, w_042_1298, w_042_1301, w_042_1302, w_042_1303, w_042_1304, w_042_1305, w_042_1306, w_042_1309, w_042_1311, w_042_1312, w_042_1313, w_042_1314, w_042_1316, w_042_1317, w_042_1320, w_042_1322, w_042_1326, w_042_1327, w_042_1331, w_042_1332, w_042_1333, w_042_1334, w_042_1336, w_042_1339, w_042_1341, w_042_1345, w_042_1346, w_042_1349, w_042_1351, w_042_1352, w_042_1353, w_042_1354, w_042_1356, w_042_1357, w_042_1358, w_042_1359, w_042_1360, w_042_1362, w_042_1368, w_042_1369, w_042_1371, w_042_1372, w_042_1373, w_042_1374, w_042_1376, w_042_1377, w_042_1380, w_042_1383, w_042_1384, w_042_1385, w_042_1387, w_042_1388, w_042_1389, w_042_1392, w_042_1393, w_042_1394, w_042_1395, w_042_1396, w_042_1397, w_042_1399, w_042_1401, w_042_1402, w_042_1403, w_042_1404, w_042_1405, w_042_1406, w_042_1410, w_042_1412, w_042_1415, w_042_1416, w_042_1417, w_042_1421, w_042_1422, w_042_1423, w_042_1426, w_042_1428, w_042_1432, w_042_1434, w_042_1435, w_042_1437, w_042_1439, w_042_1441, w_042_1442, w_042_1443, w_042_1444, w_042_1445, w_042_1446, w_042_1447, w_042_1448, w_042_1449, w_042_1451, w_042_1452, w_042_1453, w_042_1455, w_042_1456, w_042_1457, w_042_1458, w_042_1459, w_042_1460, w_042_1461, w_042_1464, w_042_1465, w_042_1466, w_042_1469, w_042_1470, w_042_1474, w_042_1478, w_042_1483, w_042_1485, w_042_1487, w_042_1489, w_042_1490, w_042_1491, w_042_1492, w_042_1494, w_042_1496, w_042_1498, w_042_1507, w_042_1508, w_042_1510, w_042_1512, w_042_1515, w_042_1518, w_042_1521, w_042_1522, w_042_1523, w_042_1524, w_042_1525, w_042_1527, w_042_1528, w_042_1529, w_042_1530, w_042_1532, w_042_1533, w_042_1535, w_042_1537, w_042_1538, w_042_1541, w_042_1543, w_042_1544, w_042_1547, w_042_1549, w_042_1550, w_042_1551, w_042_1552, w_042_1553, w_042_1555, w_042_1556, w_042_1557, w_042_1558, w_042_1561, w_042_1563, w_042_1564, w_042_1565, w_042_1567, w_042_1569, w_042_1570, w_042_1571, w_042_1574, w_042_1576, w_042_1577, w_042_1580, w_042_1582, w_042_1583, w_042_1584, w_042_1587, w_042_1589, w_042_1590, w_042_1592, w_042_1593, w_042_1595, w_042_1598, w_042_1601, w_042_1602, w_042_1603, w_042_1604, w_042_1605, w_042_1613, w_042_1615, w_042_1617, w_042_1622, w_042_1625, w_042_1627, w_042_1628, w_042_1630, w_042_1631, w_042_1632, w_042_1636, w_042_1638, w_042_1639, w_042_1640, w_042_1645, w_042_1646, w_042_1647, w_042_1648, w_042_1649, w_042_1650, w_042_1652, w_042_1653, w_042_1656, w_042_1657, w_042_1660, w_042_1665, w_042_1667, w_042_1668, w_042_1670, w_042_1672, w_042_1673, w_042_1674, w_042_1677, w_042_1679, w_042_1682, w_042_1683, w_042_1684, w_042_1687, w_042_1688, w_042_1689, w_042_1691, w_042_1695, w_042_1696, w_042_1698, w_042_1699, w_042_1700, w_042_1702, w_042_1703, w_042_1705, w_042_1706, w_042_1708, w_042_1711, w_042_1713, w_042_1715, w_042_1716, w_042_1719, w_042_1722, w_042_1723, w_042_1726, w_042_1729, w_042_1730, w_042_1731, w_042_1732, w_042_1733, w_042_1734, w_042_1737, w_042_1740, w_042_1741, w_042_1743, w_042_1744, w_042_1745, w_042_1747, w_042_1748, w_042_1749, w_042_1750, w_042_1752, w_042_1754, w_042_1758, w_042_1761, w_042_1763, w_042_1765, w_042_1766, w_042_1767, w_042_1768, w_042_1769, w_042_1772, w_042_1776, w_042_1777, w_042_1780, w_042_1781, w_042_1782, w_042_1785, w_042_1789, w_042_1793, w_042_1795, w_042_1796, w_042_1798, w_042_1800, w_042_1801, w_042_1802, w_042_1803, w_042_1804, w_042_1811, w_042_1814, w_042_1816, w_042_1818, w_042_1819, w_042_1820, w_042_1821, w_042_1822, w_042_1825, w_042_1826, w_042_1828, w_042_1829, w_042_1830, w_042_1831, w_042_1832, w_042_1836, w_042_1839, w_042_1843, w_042_1845, w_042_1846, w_042_1848, w_042_1849, w_042_1853, w_042_1854, w_042_1855, w_042_1856, w_042_1859, w_042_1862, w_042_1865, w_042_1866, w_042_1868, w_042_1870, w_042_1872, w_042_1873, w_042_1874, w_042_1875, w_042_1877, w_042_1878, w_042_1881, w_042_1882, w_042_1885, w_042_1888, w_042_1889, w_042_1890, w_042_1893, w_042_1896, w_042_1898, w_042_1899, w_042_1901, w_042_1902, w_042_1903, w_042_1906, w_042_1910, w_042_1912, w_042_1913, w_042_1914, w_042_1917, w_042_1918, w_042_1920, w_042_1921, w_042_1923, w_042_1927, w_042_1928, w_042_1930, w_042_1933, w_042_1934, w_042_1935, w_042_1936, w_042_1939, w_042_1942, w_042_1943, w_042_1945, w_042_1948, w_042_1949, w_042_1950, w_042_1951, w_042_1955, w_042_1956, w_042_1957, w_042_1958, w_042_1959, w_042_1961, w_042_1963, w_042_1964, w_042_1966, w_042_1967, w_042_1969, w_042_1971, w_042_1972, w_042_1973, w_042_1974, w_042_1979, w_042_1982, w_042_1984, w_042_1985, w_042_1986, w_042_1987, w_042_1990, w_042_1992, w_042_1993, w_042_1995, w_042_1997, w_042_1998, w_042_1999, w_042_2001, w_042_2004, w_042_2008, w_042_2010, w_042_2011, w_042_2016, w_042_2020, w_042_2023, w_042_2024, w_042_2026, w_042_2027, w_042_2028, w_042_2029, w_042_2031, w_042_2032, w_042_2036, w_042_2037, w_042_2039, w_042_2045, w_042_2049, w_042_2052, w_042_2055, w_042_2056, w_042_2057, w_042_2058, w_042_2061, w_042_2063, w_042_2064, w_042_2067, w_042_2068, w_042_2069, w_042_2070, w_042_2075, w_042_2076, w_042_2077, w_042_2082, w_042_2083, w_042_2084, w_042_2085, w_042_2087, w_042_2095, w_042_2096, w_042_2097, w_042_2098, w_042_2102, w_042_2103, w_042_2104, w_042_2106, w_042_2107, w_042_2108, w_042_2109, w_042_2110, w_042_2111, w_042_2112, w_042_2115, w_042_2116, w_042_2117, w_042_2118, w_042_2120, w_042_2121, w_042_2123, w_042_2127, w_042_2131, w_042_2132, w_042_2137, w_042_2138, w_042_2139, w_042_2140, w_042_2141, w_042_2143, w_042_2145, w_042_2146, w_042_2149, w_042_2150, w_042_2151, w_042_2152, w_042_2153, w_042_2154, w_042_2156, w_042_2157, w_042_2160, w_042_2161, w_042_2162, w_042_2163, w_042_2165, w_042_2167, w_042_2168, w_042_2171, w_042_2173, w_042_2177, w_042_2179, w_042_2181, w_042_2182, w_042_2185, w_042_2187, w_042_2188, w_042_2190, w_042_2192, w_042_2193, w_042_2194, w_042_2195, w_042_2197, w_042_2199, w_042_2202, w_042_2203, w_042_2204, w_042_2205, w_042_2206, w_042_2208, w_042_2209, w_042_2212, w_042_2215, w_042_2217, w_042_2221, w_042_2225, w_042_2231, w_042_2233, w_042_2234, w_042_2236, w_042_2237, w_042_2239, w_042_2240, w_042_2243, w_042_2244, w_042_2245, w_042_2246, w_042_2248, w_042_2250, w_042_2251, w_042_2254, w_042_2255, w_042_2258, w_042_2259, w_042_2261, w_042_2266, w_042_2272, w_042_2273, w_042_2274, w_042_2276, w_042_2278, w_042_2280, w_042_2284, w_042_2286, w_042_2290, w_042_2292, w_042_2293, w_042_2294, w_042_2295, w_042_2297, w_042_2299, w_042_2301, w_042_2303, w_042_2306, w_042_2307, w_042_2308, w_042_2309, w_042_2311, w_042_2315, w_042_2318, w_042_2321, w_042_2323, w_042_2324, w_042_2325, w_042_2326, w_042_2328, w_042_2329, w_042_2331, w_042_2333, w_042_2334, w_042_2335, w_042_2337, w_042_2338, w_042_2339, w_042_2340, w_042_2345, w_042_2346, w_042_2348, w_042_2349, w_042_2350, w_042_2352, w_042_2353, w_042_2354, w_042_2355, w_042_2356, w_042_2358, w_042_2359, w_042_2360, w_042_2361, w_042_2363, w_042_2366, w_042_2369, w_042_2372, w_042_2377, w_042_2378, w_042_2380, w_042_2382, w_042_2384, w_042_2385, w_042_2387, w_042_2388, w_042_2391, w_042_2392, w_042_2394, w_042_2396, w_042_2397, w_042_2400, w_042_2401, w_042_2403, w_042_2405, w_042_2407, w_042_2410, w_042_2411, w_042_2412, w_042_2414, w_042_2415, w_042_2416, w_042_2417, w_042_2421, w_042_2422, w_042_2423, w_042_2425, w_042_2427, w_042_2428, w_042_2430, w_042_2431, w_042_2433, w_042_2435, w_042_2437, w_042_2438, w_042_2439, w_042_2443, w_042_2445, w_042_2447, w_042_2450, w_042_2451, w_042_2453, w_042_2454, w_042_2457, w_042_2458, w_042_2460, w_042_2462, w_042_2464, w_042_2467, w_042_2469, w_042_2473, w_042_2474, w_042_2475, w_042_2477, w_042_2478, w_042_2483, w_042_2486, w_042_2487, w_042_2488, w_042_2489, w_042_2490, w_042_2491, w_042_2493, w_042_2494, w_042_2496, w_042_2497, w_042_2498, w_042_2499, w_042_2500, w_042_2502, w_042_2503, w_042_2512, w_042_2513, w_042_2514, w_042_2519, w_042_2522, w_042_2524, w_042_2528, w_042_2532, w_042_2533, w_042_2534, w_042_2540, w_042_2542, w_042_2543, w_042_2546, w_042_2548, w_042_2549, w_042_2550, w_042_2551, w_042_2552, w_042_2553, w_042_2555, w_042_2557, w_042_2558, w_042_2560, w_042_2564, w_042_2567, w_042_2569, w_042_2571, w_042_2572, w_042_2574, w_042_2576, w_042_2577, w_042_2578, w_042_2581, w_042_2582, w_042_2583, w_042_2585, w_042_2586, w_042_2587, w_042_2588, w_042_2589, w_042_2591, w_042_2595, w_042_2597, w_042_2599, w_042_2603, w_042_2605, w_042_2607, w_042_2608, w_042_2610, w_042_2611, w_042_2612, w_042_2613, w_042_2620, w_042_2621, w_042_2622, w_042_2623, w_042_2624, w_042_2626, w_042_2627, w_042_2628, w_042_2629, w_042_2630, w_042_2632, w_042_2633, w_042_2634, w_042_2636, w_042_2637, w_042_2638, w_042_2642, w_042_2647, w_042_2649, w_042_2650, w_042_2651, w_042_2653, w_042_2654, w_042_2656, w_042_2657, w_042_2658, w_042_2659, w_042_2660, w_042_2662, w_042_2663, w_042_2664, w_042_2665, w_042_2666, w_042_2667, w_042_2668, w_042_2670, w_042_2675, w_042_2676, w_042_2682, w_042_2684, w_042_2685, w_042_2686, w_042_2687, w_042_2688, w_042_2689, w_042_2692, w_042_2693, w_042_2694, w_042_2695, w_042_2696, w_042_2697, w_042_2698, w_042_2700, w_042_2701, w_042_2702, w_042_2705, w_042_2706, w_042_2707, w_042_2709, w_042_2710, w_042_2712, w_042_2713, w_042_2715, w_042_2716, w_042_2719, w_042_2720, w_042_2725, w_042_2726, w_042_2727, w_042_2728, w_042_2730, w_042_2731, w_042_2733, w_042_2734, w_042_2735, w_042_2737, w_042_2740, w_042_2741, w_042_2742, w_042_2743, w_042_2745, w_042_2746, w_042_2748, w_042_2750, w_042_2754, w_042_2755, w_042_2756, w_042_2757, w_042_2759, w_042_2761, w_042_2764, w_042_2765, w_042_2767, w_042_2768, w_042_2769, w_042_2770, w_042_2773, w_042_2775, w_042_2777, w_042_2778, w_042_2781, w_042_2782, w_042_2783, w_042_2784, w_042_2785, w_042_2787, w_042_2788, w_042_2790, w_042_2792, w_042_2793, w_042_2794, w_042_2795, w_042_2796, w_042_2797, w_042_2799, w_042_2800, w_042_2803, w_042_2804, w_042_2805, w_042_2807, w_042_2809, w_042_2810, w_042_2812, w_042_2814, w_042_2815, w_042_2816, w_042_2817, w_042_2820, w_042_2821, w_042_2822, w_042_2823, w_042_2824, w_042_2828, w_042_2830, w_042_2831, w_042_2833, w_042_2834, w_042_2835, w_042_2836, w_042_2842, w_042_2843, w_042_2844, w_042_2846, w_042_2848, w_042_2849, w_042_2850, w_042_2851, w_042_2853, w_042_2856, w_042_2857, w_042_2859, w_042_2864, w_042_2868, w_042_2869, w_042_2874, w_042_2875, w_042_2876, w_042_2879, w_042_2880, w_042_2881, w_042_2883, w_042_2884, w_042_2885, w_042_2886, w_042_2887, w_042_2888, w_042_2889, w_042_2893, w_042_2896, w_042_2897, w_042_2898, w_042_2899, w_042_2900, w_042_2901, w_042_2902, w_042_2904, w_042_2905, w_042_2906, w_042_2909, w_042_2911, w_042_2916, w_042_2917, w_042_2918, w_042_2922, w_042_2927, w_042_2930, w_042_2931, w_042_2932, w_042_2933, w_042_2934, w_042_2940, w_042_2941, w_042_2943, w_042_2944, w_042_2945, w_042_2946, w_042_2947, w_042_2948, w_042_2949, w_042_2950, w_042_2951, w_042_2954, w_042_2959, w_042_2961, w_042_2962, w_042_2964, w_042_2965, w_042_2966, w_042_2967, w_042_2968, w_042_2969, w_042_2971, w_042_2977, w_042_2979, w_042_2981, w_042_2983, w_042_2984, w_042_2987, w_042_2988, w_042_2989, w_042_2992, w_042_2994, w_042_2996, w_042_2997, w_042_2999, w_042_3001, w_042_3002, w_042_3003, w_042_3004, w_042_3005, w_042_3008, w_042_3009, w_042_3012, w_042_3013, w_042_3014, w_042_3015, w_042_3017, w_042_3018, w_042_3021, w_042_3022, w_042_3023, w_042_3029, w_042_3030, w_042_3033, w_042_3035, w_042_3038, w_042_3039, w_042_3041, w_042_3042, w_042_3044, w_042_3045, w_042_3046, w_042_3048, w_042_3050, w_042_3051, w_042_3057, w_042_3058, w_042_3061, w_042_3064, w_042_3065, w_042_3067, w_042_3068, w_042_3070, w_042_3071, w_042_3073, w_042_3074, w_042_3078, w_042_3079, w_042_3080, w_042_3081, w_042_3083, w_042_3086, w_042_3089, w_042_3091, w_042_3092, w_042_3094, w_042_3096, w_042_3098, w_042_3100, w_042_3103, w_042_3105, w_042_3107, w_042_3114, w_042_3116, w_042_3118, w_042_3119, w_042_3121, w_042_3122, w_042_3123, w_042_3124, w_042_3127, w_042_3129, w_042_3132, w_042_3133, w_042_3134, w_042_3135, w_042_3136, w_042_3141, w_042_3144, w_042_3145, w_042_3146, w_042_3147, w_042_3151, w_042_3154, w_042_3155, w_042_3156, w_042_3157, w_042_3158, w_042_3160, w_042_3164, w_042_3166, w_042_3169, w_042_3171, w_042_3172, w_042_3174, w_042_3175, w_042_3176, w_042_3177, w_042_3179, w_042_3181, w_042_3186, w_042_3187, w_042_3190, w_042_3191, w_042_3192, w_042_3194, w_042_3196, w_042_3199, w_042_3201, w_042_3203, w_042_3206, w_042_3209, w_042_3211, w_042_3214, w_042_3215, w_042_3217, w_042_3218, w_042_3220, w_042_3223, w_042_3224, w_042_3226, w_042_3228, w_042_3230, w_042_3232, w_042_3234, w_042_3238, w_042_3239, w_042_3242, w_042_3244, w_042_3245, w_042_3246, w_042_3247, w_042_3248, w_042_3250, w_042_3252, w_042_3253, w_042_3254, w_042_3255, w_042_3257, w_042_3261, w_042_3263, w_042_3265, w_042_3267, w_042_3268, w_042_3269, w_042_3270, w_042_3271, w_042_3275, w_042_3279, w_042_3280, w_042_3282, w_042_3283, w_042_3285, w_042_3288, w_042_3295, w_042_3296, w_042_3298, w_042_3299, w_042_3300, w_042_3301, w_042_3306, w_042_3308, w_042_3309, w_042_3310, w_042_3311, w_042_3313, w_042_3319, w_042_3322, w_042_3324, w_042_3325, w_042_3326, w_042_3327, w_042_3331, w_042_3332, w_042_3336, w_042_3340, w_042_3341, w_042_3343, w_042_3344, w_042_3350, w_042_3351, w_042_3353, w_042_3355, w_042_3356, w_042_3357, w_042_3359, w_042_3360, w_042_3361, w_042_3362, w_042_3364, w_042_3366, w_042_3370, w_042_3374, w_042_3377, w_042_3378, w_042_3380, w_042_3383, w_042_3384, w_042_3385, w_042_3386, w_042_3389, w_042_3390, w_042_3391, w_042_3392, w_042_3393, w_042_3394, w_042_3396, w_042_3398, w_042_3403, w_042_3406, w_042_3407, w_042_3408, w_042_3409, w_042_3410, w_042_3412, w_042_3415, w_042_3418, w_042_3419, w_042_3426, w_042_3427, w_042_3429, w_042_3430, w_042_3431, w_042_3432, w_042_3433, w_042_3434, w_042_3436, w_042_3439, w_042_3440, w_042_3441, w_042_3442, w_042_3443, w_042_3444, w_042_3445, w_042_3448, w_042_3450, w_042_3452, w_042_3454, w_042_3455, w_042_3458, w_042_3459, w_042_3460, w_042_3461, w_042_3462, w_042_3463, w_042_3464, w_042_3466, w_042_3467, w_042_3469, w_042_3470, w_042_3471, w_042_3475, w_042_3477, w_042_3481, w_042_3482, w_042_3484, w_042_3485, w_042_3493, w_042_3494, w_042_3495, w_042_3496, w_042_3498, w_042_3502, w_042_3505, w_042_3506, w_042_3507, w_042_3510, w_042_3513, w_042_3515, w_042_3516, w_042_3517, w_042_3519, w_042_3520, w_042_3523, w_042_3524, w_042_3525, w_042_3527, w_042_3529, w_042_3531, w_042_3534, w_042_3537, w_042_3538, w_042_3540, w_042_3541, w_042_3543, w_042_3544, w_042_3545, w_042_3550, w_042_3551, w_042_3555, w_042_3556, w_042_3557, w_042_3558, w_042_3559, w_042_3560, w_042_3561, w_042_3562, w_042_3565, w_042_3566, w_042_3568, w_042_3570, w_042_3571, w_042_3573, w_042_3574, w_042_3575, w_042_3577, w_042_3578, w_042_3579, w_042_3581, w_042_3583, w_042_3586, w_042_3587, w_042_3588, w_042_3589, w_042_3591, w_042_3593, w_042_3595, w_042_3596, w_042_3598, w_042_3601, w_042_3603, w_042_3606, w_042_3608, w_042_3609, w_042_3610, w_042_3611, w_042_3613, w_042_3615, w_042_3616, w_042_3622, w_042_3623, w_042_3624, w_042_3625, w_042_3627, w_042_3630, w_042_3634, w_042_3635, w_042_3636, w_042_3637, w_042_3638, w_042_3639, w_042_3641, w_042_3642, w_042_3645, w_042_3647, w_042_3649, w_042_3650, w_042_3651, w_042_3653, w_042_3654, w_042_3660, w_042_3663, w_042_3664, w_042_3665, w_042_3667, w_042_3668, w_042_3669, w_042_3671, w_042_3672, w_042_3673, w_042_3674, w_042_3675, w_042_3690, w_042_3691, w_042_3696, w_042_3697, w_042_3698, w_042_3699, w_042_3701, w_042_3702, w_042_3704, w_042_3705, w_042_3706, w_042_3707, w_042_3708, w_042_3711, w_042_3712, w_042_3713, w_042_3714, w_042_3717, w_042_3719, w_042_3721, w_042_3724, w_042_3727, w_042_3728, w_042_3731, w_042_3732, w_042_3734, w_042_3735, w_042_3738, w_042_3739, w_042_3741, w_042_3743, w_042_3744, w_042_3746, w_042_3747, w_042_3749, w_042_3751, w_042_3752, w_042_3754, w_042_3756, w_042_3758, w_042_3760, w_042_3761, w_042_3762, w_042_3763, w_042_3768, w_042_3769, w_042_3770, w_042_3771, w_042_3772, w_042_3773, w_042_3777, w_042_3779, w_042_3780, w_042_3784, w_042_3785, w_042_3787, w_042_3788, w_042_3789, w_042_3792, w_042_3793, w_042_3794, w_042_3795, w_042_3796, w_042_3799, w_042_3801, w_042_3803, w_042_3804, w_042_3806, w_042_3807, w_042_3808, w_042_3810, w_042_3812, w_042_3814, w_042_3816, w_042_3819, w_042_3820, w_042_3821, w_042_3824, w_042_3826, w_042_3829, w_042_3832, w_042_3833, w_042_3834, w_042_3835, w_042_3837, w_042_3838, w_042_3840, w_042_3842, w_042_3843, w_042_3844, w_042_3846, w_042_3849, w_042_3850, w_042_3851, w_042_3855, w_042_3856, w_042_3860, w_042_3863, w_042_3864, w_042_3866, w_042_3867, w_042_3869, w_042_3872, w_042_3876, w_042_3878, w_042_3879, w_042_3881, w_042_3886, w_042_3890, w_042_3891, w_042_3899, w_042_3901, w_042_3902, w_042_3903, w_042_3906, w_042_3907, w_042_3909, w_042_3912, w_042_3914, w_042_3915, w_042_3918, w_042_3919, w_042_3922, w_042_3923, w_042_3924, w_042_3926, w_042_3929, w_042_3930, w_042_3932, w_042_3933, w_042_3934, w_042_3935, w_042_3936, w_042_3938, w_042_3939, w_042_3940, w_042_3941, w_042_3942, w_042_3943, w_042_3944, w_042_3946, w_042_3949, w_042_3950, w_042_3951, w_042_3953, w_042_3955, w_042_3956, w_042_3957, w_042_3959, w_042_3962, w_042_3963, w_042_3964, w_042_3967, w_042_3968, w_042_3969, w_042_3970, w_042_3971, w_042_3972, w_042_3974, w_042_3975, w_042_3978, w_042_3982, w_042_3983, w_042_3984, w_042_3985, w_042_3987, w_042_3989, w_042_3991, w_042_3992, w_042_3994, w_042_3996, w_042_3998, w_042_3999, w_042_4007, w_042_4009, w_042_4013, w_042_4014, w_042_4015, w_042_4022, w_042_4024, w_042_4025, w_042_4026, w_042_4027, w_042_4028, w_042_4029, w_042_4030, w_042_4033, w_042_4035, w_042_4036, w_042_4038, w_042_4039, w_042_4040, w_042_4041, w_042_4042, w_042_4043, w_042_4045, w_042_4049, w_042_4050, w_042_4051, w_042_4052, w_042_4053, w_042_4055, w_042_4056, w_042_4058, w_042_4061, w_042_4062, w_042_4065, w_042_4067, w_042_4068, w_042_4069, w_042_4070, w_042_4073, w_042_4076, w_042_4078, w_042_4079, w_042_4082, w_042_4083, w_042_4084, w_042_4086, w_042_4087, w_042_4089, w_042_4090, w_042_4092, w_042_4093, w_042_4095, w_042_4096, w_042_4097, w_042_4100, w_042_4104, w_042_4107, w_042_4109, w_042_4110, w_042_4112, w_042_4113, w_042_4117, w_042_4118, w_042_4119, w_042_4120, w_042_4122, w_042_4123, w_042_4124, w_042_4125, w_042_4126, w_042_4127, w_042_4133, w_042_4134, w_042_4135, w_042_4136, w_042_4137, w_042_4138, w_042_4139, w_042_4140, w_042_4143, w_042_4145, w_042_4146, w_042_4147, w_042_4148, w_042_4149, w_042_4151, w_042_4154, w_042_4155, w_042_4156, w_042_4157, w_042_4160, w_042_4162, w_042_4163, w_042_4164, w_042_4166, w_042_4167, w_042_4171, w_042_4174, w_042_4176, w_042_4178, w_042_4179, w_042_4180, w_042_4183, w_042_4184, w_042_4185, w_042_4186, w_042_4189, w_042_4192, w_042_4196, w_042_4197, w_042_4198, w_042_4201, w_042_4202, w_042_4203, w_042_4206, w_042_4207, w_042_4208, w_042_4211, w_042_4212, w_042_4216, w_042_4219, w_042_4220, w_042_4221, w_042_4222, w_042_4223, w_042_4224, w_042_4225, w_042_4226, w_042_4227, w_042_4228, w_042_4229, w_042_4230, w_042_4231, w_042_4232, w_042_4233, w_042_4235, w_042_4236, w_042_4240, w_042_4243, w_042_4245, w_042_4247, w_042_4250, w_042_4251, w_042_4254, w_042_4255, w_042_4256, w_042_4257, w_042_4258, w_042_4260, w_042_4262, w_042_4264, w_042_4268, w_042_4269, w_042_4271, w_042_4273, w_042_4278, w_042_4279, w_042_4281, w_042_4282, w_042_4283, w_042_4286, w_042_4287, w_042_4288, w_042_4289, w_042_4295, w_042_4297, w_042_4298, w_042_4299, w_042_4300, w_042_4301, w_042_4302, w_042_4303, w_042_4307, w_042_4308, w_042_4309, w_042_4313, w_042_4315, w_042_4316, w_042_4318, w_042_4319, w_042_4322, w_042_4328, w_042_4329, w_042_4331, w_042_4332, w_042_4337, w_042_4338, w_042_4342, w_042_4344, w_042_4346, w_042_4349, w_042_4351, w_042_4352, w_042_4354, w_042_4356, w_042_4360, w_042_4361, w_042_4362, w_042_4364, w_042_4365, w_042_4366, w_042_4369, w_042_4371, w_042_4372, w_042_4375, w_042_4377, w_042_4378, w_042_4380, w_042_4383, w_042_4384, w_042_4387, w_042_4388, w_042_4389, w_042_4391, w_042_4392, w_042_4396, w_042_4397, w_042_4398, w_042_4402, w_042_4403, w_042_4405, w_042_4406, w_042_4407, w_042_4410, w_042_4411, w_042_4414, w_042_4415, w_042_4418, w_042_4420, w_042_4421, w_042_4424, w_042_4425, w_042_4426, w_042_4427, w_042_4428, w_042_4431, w_042_4432, w_042_4434, w_042_4435, w_042_4436, w_042_4437, w_042_4438, w_042_4442, w_042_4444, w_042_4447, w_042_4449, w_042_4450, w_042_4451, w_042_4452, w_042_4455, w_042_4456, w_042_4457, w_042_4459, w_042_4461, w_042_4465, w_042_4467, w_042_4468, w_042_4469, w_042_4475, w_042_4476, w_042_4477, w_042_4478, w_042_4479, w_042_4481, w_042_4482, w_042_4483, w_042_4485, w_042_4487, w_042_4489, w_042_4490, w_042_4493, w_042_4494, w_042_4495, w_042_4497, w_042_4498, w_042_4499, w_042_4500, w_042_4501, w_042_4504, w_042_4505, w_042_4507, w_042_4508, w_042_4510, w_042_4512, w_042_4514, w_042_4515, w_042_4517, w_042_4518, w_042_4521, w_042_4523, w_042_4525, w_042_4526, w_042_4531, w_042_4533, w_042_4535, w_042_4536, w_042_4539, w_042_4541, w_042_4544, w_042_4545, w_042_4549, w_042_4550, w_042_4551, w_042_4552, w_042_4553, w_042_4555, w_042_4556, w_042_4558, w_042_4559, w_042_4560, w_042_4563, w_042_4567, w_042_4568, w_042_4569, w_042_4570, w_042_4571, w_042_4573, w_042_4574, w_042_4577, w_042_4578, w_042_4580, w_042_4582, w_042_4588, w_042_4589, w_042_4591, w_042_4592, w_042_4594, w_042_4597, w_042_4598, w_042_4599, w_042_4601, w_042_4602, w_042_4603, w_042_4605, w_042_4606, w_042_4607, w_042_4608, w_042_4609, w_042_4610, w_042_4611, w_042_4612, w_042_4613, w_042_4614, w_042_4615, w_042_4618, w_042_4620, w_042_4625, w_042_4626, w_042_4631, w_042_4633, w_042_4634, w_042_4635, w_042_4639, w_042_4640, w_042_4645, w_042_4648, w_042_4651, w_042_4652, w_042_4653, w_042_4656, w_042_4659, w_042_4663, w_042_4664, w_042_4665, w_042_4666, w_042_4667, w_042_4669, w_042_4672;
  wire w_043_000, w_043_002, w_043_003, w_043_004, w_043_005, w_043_006, w_043_009, w_043_010, w_043_011, w_043_012, w_043_013, w_043_015, w_043_016, w_043_017, w_043_019, w_043_022, w_043_023, w_043_025, w_043_026, w_043_027, w_043_028, w_043_029, w_043_030, w_043_032, w_043_034, w_043_035, w_043_036, w_043_037, w_043_039, w_043_040, w_043_041, w_043_042, w_043_043, w_043_044, w_043_045, w_043_046, w_043_047, w_043_048, w_043_049, w_043_050, w_043_051, w_043_052, w_043_054, w_043_056, w_043_058, w_043_059, w_043_060, w_043_061, w_043_062, w_043_063, w_043_065, w_043_066, w_043_067, w_043_070, w_043_071, w_043_072, w_043_073, w_043_074, w_043_075, w_043_076, w_043_077, w_043_080, w_043_081, w_043_083, w_043_084, w_043_085, w_043_086, w_043_087, w_043_088, w_043_089, w_043_090, w_043_091, w_043_092, w_043_093, w_043_094, w_043_095, w_043_097, w_043_098, w_043_099, w_043_101, w_043_102, w_043_103, w_043_104, w_043_105, w_043_107, w_043_108, w_043_109, w_043_110, w_043_111, w_043_113, w_043_114, w_043_115, w_043_117, w_043_118, w_043_119, w_043_120, w_043_121, w_043_122, w_043_123, w_043_124, w_043_125, w_043_127, w_043_128, w_043_129, w_043_130, w_043_132, w_043_134, w_043_136, w_043_137, w_043_138, w_043_139, w_043_141, w_043_142, w_043_143, w_043_144, w_043_145, w_043_146, w_043_147, w_043_148, w_043_150, w_043_151, w_043_152, w_043_155, w_043_157, w_043_158, w_043_159, w_043_162, w_043_163, w_043_164, w_043_165, w_043_168, w_043_169, w_043_170, w_043_171, w_043_172, w_043_173, w_043_174, w_043_175, w_043_177, w_043_178, w_043_179, w_043_181, w_043_182, w_043_183, w_043_184, w_043_186, w_043_187, w_043_188, w_043_189, w_043_190, w_043_192, w_043_193, w_043_194, w_043_195, w_043_196, w_043_198, w_043_199, w_043_200, w_043_201, w_043_202, w_043_203, w_043_204, w_043_205, w_043_206, w_043_207, w_043_208, w_043_211, w_043_212, w_043_213, w_043_215, w_043_216, w_043_217, w_043_218, w_043_219, w_043_221, w_043_222, w_043_224, w_043_225, w_043_226, w_043_227, w_043_228, w_043_231, w_043_233, w_043_234, w_043_235, w_043_236, w_043_237, w_043_238, w_043_239, w_043_241, w_043_242, w_043_243, w_043_244, w_043_245, w_043_248, w_043_249, w_043_250, w_043_251, w_043_253, w_043_254, w_043_255, w_043_256, w_043_258, w_043_259, w_043_260, w_043_262, w_043_264, w_043_265, w_043_266, w_043_267, w_043_268, w_043_269, w_043_270, w_043_272, w_043_273, w_043_274, w_043_275, w_043_279, w_043_280, w_043_281, w_043_282, w_043_283, w_043_284, w_043_285, w_043_286, w_043_287, w_043_288, w_043_289, w_043_290, w_043_294, w_043_295, w_043_296, w_043_297, w_043_298, w_043_299, w_043_300, w_043_301, w_043_302, w_043_303, w_043_304, w_043_305, w_043_306, w_043_307, w_043_308, w_043_309, w_043_310, w_043_311, w_043_312, w_043_313, w_043_314, w_043_316, w_043_317, w_043_318, w_043_319, w_043_320, w_043_322, w_043_323, w_043_324, w_043_325, w_043_326, w_043_327, w_043_328, w_043_329, w_043_330, w_043_331, w_043_332, w_043_333, w_043_334, w_043_335, w_043_336, w_043_339, w_043_340, w_043_342, w_043_344, w_043_345, w_043_347, w_043_348, w_043_349, w_043_350, w_043_351, w_043_357, w_043_358, w_043_360, w_043_362, w_043_364, w_043_365, w_043_366, w_043_367, w_043_370, w_043_371, w_043_372, w_043_373, w_043_374, w_043_375, w_043_378, w_043_379, w_043_380, w_043_381, w_043_382, w_043_383, w_043_385, w_043_386, w_043_387, w_043_389, w_043_390, w_043_391, w_043_392, w_043_394, w_043_395, w_043_396, w_043_397, w_043_398, w_043_399, w_043_400, w_043_401, w_043_402, w_043_403, w_043_404, w_043_406, w_043_407, w_043_408, w_043_411, w_043_412, w_043_413, w_043_414, w_043_415, w_043_417, w_043_418, w_043_420, w_043_421, w_043_423, w_043_424, w_043_425, w_043_426, w_043_427, w_043_428, w_043_430, w_043_431, w_043_433, w_043_434, w_043_435, w_043_436, w_043_439, w_043_440, w_043_441, w_043_442, w_043_444, w_043_445, w_043_446, w_043_447, w_043_448, w_043_449, w_043_450, w_043_451, w_043_453, w_043_454, w_043_455, w_043_456, w_043_459, w_043_460, w_043_462, w_043_463, w_043_465, w_043_467, w_043_468, w_043_469, w_043_471, w_043_472, w_043_473, w_043_474, w_043_476, w_043_477, w_043_478, w_043_479, w_043_480, w_043_482, w_043_483, w_043_484, w_043_487, w_043_488, w_043_489, w_043_492, w_043_494, w_043_495, w_043_496, w_043_497, w_043_499, w_043_500, w_043_501, w_043_502, w_043_503, w_043_504, w_043_505, w_043_506, w_043_507, w_043_508, w_043_509, w_043_510, w_043_511, w_043_513, w_043_514, w_043_515, w_043_516, w_043_517, w_043_518, w_043_519, w_043_520, w_043_521, w_043_522, w_043_523, w_043_524, w_043_525, w_043_526, w_043_527, w_043_529, w_043_530, w_043_531, w_043_532, w_043_533, w_043_534, w_043_535, w_043_537, w_043_538, w_043_539, w_043_540, w_043_541, w_043_542, w_043_543, w_043_545, w_043_547, w_043_548, w_043_550, w_043_551, w_043_552, w_043_553, w_043_554, w_043_555, w_043_556, w_043_557, w_043_558, w_043_559, w_043_560, w_043_561, w_043_562, w_043_563, w_043_568, w_043_569, w_043_570, w_043_571, w_043_572, w_043_573, w_043_574, w_043_576, w_043_578, w_043_579, w_043_580, w_043_581, w_043_582, w_043_583, w_043_584, w_043_585, w_043_586, w_043_587, w_043_588, w_043_589, w_043_591, w_043_592, w_043_593, w_043_594, w_043_595, w_043_596, w_043_597, w_043_599, w_043_601, w_043_602, w_043_603, w_043_604, w_043_605, w_043_606, w_043_607, w_043_608, w_043_610, w_043_611, w_043_612, w_043_614, w_043_616, w_043_617, w_043_619, w_043_620, w_043_621, w_043_622, w_043_623, w_043_626, w_043_627, w_043_628, w_043_629, w_043_630, w_043_631, w_043_632, w_043_633, w_043_635, w_043_637, w_043_638, w_043_639, w_043_640, w_043_642, w_043_644, w_043_645, w_043_647, w_043_648, w_043_649, w_043_650, w_043_651, w_043_652, w_043_653, w_043_654, w_043_655, w_043_656, w_043_658, w_043_659, w_043_660, w_043_661, w_043_662, w_043_663, w_043_664, w_043_666, w_043_667, w_043_669, w_043_671, w_043_672, w_043_673, w_043_674, w_043_675, w_043_676, w_043_677, w_043_678, w_043_679, w_043_680, w_043_681, w_043_684, w_043_685, w_043_686, w_043_688, w_043_689, w_043_691, w_043_692, w_043_693, w_043_694, w_043_695, w_043_696, w_043_699, w_043_700, w_043_701, w_043_703, w_043_704, w_043_705, w_043_706, w_043_707, w_043_708, w_043_712, w_043_714, w_043_715, w_043_717, w_043_719, w_043_722, w_043_723, w_043_724, w_043_728, w_043_730, w_043_731, w_043_733, w_043_734, w_043_735, w_043_736, w_043_737, w_043_738, w_043_739, w_043_740, w_043_741, w_043_743, w_043_744, w_043_745, w_043_746, w_043_747, w_043_748, w_043_749, w_043_752, w_043_756, w_043_757, w_043_758, w_043_759, w_043_760, w_043_761, w_043_762, w_043_763, w_043_765, w_043_766, w_043_767, w_043_768, w_043_769, w_043_770, w_043_771, w_043_772, w_043_773, w_043_774, w_043_775, w_043_776, w_043_778, w_043_779, w_043_780, w_043_781, w_043_782, w_043_783, w_043_784, w_043_785, w_043_787, w_043_788, w_043_789, w_043_790, w_043_791, w_043_792, w_043_793, w_043_796, w_043_797, w_043_798, w_043_800, w_043_802, w_043_803, w_043_804, w_043_805, w_043_806, w_043_807, w_043_808, w_043_809, w_043_810, w_043_811, w_043_813, w_043_816, w_043_818, w_043_819, w_043_820, w_043_821, w_043_822, w_043_823, w_043_824, w_043_826, w_043_827, w_043_828, w_043_829, w_043_830, w_043_831, w_043_832, w_043_833, w_043_834, w_043_837, w_043_839, w_043_840, w_043_841, w_043_842, w_043_844, w_043_845, w_043_846, w_043_847, w_043_848, w_043_849, w_043_850, w_043_851, w_043_852, w_043_854, w_043_855, w_043_856, w_043_857, w_043_859, w_043_860, w_043_861, w_043_862, w_043_863, w_043_864, w_043_865, w_043_866, w_043_867, w_043_868, w_043_871, w_043_872, w_043_873, w_043_874, w_043_875, w_043_876, w_043_878, w_043_879, w_043_880, w_043_881, w_043_883, w_043_884, w_043_885, w_043_887, w_043_888, w_043_889, w_043_890, w_043_891, w_043_892, w_043_893, w_043_894, w_043_895, w_043_896, w_043_897, w_043_898, w_043_899, w_043_901, w_043_902, w_043_903, w_043_904, w_043_905, w_043_906, w_043_907, w_043_908, w_043_909, w_043_910, w_043_911, w_043_912, w_043_913, w_043_914, w_043_915, w_043_916, w_043_917, w_043_918, w_043_919, w_043_920, w_043_922, w_043_923, w_043_924, w_043_925, w_043_927, w_043_928, w_043_929, w_043_930, w_043_931, w_043_932, w_043_933, w_043_934, w_043_935, w_043_936, w_043_937, w_043_938, w_043_941, w_043_942, w_043_943, w_043_944, w_043_945, w_043_946, w_043_947, w_043_948, w_043_950, w_043_951, w_043_952, w_043_953, w_043_954, w_043_956, w_043_957, w_043_958, w_043_959, w_043_961, w_043_962, w_043_963, w_043_964, w_043_965, w_043_966, w_043_968, w_043_969, w_043_970, w_043_971, w_043_972, w_043_974, w_043_975, w_043_976, w_043_977, w_043_978, w_043_979, w_043_980, w_043_981, w_043_982, w_043_983, w_043_984, w_043_987, w_043_988, w_043_989, w_043_990, w_043_993, w_043_994, w_043_995, w_043_996, w_043_997, w_043_999, w_043_1000, w_043_1001, w_043_1003, w_043_1004, w_043_1007, w_043_1008, w_043_1009, w_043_1010, w_043_1011, w_043_1012, w_043_1013, w_043_1015, w_043_1016, w_043_1017, w_043_1020, w_043_1021, w_043_1022, w_043_1023, w_043_1024, w_043_1026, w_043_1028, w_043_1029, w_043_1030, w_043_1031, w_043_1032, w_043_1033, w_043_1034, w_043_1035, w_043_1037, w_043_1038, w_043_1039, w_043_1040, w_043_1041, w_043_1043, w_043_1044, w_043_1045, w_043_1046, w_043_1048, w_043_1049, w_043_1050, w_043_1051, w_043_1053, w_043_1054, w_043_1056, w_043_1057, w_043_1058, w_043_1061, w_043_1062, w_043_1064, w_043_1065, w_043_1066, w_043_1067, w_043_1069, w_043_1070, w_043_1071, w_043_1072, w_043_1073, w_043_1074, w_043_1075, w_043_1076, w_043_1077, w_043_1078, w_043_1079, w_043_1080, w_043_1081, w_043_1082, w_043_1083, w_043_1084, w_043_1085, w_043_1086, w_043_1088, w_043_1089, w_043_1090, w_043_1092, w_043_1093, w_043_1095, w_043_1098, w_043_1099, w_043_1101, w_043_1104, w_043_1107, w_043_1109, w_043_1110, w_043_1111, w_043_1112, w_043_1115, w_043_1116, w_043_1118, w_043_1119, w_043_1120, w_043_1121, w_043_1122, w_043_1124, w_043_1125, w_043_1126, w_043_1127, w_043_1128, w_043_1129, w_043_1130, w_043_1131, w_043_1132, w_043_1133, w_043_1134, w_043_1135, w_043_1136, w_043_1140, w_043_1141, w_043_1142, w_043_1143, w_043_1144, w_043_1145, w_043_1146, w_043_1147, w_043_1148, w_043_1149, w_043_1150, w_043_1151, w_043_1153, w_043_1154, w_043_1155, w_043_1156, w_043_1157, w_043_1158, w_043_1159, w_043_1160, w_043_1161, w_043_1162, w_043_1164, w_043_1165, w_043_1166, w_043_1167, w_043_1168, w_043_1169, w_043_1170, w_043_1171, w_043_1172, w_043_1174, w_043_1175, w_043_1176, w_043_1177, w_043_1178, w_043_1179, w_043_1180, w_043_1181, w_043_1182, w_043_1183, w_043_1184, w_043_1185, w_043_1186, w_043_1187, w_043_1189, w_043_1190, w_043_1191, w_043_1192, w_043_1195, w_043_1196, w_043_1197, w_043_1198, w_043_1200, w_043_1202, w_043_1203, w_043_1205, w_043_1207, w_043_1208, w_043_1209, w_043_1210, w_043_1212, w_043_1214, w_043_1215, w_043_1216, w_043_1217, w_043_1218, w_043_1219, w_043_1221, w_043_1222, w_043_1224, w_043_1225, w_043_1227, w_043_1228, w_043_1229, w_043_1230, w_043_1231, w_043_1232, w_043_1234, w_043_1235, w_043_1236, w_043_1238, w_043_1239, w_043_1240, w_043_1241, w_043_1242, w_043_1243, w_043_1245, w_043_1246, w_043_1247, w_043_1248, w_043_1249, w_043_1252, w_043_1253, w_043_1255, w_043_1256, w_043_1257, w_043_1259, w_043_1260, w_043_1261, w_043_1262, w_043_1263, w_043_1264, w_043_1265, w_043_1268, w_043_1269, w_043_1270, w_043_1271, w_043_1272, w_043_1273, w_043_1274, w_043_1275, w_043_1276, w_043_1277, w_043_1278, w_043_1279, w_043_1280, w_043_1281, w_043_1282, w_043_1283, w_043_1284, w_043_1285, w_043_1286, w_043_1288, w_043_1289, w_043_1290, w_043_1291, w_043_1292, w_043_1293, w_043_1294, w_043_1295, w_043_1296, w_043_1297, w_043_1299, w_043_1300, w_043_1302, w_043_1303, w_043_1304, w_043_1305, w_043_1306, w_043_1309, w_043_1310, w_043_1311, w_043_1312, w_043_1313, w_043_1315, w_043_1316, w_043_1317, w_043_1319, w_043_1320, w_043_1321, w_043_1323, w_043_1324, w_043_1327, w_043_1328, w_043_1329, w_043_1331, w_043_1332, w_043_1333, w_043_1334, w_043_1335, w_043_1336, w_043_1337, w_043_1338, w_043_1340, w_043_1344, w_043_1346, w_043_1347, w_043_1348, w_043_1349, w_043_1350, w_043_1351, w_043_1352, w_043_1353, w_043_1354, w_043_1355, w_043_1356, w_043_1357, w_043_1358, w_043_1359, w_043_1360, w_043_1361, w_043_1364, w_043_1366, w_043_1367, w_043_1368, w_043_1371, w_043_1372, w_043_1373, w_043_1374, w_043_1375, w_043_1376, w_043_1379, w_043_1380, w_043_1382, w_043_1384, w_043_1385, w_043_1386, w_043_1388, w_043_1389, w_043_1392, w_043_1393, w_043_1394, w_043_1395, w_043_1396, w_043_1400, w_043_1402, w_043_1403, w_043_1404, w_043_1405, w_043_1406, w_043_1407, w_043_1408, w_043_1411, w_043_1412, w_043_1413, w_043_1415, w_043_1417, w_043_1418, w_043_1419, w_043_1420, w_043_1421, w_043_1422, w_043_1423, w_043_1424, w_043_1425, w_043_1426, w_043_1428, w_043_1429, w_043_1431, w_043_1432, w_043_1435, w_043_1436, w_043_1437, w_043_1438, w_043_1439, w_043_1441, w_043_1442, w_043_1444, w_043_1445, w_043_1447, w_043_1449, w_043_1450, w_043_1451, w_043_1452, w_043_1453, w_043_1454, w_043_1456, w_043_1457, w_043_1458, w_043_1459, w_043_1461, w_043_1463, w_043_1465, w_043_1466, w_043_1467, w_043_1469, w_043_1470, w_043_1471, w_043_1472, w_043_1475, w_043_1476, w_043_1477, w_043_1478, w_043_1479, w_043_1480, w_043_1481, w_043_1482, w_043_1483, w_043_1484, w_043_1485, w_043_1486, w_043_1487, w_043_1489, w_043_1491, w_043_1492, w_043_1494, w_043_1498, w_043_1499, w_043_1500, w_043_1501, w_043_1502, w_043_1505, w_043_1506, w_043_1507, w_043_1508, w_043_1509, w_043_1511, w_043_1512, w_043_1513, w_043_1514, w_043_1515, w_043_1516, w_043_1517, w_043_1518, w_043_1519, w_043_1520, w_043_1521, w_043_1523, w_043_1525, w_043_1527, w_043_1528, w_043_1529, w_043_1530, w_043_1532, w_043_1533, w_043_1534, w_043_1535, w_043_1536, w_043_1538, w_043_1539, w_043_1540, w_043_1541, w_043_1542, w_043_1543, w_043_1544, w_043_1546, w_043_1547, w_043_1548, w_043_1549, w_043_1550, w_043_1551, w_043_1552, w_043_1553, w_043_1554, w_043_1555, w_043_1556, w_043_1557, w_043_1558, w_043_1559, w_043_1560, w_043_1561, w_043_1562, w_043_1564, w_043_1565, w_043_1566, w_043_1568, w_043_1569, w_043_1570, w_043_1571, w_043_1572, w_043_1574, w_043_1575, w_043_1576, w_043_1579, w_043_1580, w_043_1581, w_043_1582, w_043_1583, w_043_1584, w_043_1586, w_043_1588, w_043_1589, w_043_1591, w_043_1593, w_043_1594, w_043_1595, w_043_1598, w_043_1599, w_043_1600, w_043_1601, w_043_1604, w_043_1606, w_043_1607, w_043_1610, w_043_1612, w_043_1613, w_043_1614, w_043_1615, w_043_1616, w_043_1617, w_043_1618, w_043_1619, w_043_1620, w_043_1622, w_043_1623, w_043_1624, w_043_1625, w_043_1626, w_043_1627, w_043_1628, w_043_1629, w_043_1630, w_043_1632, w_043_1633, w_043_1634, w_043_1635, w_043_1636, w_043_1638, w_043_1640, w_043_1642, w_043_1643, w_043_1644, w_043_1645, w_043_1646, w_043_1648, w_043_1650, w_043_1651, w_043_1652, w_043_1653, w_043_1654, w_043_1655, w_043_1656, w_043_1657, w_043_1658, w_043_1659, w_043_1660, w_043_1661, w_043_1662, w_043_1663, w_043_1664, w_043_1665, w_043_1666, w_043_1667, w_043_1668, w_043_1669, w_043_1670, w_043_1671, w_043_1673, w_043_1674, w_043_1676, w_043_1677, w_043_1678, w_043_1679, w_043_1681, w_043_1682, w_043_1683, w_043_1685, w_043_1686, w_043_1687, w_043_1688, w_043_1689, w_043_1690, w_043_1691, w_043_1692, w_043_1693, w_043_1694, w_043_1695, w_043_1696, w_043_1697, w_043_1698, w_043_1699, w_043_1701, w_043_1702, w_043_1703, w_043_1705, w_043_1706, w_043_1707, w_043_1709, w_043_1710, w_043_1711, w_043_1712, w_043_1713, w_043_1714, w_043_1715, w_043_1716, w_043_1718, w_043_1719, w_043_1720, w_043_1721, w_043_1722, w_043_1723, w_043_1724, w_043_1725, w_043_1726, w_043_1727, w_043_1729, w_043_1730, w_043_1732, w_043_1733, w_043_1735, w_043_1736, w_043_1737, w_043_1738, w_043_1741, w_043_1742, w_043_1743, w_043_1744, w_043_1745, w_043_1746, w_043_1747, w_043_1748, w_043_1750, w_043_1751, w_043_1752, w_043_1753, w_043_1755, w_043_1756, w_043_1758, w_043_1759, w_043_1760, w_043_1762, w_043_1763, w_043_1764, w_043_1765, w_043_1766, w_043_1767, w_043_1768, w_043_1769, w_043_1770, w_043_1772, w_043_1774, w_043_1775, w_043_1776, w_043_1778, w_043_1779, w_043_1781, w_043_1782, w_043_1783, w_043_1784, w_043_1785, w_043_1786, w_043_1787, w_043_1788, w_043_1789, w_043_1791, w_043_1792, w_043_1793, w_043_1795, w_043_1796, w_043_1797, w_043_1798, w_043_1799, w_043_1800, w_043_1801, w_043_1802, w_043_1804, w_043_1807, w_043_1810, w_043_1811, w_043_1812, w_043_1813, w_043_1814, w_043_1816, w_043_1817, w_043_1819, w_043_1822, w_043_1824, w_043_1825, w_043_1826, w_043_1828, w_043_1829, w_043_1830, w_043_1831, w_043_1832, w_043_1833, w_043_1834, w_043_1835, w_043_1836, w_043_1837, w_043_1838, w_043_1839, w_043_1840, w_043_1841, w_043_1842, w_043_1843, w_043_1844, w_043_1845, w_043_1846, w_043_1847, w_043_1848, w_043_1849, w_043_1850, w_043_1851, w_043_1852, w_043_1853, w_043_1854, w_043_1855, w_043_1856, w_043_1858, w_043_1859, w_043_1860, w_043_1861, w_043_1862, w_043_1863, w_043_1864, w_043_1865, w_043_1866, w_043_1867, w_043_1871, w_043_1873, w_043_1874, w_043_1875, w_043_1877, w_043_1878, w_043_1879, w_043_1880, w_043_1881, w_043_1882, w_043_1883, w_043_1884, w_043_1888, w_043_1890, w_043_1891, w_043_1892, w_043_1893, w_043_1895, w_043_1896, w_043_1897, w_043_1899, w_043_1900, w_043_1902, w_043_1903, w_043_1904, w_043_1905, w_043_1906, w_043_1907, w_043_1908, w_043_1909, w_043_1910, w_043_1911, w_043_1912, w_043_1913, w_043_1914, w_043_1915, w_043_1916, w_043_1917, w_043_1918, w_043_1919, w_043_1920, w_043_1922, w_043_1923, w_043_1924, w_043_1925, w_043_1928, w_043_1929, w_043_1930, w_043_1931, w_043_1935, w_043_1936, w_043_1938, w_043_1939, w_043_1940, w_043_1942, w_043_1943, w_043_1944, w_043_1945, w_043_1946, w_043_1949, w_043_1950, w_043_1951, w_043_1952, w_043_1953, w_043_1954, w_043_1956, w_043_1957, w_043_1959, w_043_1960, w_043_1962, w_043_1964, w_043_1965, w_043_1966, w_043_1968, w_043_1969, w_043_1970, w_043_1971, w_043_1972, w_043_1973, w_043_1974, w_043_1975, w_043_1976, w_043_1981, w_043_1982, w_043_1983, w_043_1984, w_043_1985, w_043_1986, w_043_1987, w_043_1989, w_043_1990, w_043_1991, w_043_1992, w_043_1994, w_043_1995, w_043_1996, w_043_1997, w_043_1998, w_043_1999, w_043_2000, w_043_2001, w_043_2002, w_043_2004, w_043_2005, w_043_2006, w_043_2007, w_043_2008, w_043_2009, w_043_2010, w_043_2011, w_043_2013, w_043_2014, w_043_2015, w_043_2017, w_043_2018, w_043_2019, w_043_2020, w_043_2021, w_043_2022, w_043_2023, w_043_2024, w_043_2025, w_043_2027, w_043_2028, w_043_2030, w_043_2031, w_043_2032, w_043_2033, w_043_2034, w_043_2036, w_043_2037, w_043_2040, w_043_2041, w_043_2042, w_043_2043, w_043_2044, w_043_2045, w_043_2046, w_043_2048, w_043_2049, w_043_2050, w_043_2052, w_043_2054, w_043_2055, w_043_2056, w_043_2057, w_043_2058, w_043_2059, w_043_2060, w_043_2061, w_043_2062, w_043_2063, w_043_2064, w_043_2065, w_043_2066, w_043_2068, w_043_2069, w_043_2070, w_043_2071, w_043_2074, w_043_2075, w_043_2076, w_043_2077, w_043_2078, w_043_2079, w_043_2080, w_043_2082, w_043_2083, w_043_2084, w_043_2085, w_043_2087, w_043_2089, w_043_2091, w_043_2092, w_043_2093, w_043_2094, w_043_2095, w_043_2096, w_043_2097, w_043_2098, w_043_2102, w_043_2103, w_043_2104, w_043_2106, w_043_2107, w_043_2109, w_043_2110, w_043_2111, w_043_2112, w_043_2115, w_043_2116, w_043_2119, w_043_2120, w_043_2122, w_043_2123, w_043_2125, w_043_2127, w_043_2129, w_043_2133, w_043_2135, w_043_2136, w_043_2141, w_043_2142, w_043_2143, w_043_2144, w_043_2146, w_043_2149, w_043_2151, w_043_2152, w_043_2153, w_043_2154, w_043_2156, w_043_2157, w_043_2159, w_043_2161, w_043_2162, w_043_2164, w_043_2165, w_043_2170, w_043_2171, w_043_2175, w_043_2176, w_043_2177, w_043_2178, w_043_2179, w_043_2180, w_043_2182, w_043_2183, w_043_2186, w_043_2187, w_043_2190, w_043_2191, w_043_2192, w_043_2193, w_043_2194, w_043_2196, w_043_2197, w_043_2199, w_043_2202, w_043_2205, w_043_2208, w_043_2211, w_043_2212, w_043_2213, w_043_2214, w_043_2216, w_043_2218, w_043_2219, w_043_2220, w_043_2221, w_043_2222, w_043_2224, w_043_2230, w_043_2231, w_043_2232, w_043_2234, w_043_2235, w_043_2236, w_043_2237, w_043_2238, w_043_2240, w_043_2244, w_043_2248, w_043_2250, w_043_2251, w_043_2252, w_043_2254, w_043_2255, w_043_2256, w_043_2257, w_043_2261, w_043_2262, w_043_2264, w_043_2270, w_043_2271, w_043_2272, w_043_2274, w_043_2275, w_043_2277, w_043_2280, w_043_2281, w_043_2282, w_043_2286, w_043_2287, w_043_2293, w_043_2295, w_043_2298, w_043_2300, w_043_2303, w_043_2304, w_043_2306, w_043_2307, w_043_2308, w_043_2309, w_043_2311, w_043_2312, w_043_2313, w_043_2314, w_043_2315, w_043_2316, w_043_2317, w_043_2319, w_043_2322, w_043_2323, w_043_2324, w_043_2325, w_043_2326, w_043_2327, w_043_2333, w_043_2334, w_043_2335, w_043_2336, w_043_2337, w_043_2338, w_043_2340, w_043_2341, w_043_2342, w_043_2343, w_043_2345, w_043_2347, w_043_2348, w_043_2350, w_043_2354, w_043_2355, w_043_2356, w_043_2359, w_043_2360, w_043_2361, w_043_2363, w_043_2364, w_043_2365, w_043_2366, w_043_2367, w_043_2368, w_043_2371, w_043_2374, w_043_2377, w_043_2379, w_043_2380, w_043_2381, w_043_2382, w_043_2383, w_043_2384, w_043_2385, w_043_2386, w_043_2387, w_043_2390, w_043_2391, w_043_2392, w_043_2393, w_043_2394, w_043_2395, w_043_2396, w_043_2398, w_043_2401, w_043_2402, w_043_2403, w_043_2404, w_043_2405, w_043_2407, w_043_2410, w_043_2412, w_043_2414, w_043_2415, w_043_2417, w_043_2419, w_043_2421, w_043_2422, w_043_2423, w_043_2424, w_043_2426, w_043_2428, w_043_2429, w_043_2430, w_043_2431, w_043_2432, w_043_2437, w_043_2443, w_043_2447, w_043_2448, w_043_2450, w_043_2452, w_043_2453, w_043_2458, w_043_2459, w_043_2460, w_043_2464, w_043_2465, w_043_2466, w_043_2468, w_043_2469, w_043_2470, w_043_2473, w_043_2474, w_043_2475, w_043_2476, w_043_2479, w_043_2480, w_043_2482, w_043_2483, w_043_2484, w_043_2487, w_043_2489, w_043_2490, w_043_2491, w_043_2493, w_043_2495, w_043_2496, w_043_2497, w_043_2498, w_043_2499, w_043_2501, w_043_2503, w_043_2507, w_043_2508, w_043_2509, w_043_2510, w_043_2511, w_043_2512, w_043_2513, w_043_2516, w_043_2520, w_043_2525, w_043_2526, w_043_2527, w_043_2528, w_043_2529, w_043_2530, w_043_2531, w_043_2533, w_043_2534, w_043_2535, w_043_2536, w_043_2539, w_043_2544, w_043_2545, w_043_2547, w_043_2551, w_043_2552, w_043_2555, w_043_2556, w_043_2558, w_043_2559, w_043_2560, w_043_2561, w_043_2563, w_043_2565, w_043_2566, w_043_2567, w_043_2569, w_043_2570, w_043_2571, w_043_2572, w_043_2573, w_043_2576, w_043_2578, w_043_2579, w_043_2580, w_043_2581, w_043_2582, w_043_2583, w_043_2585, w_043_2587, w_043_2588, w_043_2589, w_043_2590, w_043_2593, w_043_2594, w_043_2598, w_043_2599, w_043_2600, w_043_2601, w_043_2602, w_043_2604, w_043_2609, w_043_2610, w_043_2611, w_043_2613, w_043_2615, w_043_2617, w_043_2618, w_043_2623, w_043_2624, w_043_2625, w_043_2627, w_043_2629, w_043_2630, w_043_2632, w_043_2635, w_043_2636, w_043_2638, w_043_2639, w_043_2641, w_043_2644, w_043_2645, w_043_2647, w_043_2648, w_043_2649, w_043_2651, w_043_2652, w_043_2653, w_043_2654, w_043_2656, w_043_2657, w_043_2658, w_043_2666, w_043_2667, w_043_2668, w_043_2670, w_043_2674, w_043_2676, w_043_2680, w_043_2684, w_043_2687, w_043_2688, w_043_2689, w_043_2691, w_043_2692, w_043_2695, w_043_2696, w_043_2698, w_043_2702, w_043_2705, w_043_2707, w_043_2711, w_043_2712, w_043_2714, w_043_2717, w_043_2718, w_043_2719, w_043_2720, w_043_2721, w_043_2722, w_043_2723, w_043_2725, w_043_2727, w_043_2728, w_043_2730, w_043_2735, w_043_2736, w_043_2737, w_043_2740, w_043_2741, w_043_2742, w_043_2743, w_043_2745, w_043_2747, w_043_2750, w_043_2752, w_043_2755, w_043_2756, w_043_2759, w_043_2760, w_043_2762, w_043_2763, w_043_2764, w_043_2766, w_043_2767, w_043_2770, w_043_2774, w_043_2776, w_043_2777, w_043_2778, w_043_2781, w_043_2785, w_043_2786, w_043_2788, w_043_2789, w_043_2790, w_043_2791, w_043_2794, w_043_2795, w_043_2796, w_043_2797, w_043_2798, w_043_2802, w_043_2803, w_043_2804, w_043_2806, w_043_2808, w_043_2809, w_043_2812, w_043_2813, w_043_2815, w_043_2816, w_043_2817, w_043_2820, w_043_2821, w_043_2823, w_043_2825, w_043_2826, w_043_2827, w_043_2828, w_043_2829, w_043_2830, w_043_2833, w_043_2835, w_043_2836, w_043_2837, w_043_2841, w_043_2842, w_043_2843, w_043_2844, w_043_2845, w_043_2849, w_043_2850, w_043_2852, w_043_2854, w_043_2855, w_043_2857, w_043_2860, w_043_2861, w_043_2862, w_043_2864, w_043_2865, w_043_2869, w_043_2873, w_043_2876, w_043_2879, w_043_2880, w_043_2881, w_043_2882;
  wire w_044_002, w_044_003, w_044_004, w_044_005, w_044_006, w_044_008, w_044_009, w_044_011, w_044_012, w_044_013, w_044_014, w_044_017, w_044_018, w_044_019, w_044_020, w_044_021, w_044_022, w_044_023, w_044_026, w_044_027, w_044_028, w_044_029, w_044_030, w_044_031, w_044_032, w_044_033, w_044_034, w_044_037, w_044_038, w_044_039, w_044_040, w_044_043, w_044_044, w_044_045, w_044_046, w_044_047, w_044_048, w_044_049, w_044_050, w_044_051, w_044_052, w_044_053, w_044_054, w_044_055, w_044_056, w_044_057, w_044_058, w_044_059, w_044_060, w_044_061, w_044_062, w_044_063, w_044_064, w_044_065, w_044_066, w_044_067, w_044_068, w_044_070, w_044_073, w_044_074, w_044_076, w_044_078, w_044_079, w_044_082, w_044_083, w_044_084, w_044_085, w_044_086, w_044_088, w_044_090, w_044_091, w_044_092, w_044_093, w_044_094, w_044_095, w_044_098, w_044_104, w_044_105, w_044_106, w_044_107, w_044_108, w_044_109, w_044_110, w_044_111, w_044_112, w_044_113, w_044_116, w_044_120, w_044_121, w_044_123, w_044_124, w_044_126, w_044_128, w_044_131, w_044_132, w_044_136, w_044_140, w_044_141, w_044_142, w_044_143, w_044_144, w_044_145, w_044_147, w_044_148, w_044_151, w_044_154, w_044_157, w_044_158, w_044_159, w_044_160, w_044_161, w_044_162, w_044_163, w_044_167, w_044_168, w_044_171, w_044_172, w_044_174, w_044_175, w_044_176, w_044_183, w_044_184, w_044_185, w_044_187, w_044_190, w_044_191, w_044_193, w_044_196, w_044_199, w_044_202, w_044_203, w_044_206, w_044_208, w_044_209, w_044_213, w_044_215, w_044_216, w_044_217, w_044_223, w_044_224, w_044_225, w_044_226, w_044_228, w_044_230, w_044_231, w_044_234, w_044_235, w_044_237, w_044_241, w_044_244, w_044_245, w_044_249, w_044_251, w_044_252, w_044_253, w_044_255, w_044_257, w_044_259, w_044_260, w_044_261, w_044_263, w_044_264, w_044_265, w_044_267, w_044_270, w_044_271, w_044_272, w_044_273, w_044_274, w_044_275, w_044_277, w_044_282, w_044_284, w_044_287, w_044_288, w_044_289, w_044_293, w_044_297, w_044_298, w_044_300, w_044_305, w_044_307, w_044_310, w_044_313, w_044_314, w_044_315, w_044_316, w_044_318, w_044_320, w_044_326, w_044_329, w_044_331, w_044_333, w_044_334, w_044_335, w_044_338, w_044_340, w_044_342, w_044_343, w_044_344, w_044_346, w_044_349, w_044_350, w_044_353, w_044_354, w_044_357, w_044_362, w_044_364, w_044_367, w_044_370, w_044_377, w_044_378, w_044_379, w_044_381, w_044_382, w_044_383, w_044_384, w_044_385, w_044_389, w_044_391, w_044_393, w_044_394, w_044_397, w_044_403, w_044_405, w_044_406, w_044_408, w_044_410, w_044_412, w_044_413, w_044_414, w_044_416, w_044_417, w_044_420, w_044_421, w_044_422, w_044_429, w_044_431, w_044_432, w_044_439, w_044_441, w_044_443, w_044_444, w_044_445, w_044_446, w_044_449, w_044_451, w_044_456, w_044_458, w_044_459, w_044_461, w_044_463, w_044_468, w_044_471, w_044_472, w_044_475, w_044_478, w_044_482, w_044_487, w_044_490, w_044_493, w_044_495, w_044_496, w_044_499, w_044_502, w_044_504, w_044_506, w_044_508, w_044_509, w_044_511, w_044_512, w_044_516, w_044_517, w_044_520, w_044_523, w_044_525, w_044_528, w_044_529, w_044_532, w_044_533, w_044_536, w_044_537, w_044_538, w_044_540, w_044_541, w_044_543, w_044_544, w_044_548, w_044_549, w_044_551, w_044_552, w_044_553, w_044_554, w_044_555, w_044_557, w_044_561, w_044_564, w_044_570, w_044_575, w_044_580, w_044_584, w_044_587, w_044_588, w_044_590, w_044_593, w_044_594, w_044_606, w_044_607, w_044_609, w_044_614, w_044_615, w_044_620, w_044_624, w_044_625, w_044_626, w_044_635, w_044_636, w_044_637, w_044_641, w_044_643, w_044_645, w_044_646, w_044_647, w_044_648, w_044_652, w_044_654, w_044_656, w_044_657, w_044_659, w_044_660, w_044_661, w_044_662, w_044_663, w_044_666, w_044_667, w_044_668, w_044_669, w_044_673, w_044_675, w_044_677, w_044_680, w_044_681, w_044_682, w_044_683, w_044_684, w_044_687, w_044_688, w_044_690, w_044_691, w_044_693, w_044_695, w_044_697, w_044_698, w_044_699, w_044_702, w_044_704, w_044_705, w_044_706, w_044_707, w_044_708, w_044_709, w_044_711, w_044_712, w_044_713, w_044_714, w_044_715, w_044_717, w_044_718, w_044_719, w_044_722, w_044_724, w_044_726, w_044_727, w_044_728, w_044_729, w_044_733, w_044_734, w_044_736, w_044_737, w_044_738, w_044_740, w_044_743, w_044_745, w_044_746, w_044_748, w_044_749, w_044_752, w_044_753, w_044_754, w_044_756, w_044_758, w_044_760, w_044_761, w_044_764, w_044_768, w_044_769, w_044_772, w_044_774, w_044_775, w_044_777, w_044_779, w_044_780, w_044_781, w_044_783, w_044_785, w_044_786, w_044_787, w_044_788, w_044_790, w_044_797, w_044_800, w_044_802, w_044_804, w_044_805, w_044_807, w_044_808, w_044_811, w_044_812, w_044_815, w_044_816, w_044_817, w_044_818, w_044_819, w_044_820, w_044_822, w_044_824, w_044_826, w_044_833, w_044_834, w_044_835, w_044_837, w_044_840, w_044_841, w_044_845, w_044_846, w_044_851, w_044_853, w_044_854, w_044_855, w_044_862, w_044_863, w_044_866, w_044_867, w_044_868, w_044_870, w_044_874, w_044_875, w_044_878, w_044_879, w_044_880, w_044_883, w_044_885, w_044_887, w_044_888, w_044_889, w_044_894, w_044_898, w_044_900, w_044_903, w_044_905, w_044_906, w_044_907, w_044_908, w_044_909, w_044_910, w_044_920, w_044_921, w_044_924, w_044_928, w_044_931, w_044_932, w_044_933, w_044_935, w_044_936, w_044_938, w_044_939, w_044_940, w_044_941, w_044_942, w_044_943, w_044_944, w_044_945, w_044_946, w_044_948, w_044_953, w_044_957, w_044_958, w_044_960, w_044_963, w_044_964, w_044_965, w_044_968, w_044_970, w_044_972, w_044_973, w_044_976, w_044_978, w_044_979, w_044_980, w_044_981, w_044_982, w_044_984, w_044_985, w_044_986, w_044_988, w_044_990, w_044_991, w_044_992, w_044_993, w_044_996, w_044_997, w_044_999, w_044_1000, w_044_1001, w_044_1002, w_044_1006, w_044_1008, w_044_1010, w_044_1011, w_044_1012, w_044_1014, w_044_1017, w_044_1018, w_044_1019, w_044_1022, w_044_1024, w_044_1027, w_044_1028, w_044_1032, w_044_1034, w_044_1036, w_044_1037, w_044_1039, w_044_1040, w_044_1041, w_044_1049, w_044_1053, w_044_1055, w_044_1056, w_044_1057, w_044_1058, w_044_1060, w_044_1061, w_044_1062, w_044_1063, w_044_1064, w_044_1065, w_044_1069, w_044_1070, w_044_1073, w_044_1074, w_044_1075, w_044_1076, w_044_1077, w_044_1078, w_044_1082, w_044_1084, w_044_1088, w_044_1089, w_044_1091, w_044_1092, w_044_1096, w_044_1097, w_044_1099, w_044_1104, w_044_1105, w_044_1106, w_044_1108, w_044_1110, w_044_1112, w_044_1116, w_044_1118, w_044_1119, w_044_1120, w_044_1124, w_044_1126, w_044_1129, w_044_1131, w_044_1132, w_044_1133, w_044_1134, w_044_1135, w_044_1136, w_044_1138, w_044_1139, w_044_1140, w_044_1142, w_044_1144, w_044_1145, w_044_1146, w_044_1149, w_044_1151, w_044_1152, w_044_1157, w_044_1160, w_044_1161, w_044_1162, w_044_1164, w_044_1167, w_044_1171, w_044_1172, w_044_1175, w_044_1176, w_044_1180, w_044_1183, w_044_1186, w_044_1187, w_044_1188, w_044_1191, w_044_1192, w_044_1195, w_044_1196, w_044_1197, w_044_1198, w_044_1199, w_044_1200, w_044_1203, w_044_1205, w_044_1206, w_044_1208, w_044_1209, w_044_1212, w_044_1213, w_044_1215, w_044_1216, w_044_1217, w_044_1221, w_044_1223, w_044_1225, w_044_1226, w_044_1227, w_044_1228, w_044_1229, w_044_1230, w_044_1233, w_044_1234, w_044_1236, w_044_1237, w_044_1241, w_044_1242, w_044_1244, w_044_1245, w_044_1246, w_044_1247, w_044_1252, w_044_1254, w_044_1258, w_044_1263, w_044_1267, w_044_1269, w_044_1273, w_044_1275, w_044_1282, w_044_1283, w_044_1284, w_044_1288, w_044_1290, w_044_1293, w_044_1295, w_044_1296, w_044_1297, w_044_1298, w_044_1299, w_044_1305, w_044_1307, w_044_1309, w_044_1310, w_044_1312, w_044_1316, w_044_1318, w_044_1321, w_044_1322, w_044_1324, w_044_1325, w_044_1329, w_044_1332, w_044_1333, w_044_1341, w_044_1342, w_044_1343, w_044_1344, w_044_1345, w_044_1347, w_044_1349, w_044_1350, w_044_1351, w_044_1352, w_044_1353, w_044_1354, w_044_1357, w_044_1363, w_044_1364, w_044_1365, w_044_1366, w_044_1367, w_044_1368, w_044_1369, w_044_1371, w_044_1373, w_044_1374, w_044_1377, w_044_1378, w_044_1380, w_044_1386, w_044_1387, w_044_1394, w_044_1396, w_044_1397, w_044_1399, w_044_1402, w_044_1407, w_044_1409, w_044_1410, w_044_1412, w_044_1413, w_044_1414, w_044_1416, w_044_1417, w_044_1419, w_044_1420, w_044_1422, w_044_1423, w_044_1424, w_044_1425, w_044_1426, w_044_1430, w_044_1432, w_044_1436, w_044_1437, w_044_1439, w_044_1440, w_044_1441, w_044_1442, w_044_1444, w_044_1445, w_044_1447, w_044_1448, w_044_1450, w_044_1452, w_044_1453, w_044_1455, w_044_1456, w_044_1457, w_044_1458, w_044_1461, w_044_1466, w_044_1467, w_044_1468, w_044_1469, w_044_1471, w_044_1472, w_044_1473, w_044_1474, w_044_1475, w_044_1477, w_044_1481, w_044_1483, w_044_1485, w_044_1486, w_044_1487, w_044_1488, w_044_1491, w_044_1492, w_044_1493, w_044_1495, w_044_1497, w_044_1500, w_044_1504, w_044_1508, w_044_1511, w_044_1512, w_044_1513, w_044_1515, w_044_1516, w_044_1517, w_044_1518, w_044_1523, w_044_1525, w_044_1527, w_044_1528, w_044_1531, w_044_1532, w_044_1534, w_044_1537, w_044_1538, w_044_1540, w_044_1544, w_044_1545, w_044_1546, w_044_1547, w_044_1549, w_044_1550, w_044_1553, w_044_1559, w_044_1566, w_044_1572, w_044_1573, w_044_1574, w_044_1580, w_044_1583, w_044_1584, w_044_1587, w_044_1589, w_044_1591, w_044_1592, w_044_1593, w_044_1594, w_044_1596, w_044_1597, w_044_1598, w_044_1604, w_044_1606, w_044_1608, w_044_1617, w_044_1618, w_044_1619, w_044_1620, w_044_1625, w_044_1627, w_044_1629, w_044_1631, w_044_1632, w_044_1633, w_044_1636, w_044_1637, w_044_1643, w_044_1644, w_044_1645, w_044_1646, w_044_1647, w_044_1648, w_044_1650, w_044_1653, w_044_1655, w_044_1662, w_044_1664, w_044_1665, w_044_1666, w_044_1667, w_044_1668, w_044_1670, w_044_1671, w_044_1672, w_044_1673, w_044_1675, w_044_1677, w_044_1678, w_044_1679, w_044_1681, w_044_1684, w_044_1685, w_044_1688, w_044_1694, w_044_1699, w_044_1701, w_044_1703, w_044_1705, w_044_1710, w_044_1713, w_044_1715, w_044_1716, w_044_1719, w_044_1720, w_044_1721, w_044_1722, w_044_1724, w_044_1728, w_044_1729, w_044_1731, w_044_1734, w_044_1738, w_044_1740, w_044_1741, w_044_1742, w_044_1743, w_044_1745, w_044_1746, w_044_1748, w_044_1749, w_044_1750, w_044_1751, w_044_1752, w_044_1754, w_044_1755, w_044_1757, w_044_1762, w_044_1763, w_044_1767, w_044_1769, w_044_1770, w_044_1774, w_044_1775, w_044_1777, w_044_1778, w_044_1779, w_044_1780, w_044_1782, w_044_1783, w_044_1784, w_044_1786, w_044_1787, w_044_1789, w_044_1791, w_044_1792, w_044_1793, w_044_1794, w_044_1795, w_044_1796, w_044_1797, w_044_1798, w_044_1802, w_044_1804, w_044_1808, w_044_1809, w_044_1812, w_044_1816, w_044_1818, w_044_1819, w_044_1821, w_044_1822, w_044_1823, w_044_1824, w_044_1825, w_044_1826, w_044_1833, w_044_1834, w_044_1835, w_044_1838, w_044_1839, w_044_1840, w_044_1841, w_044_1842, w_044_1843, w_044_1844, w_044_1847, w_044_1848, w_044_1850, w_044_1851, w_044_1854, w_044_1855, w_044_1857, w_044_1858, w_044_1862, w_044_1863, w_044_1866, w_044_1869, w_044_1870, w_044_1871, w_044_1872, w_044_1873, w_044_1875, w_044_1876, w_044_1877, w_044_1878, w_044_1879, w_044_1883, w_044_1884, w_044_1887, w_044_1891, w_044_1892, w_044_1894, w_044_1895, w_044_1896, w_044_1897, w_044_1900, w_044_1903, w_044_1905, w_044_1906, w_044_1907, w_044_1910, w_044_1911, w_044_1913, w_044_1915, w_044_1917, w_044_1919, w_044_1923, w_044_1924, w_044_1926, w_044_1927, w_044_1928, w_044_1930, w_044_1933, w_044_1936, w_044_1940, w_044_1941, w_044_1944, w_044_1947, w_044_1949, w_044_1950, w_044_1953, w_044_1954, w_044_1956, w_044_1958, w_044_1961, w_044_1962, w_044_1963, w_044_1965, w_044_1966, w_044_1968, w_044_1969, w_044_1970, w_044_1971, w_044_1972, w_044_1973, w_044_1974, w_044_1975, w_044_1976, w_044_1980, w_044_1983, w_044_1985, w_044_1987, w_044_1989, w_044_1991, w_044_1992, w_044_1994, w_044_1995, w_044_1999, w_044_2001, w_044_2002, w_044_2003, w_044_2006, w_044_2008, w_044_2009, w_044_2011, w_044_2013, w_044_2014, w_044_2018, w_044_2019, w_044_2020, w_044_2023, w_044_2024, w_044_2026, w_044_2027, w_044_2035, w_044_2036, w_044_2037, w_044_2038, w_044_2040, w_044_2041, w_044_2042, w_044_2043, w_044_2044, w_044_2047, w_044_2049, w_044_2050, w_044_2051, w_044_2055, w_044_2056, w_044_2057, w_044_2060, w_044_2063, w_044_2064, w_044_2066, w_044_2067, w_044_2068, w_044_2070, w_044_2071, w_044_2073, w_044_2074, w_044_2075, w_044_2076, w_044_2080, w_044_2081, w_044_2083, w_044_2085, w_044_2086, w_044_2087, w_044_2090, w_044_2093, w_044_2094, w_044_2096, w_044_2098, w_044_2101, w_044_2104, w_044_2105, w_044_2107, w_044_2108, w_044_2113, w_044_2115, w_044_2116, w_044_2117, w_044_2118, w_044_2119, w_044_2124, w_044_2125, w_044_2126, w_044_2127, w_044_2129, w_044_2130, w_044_2131, w_044_2132, w_044_2133, w_044_2134, w_044_2136, w_044_2138, w_044_2140, w_044_2141, w_044_2144, w_044_2145, w_044_2150, w_044_2153, w_044_2154, w_044_2157, w_044_2158, w_044_2159, w_044_2162, w_044_2163, w_044_2165, w_044_2166, w_044_2167, w_044_2169, w_044_2173, w_044_2175, w_044_2176, w_044_2177, w_044_2178, w_044_2179, w_044_2180, w_044_2181, w_044_2182, w_044_2183, w_044_2186, w_044_2188, w_044_2189, w_044_2190, w_044_2191, w_044_2193, w_044_2195, w_044_2196, w_044_2197, w_044_2198, w_044_2199, w_044_2200, w_044_2201, w_044_2203, w_044_2207, w_044_2208, w_044_2212, w_044_2213, w_044_2214, w_044_2216, w_044_2217, w_044_2218, w_044_2219, w_044_2220, w_044_2221, w_044_2222, w_044_2223, w_044_2226, w_044_2232, w_044_2233, w_044_2235, w_044_2237, w_044_2239, w_044_2245, w_044_2246, w_044_2248, w_044_2250, w_044_2251, w_044_2256, w_044_2257, w_044_2260, w_044_2261, w_044_2262, w_044_2264, w_044_2268, w_044_2270, w_044_2272, w_044_2274, w_044_2275, w_044_2276, w_044_2278, w_044_2285, w_044_2287, w_044_2291, w_044_2292, w_044_2294, w_044_2297, w_044_2298, w_044_2299, w_044_2304, w_044_2305, w_044_2306, w_044_2308, w_044_2309, w_044_2310, w_044_2311, w_044_2312, w_044_2314, w_044_2316, w_044_2318, w_044_2320, w_044_2321, w_044_2322, w_044_2324, w_044_2325, w_044_2326, w_044_2329, w_044_2330, w_044_2332, w_044_2334, w_044_2335, w_044_2337, w_044_2340, w_044_2342, w_044_2343, w_044_2348, w_044_2349, w_044_2350, w_044_2351, w_044_2352, w_044_2353, w_044_2355, w_044_2356, w_044_2358, w_044_2359, w_044_2360, w_044_2363, w_044_2365, w_044_2367, w_044_2368, w_044_2371, w_044_2372, w_044_2378, w_044_2379, w_044_2380, w_044_2381, w_044_2384, w_044_2386, w_044_2387, w_044_2388, w_044_2390, w_044_2391, w_044_2392, w_044_2394, w_044_2397, w_044_2399, w_044_2400, w_044_2402, w_044_2403, w_044_2406, w_044_2407, w_044_2408, w_044_2409, w_044_2411, w_044_2412, w_044_2413, w_044_2414, w_044_2415, w_044_2416, w_044_2417, w_044_2418, w_044_2419, w_044_2420, w_044_2421, w_044_2423, w_044_2424, w_044_2425, w_044_2428, w_044_2433, w_044_2434, w_044_2437, w_044_2441, w_044_2442, w_044_2443, w_044_2445, w_044_2446, w_044_2450, w_044_2451, w_044_2457, w_044_2459, w_044_2461, w_044_2464, w_044_2467, w_044_2469, w_044_2470, w_044_2471, w_044_2472, w_044_2473, w_044_2474, w_044_2475, w_044_2481, w_044_2482, w_044_2484, w_044_2485, w_044_2487, w_044_2488, w_044_2490, w_044_2491, w_044_2493, w_044_2496, w_044_2497, w_044_2498, w_044_2499, w_044_2501, w_044_2502, w_044_2506, w_044_2508, w_044_2509, w_044_2513, w_044_2515, w_044_2516, w_044_2522, w_044_2523, w_044_2528, w_044_2530, w_044_2533, w_044_2535, w_044_2537, w_044_2540, w_044_2542, w_044_2543, w_044_2547, w_044_2549, w_044_2550, w_044_2552, w_044_2554, w_044_2555, w_044_2558, w_044_2560, w_044_2561, w_044_2564, w_044_2565, w_044_2566, w_044_2567, w_044_2568, w_044_2569, w_044_2571, w_044_2572, w_044_2573, w_044_2574, w_044_2576, w_044_2577, w_044_2580, w_044_2581, w_044_2582, w_044_2583, w_044_2584, w_044_2585, w_044_2586, w_044_2590, w_044_2595, w_044_2597, w_044_2599, w_044_2602, w_044_2604, w_044_2606, w_044_2607, w_044_2608, w_044_2609, w_044_2610, w_044_2615, w_044_2617, w_044_2618, w_044_2619, w_044_2620, w_044_2622, w_044_2623, w_044_2624, w_044_2627, w_044_2628, w_044_2632, w_044_2633, w_044_2635, w_044_2636, w_044_2638, w_044_2639, w_044_2641, w_044_2644, w_044_2647, w_044_2652, w_044_2654, w_044_2657, w_044_2659, w_044_2660, w_044_2662, w_044_2664, w_044_2668, w_044_2669, w_044_2670, w_044_2671, w_044_2672, w_044_2674, w_044_2677, w_044_2681, w_044_2682, w_044_2683, w_044_2684, w_044_2686, w_044_2687, w_044_2688, w_044_2695, w_044_2697, w_044_2698, w_044_2702, w_044_2705, w_044_2707, w_044_2708, w_044_2711, w_044_2712, w_044_2714, w_044_2716, w_044_2719, w_044_2720, w_044_2722, w_044_2724, w_044_2725, w_044_2726, w_044_2730, w_044_2731, w_044_2732, w_044_2733, w_044_2734, w_044_2735, w_044_2736, w_044_2737, w_044_2739, w_044_2742, w_044_2746, w_044_2751, w_044_2753, w_044_2756, w_044_2757, w_044_2759, w_044_2760, w_044_2762, w_044_2763, w_044_2765, w_044_2768, w_044_2769, w_044_2772, w_044_2773, w_044_2774, w_044_2775, w_044_2776, w_044_2793, w_044_2796, w_044_2797, w_044_2800, w_044_2802, w_044_2803, w_044_2805, w_044_2806, w_044_2807, w_044_2808, w_044_2809, w_044_2813, w_044_2814, w_044_2815, w_044_2816, w_044_2820, w_044_2823, w_044_2824, w_044_2825, w_044_2826, w_044_2827, w_044_2829, w_044_2832, w_044_2833, w_044_2835, w_044_2836, w_044_2843, w_044_2844, w_044_2846, w_044_2848, w_044_2851, w_044_2852, w_044_2854, w_044_2855, w_044_2856, w_044_2858, w_044_2860, w_044_2861, w_044_2862, w_044_2863, w_044_2864, w_044_2865, w_044_2866, w_044_2872, w_044_2875, w_044_2876, w_044_2878, w_044_2885, w_044_2886, w_044_2889, w_044_2894, w_044_2895, w_044_2899, w_044_2902, w_044_2904, w_044_2906, w_044_2907, w_044_2908, w_044_2911, w_044_2913, w_044_2915, w_044_2916, w_044_2918, w_044_2920, w_044_2923, w_044_2924, w_044_2925, w_044_2927, w_044_2930, w_044_2931, w_044_2932, w_044_2934, w_044_2939, w_044_2940, w_044_2944, w_044_2945, w_044_2946, w_044_2948, w_044_2950, w_044_2954, w_044_2955, w_044_2956, w_044_2958, w_044_2959, w_044_2962, w_044_2964, w_044_2965, w_044_2968, w_044_2970, w_044_2971, w_044_2972, w_044_2975, w_044_2976, w_044_2978, w_044_2979, w_044_2981, w_044_2982, w_044_2983, w_044_2984, w_044_2985, w_044_2987, w_044_2988, w_044_2990, w_044_2992, w_044_2993, w_044_2994, w_044_2995, w_044_2996, w_044_2999, w_044_3000, w_044_3001, w_044_3005, w_044_3006, w_044_3007, w_044_3008, w_044_3010, w_044_3012, w_044_3013, w_044_3014, w_044_3015, w_044_3017, w_044_3019, w_044_3020, w_044_3021, w_044_3024, w_044_3029, w_044_3035, w_044_3036, w_044_3038, w_044_3039, w_044_3040, w_044_3042, w_044_3045, w_044_3047, w_044_3048, w_044_3049, w_044_3050, w_044_3055, w_044_3056, w_044_3057, w_044_3058, w_044_3063, w_044_3065, w_044_3068, w_044_3069, w_044_3070, w_044_3071, w_044_3072, w_044_3073, w_044_3074, w_044_3075, w_044_3077, w_044_3078, w_044_3080, w_044_3081, w_044_3084, w_044_3086, w_044_3089, w_044_3093, w_044_3095, w_044_3098, w_044_3102, w_044_3104, w_044_3105, w_044_3108, w_044_3109, w_044_3111, w_044_3118, w_044_3119, w_044_3123, w_044_3126, w_044_3133, w_044_3134, w_044_3135, w_044_3136, w_044_3137, w_044_3143, w_044_3144, w_044_3145, w_044_3146, w_044_3147, w_044_3148, w_044_3149, w_044_3150, w_044_3151, w_044_3153, w_044_3154, w_044_3155, w_044_3157, w_044_3158, w_044_3159, w_044_3162, w_044_3163, w_044_3164, w_044_3165, w_044_3166, w_044_3169, w_044_3171, w_044_3174, w_044_3176, w_044_3177, w_044_3179, w_044_3181, w_044_3182, w_044_3184, w_044_3186, w_044_3187, w_044_3188, w_044_3189, w_044_3190, w_044_3196, w_044_3201, w_044_3202, w_044_3206, w_044_3209, w_044_3210, w_044_3211, w_044_3212, w_044_3214, w_044_3216, w_044_3218, w_044_3219, w_044_3220, w_044_3223, w_044_3224, w_044_3228, w_044_3229, w_044_3230, w_044_3232, w_044_3234, w_044_3235, w_044_3236, w_044_3238, w_044_3242, w_044_3243, w_044_3244, w_044_3246, w_044_3247, w_044_3249, w_044_3251, w_044_3253, w_044_3255, w_044_3260, w_044_3264, w_044_3265, w_044_3267, w_044_3268, w_044_3271, w_044_3272, w_044_3273, w_044_3277, w_044_3279, w_044_3282, w_044_3283, w_044_3286, w_044_3288, w_044_3290, w_044_3293, w_044_3295, w_044_3296, w_044_3297, w_044_3302, w_044_3308, w_044_3309, w_044_3311, w_044_3312, w_044_3315, w_044_3320, w_044_3326, w_044_3327, w_044_3330, w_044_3331, w_044_3332, w_044_3333, w_044_3336, w_044_3337, w_044_3338, w_044_3339, w_044_3345, w_044_3346, w_044_3349, w_044_3350, w_044_3351, w_044_3352, w_044_3354, w_044_3355, w_044_3358, w_044_3359, w_044_3362, w_044_3363, w_044_3365, w_044_3366, w_044_3370, w_044_3371, w_044_3372, w_044_3373, w_044_3376, w_044_3377, w_044_3379, w_044_3380, w_044_3385, w_044_3387, w_044_3388, w_044_3393, w_044_3394, w_044_3397, w_044_3399, w_044_3402, w_044_3403, w_044_3406, w_044_3407, w_044_3408, w_044_3409, w_044_3410, w_044_3415, w_044_3417, w_044_3418, w_044_3419, w_044_3421, w_044_3422, w_044_3424, w_044_3428, w_044_3429, w_044_3430, w_044_3431, w_044_3433, w_044_3435, w_044_3437, w_044_3439, w_044_3440, w_044_3442, w_044_3444, w_044_3446, w_044_3447, w_044_3448, w_044_3453, w_044_3457, w_044_3458, w_044_3463, w_044_3464, w_044_3465, w_044_3466, w_044_3467, w_044_3469, w_044_3470, w_044_3471, w_044_3472, w_044_3473, w_044_3475, w_044_3476, w_044_3479, w_044_3480, w_044_3486, w_044_3487, w_044_3492, w_044_3494, w_044_3501, w_044_3502, w_044_3503, w_044_3504, w_044_3505, w_044_3506, w_044_3508, w_044_3509, w_044_3511, w_044_3513, w_044_3514, w_044_3515, w_044_3516, w_044_3517, w_044_3518, w_044_3525, w_044_3527, w_044_3528, w_044_3529, w_044_3530, w_044_3531, w_044_3532, w_044_3535, w_044_3538, w_044_3539, w_044_3540, w_044_3543, w_044_3545, w_044_3546, w_044_3548, w_044_3549, w_044_3550, w_044_3551, w_044_3553, w_044_3555, w_044_3556, w_044_3558, w_044_3560, w_044_3562, w_044_3565, w_044_3566, w_044_3570, w_044_3572, w_044_3574, w_044_3575, w_044_3579, w_044_3582, w_044_3584, w_044_3586, w_044_3587, w_044_3588, w_044_3592, w_044_3593, w_044_3594, w_044_3599, w_044_3600, w_044_3601, w_044_3605, w_044_3606, w_044_3607, w_044_3608, w_044_3609, w_044_3610, w_044_3616, w_044_3617, w_044_3618, w_044_3619, w_044_3621, w_044_3622, w_044_3623, w_044_3625, w_044_3634, w_044_3636, w_044_3637, w_044_3638, w_044_3640, w_044_3646, w_044_3649, w_044_3653, w_044_3655, w_044_3658, w_044_3660, w_044_3663, w_044_3664, w_044_3666, w_044_3668, w_044_3675, w_044_3676, w_044_3677, w_044_3679, w_044_3681, w_044_3682, w_044_3685, w_044_3688, w_044_3689, w_044_3690, w_044_3691, w_044_3694, w_044_3695, w_044_3696, w_044_3698, w_044_3700, w_044_3701, w_044_3703, w_044_3707, w_044_3708, w_044_3709, w_044_3713, w_044_3715, w_044_3716, w_044_3718, w_044_3721, w_044_3722, w_044_3723, w_044_3725, w_044_3726, w_044_3727, w_044_3729, w_044_3730, w_044_3731, w_044_3735, w_044_3736, w_044_3738, w_044_3739, w_044_3742, w_044_3743, w_044_3745, w_044_3748, w_044_3749, w_044_3755, w_044_3758, w_044_3759, w_044_3765, w_044_3766, w_044_3769, w_044_3771, w_044_3772, w_044_3773, w_044_3774, w_044_3775, w_044_3776, w_044_3780, w_044_3781, w_044_3785, w_044_3786, w_044_3788, w_044_3789, w_044_3790, w_044_3792, w_044_3793, w_044_3794, w_044_3795, w_044_3796, w_044_3798, w_044_3799, w_044_3800, w_044_3801, w_044_3804, w_044_3806, w_044_3807, w_044_3810, w_044_3813, w_044_3814, w_044_3815, w_044_3816, w_044_3817, w_044_3819, w_044_3822, w_044_3824, w_044_3827, w_044_3828, w_044_3832, w_044_3833, w_044_3834, w_044_3839, w_044_3840, w_044_3843, w_044_3844, w_044_3846, w_044_3850, w_044_3851, w_044_3855, w_044_3858, w_044_3861, w_044_3862, w_044_3864, w_044_3865, w_044_3866, w_044_3868, w_044_3869, w_044_3871, w_044_3873, w_044_3874, w_044_3876, w_044_3877, w_044_3879, w_044_3880, w_044_3881, w_044_3884, w_044_3886, w_044_3887, w_044_3888, w_044_3889, w_044_3891, w_044_3892, w_044_3894, w_044_3895, w_044_3897, w_044_3898, w_044_3900, w_044_3901, w_044_3902, w_044_3903, w_044_3904, w_044_3905, w_044_3906, w_044_3910, w_044_3911, w_044_3912, w_044_3913, w_044_3916, w_044_3920, w_044_3921, w_044_3925, w_044_3926, w_044_3927, w_044_3928, w_044_3930, w_044_3932, w_044_3933, w_044_3936, w_044_3937, w_044_3938, w_044_3939, w_044_3941, w_044_3942, w_044_3943, w_044_3945, w_044_3948, w_044_3949, w_044_3952, w_044_3954, w_044_3957, w_044_3959, w_044_3963, w_044_3964, w_044_3967, w_044_3968, w_044_3970, w_044_3977, w_044_3978, w_044_3979, w_044_3981, w_044_3985, w_044_3987, w_044_3990, w_044_3991, w_044_3992, w_044_3997, w_044_3998, w_044_3999, w_044_4001, w_044_4005, w_044_4006, w_044_4012, w_044_4013, w_044_4014, w_044_4015, w_044_4017, w_044_4018, w_044_4019, w_044_4020, w_044_4021, w_044_4026, w_044_4027, w_044_4028, w_044_4029, w_044_4033, w_044_4034, w_044_4035, w_044_4036, w_044_4039, w_044_4040, w_044_4045, w_044_4048, w_044_4049, w_044_4056, w_044_4057, w_044_4058, w_044_4059, w_044_4060, w_044_4061, w_044_4063, w_044_4067, w_044_4068, w_044_4069, w_044_4072, w_044_4075, w_044_4076, w_044_4079, w_044_4080, w_044_4082, w_044_4085, w_044_4087, w_044_4090, w_044_4092, w_044_4093, w_044_4095, w_044_4096, w_044_4098, w_044_4100, w_044_4102, w_044_4103, w_044_4104, w_044_4105, w_044_4107, w_044_4108, w_044_4110, w_044_4111, w_044_4112, w_044_4113, w_044_4114, w_044_4115, w_044_4117, w_044_4118, w_044_4120, w_044_4122, w_044_4124, w_044_4128, w_044_4129, w_044_4133, w_044_4134, w_044_4137, w_044_4142, w_044_4144, w_044_4145, w_044_4148, w_044_4150, w_044_4152, w_044_4153, w_044_4155, w_044_4157, w_044_4162, w_044_4163, w_044_4164, w_044_4165, w_044_4166, w_044_4168, w_044_4169, w_044_4170, w_044_4171, w_044_4172, w_044_4173, w_044_4174, w_044_4178, w_044_4182, w_044_4184, w_044_4185, w_044_4187, w_044_4188, w_044_4189, w_044_4190, w_044_4191, w_044_4192, w_044_4195, w_044_4196, w_044_4198, w_044_4199, w_044_4203, w_044_4204, w_044_4206, w_044_4207, w_044_4211, w_044_4213, w_044_4214, w_044_4216, w_044_4217, w_044_4218, w_044_4219, w_044_4221, w_044_4223, w_044_4225, w_044_4226, w_044_4229, w_044_4230, w_044_4232, w_044_4235, w_044_4237, w_044_4238, w_044_4243, w_044_4244, w_044_4247, w_044_4249, w_044_4250, w_044_4251, w_044_4253, w_044_4254, w_044_4255, w_044_4257, w_044_4261, w_044_4262, w_044_4268, w_044_4269, w_044_4272, w_044_4273, w_044_4276, w_044_4281, w_044_4282, w_044_4287, w_044_4288, w_044_4290, w_044_4291, w_044_4292, w_044_4294, w_044_4295, w_044_4297, w_044_4299, w_044_4301, w_044_4303, w_044_4304, w_044_4310, w_044_4311, w_044_4314, w_044_4315, w_044_4316, w_044_4317, w_044_4319, w_044_4320, w_044_4321, w_044_4322, w_044_4323, w_044_4328, w_044_4330, w_044_4333, w_044_4335, w_044_4337, w_044_4338, w_044_4339, w_044_4340, w_044_4341, w_044_4343, w_044_4344, w_044_4346, w_044_4349, w_044_4350, w_044_4351, w_044_4360, w_044_4361, w_044_4363, w_044_4364, w_044_4365, w_044_4367, w_044_4368, w_044_4369, w_044_4370, w_044_4371, w_044_4373, w_044_4374, w_044_4375, w_044_4376, w_044_4377, w_044_4380, w_044_4382, w_044_4384, w_044_4385, w_044_4390, w_044_4396, w_044_4397, w_044_4398, w_044_4401, w_044_4403, w_044_4407, w_044_4408, w_044_4410, w_044_4411, w_044_4414, w_044_4415, w_044_4417, w_044_4422, w_044_4423, w_044_4426, w_044_4427, w_044_4428, w_044_4430, w_044_4435, w_044_4437, w_044_4438, w_044_4440, w_044_4442, w_044_4443, w_044_4444, w_044_4445, w_044_4446, w_044_4448, w_044_4452, w_044_4453, w_044_4454, w_044_4456, w_044_4457, w_044_4458, w_044_4460, w_044_4467, w_044_4471, w_044_4472, w_044_4474, w_044_4476, w_044_4478, w_044_4479, w_044_4480, w_044_4486, w_044_4487, w_044_4490, w_044_4492, w_044_4494, w_044_4495, w_044_4496, w_044_4498, w_044_4501, w_044_4502, w_044_4503, w_044_4506, w_044_4509, w_044_4511, w_044_4512, w_044_4513, w_044_4515, w_044_4516, w_044_4517, w_044_4519, w_044_4520, w_044_4522, w_044_4524, w_044_4525, w_044_4526, w_044_4527, w_044_4529, w_044_4532, w_044_4533, w_044_4534, w_044_4535, w_044_4537, w_044_4538, w_044_4539, w_044_4540, w_044_4543, w_044_4547, w_044_4548, w_044_4549, w_044_4550, w_044_4554, w_044_4556, w_044_4559, w_044_4560, w_044_4561, w_044_4562, w_044_4570, w_044_4571, w_044_4572, w_044_4573, w_044_4574, w_044_4578, w_044_4584, w_044_4586, w_044_4588, w_044_4589, w_044_4590, w_044_4595, w_044_4598, w_044_4599, w_044_4600, w_044_4602, w_044_4607, w_044_4608, w_044_4609, w_044_4610, w_044_4613, w_044_4618, w_044_4619, w_044_4621, w_044_4622, w_044_4624, w_044_4628, w_044_4630, w_044_4631, w_044_4632, w_044_4634, w_044_4636, w_044_4637, w_044_4638, w_044_4639, w_044_4642, w_044_4643, w_044_4644, w_044_4645, w_044_4647, w_044_4648, w_044_4650, w_044_4652, w_044_4654, w_044_4662, w_044_4663, w_044_4665, w_044_4667, w_044_4670, w_044_4674, w_044_4675, w_044_4676, w_044_4679, w_044_4681, w_044_4683, w_044_4685, w_044_4687, w_044_4688, w_044_4697, w_044_4700, w_044_4702, w_044_4703, w_044_4704, w_044_4706, w_044_4708, w_044_4709, w_044_4713, w_044_4719, w_044_4720, w_044_4721, w_044_4722, w_044_4724, w_044_4725, w_044_4726, w_044_4729, w_044_4730, w_044_4731, w_044_4733, w_044_4735, w_044_4737, w_044_4738, w_044_4739, w_044_4740, w_044_4743, w_044_4744, w_044_4745, w_044_4748, w_044_4751, w_044_4752, w_044_4754, w_044_4756, w_044_4757, w_044_4758, w_044_4759, w_044_4761, w_044_4762, w_044_4763, w_044_4764, w_044_4766, w_044_4767, w_044_4768, w_044_4770, w_044_4771, w_044_4773, w_044_4774, w_044_4777, w_044_4780, w_044_4782, w_044_4784, w_044_4791, w_044_4793, w_044_4794, w_044_4797, w_044_4798, w_044_4800, w_044_4802, w_044_4805, w_044_4807, w_044_4810, w_044_4811, w_044_4812, w_044_4815, w_044_4816, w_044_4822, w_044_4823, w_044_4827, w_044_4828, w_044_4830, w_044_4831, w_044_4834, w_044_4838, w_044_4839, w_044_4840, w_044_4841, w_044_4842, w_044_4846, w_044_4850, w_044_4851, w_044_4852, w_044_4853, w_044_4854, w_044_4855, w_044_4857, w_044_4859, w_044_4860, w_044_4861, w_044_4863, w_044_4865, w_044_4867, w_044_4868, w_044_4870, w_044_4871, w_044_4873, w_044_4874, w_044_4883, w_044_4886, w_044_4888, w_044_4890, w_044_4891, w_044_4892, w_044_4893, w_044_4896, w_044_4899, w_044_4903, w_044_4906, w_044_4907, w_044_4908, w_044_4909, w_044_4911, w_044_4914, w_044_4915, w_044_4917, w_044_4920, w_044_4921, w_044_4922, w_044_4923, w_044_4924, w_044_4925, w_044_4927, w_044_4928, w_044_4931, w_044_4932, w_044_4933, w_044_4934, w_044_4935, w_044_4936, w_044_4937, w_044_4938, w_044_4939, w_044_4940, w_044_4941, w_044_4943, w_044_4945, w_044_4946, w_044_4947, w_044_4948, w_044_4949, w_044_4950, w_044_4951, w_044_4952, w_044_4954, w_044_4956, w_044_4957, w_044_4958, w_044_4959, w_044_4961, w_044_4963, w_044_4964, w_044_4965, w_044_4966, w_044_4967, w_044_4968, w_044_4969, w_044_4970, w_044_4971, w_044_4973, w_044_4975, w_044_4976, w_044_4977, w_044_4978, w_044_4979, w_044_4980, w_044_4981, w_044_4982, w_044_4983, w_044_4984, w_044_4986;
  wire w_045_000, w_045_001, w_045_002, w_045_003, w_045_004, w_045_005, w_045_006, w_045_009, w_045_010, w_045_011, w_045_012, w_045_013, w_045_014, w_045_015, w_045_016, w_045_017, w_045_018, w_045_021, w_045_022, w_045_023, w_045_024, w_045_025, w_045_026, w_045_027, w_045_028, w_045_029, w_045_030, w_045_031, w_045_032, w_045_034, w_045_035, w_045_036, w_045_037, w_045_039, w_045_040, w_045_041, w_045_042, w_045_043, w_045_044, w_045_045, w_045_046, w_045_047, w_045_048, w_045_049, w_045_050, w_045_051, w_045_052, w_045_053, w_045_054, w_045_055, w_045_056, w_045_057, w_045_058, w_045_060, w_045_061, w_045_062, w_045_063, w_045_064, w_045_065, w_045_066, w_045_067, w_045_068, w_045_069, w_045_070, w_045_071, w_045_072, w_045_073, w_045_074, w_045_075, w_045_076, w_045_077, w_045_078, w_045_079, w_045_080, w_045_083, w_045_084, w_045_085, w_045_086, w_045_087, w_045_088, w_045_089, w_045_090, w_045_091, w_045_092, w_045_093, w_045_094, w_045_095, w_045_096, w_045_097, w_045_098, w_045_099, w_045_100, w_045_101, w_045_103, w_045_104, w_045_105, w_045_106, w_045_107, w_045_108, w_045_109, w_045_110, w_045_111, w_045_112, w_045_113, w_045_114, w_045_115, w_045_116, w_045_117, w_045_118, w_045_119, w_045_120, w_045_121, w_045_122, w_045_123, w_045_124, w_045_125, w_045_126, w_045_127, w_045_128, w_045_129, w_045_131, w_045_132, w_045_133, w_045_134, w_045_136, w_045_137, w_045_138, w_045_139, w_045_140, w_045_141, w_045_143, w_045_144, w_045_145, w_045_146, w_045_147, w_045_148, w_045_149, w_045_150, w_045_151, w_045_152, w_045_153, w_045_154, w_045_156, w_045_157, w_045_158, w_045_159, w_045_161, w_045_162, w_045_163, w_045_166, w_045_167, w_045_169, w_045_170, w_045_171, w_045_172, w_045_173, w_045_174, w_045_175, w_045_176, w_045_177, w_045_178, w_045_179, w_045_180, w_045_181, w_045_182, w_045_183, w_045_184, w_045_186, w_045_188, w_045_189, w_045_190, w_045_192, w_045_193, w_045_194, w_045_195, w_045_196, w_045_197, w_045_199, w_045_200, w_045_201, w_045_202, w_045_203, w_045_204, w_045_205, w_045_206, w_045_207, w_045_208, w_045_209, w_045_210, w_045_211, w_045_212, w_045_213, w_045_214, w_045_215, w_045_216, w_045_217, w_045_218, w_045_219, w_045_220, w_045_221, w_045_222, w_045_223, w_045_224, w_045_225, w_045_226, w_045_227, w_045_228, w_045_229, w_045_230, w_045_232, w_045_235, w_045_236, w_045_237, w_045_238, w_045_239, w_045_240, w_045_241, w_045_242, w_045_243, w_045_244, w_045_245, w_045_246, w_045_247, w_045_248, w_045_249, w_045_250, w_045_251, w_045_252, w_045_253, w_045_254, w_045_255, w_045_256, w_045_257, w_045_260, w_045_261, w_045_262, w_045_263, w_045_264, w_045_265, w_045_266, w_045_267, w_045_268, w_045_269, w_045_270, w_045_271, w_045_272, w_045_273, w_045_274, w_045_275, w_045_276, w_045_277, w_045_278, w_045_279, w_045_281, w_045_282, w_045_283, w_045_284, w_045_285, w_045_286, w_045_287, w_045_288, w_045_289, w_045_290, w_045_291, w_045_292, w_045_293, w_045_294, w_045_295, w_045_296, w_045_297, w_045_298, w_045_299, w_045_300, w_045_301, w_045_302, w_045_303, w_045_304, w_045_305, w_045_306, w_045_307, w_045_308, w_045_309, w_045_310, w_045_311, w_045_312, w_045_313, w_045_314, w_045_316, w_045_317, w_045_318, w_045_319, w_045_320, w_045_322, w_045_323, w_045_324, w_045_325, w_045_326, w_045_327, w_045_328, w_045_329, w_045_330, w_045_331, w_045_333, w_045_334, w_045_335, w_045_336, w_045_337, w_045_338, w_045_339, w_045_340, w_045_342, w_045_343, w_045_345, w_045_346, w_045_347, w_045_348, w_045_349, w_045_350, w_045_351, w_045_352, w_045_353, w_045_354, w_045_355, w_045_356, w_045_357, w_045_358, w_045_360, w_045_361, w_045_362, w_045_363, w_045_364, w_045_365, w_045_367, w_045_368, w_045_369, w_045_370, w_045_371, w_045_372, w_045_373, w_045_374, w_045_375, w_045_376, w_045_377, w_045_378, w_045_379, w_045_380, w_045_381, w_045_382, w_045_383, w_045_384, w_045_387, w_045_388, w_045_389, w_045_390, w_045_391, w_045_392, w_045_393, w_045_394, w_045_395, w_045_396, w_045_397, w_045_398, w_045_399, w_045_400, w_045_401, w_045_402, w_045_403, w_045_404, w_045_405, w_045_406, w_045_407, w_045_408, w_045_409, w_045_410, w_045_411, w_045_412, w_045_413, w_045_415, w_045_416, w_045_417, w_045_418, w_045_419, w_045_420, w_045_421, w_045_422, w_045_423, w_045_424, w_045_426, w_045_427, w_045_428, w_045_429, w_045_430, w_045_431, w_045_432, w_045_433, w_045_435, w_045_436, w_045_437, w_045_438, w_045_439, w_045_440, w_045_442, w_045_443, w_045_444, w_045_445, w_045_446, w_045_448, w_045_449, w_045_450, w_045_451, w_045_452, w_045_453, w_045_454, w_045_455, w_045_456, w_045_457, w_045_458, w_045_459, w_045_460, w_045_461, w_045_462, w_045_463, w_045_464, w_045_465, w_045_466, w_045_467, w_045_468, w_045_469, w_045_471, w_045_472, w_045_473, w_045_474, w_045_475, w_045_476, w_045_477, w_045_478, w_045_479, w_045_480, w_045_481, w_045_483, w_045_484, w_045_485, w_045_486, w_045_489, w_045_490, w_045_491, w_045_492, w_045_493, w_045_494, w_045_495, w_045_496, w_045_497, w_045_498, w_045_500, w_045_501, w_045_502, w_045_503, w_045_504, w_045_505, w_045_506, w_045_508, w_045_509, w_045_510, w_045_511, w_045_512, w_045_515, w_045_516, w_045_517, w_045_518, w_045_519, w_045_520, w_045_521, w_045_523, w_045_524, w_045_528, w_045_529, w_045_530, w_045_531, w_045_532, w_045_533, w_045_534, w_045_535, w_045_536, w_045_537, w_045_538, w_045_539, w_045_540, w_045_541, w_045_542, w_045_543, w_045_544, w_045_545, w_045_546, w_045_547, w_045_548, w_045_549, w_045_550, w_045_551, w_045_552, w_045_553, w_045_554, w_045_555, w_045_556, w_045_557, w_045_558, w_045_559, w_045_560, w_045_561, w_045_562, w_045_563, w_045_564, w_045_565, w_045_566, w_045_567, w_045_568, w_045_569, w_045_570, w_045_571, w_045_572, w_045_574, w_045_575, w_045_576, w_045_577, w_045_578, w_045_579, w_045_580, w_045_582, w_045_583, w_045_584, w_045_585, w_045_586, w_045_587, w_045_588, w_045_589, w_045_591, w_045_592, w_045_593, w_045_594, w_045_595, w_045_596, w_045_597, w_045_598, w_045_599, w_045_600, w_045_601, w_045_602, w_045_603, w_045_604, w_045_605, w_045_606, w_045_607, w_045_608, w_045_609, w_045_610, w_045_611, w_045_612, w_045_613, w_045_614, w_045_615, w_045_618, w_045_619, w_045_620, w_045_621, w_045_622, w_045_623, w_045_624, w_045_625, w_045_626, w_045_628, w_045_629, w_045_630, w_045_632, w_045_633, w_045_634, w_045_635, w_045_637, w_045_638, w_045_639, w_045_640, w_045_641, w_045_642, w_045_643, w_045_644, w_045_645, w_045_646, w_045_647, w_045_648, w_045_649, w_045_650, w_045_651, w_045_653, w_045_654, w_045_656, w_045_659, w_045_660, w_045_661, w_045_662, w_045_663, w_045_664, w_045_667, w_045_668, w_045_669, w_045_670, w_045_671, w_045_673, w_045_674, w_045_676, w_045_678, w_045_680, w_045_681, w_045_682, w_045_683, w_045_684, w_045_687, w_045_688, w_045_689, w_045_690, w_045_692, w_045_693, w_045_696, w_045_698, w_045_699, w_045_700, w_045_701, w_045_703, w_045_704, w_045_707, w_045_708, w_045_710, w_045_713, w_045_714, w_045_716, w_045_717, w_045_718, w_045_722, w_045_723, w_045_724, w_045_725, w_045_726, w_045_727, w_045_728, w_045_731, w_045_732, w_045_734, w_045_735, w_045_736, w_045_737, w_045_738, w_045_739, w_045_740, w_045_741, w_045_742, w_045_744, w_045_745, w_045_747, w_045_748, w_045_749, w_045_750, w_045_751, w_045_753, w_045_754, w_045_755, w_045_756, w_045_759, w_045_762, w_045_763, w_045_765, w_045_766, w_045_767, w_045_769, w_045_770, w_045_771, w_045_772, w_045_774, w_045_775, w_045_777, w_045_778, w_045_779, w_045_781, w_045_782, w_045_783, w_045_784, w_045_785, w_045_788, w_045_789, w_045_791, w_045_792, w_045_795, w_045_796, w_045_798, w_045_799, w_045_800, w_045_801, w_045_802, w_045_803, w_045_804, w_045_805, w_045_806, w_045_807, w_045_808, w_045_812, w_045_813, w_045_814, w_045_815, w_045_816, w_045_817, w_045_819, w_045_820, w_045_821, w_045_822, w_045_824, w_045_825, w_045_827, w_045_828, w_045_829, w_045_830, w_045_831, w_045_832, w_045_833, w_045_834, w_045_835, w_045_836, w_045_837, w_045_838, w_045_841, w_045_842, w_045_844, w_045_846, w_045_848, w_045_849, w_045_853, w_045_854, w_045_855, w_045_856, w_045_857, w_045_858, w_045_859, w_045_861, w_045_862, w_045_864, w_045_865, w_045_866, w_045_867, w_045_868, w_045_870, w_045_871, w_045_872, w_045_873, w_045_874, w_045_875, w_045_877, w_045_878, w_045_879, w_045_880, w_045_881, w_045_882, w_045_884, w_045_885, w_045_886, w_045_887, w_045_888, w_045_890, w_045_891, w_045_895, w_045_896, w_045_897, w_045_898, w_045_899, w_045_900, w_045_901, w_045_903, w_045_905, w_045_906, w_045_912, w_045_913, w_045_914, w_045_915, w_045_916, w_045_917, w_045_919, w_045_920, w_045_921, w_045_923, w_045_925, w_045_926, w_045_927, w_045_929, w_045_930, w_045_931, w_045_932, w_045_933, w_045_934, w_045_936, w_045_938, w_045_939, w_045_940, w_045_942, w_045_943, w_045_944, w_045_947, w_045_948, w_045_950, w_045_952, w_045_953, w_045_955, w_045_956, w_045_957, w_045_958, w_045_960, w_045_961, w_045_962, w_045_963, w_045_964, w_045_965, w_045_966, w_045_967, w_045_969, w_045_970, w_045_971, w_045_972, w_045_975, w_045_976, w_045_977, w_045_979, w_045_981, w_045_982, w_045_983, w_045_985, w_045_986, w_045_988, w_045_989, w_045_990, w_045_992, w_045_993, w_045_994, w_045_996, w_045_998, w_045_999, w_045_1000, w_045_1002, w_045_1003, w_045_1005, w_045_1007, w_045_1009, w_045_1013, w_045_1014, w_045_1015, w_045_1016, w_045_1018, w_045_1021, w_045_1022, w_045_1024, w_045_1025, w_045_1026, w_045_1027, w_045_1030, w_045_1031, w_045_1032, w_045_1033, w_045_1036, w_045_1038, w_045_1039, w_045_1040, w_045_1041, w_045_1043, w_045_1044, w_045_1045, w_045_1047, w_045_1050, w_045_1051, w_045_1052, w_045_1054, w_045_1056, w_045_1057, w_045_1059, w_045_1060, w_045_1061, w_045_1062, w_045_1063, w_045_1065, w_045_1066, w_045_1067, w_045_1073, w_045_1074, w_045_1075, w_045_1076, w_045_1077, w_045_1078, w_045_1079, w_045_1080, w_045_1081, w_045_1082, w_045_1083, w_045_1086, w_045_1087, w_045_1088, w_045_1089, w_045_1090, w_045_1091, w_045_1092, w_045_1094, w_045_1096, w_045_1097, w_045_1099, w_045_1100, w_045_1101, w_045_1102, w_045_1103, w_045_1105, w_045_1106, w_045_1107, w_045_1108, w_045_1112, w_045_1113, w_045_1114, w_045_1115, w_045_1116, w_045_1117, w_045_1119, w_045_1120, w_045_1121, w_045_1122, w_045_1123, w_045_1124, w_045_1125, w_045_1127, w_045_1128, w_045_1129, w_045_1130, w_045_1131, w_045_1132, w_045_1134, w_045_1135, w_045_1136, w_045_1137, w_045_1138, w_045_1139, w_045_1140, w_045_1141, w_045_1145, w_045_1146, w_045_1148, w_045_1149, w_045_1151, w_045_1152, w_045_1153, w_045_1154, w_045_1155, w_045_1156, w_045_1157, w_045_1158, w_045_1160, w_045_1161, w_045_1164, w_045_1166, w_045_1167, w_045_1169, w_045_1170, w_045_1171, w_045_1173, w_045_1174, w_045_1175, w_045_1176, w_045_1177, w_045_1178, w_045_1179, w_045_1180, w_045_1182, w_045_1183, w_045_1184, w_045_1186, w_045_1187, w_045_1188, w_045_1189, w_045_1190, w_045_1191, w_045_1192, w_045_1193, w_045_1197, w_045_1198, w_045_1199, w_045_1200, w_045_1201, w_045_1203, w_045_1205, w_045_1207, w_045_1208, w_045_1209, w_045_1211, w_045_1212, w_045_1213, w_045_1214, w_045_1216, w_045_1217, w_045_1218, w_045_1219, w_045_1221, w_045_1223, w_045_1224, w_045_1225, w_045_1227, w_045_1231, w_045_1234, w_045_1235, w_045_1236, w_045_1237, w_045_1238, w_045_1240, w_045_1241, w_045_1242, w_045_1244, w_045_1245, w_045_1246, w_045_1247, w_045_1248, w_045_1249, w_045_1250, w_045_1251, w_045_1253, w_045_1254, w_045_1255, w_045_1256, w_045_1257, w_045_1258, w_045_1259, w_045_1260, w_045_1261, w_045_1262, w_045_1263, w_045_1264, w_045_1265, w_045_1266, w_045_1267, w_045_1268, w_045_1270, w_045_1271, w_045_1272, w_045_1273, w_045_1274, w_045_1275, w_045_1276, w_045_1277, w_045_1278, w_045_1279, w_045_1280, w_045_1281, w_045_1284, w_045_1285, w_045_1288, w_045_1289, w_045_1290, w_045_1291, w_045_1292, w_045_1293, w_045_1296, w_045_1298, w_045_1299, w_045_1300, w_045_1301, w_045_1302, w_045_1304, w_045_1305, w_045_1306, w_045_1307, w_045_1309, w_045_1310, w_045_1311, w_045_1312, w_045_1315, w_045_1316, w_045_1318, w_045_1319, w_045_1321, w_045_1322, w_045_1323, w_045_1324, w_045_1327, w_045_1328, w_045_1329, w_045_1330, w_045_1331, w_045_1332, w_045_1333, w_045_1334, w_045_1335, w_045_1336, w_045_1338, w_045_1340, w_045_1341, w_045_1343, w_045_1344, w_045_1345, w_045_1346, w_045_1348, w_045_1349, w_045_1352, w_045_1353, w_045_1354, w_045_1355, w_045_1356, w_045_1357, w_045_1358, w_045_1359, w_045_1362, w_045_1363, w_045_1365, w_045_1366, w_045_1367, w_045_1368, w_045_1370, w_045_1371, w_045_1375, w_045_1376, w_045_1378, w_045_1379, w_045_1380, w_045_1381, w_045_1382, w_045_1383, w_045_1384, w_045_1385, w_045_1386, w_045_1387, w_045_1388, w_045_1389, w_045_1390, w_045_1391, w_045_1392, w_045_1393, w_045_1394, w_045_1395, w_045_1396, w_045_1398, w_045_1401, w_045_1402, w_045_1403, w_045_1404, w_045_1405, w_045_1406, w_045_1407, w_045_1408, w_045_1409, w_045_1410, w_045_1411, w_045_1412, w_045_1413, w_045_1414, w_045_1415, w_045_1416, w_045_1417, w_045_1418, w_045_1419, w_045_1420, w_045_1422, w_045_1423, w_045_1424, w_045_1425, w_045_1426, w_045_1427, w_045_1432, w_045_1434, w_045_1435, w_045_1438, w_045_1439, w_045_1440, w_045_1441, w_045_1442, w_045_1443, w_045_1444, w_045_1445, w_045_1446, w_045_1447, w_045_1448, w_045_1450, w_045_1451, w_045_1453, w_045_1454, w_045_1456, w_045_1457, w_045_1458, w_045_1459, w_045_1462, w_045_1463, w_045_1464, w_045_1468, w_045_1472, w_045_1474, w_045_1475, w_045_1476, w_045_1477, w_045_1478, w_045_1479, w_045_1480, w_045_1481, w_045_1482, w_045_1483, w_045_1484, w_045_1487, w_045_1488, w_045_1489, w_045_1490, w_045_1491, w_045_1492, w_045_1493, w_045_1497, w_045_1498, w_045_1499, w_045_1500, w_045_1504, w_045_1505, w_045_1506, w_045_1507, w_045_1509, w_045_1510, w_045_1511, w_045_1512, w_045_1513, w_045_1514, w_045_1515, w_045_1516, w_045_1519, w_045_1520, w_045_1521, w_045_1523, w_045_1525, w_045_1528, w_045_1529, w_045_1530, w_045_1532, w_045_1533, w_045_1534, w_045_1535, w_045_1537, w_045_1538, w_045_1539, w_045_1541, w_045_1543, w_045_1544, w_045_1546, w_045_1547, w_045_1548, w_045_1550, w_045_1551, w_045_1552, w_045_1556, w_045_1557, w_045_1559, w_045_1562, w_045_1563, w_045_1564, w_045_1565, w_045_1567, w_045_1568, w_045_1569, w_045_1571, w_045_1572, w_045_1573, w_045_1574, w_045_1575, w_045_1576, w_045_1577, w_045_1578, w_045_1579, w_045_1580, w_045_1581, w_045_1582, w_045_1583, w_045_1584, w_045_1585, w_045_1587, w_045_1589, w_045_1590, w_045_1591, w_045_1592, w_045_1593, w_045_1594, w_045_1595, w_045_1596, w_045_1597, w_045_1598, w_045_1599, w_045_1600, w_045_1601, w_045_1602, w_045_1603, w_045_1605, w_045_1607, w_045_1608, w_045_1609, w_045_1610, w_045_1611, w_045_1612, w_045_1615, w_045_1616, w_045_1617, w_045_1619, w_045_1620, w_045_1622, w_045_1623, w_045_1624, w_045_1625, w_045_1626, w_045_1627, w_045_1628, w_045_1629, w_045_1630, w_045_1631, w_045_1632, w_045_1634, w_045_1635, w_045_1636, w_045_1638, w_045_1639, w_045_1640, w_045_1641, w_045_1643, w_045_1644, w_045_1645, w_045_1646, w_045_1647, w_045_1649, w_045_1650, w_045_1651, w_045_1652, w_045_1654, w_045_1655, w_045_1656, w_045_1657, w_045_1659, w_045_1660, w_045_1661, w_045_1662, w_045_1665, w_045_1666, w_045_1669, w_045_1671, w_045_1672, w_045_1673, w_045_1675, w_045_1677, w_045_1678, w_045_1679, w_045_1681, w_045_1683, w_045_1685, w_045_1686, w_045_1688, w_045_1690, w_045_1691, w_045_1694, w_045_1695, w_045_1696, w_045_1697, w_045_1698, w_045_1699, w_045_1700, w_045_1701, w_045_1702, w_045_1703, w_045_1704, w_045_1705, w_045_1707, w_045_1708, w_045_1709, w_045_1711, w_045_1712, w_045_1713, w_045_1714, w_045_1715, w_045_1716, w_045_1717, w_045_1719, w_045_1720, w_045_1721, w_045_1722, w_045_1723, w_045_1725, w_045_1727, w_045_1728, w_045_1729, w_045_1730, w_045_1731, w_045_1732, w_045_1733, w_045_1735, w_045_1736, w_045_1739, w_045_1740, w_045_1741, w_045_1742, w_045_1743, w_045_1744, w_045_1746, w_045_1747, w_045_1748, w_045_1749, w_045_1750, w_045_1751, w_045_1752, w_045_1754, w_045_1755, w_045_1756, w_045_1757, w_045_1758, w_045_1759, w_045_1760, w_045_1762, w_045_1763, w_045_1765, w_045_1766, w_045_1768, w_045_1769, w_045_1770, w_045_1771, w_045_1774, w_045_1775, w_045_1777, w_045_1778, w_045_1779, w_045_1781, w_045_1784, w_045_1785, w_045_1786, w_045_1787, w_045_1788, w_045_1789, w_045_1790, w_045_1791, w_045_1792, w_045_1793, w_045_1794, w_045_1795, w_045_1796, w_045_1797, w_045_1798, w_045_1800, w_045_1801, w_045_1802, w_045_1803, w_045_1804, w_045_1806, w_045_1807, w_045_1809, w_045_1810, w_045_1811, w_045_1813, w_045_1814, w_045_1815, w_045_1816, w_045_1817, w_045_1818, w_045_1819, w_045_1820, w_045_1821, w_045_1822, w_045_1824, w_045_1825, w_045_1826, w_045_1828, w_045_1829, w_045_1830, w_045_1831, w_045_1832, w_045_1833, w_045_1834, w_045_1835, w_045_1836, w_045_1837, w_045_1840, w_045_1841, w_045_1842, w_045_1843, w_045_1844, w_045_1846, w_045_1847, w_045_1848, w_045_1849, w_045_1850, w_045_1853, w_045_1856, w_045_1857, w_045_1858, w_045_1859, w_045_1860, w_045_1863, w_045_1865, w_045_1867, w_045_1868, w_045_1869, w_045_1872, w_045_1873, w_045_1876, w_045_1877, w_045_1878, w_045_1879, w_045_1880, w_045_1881, w_045_1882, w_045_1884, w_045_1885, w_045_1886, w_045_1889, w_045_1890, w_045_1892, w_045_1893, w_045_1894, w_045_1895, w_045_1896, w_045_1897, w_045_1898, w_045_1899, w_045_1900, w_045_1901, w_045_1903, w_045_1904, w_045_1905, w_045_1906, w_045_1907, w_045_1908, w_045_1910, w_045_1912, w_045_1913, w_045_1914, w_045_1915, w_045_1916, w_045_1917, w_045_1918, w_045_1919, w_045_1920, w_045_1921, w_045_1923, w_045_1924, w_045_1925, w_045_1926, w_045_1927, w_045_1928, w_045_1929, w_045_1930, w_045_1931, w_045_1932, w_045_1933, w_045_1934, w_045_1937, w_045_1939, w_045_1941, w_045_1942, w_045_1943, w_045_1944, w_045_1947, w_045_1948, w_045_1950, w_045_1951, w_045_1952, w_045_1953, w_045_1955, w_045_1957, w_045_1958, w_045_1959, w_045_1960, w_045_1962, w_045_1964, w_045_1966, w_045_1967, w_045_1969, w_045_1970, w_045_1971, w_045_1972, w_045_1974, w_045_1975, w_045_1978, w_045_1980, w_045_1981, w_045_1982, w_045_1983, w_045_1984, w_045_1985, w_045_1986, w_045_1990, w_045_1991, w_045_1992, w_045_1993, w_045_1994, w_045_1995, w_045_1996, w_045_1997, w_045_1998, w_045_1999, w_045_2000, w_045_2002, w_045_2003, w_045_2004, w_045_2009, w_045_2010, w_045_2011, w_045_2012, w_045_2013, w_045_2015, w_045_2017, w_045_2018, w_045_2021, w_045_2022, w_045_2023, w_045_2024, w_045_2025, w_045_2026, w_045_2027, w_045_2028, w_045_2030, w_045_2032, w_045_2033, w_045_2034, w_045_2036, w_045_2037, w_045_2038, w_045_2039, w_045_2040, w_045_2041, w_045_2042, w_045_2043, w_045_2045, w_045_2046, w_045_2047, w_045_2049, w_045_2052, w_045_2053, w_045_2055, w_045_2056, w_045_2057, w_045_2060, w_045_2061, w_045_2062, w_045_2064, w_045_2065, w_045_2066, w_045_2068, w_045_2069, w_045_2070, w_045_2071, w_045_2072, w_045_2073, w_045_2074, w_045_2076, w_045_2079, w_045_2080, w_045_2081, w_045_2082, w_045_2083, w_045_2084, w_045_2085, w_045_2086, w_045_2087, w_045_2088, w_045_2090, w_045_2091, w_045_2093, w_045_2094, w_045_2095, w_045_2097, w_045_2098, w_045_2099, w_045_2100, w_045_2101, w_045_2102, w_045_2103, w_045_2104, w_045_2105, w_045_2106, w_045_2107, w_045_2108, w_045_2110, w_045_2111, w_045_2112, w_045_2113, w_045_2114, w_045_2115, w_045_2116, w_045_2117, w_045_2119, w_045_2120, w_045_2122, w_045_2124, w_045_2125, w_045_2126, w_045_2130, w_045_2132, w_045_2133, w_045_2134, w_045_2135, w_045_2136, w_045_2138, w_045_2140, w_045_2141, w_045_2142, w_045_2143, w_045_2144, w_045_2145, w_045_2146, w_045_2147, w_045_2149, w_045_2151, w_045_2152, w_045_2153, w_045_2154, w_045_2155, w_045_2156, w_045_2157, w_045_2159, w_045_2161, w_045_2162, w_045_2163, w_045_2166, w_045_2167, w_045_2168, w_045_2169, w_045_2170, w_045_2171;
  wire w_046_001, w_046_002, w_046_003, w_046_005, w_046_007, w_046_008, w_046_009, w_046_011, w_046_012, w_046_013, w_046_014, w_046_015, w_046_016, w_046_018, w_046_019, w_046_020, w_046_022, w_046_023, w_046_025, w_046_026, w_046_027, w_046_028, w_046_029, w_046_031, w_046_032, w_046_035, w_046_036, w_046_038, w_046_040, w_046_041, w_046_042, w_046_044, w_046_045, w_046_046, w_046_047, w_046_049, w_046_050, w_046_053, w_046_055, w_046_056, w_046_057, w_046_058, w_046_059, w_046_060, w_046_061, w_046_063, w_046_065, w_046_066, w_046_067, w_046_068, w_046_069, w_046_070, w_046_071, w_046_072, w_046_073, w_046_074, w_046_075, w_046_076, w_046_077, w_046_078, w_046_079, w_046_080, w_046_083, w_046_084, w_046_085, w_046_086, w_046_087, w_046_088, w_046_089, w_046_091, w_046_092, w_046_093, w_046_094, w_046_096, w_046_098, w_046_099, w_046_100, w_046_101, w_046_102, w_046_103, w_046_104, w_046_105, w_046_107, w_046_108, w_046_110, w_046_111, w_046_112, w_046_114, w_046_115, w_046_117, w_046_118, w_046_119, w_046_120, w_046_121, w_046_122, w_046_123, w_046_124, w_046_126, w_046_127, w_046_128, w_046_129, w_046_130, w_046_131, w_046_132, w_046_133, w_046_134, w_046_135, w_046_136, w_046_137, w_046_138, w_046_139, w_046_140, w_046_141, w_046_143, w_046_144, w_046_146, w_046_147, w_046_148, w_046_149, w_046_152, w_046_154, w_046_155, w_046_157, w_046_159, w_046_162, w_046_163, w_046_164, w_046_165, w_046_166, w_046_167, w_046_168, w_046_169, w_046_170, w_046_171, w_046_172, w_046_173, w_046_174, w_046_177, w_046_178, w_046_180, w_046_181, w_046_183, w_046_184, w_046_185, w_046_187, w_046_188, w_046_189, w_046_191, w_046_192, w_046_193, w_046_194, w_046_195, w_046_199, w_046_200, w_046_201, w_046_204, w_046_205, w_046_207, w_046_209, w_046_210, w_046_213, w_046_214, w_046_216, w_046_217, w_046_218, w_046_219, w_046_220, w_046_222, w_046_223, w_046_227, w_046_229, w_046_231, w_046_232, w_046_234, w_046_235, w_046_236, w_046_237, w_046_238, w_046_239, w_046_241, w_046_242, w_046_244, w_046_246, w_046_247, w_046_248, w_046_249, w_046_250, w_046_252, w_046_254, w_046_255, w_046_256, w_046_257, w_046_258, w_046_262, w_046_264, w_046_265, w_046_266, w_046_268, w_046_269, w_046_270, w_046_271, w_046_272, w_046_275, w_046_276, w_046_279, w_046_280, w_046_281, w_046_284, w_046_285, w_046_286, w_046_287, w_046_288, w_046_292, w_046_293, w_046_294, w_046_296, w_046_298, w_046_299, w_046_300, w_046_301, w_046_302, w_046_303, w_046_304, w_046_305, w_046_306, w_046_307, w_046_311, w_046_312, w_046_314, w_046_315, w_046_316, w_046_317, w_046_319, w_046_320, w_046_321, w_046_325, w_046_326, w_046_327, w_046_329, w_046_330, w_046_331, w_046_333, w_046_335, w_046_336, w_046_337, w_046_338, w_046_340, w_046_341, w_046_342, w_046_343, w_046_345, w_046_346, w_046_347, w_046_348, w_046_349, w_046_350, w_046_351, w_046_352, w_046_353, w_046_355, w_046_356, w_046_359, w_046_360, w_046_361, w_046_362, w_046_363, w_046_364, w_046_365, w_046_366, w_046_367, w_046_368, w_046_369, w_046_371, w_046_372, w_046_375, w_046_376, w_046_378, w_046_379, w_046_380, w_046_382, w_046_383, w_046_384, w_046_385, w_046_386, w_046_387, w_046_388, w_046_389, w_046_390, w_046_391, w_046_392, w_046_393, w_046_395, w_046_398, w_046_400, w_046_401, w_046_403, w_046_404, w_046_405, w_046_406, w_046_407, w_046_409, w_046_410, w_046_411, w_046_412, w_046_413, w_046_414, w_046_415, w_046_416, w_046_417, w_046_419, w_046_420, w_046_421, w_046_422, w_046_423, w_046_424, w_046_425, w_046_426, w_046_427, w_046_429, w_046_432, w_046_434, w_046_435, w_046_436, w_046_437, w_046_438, w_046_440, w_046_445, w_046_446, w_046_447, w_046_451, w_046_456, w_046_458, w_046_459, w_046_461, w_046_463, w_046_464, w_046_465, w_046_466, w_046_467, w_046_468, w_046_469, w_046_470, w_046_471, w_046_473, w_046_474, w_046_475, w_046_477, w_046_479, w_046_480, w_046_481, w_046_482, w_046_483, w_046_484, w_046_485, w_046_487, w_046_489, w_046_490, w_046_491, w_046_492, w_046_493, w_046_494, w_046_495, w_046_496, w_046_497, w_046_498, w_046_499, w_046_500, w_046_501, w_046_502, w_046_504, w_046_506, w_046_507, w_046_509, w_046_510, w_046_511, w_046_512, w_046_513, w_046_514, w_046_515, w_046_517, w_046_518, w_046_520, w_046_521, w_046_522, w_046_523, w_046_524, w_046_525, w_046_526, w_046_527, w_046_528, w_046_529, w_046_530, w_046_531, w_046_532, w_046_533, w_046_534, w_046_535, w_046_537, w_046_538, w_046_539, w_046_540, w_046_541, w_046_542, w_046_545, w_046_547, w_046_548, w_046_549, w_046_551, w_046_552, w_046_553, w_046_554, w_046_556, w_046_557, w_046_558, w_046_559, w_046_560, w_046_561, w_046_562, w_046_563, w_046_564, w_046_566, w_046_569, w_046_570, w_046_571, w_046_573, w_046_574, w_046_577, w_046_581, w_046_582, w_046_583, w_046_584, w_046_586, w_046_587, w_046_588, w_046_589, w_046_593, w_046_595, w_046_596, w_046_597, w_046_598, w_046_599, w_046_600, w_046_604, w_046_605, w_046_606, w_046_608, w_046_609, w_046_610, w_046_611, w_046_612, w_046_613, w_046_614, w_046_615, w_046_617, w_046_618, w_046_619, w_046_620, w_046_621, w_046_622, w_046_624, w_046_625, w_046_628, w_046_629, w_046_630, w_046_631, w_046_632, w_046_633, w_046_634, w_046_635, w_046_636, w_046_638, w_046_639, w_046_640, w_046_641, w_046_645, w_046_646, w_046_647, w_046_648, w_046_649, w_046_650, w_046_651, w_046_654, w_046_656, w_046_657, w_046_659, w_046_660, w_046_662, w_046_664, w_046_665, w_046_667, w_046_668, w_046_670, w_046_671, w_046_672, w_046_673, w_046_674, w_046_675, w_046_676, w_046_677, w_046_678, w_046_680, w_046_682, w_046_683, w_046_685, w_046_686, w_046_687, w_046_688, w_046_689, w_046_690, w_046_691, w_046_692, w_046_693, w_046_695, w_046_696, w_046_697, w_046_698, w_046_700, w_046_701, w_046_702, w_046_703, w_046_704, w_046_706, w_046_707, w_046_708, w_046_709, w_046_711, w_046_713, w_046_714, w_046_715, w_046_716, w_046_717, w_046_718, w_046_719, w_046_720, w_046_721, w_046_722, w_046_723, w_046_724, w_046_726, w_046_727, w_046_728, w_046_729, w_046_730, w_046_731, w_046_734, w_046_735, w_046_736, w_046_737, w_046_739, w_046_740, w_046_742, w_046_743, w_046_744, w_046_745, w_046_746, w_046_747, w_046_748, w_046_750, w_046_751, w_046_752, w_046_754, w_046_756, w_046_757, w_046_758, w_046_760, w_046_762, w_046_763, w_046_764, w_046_765, w_046_766, w_046_767, w_046_768, w_046_769, w_046_771, w_046_772, w_046_773, w_046_774, w_046_775, w_046_776, w_046_778, w_046_781, w_046_783, w_046_784, w_046_787, w_046_788, w_046_789, w_046_791, w_046_792, w_046_793, w_046_794, w_046_796, w_046_797, w_046_798, w_046_799, w_046_800, w_046_801, w_046_804, w_046_805, w_046_806, w_046_807, w_046_808, w_046_809, w_046_810, w_046_812, w_046_813, w_046_814, w_046_815, w_046_816, w_046_817, w_046_819, w_046_820, w_046_821, w_046_822, w_046_823, w_046_824, w_046_825, w_046_826, w_046_827, w_046_828, w_046_830, w_046_831, w_046_833, w_046_834, w_046_835, w_046_837, w_046_838, w_046_839, w_046_840, w_046_841, w_046_843, w_046_844, w_046_846, w_046_849, w_046_850, w_046_851, w_046_852, w_046_853, w_046_854, w_046_855, w_046_857, w_046_858, w_046_860, w_046_861, w_046_864, w_046_865, w_046_866, w_046_868, w_046_869, w_046_871, w_046_872, w_046_873, w_046_874, w_046_875, w_046_877, w_046_879, w_046_880, w_046_881, w_046_882, w_046_883, w_046_884, w_046_885, w_046_886, w_046_889, w_046_890, w_046_891, w_046_892, w_046_894, w_046_897, w_046_898, w_046_900, w_046_901, w_046_904, w_046_905, w_046_906, w_046_909, w_046_910, w_046_911, w_046_912, w_046_913, w_046_914, w_046_916, w_046_918, w_046_919, w_046_920, w_046_921, w_046_922, w_046_923, w_046_924, w_046_925, w_046_926, w_046_927, w_046_928, w_046_929, w_046_930, w_046_931, w_046_932, w_046_933, w_046_934, w_046_936, w_046_937, w_046_938, w_046_939, w_046_940, w_046_941, w_046_942, w_046_943, w_046_946, w_046_949, w_046_953, w_046_956, w_046_957, w_046_959, w_046_960, w_046_961, w_046_962, w_046_965, w_046_966, w_046_967, w_046_969, w_046_971, w_046_972, w_046_973, w_046_974, w_046_975, w_046_977, w_046_979, w_046_981, w_046_984, w_046_985, w_046_986, w_046_987, w_046_988, w_046_991, w_046_992, w_046_993, w_046_994, w_046_995, w_046_997, w_046_1000, w_046_1002, w_046_1003, w_046_1004, w_046_1005, w_046_1006, w_046_1007, w_046_1008, w_046_1011, w_046_1012, w_046_1013, w_046_1014, w_046_1017, w_046_1020, w_046_1021, w_046_1023, w_046_1026, w_046_1027, w_046_1028, w_046_1029, w_046_1030, w_046_1031, w_046_1032, w_046_1033, w_046_1034, w_046_1035, w_046_1036, w_046_1038, w_046_1040, w_046_1041, w_046_1042, w_046_1044, w_046_1045, w_046_1048, w_046_1049, w_046_1050, w_046_1051, w_046_1053, w_046_1054, w_046_1055, w_046_1056, w_046_1057, w_046_1058, w_046_1059, w_046_1060, w_046_1061, w_046_1062, w_046_1063, w_046_1064, w_046_1067, w_046_1068, w_046_1069, w_046_1070, w_046_1071, w_046_1072, w_046_1074, w_046_1075, w_046_1076, w_046_1077, w_046_1078, w_046_1079, w_046_1081, w_046_1082, w_046_1083, w_046_1084, w_046_1085, w_046_1087, w_046_1088, w_046_1090, w_046_1091, w_046_1092, w_046_1093, w_046_1094, w_046_1097, w_046_1098, w_046_1099, w_046_1101, w_046_1103, w_046_1104, w_046_1106, w_046_1107, w_046_1109, w_046_1110, w_046_1111, w_046_1112, w_046_1113, w_046_1116, w_046_1118, w_046_1119, w_046_1120, w_046_1121, w_046_1123, w_046_1124, w_046_1125, w_046_1126, w_046_1128, w_046_1130, w_046_1131, w_046_1132, w_046_1133, w_046_1136, w_046_1137, w_046_1138, w_046_1139, w_046_1140, w_046_1144, w_046_1145, w_046_1146, w_046_1147, w_046_1148, w_046_1150, w_046_1152, w_046_1153, w_046_1154, w_046_1155, w_046_1156, w_046_1157, w_046_1158, w_046_1159, w_046_1160, w_046_1161, w_046_1162, w_046_1163, w_046_1164, w_046_1166, w_046_1167, w_046_1168, w_046_1169, w_046_1170, w_046_1171, w_046_1172, w_046_1174, w_046_1175, w_046_1177, w_046_1178, w_046_1179, w_046_1180, w_046_1181, w_046_1182, w_046_1183, w_046_1184, w_046_1185, w_046_1186, w_046_1187, w_046_1188, w_046_1191, w_046_1192, w_046_1193, w_046_1194, w_046_1197, w_046_1198, w_046_1199, w_046_1201, w_046_1202, w_046_1203, w_046_1204, w_046_1205, w_046_1206, w_046_1207, w_046_1208, w_046_1209, w_046_1210, w_046_1213, w_046_1214, w_046_1217, w_046_1218, w_046_1219, w_046_1220, w_046_1222, w_046_1223, w_046_1224, w_046_1225, w_046_1227, w_046_1228, w_046_1229, w_046_1231, w_046_1233, w_046_1234, w_046_1236, w_046_1237, w_046_1238, w_046_1239, w_046_1240, w_046_1241, w_046_1242, w_046_1243, w_046_1246, w_046_1247, w_046_1248, w_046_1249, w_046_1251, w_046_1252, w_046_1253, w_046_1255, w_046_1261, w_046_1262, w_046_1265, w_046_1266, w_046_1267, w_046_1268, w_046_1270, w_046_1271, w_046_1272, w_046_1273, w_046_1274, w_046_1275, w_046_1276, w_046_1277, w_046_1278, w_046_1279, w_046_1282, w_046_1283, w_046_1284, w_046_1285, w_046_1286, w_046_1287, w_046_1288, w_046_1290, w_046_1291, w_046_1292, w_046_1293, w_046_1297, w_046_1298, w_046_1299, w_046_1300, w_046_1301, w_046_1302, w_046_1303, w_046_1307, w_046_1309, w_046_1310, w_046_1311, w_046_1312, w_046_1313, w_046_1314, w_046_1315, w_046_1316, w_046_1317, w_046_1320, w_046_1323, w_046_1324, w_046_1325, w_046_1326, w_046_1327, w_046_1329, w_046_1330, w_046_1332, w_046_1333, w_046_1335, w_046_1338, w_046_1339, w_046_1340, w_046_1341, w_046_1343, w_046_1347, w_046_1348, w_046_1349, w_046_1350, w_046_1351, w_046_1352, w_046_1354, w_046_1355, w_046_1357, w_046_1358, w_046_1359, w_046_1360, w_046_1361, w_046_1362, w_046_1363, w_046_1364, w_046_1367, w_046_1368, w_046_1370, w_046_1372, w_046_1374, w_046_1375, w_046_1376, w_046_1377, w_046_1378, w_046_1379, w_046_1381, w_046_1382, w_046_1383, w_046_1384, w_046_1386, w_046_1387, w_046_1388, w_046_1390, w_046_1391, w_046_1392, w_046_1393, w_046_1394, w_046_1395, w_046_1396, w_046_1397, w_046_1399, w_046_1400, w_046_1401, w_046_1402, w_046_1404, w_046_1405, w_046_1406, w_046_1407, w_046_1408, w_046_1410, w_046_1411, w_046_1412, w_046_1414, w_046_1418, w_046_1419, w_046_1420, w_046_1421, w_046_1423, w_046_1425, w_046_1427, w_046_1428, w_046_1429, w_046_1431, w_046_1432, w_046_1433, w_046_1434, w_046_1436, w_046_1438, w_046_1439, w_046_1440, w_046_1441, w_046_1442, w_046_1443, w_046_1444, w_046_1447, w_046_1448, w_046_1449, w_046_1450, w_046_1451, w_046_1452, w_046_1453, w_046_1454, w_046_1455, w_046_1456, w_046_1457, w_046_1459, w_046_1460, w_046_1461, w_046_1463, w_046_1464, w_046_1465, w_046_1466, w_046_1467, w_046_1468, w_046_1469, w_046_1470, w_046_1471, w_046_1472, w_046_1473, w_046_1474, w_046_1477, w_046_1478, w_046_1479, w_046_1480, w_046_1481, w_046_1482, w_046_1483, w_046_1486, w_046_1487, w_046_1488, w_046_1489, w_046_1490, w_046_1491, w_046_1495, w_046_1496, w_046_1497, w_046_1498, w_046_1499, w_046_1500, w_046_1501, w_046_1502, w_046_1504, w_046_1505, w_046_1506, w_046_1507, w_046_1511, w_046_1512, w_046_1513, w_046_1515, w_046_1517, w_046_1519, w_046_1524, w_046_1525, w_046_1527, w_046_1528, w_046_1529, w_046_1530, w_046_1531, w_046_1532, w_046_1533, w_046_1534, w_046_1536, w_046_1537, w_046_1539, w_046_1540, w_046_1541, w_046_1542, w_046_1544, w_046_1546, w_046_1547, w_046_1548, w_046_1549, w_046_1550, w_046_1551, w_046_1553, w_046_1554, w_046_1556, w_046_1557, w_046_1558, w_046_1559, w_046_1561, w_046_1562, w_046_1564, w_046_1565, w_046_1567, w_046_1568, w_046_1569, w_046_1572, w_046_1573, w_046_1574, w_046_1575, w_046_1577, w_046_1580, w_046_1581, w_046_1582, w_046_1584, w_046_1585, w_046_1586, w_046_1587, w_046_1589, w_046_1591, w_046_1592, w_046_1594, w_046_1595, w_046_1596, w_046_1597, w_046_1598, w_046_1599, w_046_1601, w_046_1602, w_046_1603, w_046_1609, w_046_1610, w_046_1613, w_046_1614, w_046_1615, w_046_1616, w_046_1618, w_046_1619, w_046_1622, w_046_1623, w_046_1625, w_046_1627, w_046_1628, w_046_1631, w_046_1634, w_046_1635, w_046_1638, w_046_1640, w_046_1645, w_046_1647, w_046_1648, w_046_1649, w_046_1651, w_046_1652, w_046_1654, w_046_1655, w_046_1656, w_046_1661, w_046_1665, w_046_1666, w_046_1668, w_046_1669, w_046_1672, w_046_1673, w_046_1674, w_046_1675, w_046_1676, w_046_1679, w_046_1680, w_046_1681, w_046_1683, w_046_1692, w_046_1695, w_046_1696, w_046_1699, w_046_1700, w_046_1701, w_046_1703, w_046_1706, w_046_1709, w_046_1712, w_046_1714, w_046_1715, w_046_1718, w_046_1719, w_046_1721, w_046_1724, w_046_1725, w_046_1726, w_046_1730, w_046_1733, w_046_1736, w_046_1738, w_046_1739, w_046_1744, w_046_1746, w_046_1747, w_046_1750, w_046_1752, w_046_1753, w_046_1754, w_046_1762, w_046_1765, w_046_1766, w_046_1769, w_046_1770, w_046_1771, w_046_1772, w_046_1775, w_046_1777, w_046_1778, w_046_1784, w_046_1787, w_046_1789, w_046_1792, w_046_1793, w_046_1798, w_046_1803, w_046_1805, w_046_1806, w_046_1808, w_046_1809, w_046_1812, w_046_1814, w_046_1815, w_046_1819, w_046_1820, w_046_1821, w_046_1822, w_046_1823, w_046_1824, w_046_1827, w_046_1828, w_046_1829, w_046_1830, w_046_1833, w_046_1842, w_046_1843, w_046_1847, w_046_1848, w_046_1850, w_046_1851, w_046_1857, w_046_1859, w_046_1863, w_046_1865, w_046_1867, w_046_1868, w_046_1870, w_046_1871, w_046_1874, w_046_1878, w_046_1884, w_046_1885, w_046_1890, w_046_1891, w_046_1892, w_046_1893, w_046_1895, w_046_1899, w_046_1906, w_046_1907, w_046_1908, w_046_1909, w_046_1910, w_046_1912, w_046_1913, w_046_1915, w_046_1916, w_046_1918, w_046_1923, w_046_1931, w_046_1932, w_046_1933, w_046_1935, w_046_1940, w_046_1941, w_046_1942, w_046_1944, w_046_1945, w_046_1946, w_046_1947, w_046_1952, w_046_1954, w_046_1956, w_046_1958, w_046_1959, w_046_1960, w_046_1964, w_046_1965, w_046_1967, w_046_1969, w_046_1970, w_046_1972, w_046_1973, w_046_1976, w_046_1979, w_046_1980, w_046_1981, w_046_1983, w_046_1984, w_046_1986, w_046_1988, w_046_1989, w_046_1991, w_046_1992, w_046_1993, w_046_1994, w_046_1998, w_046_1999, w_046_2002, w_046_2003, w_046_2005, w_046_2006, w_046_2008, w_046_2009, w_046_2010, w_046_2012, w_046_2013, w_046_2014, w_046_2015, w_046_2017, w_046_2020, w_046_2023, w_046_2026, w_046_2027, w_046_2028, w_046_2030, w_046_2034, w_046_2035, w_046_2037, w_046_2041, w_046_2042, w_046_2045, w_046_2048, w_046_2050, w_046_2051, w_046_2052, w_046_2053, w_046_2054, w_046_2059, w_046_2064, w_046_2065, w_046_2066, w_046_2069, w_046_2071, w_046_2074, w_046_2076, w_046_2080, w_046_2081, w_046_2082, w_046_2086, w_046_2087, w_046_2089, w_046_2090, w_046_2091, w_046_2094, w_046_2095, w_046_2096, w_046_2098, w_046_2100, w_046_2101, w_046_2103, w_046_2105, w_046_2107, w_046_2110, w_046_2112, w_046_2117, w_046_2119, w_046_2120, w_046_2121, w_046_2122, w_046_2123, w_046_2127, w_046_2128, w_046_2129, w_046_2131, w_046_2133, w_046_2134, w_046_2135, w_046_2137, w_046_2139, w_046_2140, w_046_2141, w_046_2142, w_046_2145, w_046_2148, w_046_2152, w_046_2153, w_046_2154, w_046_2157, w_046_2158, w_046_2159, w_046_2160, w_046_2161, w_046_2164, w_046_2165, w_046_2168, w_046_2173, w_046_2175, w_046_2180, w_046_2182, w_046_2186, w_046_2187, w_046_2189, w_046_2190, w_046_2191, w_046_2194, w_046_2195, w_046_2196, w_046_2197, w_046_2198, w_046_2200, w_046_2201, w_046_2203, w_046_2205, w_046_2206, w_046_2207, w_046_2208, w_046_2210, w_046_2212, w_046_2215, w_046_2217, w_046_2219, w_046_2220, w_046_2221, w_046_2223, w_046_2224, w_046_2226, w_046_2228, w_046_2229, w_046_2230, w_046_2234, w_046_2235, w_046_2236, w_046_2239, w_046_2240, w_046_2241, w_046_2242, w_046_2243, w_046_2245, w_046_2246, w_046_2248, w_046_2249, w_046_2250, w_046_2251, w_046_2252, w_046_2253, w_046_2254, w_046_2260, w_046_2264, w_046_2265, w_046_2266, w_046_2267, w_046_2268, w_046_2269, w_046_2277, w_046_2280, w_046_2281, w_046_2289, w_046_2291, w_046_2292, w_046_2294, w_046_2296, w_046_2297, w_046_2298, w_046_2300, w_046_2303, w_046_2304, w_046_2306, w_046_2307, w_046_2309, w_046_2310, w_046_2312, w_046_2314, w_046_2315, w_046_2319, w_046_2321, w_046_2323, w_046_2324, w_046_2325, w_046_2327, w_046_2330, w_046_2331, w_046_2333, w_046_2335, w_046_2336, w_046_2337, w_046_2338, w_046_2339, w_046_2341, w_046_2342, w_046_2343, w_046_2344, w_046_2346, w_046_2347, w_046_2348, w_046_2349, w_046_2351, w_046_2352, w_046_2354, w_046_2357, w_046_2363, w_046_2364, w_046_2366, w_046_2368, w_046_2372, w_046_2374, w_046_2375, w_046_2376, w_046_2377, w_046_2384, w_046_2386, w_046_2388, w_046_2391, w_046_2392, w_046_2393, w_046_2396, w_046_2399, w_046_2400, w_046_2401, w_046_2402, w_046_2403, w_046_2404, w_046_2406, w_046_2411, w_046_2413, w_046_2414, w_046_2415, w_046_2417, w_046_2418, w_046_2419, w_046_2420, w_046_2422, w_046_2423, w_046_2425, w_046_2427, w_046_2428, w_046_2430, w_046_2431, w_046_2435, w_046_2436, w_046_2437, w_046_2440, w_046_2441, w_046_2443, w_046_2444, w_046_2445, w_046_2449, w_046_2451, w_046_2453, w_046_2455, w_046_2456, w_046_2457, w_046_2458, w_046_2459, w_046_2460, w_046_2461, w_046_2466, w_046_2467, w_046_2468, w_046_2473, w_046_2475, w_046_2476, w_046_2480, w_046_2481, w_046_2482, w_046_2484, w_046_2485, w_046_2486, w_046_2493, w_046_2494, w_046_2499, w_046_2503, w_046_2506, w_046_2507, w_046_2508, w_046_2509, w_046_2510, w_046_2511, w_046_2512, w_046_2514, w_046_2516, w_046_2518, w_046_2519, w_046_2520, w_046_2523, w_046_2529, w_046_2530, w_046_2532, w_046_2533, w_046_2534, w_046_2535, w_046_2537, w_046_2540, w_046_2541, w_046_2542, w_046_2543, w_046_2546, w_046_2547, w_046_2550, w_046_2552, w_046_2553, w_046_2556, w_046_2557, w_046_2558, w_046_2561, w_046_2563, w_046_2565, w_046_2566, w_046_2575, w_046_2577, w_046_2579, w_046_2580, w_046_2581, w_046_2582, w_046_2584, w_046_2587, w_046_2592, w_046_2596, w_046_2598, w_046_2599, w_046_2600, w_046_2602, w_046_2610, w_046_2612, w_046_2613, w_046_2614, w_046_2615, w_046_2616, w_046_2620, w_046_2624, w_046_2628, w_046_2630, w_046_2632, w_046_2634, w_046_2635, w_046_2637, w_046_2642, w_046_2643, w_046_2644, w_046_2645, w_046_2646, w_046_2647, w_046_2649, w_046_2650, w_046_2652, w_046_2654, w_046_2656, w_046_2657, w_046_2659, w_046_2661, w_046_2662, w_046_2665, w_046_2666, w_046_2667, w_046_2671, w_046_2672, w_046_2673, w_046_2674, w_046_2675, w_046_2677, w_046_2678, w_046_2680, w_046_2681, w_046_2683, w_046_2686, w_046_2689, w_046_2691, w_046_2692, w_046_2696, w_046_2698, w_046_2701, w_046_2702, w_046_2703, w_046_2705, w_046_2710, w_046_2712, w_046_2713, w_046_2714, w_046_2716, w_046_2718, w_046_2721, w_046_2722, w_046_2725, w_046_2726, w_046_2728, w_046_2731, w_046_2733, w_046_2734, w_046_2739, w_046_2742, w_046_2743, w_046_2745, w_046_2746, w_046_2747, w_046_2748, w_046_2753, w_046_2757, w_046_2761, w_046_2762, w_046_2764, w_046_2773, w_046_2774, w_046_2775, w_046_2776, w_046_2780, w_046_2781, w_046_2782, w_046_2786, w_046_2787, w_046_2792, w_046_2795, w_046_2797, w_046_2798, w_046_2801, w_046_2803, w_046_2805, w_046_2806, w_046_2808, w_046_2809, w_046_2812, w_046_2813, w_046_2815, w_046_2816, w_046_2817, w_046_2818, w_046_2819, w_046_2820, w_046_2826, w_046_2827, w_046_2830, w_046_2832, w_046_2834, w_046_2836, w_046_2837, w_046_2838, w_046_2840, w_046_2842, w_046_2845, w_046_2846, w_046_2847, w_046_2849, w_046_2850, w_046_2851, w_046_2855, w_046_2856, w_046_2857, w_046_2858, w_046_2864, w_046_2866, w_046_2867, w_046_2868, w_046_2871, w_046_2873, w_046_2876, w_046_2879, w_046_2880, w_046_2884, w_046_2886, w_046_2887, w_046_2888, w_046_2889, w_046_2890, w_046_2892, w_046_2895, w_046_2897, w_046_2898, w_046_2899, w_046_2900, w_046_2902, w_046_2903, w_046_2904, w_046_2905, w_046_2906, w_046_2907, w_046_2909, w_046_2914, w_046_2915, w_046_2921, w_046_2923, w_046_2924, w_046_2925, w_046_2926, w_046_2928, w_046_2930, w_046_2932, w_046_2933, w_046_2934, w_046_2936, w_046_2937, w_046_2938, w_046_2939, w_046_2940, w_046_2941, w_046_2942, w_046_2943, w_046_2944, w_046_2946, w_046_2947, w_046_2953, w_046_2954, w_046_2956, w_046_2957, w_046_2958, w_046_2960, w_046_2963, w_046_2964, w_046_2966, w_046_2968, w_046_2969, w_046_2972, w_046_2973, w_046_2980, w_046_2982, w_046_2984, w_046_2986, w_046_2987, w_046_2988, w_046_2990, w_046_2991, w_046_2992, w_046_2993, w_046_2997, w_046_2999, w_046_3000, w_046_3002, w_046_3003, w_046_3004, w_046_3008, w_046_3009, w_046_3013, w_046_3016, w_046_3017, w_046_3018, w_046_3021, w_046_3023, w_046_3025, w_046_3027, w_046_3029, w_046_3033, w_046_3036, w_046_3040, w_046_3043, w_046_3044, w_046_3045, w_046_3050, w_046_3051, w_046_3053, w_046_3054, w_046_3056, w_046_3060, w_046_3061, w_046_3062, w_046_3063, w_046_3066, w_046_3067, w_046_3072, w_046_3073, w_046_3074, w_046_3076, w_046_3077, w_046_3078, w_046_3079, w_046_3081, w_046_3082, w_046_3085, w_046_3086, w_046_3092, w_046_3093, w_046_3094, w_046_3095, w_046_3097, w_046_3099, w_046_3100, w_046_3103, w_046_3105, w_046_3107, w_046_3110, w_046_3112, w_046_3117, w_046_3118, w_046_3119, w_046_3121, w_046_3122, w_046_3127, w_046_3129, w_046_3130, w_046_3132, w_046_3134, w_046_3136, w_046_3138, w_046_3142, w_046_3144, w_046_3145, w_046_3147, w_046_3148, w_046_3152, w_046_3154, w_046_3157, w_046_3158, w_046_3160, w_046_3161, w_046_3166, w_046_3167, w_046_3168, w_046_3169, w_046_3170, w_046_3172, w_046_3173, w_046_3176, w_046_3177, w_046_3178, w_046_3179, w_046_3180, w_046_3182, w_046_3186, w_046_3187, w_046_3189, w_046_3191, w_046_3192, w_046_3196, w_046_3201, w_046_3202, w_046_3209, w_046_3210, w_046_3211, w_046_3212, w_046_3213, w_046_3216, w_046_3220, w_046_3222, w_046_3223, w_046_3224, w_046_3226, w_046_3228, w_046_3229, w_046_3230, w_046_3234, w_046_3235, w_046_3237, w_046_3239, w_046_3240, w_046_3244, w_046_3245, w_046_3248, w_046_3249, w_046_3250, w_046_3252, w_046_3254, w_046_3259, w_046_3262, w_046_3264, w_046_3268, w_046_3270, w_046_3272, w_046_3273, w_046_3277, w_046_3278, w_046_3279, w_046_3280, w_046_3281, w_046_3282, w_046_3285, w_046_3287, w_046_3288, w_046_3289, w_046_3291, w_046_3292, w_046_3294, w_046_3295, w_046_3296, w_046_3297, w_046_3298, w_046_3300, w_046_3304, w_046_3306, w_046_3307, w_046_3308, w_046_3315, w_046_3316, w_046_3317, w_046_3319, w_046_3320, w_046_3321, w_046_3322, w_046_3325, w_046_3327, w_046_3328, w_046_3329, w_046_3334, w_046_3335, w_046_3336, w_046_3339, w_046_3341, w_046_3342, w_046_3343, w_046_3345, w_046_3348, w_046_3352, w_046_3353, w_046_3354, w_046_3356, w_046_3357, w_046_3358, w_046_3360, w_046_3361, w_046_3362, w_046_3363, w_046_3365, w_046_3372, w_046_3378, w_046_3379, w_046_3380, w_046_3382;
  wire w_047_000, w_047_001, w_047_002, w_047_003, w_047_005, w_047_006, w_047_008, w_047_009, w_047_010, w_047_011, w_047_012, w_047_013, w_047_014, w_047_015, w_047_016, w_047_017, w_047_018, w_047_019, w_047_020, w_047_021, w_047_022, w_047_023, w_047_025, w_047_026, w_047_027, w_047_028, w_047_029, w_047_030, w_047_031, w_047_032, w_047_034, w_047_035, w_047_036, w_047_037, w_047_039, w_047_040, w_047_041, w_047_042, w_047_043, w_047_044, w_047_045, w_047_046, w_047_047, w_047_048, w_047_049, w_047_050, w_047_051, w_047_052, w_047_053, w_047_054, w_047_055, w_047_056, w_047_057, w_047_058, w_047_059, w_047_060, w_047_061, w_047_062, w_047_063, w_047_064, w_047_065, w_047_066, w_047_067, w_047_068, w_047_069, w_047_070, w_047_071, w_047_072, w_047_073, w_047_074, w_047_075, w_047_076, w_047_077, w_047_078, w_047_079, w_047_080, w_047_081, w_047_082, w_047_083, w_047_084, w_047_085, w_047_086, w_047_087, w_047_088, w_047_089, w_047_090, w_047_091, w_047_092, w_047_093, w_047_094, w_047_095, w_047_096, w_047_098, w_047_099, w_047_100, w_047_101, w_047_102, w_047_103, w_047_104, w_047_105, w_047_106, w_047_107, w_047_108, w_047_109, w_047_110, w_047_111, w_047_112, w_047_113, w_047_114, w_047_115, w_047_116, w_047_117, w_047_118, w_047_119, w_047_120, w_047_121, w_047_122, w_047_124, w_047_125, w_047_126, w_047_127, w_047_128, w_047_129, w_047_130, w_047_131, w_047_132, w_047_133, w_047_134, w_047_135, w_047_136, w_047_137, w_047_138, w_047_139, w_047_140, w_047_141, w_047_142, w_047_143, w_047_144, w_047_145, w_047_146, w_047_147, w_047_149, w_047_150, w_047_151, w_047_152, w_047_153, w_047_154, w_047_155, w_047_156, w_047_157, w_047_158, w_047_159, w_047_160, w_047_161, w_047_162, w_047_163, w_047_164, w_047_165, w_047_166, w_047_167, w_047_168, w_047_169, w_047_171, w_047_174, w_047_175, w_047_176, w_047_177, w_047_178, w_047_179, w_047_180, w_047_181, w_047_182, w_047_183, w_047_185, w_047_186, w_047_187, w_047_188, w_047_190, w_047_191, w_047_192, w_047_193, w_047_194, w_047_195, w_047_196, w_047_197, w_047_198, w_047_199, w_047_200, w_047_201, w_047_202, w_047_203, w_047_204, w_047_205, w_047_206, w_047_207, w_047_208, w_047_209, w_047_210, w_047_211, w_047_212, w_047_213, w_047_214, w_047_216, w_047_217, w_047_218, w_047_219, w_047_221, w_047_222, w_047_223, w_047_224, w_047_225, w_047_226, w_047_227, w_047_230, w_047_231, w_047_232, w_047_233, w_047_234, w_047_235, w_047_236, w_047_237, w_047_238, w_047_239, w_047_240, w_047_241, w_047_243, w_047_244, w_047_245, w_047_246, w_047_247, w_047_248, w_047_249, w_047_250, w_047_251, w_047_252, w_047_253, w_047_254, w_047_255, w_047_256, w_047_257, w_047_258, w_047_259, w_047_260, w_047_261, w_047_262, w_047_263, w_047_264, w_047_265, w_047_266, w_047_267, w_047_268, w_047_269, w_047_270, w_047_271, w_047_272, w_047_273, w_047_274, w_047_275, w_047_276, w_047_277, w_047_278, w_047_279, w_047_280, w_047_281, w_047_282, w_047_283, w_047_284, w_047_285, w_047_286, w_047_287, w_047_288, w_047_289, w_047_290, w_047_291, w_047_292, w_047_294, w_047_296, w_047_297, w_047_298, w_047_299, w_047_300, w_047_301, w_047_302, w_047_304, w_047_305, w_047_306, w_047_307, w_047_308, w_047_309, w_047_310, w_047_311, w_047_312, w_047_313, w_047_314, w_047_315, w_047_316, w_047_317, w_047_318, w_047_319, w_047_320, w_047_321, w_047_323, w_047_324, w_047_325, w_047_326, w_047_327, w_047_328, w_047_329, w_047_330, w_047_331, w_047_332, w_047_333, w_047_334, w_047_335, w_047_336, w_047_337, w_047_338, w_047_339, w_047_340, w_047_341, w_047_342, w_047_343, w_047_344, w_047_345, w_047_346, w_047_347, w_047_348, w_047_349, w_047_350, w_047_351, w_047_352, w_047_353, w_047_354, w_047_355, w_047_356, w_047_357, w_047_358, w_047_359, w_047_360, w_047_361, w_047_362, w_047_364, w_047_365, w_047_367, w_047_368, w_047_370, w_047_371, w_047_372, w_047_373, w_047_374, w_047_376, w_047_377, w_047_378, w_047_380, w_047_381, w_047_382, w_047_383, w_047_384, w_047_385, w_047_386, w_047_387, w_047_388, w_047_389, w_047_390, w_047_391, w_047_393, w_047_394, w_047_395, w_047_396, w_047_397, w_047_398, w_047_399, w_047_400, w_047_401, w_047_402, w_047_403, w_047_404, w_047_405, w_047_406, w_047_407, w_047_408, w_047_409, w_047_410, w_047_411, w_047_412, w_047_413, w_047_414, w_047_415, w_047_416, w_047_417, w_047_418, w_047_419, w_047_420, w_047_421, w_047_422, w_047_423, w_047_426, w_047_427, w_047_428, w_047_429, w_047_430, w_047_431, w_047_432, w_047_433, w_047_434, w_047_435, w_047_436, w_047_437, w_047_438, w_047_439, w_047_441, w_047_442, w_047_443, w_047_444, w_047_445, w_047_446, w_047_448, w_047_449, w_047_450, w_047_451, w_047_452, w_047_453, w_047_454, w_047_455, w_047_456, w_047_457, w_047_458, w_047_459, w_047_460, w_047_461, w_047_462, w_047_463, w_047_464, w_047_465, w_047_466, w_047_467, w_047_468, w_047_469, w_047_470, w_047_471, w_047_472, w_047_474, w_047_475, w_047_476, w_047_478, w_047_479, w_047_480, w_047_481, w_047_482, w_047_483, w_047_484, w_047_485, w_047_486, w_047_487, w_047_488, w_047_489, w_047_490, w_047_491, w_047_492, w_047_493, w_047_494, w_047_495, w_047_496, w_047_497, w_047_498, w_047_499, w_047_500, w_047_501, w_047_502, w_047_503, w_047_504, w_047_505, w_047_506, w_047_507, w_047_509, w_047_510, w_047_511, w_047_512, w_047_513, w_047_514, w_047_515, w_047_516, w_047_517, w_047_518, w_047_519, w_047_520, w_047_521, w_047_522, w_047_523, w_047_524, w_047_525, w_047_526, w_047_527, w_047_528, w_047_530, w_047_531, w_047_532, w_047_533, w_047_535, w_047_536, w_047_537, w_047_538, w_047_539, w_047_540, w_047_541, w_047_542, w_047_543, w_047_544, w_047_545, w_047_547, w_047_548, w_047_549, w_047_550, w_047_551, w_047_552, w_047_554, w_047_555, w_047_556, w_047_557, w_047_559, w_047_560, w_047_561, w_047_562, w_047_563, w_047_564, w_047_565, w_047_566, w_047_567, w_047_568, w_047_569, w_047_570, w_047_571, w_047_573, w_047_574, w_047_575, w_047_576, w_047_577, w_047_578, w_047_579, w_047_580, w_047_581, w_047_582, w_047_583, w_047_584, w_047_585, w_047_586, w_047_587, w_047_589, w_047_591, w_047_592, w_047_593, w_047_594, w_047_597, w_047_598, w_047_599, w_047_600, w_047_601, w_047_602, w_047_604, w_047_606, w_047_608, w_047_609, w_047_610, w_047_611, w_047_612, w_047_613, w_047_614, w_047_615, w_047_617, w_047_618, w_047_619, w_047_620, w_047_621, w_047_622, w_047_623, w_047_624, w_047_625, w_047_626, w_047_627, w_047_628, w_047_629, w_047_630, w_047_631, w_047_632, w_047_633, w_047_634, w_047_636, w_047_637, w_047_638, w_047_639, w_047_640, w_047_641, w_047_642, w_047_646, w_047_647, w_047_648, w_047_649, w_047_650, w_047_652, w_047_653, w_047_655, w_047_656, w_047_657, w_047_658, w_047_659, w_047_660, w_047_661, w_047_662, w_047_663, w_047_664, w_047_665, w_047_666, w_047_669, w_047_670, w_047_671, w_047_672, w_047_673, w_047_674, w_047_675, w_047_676, w_047_678, w_047_679, w_047_680, w_047_681, w_047_682, w_047_683, w_047_684, w_047_685, w_047_687, w_047_689, w_047_690, w_047_691, w_047_692, w_047_693, w_047_694, w_047_695, w_047_696, w_047_697, w_047_699, w_047_700, w_047_701, w_047_702, w_047_703, w_047_704, w_047_705, w_047_706, w_047_707, w_047_709, w_047_710, w_047_711, w_047_712, w_047_713, w_047_714, w_047_715, w_047_716, w_047_718, w_047_719, w_047_720, w_047_721, w_047_722, w_047_724, w_047_726, w_047_727, w_047_728, w_047_729, w_047_730, w_047_731, w_047_732, w_047_734, w_047_735, w_047_736, w_047_737, w_047_738, w_047_739, w_047_740, w_047_741, w_047_742, w_047_743, w_047_744, w_047_745, w_047_746, w_047_747, w_047_748, w_047_749, w_047_750, w_047_752, w_047_753, w_047_754, w_047_755, w_047_756, w_047_758, w_047_759, w_047_760, w_047_761, w_047_763, w_047_764, w_047_766, w_047_768, w_047_769, w_047_770, w_047_771, w_047_772, w_047_773, w_047_774, w_047_775, w_047_776, w_047_777, w_047_778, w_047_779, w_047_780, w_047_781, w_047_782, w_047_783, w_047_784, w_047_785, w_047_786, w_047_788, w_047_789, w_047_790, w_047_791, w_047_792, w_047_793, w_047_794, w_047_795, w_047_797, w_047_799, w_047_801, w_047_802, w_047_803, w_047_804, w_047_805, w_047_807, w_047_808, w_047_809, w_047_810, w_047_811, w_047_812, w_047_813, w_047_815, w_047_816, w_047_817, w_047_818, w_047_819, w_047_820, w_047_821, w_047_822, w_047_823, w_047_824, w_047_825, w_047_826, w_047_827, w_047_828, w_047_829, w_047_830, w_047_831, w_047_832, w_047_833, w_047_834, w_047_835, w_047_836, w_047_837, w_047_838, w_047_839, w_047_840, w_047_841, w_047_842, w_047_844, w_047_845, w_047_846, w_047_847, w_047_848, w_047_849, w_047_850, w_047_851, w_047_852, w_047_853, w_047_854, w_047_855, w_047_856, w_047_857, w_047_858, w_047_860, w_047_861, w_047_862, w_047_863, w_047_864, w_047_865, w_047_866, w_047_867, w_047_868, w_047_869, w_047_870, w_047_871, w_047_872, w_047_873, w_047_874, w_047_875, w_047_876, w_047_877, w_047_878, w_047_879, w_047_880, w_047_881, w_047_882, w_047_883, w_047_884, w_047_885, w_047_886, w_047_887, w_047_888, w_047_889, w_047_890, w_047_891, w_047_892, w_047_893, w_047_894, w_047_895, w_047_896, w_047_897, w_047_898, w_047_900, w_047_902, w_047_903, w_047_904, w_047_905, w_047_906, w_047_907, w_047_910, w_047_911, w_047_912, w_047_913, w_047_914, w_047_915, w_047_916, w_047_917, w_047_918, w_047_919, w_047_920, w_047_921, w_047_922, w_047_923, w_047_924, w_047_925, w_047_926, w_047_927, w_047_928, w_047_929, w_047_930, w_047_931, w_047_932, w_047_934, w_047_935, w_047_936, w_047_937, w_047_939, w_047_940, w_047_941, w_047_942, w_047_944, w_047_945, w_047_947, w_047_948, w_047_949, w_047_950, w_047_951, w_047_953, w_047_954, w_047_955, w_047_956, w_047_957, w_047_958, w_047_959, w_047_960, w_047_961, w_047_962, w_047_963, w_047_964, w_047_965, w_047_966, w_047_967, w_047_968, w_047_969, w_047_970, w_047_971, w_047_972, w_047_973, w_047_974, w_047_975, w_047_976, w_047_977, w_047_978, w_047_979, w_047_980, w_047_981, w_047_982, w_047_983, w_047_984, w_047_985, w_047_986, w_047_987, w_047_988, w_047_989, w_047_991, w_047_992, w_047_993, w_047_994, w_047_995, w_047_996, w_047_997, w_047_998, w_047_999, w_047_1000, w_047_1001, w_047_1002, w_047_1003, w_047_1004, w_047_1006, w_047_1007, w_047_1008, w_047_1009, w_047_1010, w_047_1011, w_047_1012, w_047_1013, w_047_1014, w_047_1015, w_047_1016, w_047_1017, w_047_1018, w_047_1019, w_047_1020, w_047_1021, w_047_1022, w_047_1024, w_047_1025, w_047_1027, w_047_1028, w_047_1029, w_047_1031, w_047_1032, w_047_1033, w_047_1034, w_047_1035, w_047_1036, w_047_1037, w_047_1042, w_047_1043, w_047_1045, w_047_1046, w_047_1047, w_047_1048, w_047_1049, w_047_1050, w_047_1051, w_047_1052, w_047_1053, w_047_1054, w_047_1055, w_047_1056, w_047_1057, w_047_1059, w_047_1060, w_047_1061, w_047_1062, w_047_1063, w_047_1064, w_047_1065, w_047_1066, w_047_1067, w_047_1068, w_047_1069, w_047_1070, w_047_1071, w_047_1072, w_047_1073, w_047_1074, w_047_1075, w_047_1076, w_047_1077, w_047_1078, w_047_1079, w_047_1080, w_047_1082, w_047_1084, w_047_1086, w_047_1087, w_047_1088, w_047_1089, w_047_1090, w_047_1091, w_047_1092, w_047_1093, w_047_1094, w_047_1095, w_047_1096, w_047_1097, w_047_1098, w_047_1099, w_047_1100, w_047_1101, w_047_1102, w_047_1103, w_047_1104, w_047_1105, w_047_1106, w_047_1107, w_047_1108, w_047_1109, w_047_1110, w_047_1111, w_047_1112, w_047_1113, w_047_1114, w_047_1115, w_047_1116, w_047_1118, w_047_1121, w_047_1122, w_047_1124, w_047_1125, w_047_1126, w_047_1127, w_047_1128, w_047_1130, w_047_1131, w_047_1132, w_047_1133, w_047_1134, w_047_1135, w_047_1136, w_047_1138, w_047_1139, w_047_1140, w_047_1141, w_047_1142, w_047_1143, w_047_1144, w_047_1145, w_047_1146, w_047_1147, w_047_1148, w_047_1149, w_047_1151, w_047_1152, w_047_1154, w_047_1155, w_047_1156, w_047_1157, w_047_1158, w_047_1159, w_047_1160, w_047_1161, w_047_1162, w_047_1163, w_047_1164, w_047_1165, w_047_1166, w_047_1167, w_047_1168, w_047_1169, w_047_1170, w_047_1171, w_047_1172, w_047_1174, w_047_1175, w_047_1176, w_047_1177, w_047_1178, w_047_1180, w_047_1181, w_047_1183, w_047_1184, w_047_1185, w_047_1186, w_047_1187, w_047_1188, w_047_1189, w_047_1190, w_047_1191, w_047_1192, w_047_1193, w_047_1194, w_047_1195, w_047_1197, w_047_1198, w_047_1199, w_047_1200, w_047_1201, w_047_1202, w_047_1203, w_047_1204, w_047_1206, w_047_1207, w_047_1208, w_047_1210, w_047_1211, w_047_1213, w_047_1214, w_047_1215, w_047_1217, w_047_1218, w_047_1219, w_047_1221, w_047_1222, w_047_1224, w_047_1225, w_047_1226, w_047_1227, w_047_1229, w_047_1231, w_047_1232, w_047_1234, w_047_1235, w_047_1236, w_047_1237, w_047_1238, w_047_1241, w_047_1242, w_047_1243, w_047_1244, w_047_1246, w_047_1247, w_047_1248, w_047_1249, w_047_1250, w_047_1251, w_047_1252, w_047_1253, w_047_1254, w_047_1256, w_047_1257, w_047_1258, w_047_1259, w_047_1260, w_047_1261, w_047_1262, w_047_1263, w_047_1264, w_047_1265, w_047_1266, w_047_1267, w_047_1268, w_047_1269, w_047_1270, w_047_1271, w_047_1272, w_047_1273, w_047_1274, w_047_1275, w_047_1276, w_047_1278, w_047_1279, w_047_1281, w_047_1282, w_047_1283, w_047_1285, w_047_1286, w_047_1287, w_047_1288, w_047_1289, w_047_1290, w_047_1291, w_047_1292, w_047_1293, w_047_1295, w_047_1296, w_047_1297, w_047_1298, w_047_1300, w_047_1302, w_047_1303, w_047_1305, w_047_1307, w_047_1308, w_047_1309, w_047_1310, w_047_1311, w_047_1312, w_047_1313, w_047_1314, w_047_1315, w_047_1316, w_047_1317, w_047_1318, w_047_1319, w_047_1320, w_047_1321, w_047_1322, w_047_1323, w_047_1324, w_047_1326, w_047_1328, w_047_1329, w_047_1330, w_047_1331, w_047_1333, w_047_1334, w_047_1335, w_047_1337, w_047_1338, w_047_1339, w_047_1340, w_047_1341, w_047_1342, w_047_1343, w_047_1345, w_047_1346, w_047_1347, w_047_1348, w_047_1349, w_047_1350, w_047_1351, w_047_1352, w_047_1353, w_047_1354, w_047_1355, w_047_1356, w_047_1357, w_047_1358, w_047_1359, w_047_1360, w_047_1362, w_047_1363, w_047_1364, w_047_1365, w_047_1366, w_047_1368, w_047_1369, w_047_1370, w_047_1371, w_047_1372, w_047_1373, w_047_1374, w_047_1375, w_047_1376, w_047_1377, w_047_1378, w_047_1379, w_047_1380, w_047_1381, w_047_1382, w_047_1383, w_047_1384, w_047_1385, w_047_1386, w_047_1387, w_047_1388, w_047_1389, w_047_1390, w_047_1391, w_047_1392, w_047_1393, w_047_1394, w_047_1395, w_047_1396, w_047_1398, w_047_1399, w_047_1400, w_047_1401, w_047_1402, w_047_1403, w_047_1404, w_047_1405, w_047_1406, w_047_1407, w_047_1408, w_047_1409, w_047_1410, w_047_1411, w_047_1412, w_047_1413, w_047_1416, w_047_1417, w_047_1418, w_047_1419, w_047_1420, w_047_1421, w_047_1422, w_047_1423, w_047_1424, w_047_1425, w_047_1426, w_047_1427, w_047_1428, w_047_1429, w_047_1430, w_047_1431, w_047_1432, w_047_1433, w_047_1434, w_047_1435, w_047_1437, w_047_1438, w_047_1439, w_047_1440, w_047_1441, w_047_1443, w_047_1444, w_047_1445, w_047_1446, w_047_1447, w_047_1448, w_047_1449, w_047_1450, w_047_1451, w_047_1453, w_047_1455, w_047_1456, w_047_1457, w_047_1459, w_047_1460, w_047_1461, w_047_1462, w_047_1463, w_047_1464, w_047_1465, w_047_1466, w_047_1467, w_047_1469, w_047_1470, w_047_1471, w_047_1472, w_047_1473, w_047_1474, w_047_1476, w_047_1477, w_047_1478, w_047_1479, w_047_1480, w_047_1481, w_047_1482, w_047_1483, w_047_1484, w_047_1485, w_047_1486, w_047_1488, w_047_1490, w_047_1491, w_047_1492, w_047_1493, w_047_1494, w_047_1496;
  wire w_048_001, w_048_002, w_048_003, w_048_004, w_048_006, w_048_007, w_048_008, w_048_009, w_048_010, w_048_011, w_048_012, w_048_013, w_048_014, w_048_015, w_048_017, w_048_019, w_048_021, w_048_022, w_048_023, w_048_024, w_048_025, w_048_027, w_048_028, w_048_029, w_048_030, w_048_031, w_048_032, w_048_033, w_048_036, w_048_037, w_048_038, w_048_039, w_048_040, w_048_041, w_048_042, w_048_043, w_048_044, w_048_045, w_048_046, w_048_047, w_048_049, w_048_050, w_048_052, w_048_053, w_048_054, w_048_055, w_048_056, w_048_057, w_048_059, w_048_060, w_048_061, w_048_062, w_048_063, w_048_067, w_048_069, w_048_070, w_048_071, w_048_073, w_048_074, w_048_075, w_048_076, w_048_078, w_048_079, w_048_080, w_048_081, w_048_082, w_048_083, w_048_084, w_048_085, w_048_086, w_048_089, w_048_090, w_048_091, w_048_092, w_048_093, w_048_095, w_048_096, w_048_097, w_048_098, w_048_099, w_048_103, w_048_104, w_048_105, w_048_106, w_048_107, w_048_108, w_048_110, w_048_111, w_048_112, w_048_114, w_048_115, w_048_116, w_048_117, w_048_118, w_048_119, w_048_120, w_048_121, w_048_122, w_048_123, w_048_124, w_048_126, w_048_127, w_048_128, w_048_129, w_048_131, w_048_132, w_048_133, w_048_134, w_048_135, w_048_137, w_048_138, w_048_139, w_048_141, w_048_144, w_048_145, w_048_146, w_048_147, w_048_148, w_048_149, w_048_150, w_048_151, w_048_152, w_048_153, w_048_154, w_048_155, w_048_156, w_048_158, w_048_160, w_048_161, w_048_162, w_048_163, w_048_164, w_048_166, w_048_167, w_048_168, w_048_169, w_048_170, w_048_172, w_048_173, w_048_174, w_048_176, w_048_177, w_048_179, w_048_180, w_048_181, w_048_182, w_048_183, w_048_185, w_048_186, w_048_187, w_048_189, w_048_190, w_048_191, w_048_192, w_048_195, w_048_197, w_048_198, w_048_199, w_048_200, w_048_202, w_048_203, w_048_204, w_048_206, w_048_209, w_048_210, w_048_211, w_048_212, w_048_213, w_048_214, w_048_216, w_048_217, w_048_219, w_048_221, w_048_223, w_048_224, w_048_225, w_048_226, w_048_227, w_048_228, w_048_229, w_048_230, w_048_231, w_048_232, w_048_233, w_048_237, w_048_238, w_048_239, w_048_240, w_048_241, w_048_242, w_048_243, w_048_244, w_048_246, w_048_247, w_048_248, w_048_250, w_048_251, w_048_253, w_048_255, w_048_256, w_048_258, w_048_259, w_048_262, w_048_263, w_048_265, w_048_267, w_048_269, w_048_270, w_048_271, w_048_273, w_048_274, w_048_275, w_048_276, w_048_278, w_048_279, w_048_280, w_048_281, w_048_282, w_048_283, w_048_284, w_048_285, w_048_287, w_048_289, w_048_290, w_048_291, w_048_292, w_048_294, w_048_296, w_048_298, w_048_299, w_048_300, w_048_304, w_048_305, w_048_306, w_048_307, w_048_308, w_048_309, w_048_310, w_048_312, w_048_313, w_048_314, w_048_315, w_048_317, w_048_318, w_048_319, w_048_321, w_048_322, w_048_323, w_048_324, w_048_325, w_048_326, w_048_327, w_048_328, w_048_330, w_048_331, w_048_332, w_048_334, w_048_335, w_048_336, w_048_339, w_048_341, w_048_342, w_048_343, w_048_344, w_048_347, w_048_348, w_048_349, w_048_350, w_048_351, w_048_353, w_048_354, w_048_355, w_048_356, w_048_357, w_048_358, w_048_359, w_048_361, w_048_362, w_048_363, w_048_364, w_048_365, w_048_366, w_048_367, w_048_371, w_048_374, w_048_375, w_048_377, w_048_378, w_048_380, w_048_381, w_048_382, w_048_385, w_048_390, w_048_391, w_048_392, w_048_393, w_048_395, w_048_397, w_048_398, w_048_399, w_048_400, w_048_401, w_048_402, w_048_403, w_048_406, w_048_407, w_048_408, w_048_409, w_048_410, w_048_411, w_048_413, w_048_414, w_048_415, w_048_416, w_048_417, w_048_418, w_048_419, w_048_420, w_048_422, w_048_425, w_048_427, w_048_428, w_048_429, w_048_430, w_048_432, w_048_436, w_048_438, w_048_443, w_048_444, w_048_450, w_048_452, w_048_454, w_048_455, w_048_460, w_048_461, w_048_463, w_048_465, w_048_466, w_048_467, w_048_469, w_048_475, w_048_479, w_048_480, w_048_483, w_048_484, w_048_488, w_048_489, w_048_490, w_048_491, w_048_492, w_048_493, w_048_496, w_048_498, w_048_500, w_048_506, w_048_511, w_048_512, w_048_513, w_048_515, w_048_516, w_048_518, w_048_519, w_048_520, w_048_521, w_048_523, w_048_526, w_048_528, w_048_531, w_048_533, w_048_535, w_048_536, w_048_537, w_048_538, w_048_542, w_048_546, w_048_551, w_048_553, w_048_554, w_048_555, w_048_557, w_048_561, w_048_563, w_048_566, w_048_567, w_048_569, w_048_573, w_048_575, w_048_577, w_048_580, w_048_581, w_048_582, w_048_584, w_048_587, w_048_588, w_048_590, w_048_592, w_048_593, w_048_594, w_048_595, w_048_596, w_048_599, w_048_601, w_048_603, w_048_604, w_048_606, w_048_608, w_048_609, w_048_613, w_048_615, w_048_619, w_048_620, w_048_621, w_048_623, w_048_624, w_048_627, w_048_632, w_048_633, w_048_636, w_048_637, w_048_639, w_048_640, w_048_641, w_048_643, w_048_644, w_048_645, w_048_651, w_048_652, w_048_653, w_048_659, w_048_660, w_048_661, w_048_663, w_048_664, w_048_666, w_048_667, w_048_669, w_048_671, w_048_676, w_048_677, w_048_678, w_048_679, w_048_680, w_048_681, w_048_684, w_048_687, w_048_690, w_048_692, w_048_693, w_048_698, w_048_700, w_048_705, w_048_706, w_048_709, w_048_710, w_048_711, w_048_714, w_048_715, w_048_716, w_048_718, w_048_719, w_048_720, w_048_722, w_048_723, w_048_724, w_048_725, w_048_728, w_048_729, w_048_732, w_048_734, w_048_735, w_048_736, w_048_738, w_048_739, w_048_740, w_048_747, w_048_748, w_048_750, w_048_752, w_048_754, w_048_755, w_048_756, w_048_758, w_048_759, w_048_765, w_048_768, w_048_771, w_048_772, w_048_776, w_048_779, w_048_781, w_048_782, w_048_785, w_048_788, w_048_789, w_048_790, w_048_792, w_048_796, w_048_797, w_048_798, w_048_799, w_048_800, w_048_801, w_048_802, w_048_804, w_048_805, w_048_806, w_048_808, w_048_810, w_048_812, w_048_813, w_048_815, w_048_819, w_048_821, w_048_822, w_048_824, w_048_825, w_048_831, w_048_832, w_048_834, w_048_838, w_048_841, w_048_842, w_048_843, w_048_846, w_048_847, w_048_849, w_048_851, w_048_852, w_048_853, w_048_854, w_048_855, w_048_856, w_048_858, w_048_860, w_048_864, w_048_868, w_048_869, w_048_870, w_048_871, w_048_873, w_048_877, w_048_879, w_048_881, w_048_883, w_048_884, w_048_885, w_048_886, w_048_889, w_048_891, w_048_892, w_048_893, w_048_895, w_048_899, w_048_902, w_048_903, w_048_905, w_048_910, w_048_911, w_048_912, w_048_914, w_048_915, w_048_916, w_048_917, w_048_918, w_048_920, w_048_922, w_048_926, w_048_927, w_048_929, w_048_930, w_048_936, w_048_939, w_048_940, w_048_941, w_048_942, w_048_944, w_048_946, w_048_950, w_048_951, w_048_954, w_048_958, w_048_960, w_048_962, w_048_965, w_048_966, w_048_967, w_048_968, w_048_969, w_048_971, w_048_972, w_048_973, w_048_974, w_048_976, w_048_978, w_048_979, w_048_981, w_048_982, w_048_985, w_048_986, w_048_988, w_048_989, w_048_990, w_048_992, w_048_993, w_048_994, w_048_995, w_048_996, w_048_999, w_048_1002, w_048_1003, w_048_1006, w_048_1008, w_048_1012, w_048_1013, w_048_1014, w_048_1015, w_048_1016, w_048_1021, w_048_1022, w_048_1023, w_048_1024, w_048_1025, w_048_1031, w_048_1032, w_048_1034, w_048_1041, w_048_1042, w_048_1045, w_048_1046, w_048_1048, w_048_1049, w_048_1050, w_048_1052, w_048_1053, w_048_1055, w_048_1059, w_048_1060, w_048_1065, w_048_1066, w_048_1067, w_048_1068, w_048_1072, w_048_1075, w_048_1077, w_048_1078, w_048_1080, w_048_1085, w_048_1086, w_048_1087, w_048_1088, w_048_1089, w_048_1091, w_048_1093, w_048_1094, w_048_1095, w_048_1096, w_048_1099, w_048_1101, w_048_1103, w_048_1104, w_048_1106, w_048_1107, w_048_1108, w_048_1110, w_048_1111, w_048_1112, w_048_1113, w_048_1115, w_048_1116, w_048_1118, w_048_1120, w_048_1121, w_048_1122, w_048_1128, w_048_1129, w_048_1131, w_048_1132, w_048_1134, w_048_1135, w_048_1139, w_048_1140, w_048_1143, w_048_1145, w_048_1146, w_048_1148, w_048_1149, w_048_1150, w_048_1153, w_048_1154, w_048_1156, w_048_1158, w_048_1160, w_048_1162, w_048_1164, w_048_1165, w_048_1167, w_048_1168, w_048_1169, w_048_1172, w_048_1176, w_048_1178, w_048_1182, w_048_1187, w_048_1188, w_048_1189, w_048_1190, w_048_1191, w_048_1194, w_048_1196, w_048_1205, w_048_1206, w_048_1209, w_048_1210, w_048_1211, w_048_1212, w_048_1219, w_048_1221, w_048_1226, w_048_1227, w_048_1228, w_048_1230, w_048_1233, w_048_1235, w_048_1236, w_048_1239, w_048_1242, w_048_1245, w_048_1246, w_048_1247, w_048_1249, w_048_1250, w_048_1252, w_048_1254, w_048_1255, w_048_1256, w_048_1257, w_048_1259, w_048_1261, w_048_1262, w_048_1264, w_048_1265, w_048_1271, w_048_1272, w_048_1274, w_048_1276, w_048_1277, w_048_1281, w_048_1282, w_048_1283, w_048_1286, w_048_1287, w_048_1289, w_048_1290, w_048_1291, w_048_1292, w_048_1293, w_048_1297, w_048_1300, w_048_1301, w_048_1306, w_048_1308, w_048_1313, w_048_1315, w_048_1316, w_048_1318, w_048_1325, w_048_1326, w_048_1329, w_048_1331, w_048_1332, w_048_1336, w_048_1337, w_048_1338, w_048_1341, w_048_1344, w_048_1349, w_048_1351, w_048_1353, w_048_1356, w_048_1357, w_048_1359, w_048_1362, w_048_1364, w_048_1365, w_048_1366, w_048_1368, w_048_1369, w_048_1374, w_048_1375, w_048_1378, w_048_1380, w_048_1381, w_048_1385, w_048_1387, w_048_1389, w_048_1390, w_048_1391, w_048_1392, w_048_1393, w_048_1394, w_048_1398, w_048_1399, w_048_1403, w_048_1407, w_048_1408, w_048_1409, w_048_1412, w_048_1415, w_048_1417, w_048_1418, w_048_1419, w_048_1420, w_048_1421, w_048_1424, w_048_1427, w_048_1428, w_048_1430, w_048_1431, w_048_1436, w_048_1437, w_048_1439, w_048_1443, w_048_1444, w_048_1445, w_048_1447, w_048_1451, w_048_1452, w_048_1453, w_048_1454, w_048_1455, w_048_1456, w_048_1458, w_048_1460, w_048_1463, w_048_1464, w_048_1467, w_048_1468, w_048_1470, w_048_1471, w_048_1472, w_048_1478, w_048_1479, w_048_1482, w_048_1483, w_048_1484, w_048_1486, w_048_1487, w_048_1492, w_048_1496, w_048_1498, w_048_1499, w_048_1502, w_048_1503, w_048_1505, w_048_1506, w_048_1507, w_048_1508, w_048_1510, w_048_1511, w_048_1512, w_048_1513, w_048_1517, w_048_1518, w_048_1522, w_048_1526, w_048_1529, w_048_1532, w_048_1535, w_048_1537, w_048_1538, w_048_1541, w_048_1543, w_048_1545, w_048_1547, w_048_1548, w_048_1550, w_048_1553, w_048_1554, w_048_1555, w_048_1556, w_048_1557, w_048_1558, w_048_1559, w_048_1560, w_048_1561, w_048_1563, w_048_1564, w_048_1569, w_048_1570, w_048_1571, w_048_1572, w_048_1573, w_048_1575, w_048_1577, w_048_1580, w_048_1582, w_048_1583, w_048_1584, w_048_1587, w_048_1588, w_048_1589, w_048_1591, w_048_1595, w_048_1598, w_048_1599, w_048_1601, w_048_1602, w_048_1603, w_048_1607, w_048_1608, w_048_1609, w_048_1613, w_048_1614, w_048_1615, w_048_1616, w_048_1617, w_048_1619, w_048_1620, w_048_1622, w_048_1624, w_048_1626, w_048_1627, w_048_1628, w_048_1629, w_048_1631, w_048_1634, w_048_1635, w_048_1636, w_048_1637, w_048_1638, w_048_1639, w_048_1640, w_048_1641, w_048_1645, w_048_1646, w_048_1648, w_048_1650, w_048_1653, w_048_1654, w_048_1656, w_048_1658, w_048_1661, w_048_1666, w_048_1669, w_048_1673, w_048_1674, w_048_1676, w_048_1677, w_048_1678, w_048_1679, w_048_1685, w_048_1687, w_048_1692, w_048_1694, w_048_1695, w_048_1696, w_048_1697, w_048_1698, w_048_1701, w_048_1702, w_048_1703, w_048_1706, w_048_1708, w_048_1710, w_048_1711, w_048_1712, w_048_1713, w_048_1714, w_048_1715, w_048_1716, w_048_1717, w_048_1722, w_048_1725, w_048_1729, w_048_1730, w_048_1731, w_048_1733, w_048_1734, w_048_1736, w_048_1737, w_048_1738, w_048_1739, w_048_1743, w_048_1744, w_048_1745, w_048_1747, w_048_1748, w_048_1749, w_048_1751, w_048_1753, w_048_1754, w_048_1755, w_048_1756, w_048_1759, w_048_1760, w_048_1761, w_048_1762, w_048_1764, w_048_1765, w_048_1766, w_048_1767, w_048_1778, w_048_1779, w_048_1780, w_048_1783, w_048_1784, w_048_1786, w_048_1787, w_048_1788, w_048_1791, w_048_1794, w_048_1797, w_048_1799, w_048_1800, w_048_1801, w_048_1802, w_048_1803, w_048_1804, w_048_1806, w_048_1807, w_048_1809, w_048_1810, w_048_1812, w_048_1813, w_048_1814, w_048_1815, w_048_1816, w_048_1820, w_048_1821, w_048_1823, w_048_1824, w_048_1827, w_048_1831, w_048_1835, w_048_1836, w_048_1840, w_048_1841, w_048_1847, w_048_1850, w_048_1854, w_048_1855, w_048_1856, w_048_1857, w_048_1858, w_048_1861, w_048_1862, w_048_1864, w_048_1865, w_048_1870, w_048_1871, w_048_1872, w_048_1873, w_048_1874, w_048_1875, w_048_1877, w_048_1879, w_048_1881, w_048_1883, w_048_1887, w_048_1888, w_048_1890, w_048_1892, w_048_1893, w_048_1895, w_048_1896, w_048_1897, w_048_1898, w_048_1899, w_048_1900, w_048_1904, w_048_1906, w_048_1907, w_048_1908, w_048_1909, w_048_1910, w_048_1914, w_048_1916, w_048_1919, w_048_1922, w_048_1923, w_048_1924, w_048_1927, w_048_1929, w_048_1935, w_048_1936, w_048_1943, w_048_1944, w_048_1945, w_048_1947, w_048_1948, w_048_1951, w_048_1952, w_048_1953, w_048_1954, w_048_1961, w_048_1964, w_048_1967, w_048_1970, w_048_1971, w_048_1972, w_048_1973, w_048_1977, w_048_1980, w_048_1983, w_048_1985, w_048_1986, w_048_1987, w_048_1988, w_048_1989, w_048_1990, w_048_1991, w_048_1996, w_048_1997, w_048_2001, w_048_2002, w_048_2003, w_048_2004, w_048_2005, w_048_2007, w_048_2008, w_048_2009, w_048_2012, w_048_2013, w_048_2015, w_048_2016, w_048_2018, w_048_2022, w_048_2026, w_048_2027, w_048_2030, w_048_2031, w_048_2033, w_048_2034, w_048_2035, w_048_2036, w_048_2037, w_048_2038, w_048_2039, w_048_2041, w_048_2043, w_048_2046, w_048_2048, w_048_2050, w_048_2051, w_048_2052, w_048_2054, w_048_2057, w_048_2059, w_048_2060, w_048_2061, w_048_2063, w_048_2064, w_048_2066, w_048_2068, w_048_2069, w_048_2072, w_048_2074, w_048_2076, w_048_2078, w_048_2082, w_048_2084, w_048_2085, w_048_2086, w_048_2087, w_048_2089, w_048_2091, w_048_2093, w_048_2094, w_048_2102, w_048_2104, w_048_2106, w_048_2109, w_048_2110, w_048_2113, w_048_2114, w_048_2115, w_048_2117, w_048_2119, w_048_2121, w_048_2122, w_048_2123, w_048_2124, w_048_2130, w_048_2131, w_048_2133, w_048_2134, w_048_2141, w_048_2142, w_048_2145, w_048_2146, w_048_2150, w_048_2152, w_048_2153, w_048_2155, w_048_2157, w_048_2158, w_048_2159, w_048_2160, w_048_2161, w_048_2163, w_048_2164, w_048_2166, w_048_2167, w_048_2168, w_048_2169, w_048_2170, w_048_2171, w_048_2172, w_048_2173, w_048_2174, w_048_2179, w_048_2185, w_048_2187, w_048_2191, w_048_2192, w_048_2196, w_048_2197, w_048_2199, w_048_2202, w_048_2204, w_048_2207, w_048_2211, w_048_2212, w_048_2214, w_048_2215, w_048_2217, w_048_2218, w_048_2219, w_048_2221, w_048_2223, w_048_2224, w_048_2225, w_048_2228, w_048_2229, w_048_2231, w_048_2233, w_048_2234, w_048_2240, w_048_2241, w_048_2242, w_048_2244, w_048_2245, w_048_2246, w_048_2248, w_048_2249, w_048_2250, w_048_2251, w_048_2252, w_048_2256, w_048_2257, w_048_2258, w_048_2259, w_048_2260, w_048_2262, w_048_2272, w_048_2273, w_048_2274, w_048_2275, w_048_2277, w_048_2280, w_048_2281, w_048_2283, w_048_2285, w_048_2290, w_048_2292, w_048_2293, w_048_2296, w_048_2297, w_048_2298, w_048_2301, w_048_2309, w_048_2311, w_048_2312, w_048_2317, w_048_2318, w_048_2320, w_048_2323, w_048_2324, w_048_2326, w_048_2328, w_048_2329, w_048_2330, w_048_2331, w_048_2333, w_048_2335, w_048_2336, w_048_2338, w_048_2339, w_048_2340, w_048_2341, w_048_2343, w_048_2345, w_048_2347, w_048_2348, w_048_2349, w_048_2350, w_048_2352, w_048_2353, w_048_2355, w_048_2357, w_048_2358, w_048_2359, w_048_2362, w_048_2364, w_048_2369, w_048_2372, w_048_2373, w_048_2374, w_048_2376, w_048_2379, w_048_2380, w_048_2381, w_048_2382, w_048_2383, w_048_2387, w_048_2389, w_048_2391, w_048_2393, w_048_2394, w_048_2395, w_048_2396, w_048_2397, w_048_2400, w_048_2401, w_048_2402, w_048_2404, w_048_2406, w_048_2407, w_048_2408, w_048_2411, w_048_2414, w_048_2415, w_048_2416, w_048_2418, w_048_2420, w_048_2422, w_048_2425, w_048_2426, w_048_2428, w_048_2430, w_048_2436, w_048_2437, w_048_2438, w_048_2439, w_048_2446, w_048_2449, w_048_2452, w_048_2455, w_048_2456, w_048_2457, w_048_2458, w_048_2460, w_048_2461, w_048_2464, w_048_2465, w_048_2468, w_048_2469, w_048_2470, w_048_2471, w_048_2473, w_048_2474, w_048_2476, w_048_2477, w_048_2479, w_048_2480, w_048_2488, w_048_2489, w_048_2492, w_048_2495, w_048_2496, w_048_2497, w_048_2498, w_048_2501, w_048_2503, w_048_2504, w_048_2506, w_048_2507, w_048_2508, w_048_2511, w_048_2512, w_048_2514, w_048_2516, w_048_2517, w_048_2519, w_048_2521, w_048_2522, w_048_2523, w_048_2524, w_048_2525, w_048_2526, w_048_2533, w_048_2536, w_048_2537, w_048_2541, w_048_2545, w_048_2547, w_048_2548, w_048_2550, w_048_2551, w_048_2553, w_048_2555, w_048_2556, w_048_2561, w_048_2562, w_048_2563, w_048_2568, w_048_2571, w_048_2574, w_048_2580, w_048_2581, w_048_2585, w_048_2587, w_048_2590, w_048_2595, w_048_2596, w_048_2597, w_048_2598, w_048_2599, w_048_2600, w_048_2601, w_048_2603, w_048_2604, w_048_2608, w_048_2609, w_048_2610, w_048_2611, w_048_2613, w_048_2614, w_048_2615, w_048_2616, w_048_2621, w_048_2626, w_048_2628, w_048_2635, w_048_2636, w_048_2639, w_048_2640, w_048_2643, w_048_2644, w_048_2645, w_048_2650, w_048_2652, w_048_2656, w_048_2657, w_048_2658, w_048_2659, w_048_2661, w_048_2665, w_048_2674, w_048_2675, w_048_2679, w_048_2681, w_048_2683, w_048_2687, w_048_2691, w_048_2692, w_048_2693, w_048_2698, w_048_2699, w_048_2704, w_048_2706, w_048_2708, w_048_2711, w_048_2715, w_048_2717, w_048_2718, w_048_2719, w_048_2720, w_048_2721, w_048_2723, w_048_2724, w_048_2727, w_048_2731, w_048_2733, w_048_2734, w_048_2735, w_048_2737, w_048_2739, w_048_2742, w_048_2745, w_048_2747, w_048_2748, w_048_2749, w_048_2752, w_048_2755, w_048_2758, w_048_2764, w_048_2765, w_048_2766, w_048_2767, w_048_2773, w_048_2775, w_048_2777, w_048_2782, w_048_2785, w_048_2786, w_048_2788, w_048_2792, w_048_2793, w_048_2798, w_048_2799, w_048_2801, w_048_2803, w_048_2804, w_048_2805, w_048_2806, w_048_2807, w_048_2811, w_048_2812, w_048_2817, w_048_2818, w_048_2820, w_048_2821, w_048_2823, w_048_2824, w_048_2827, w_048_2828, w_048_2830, w_048_2833, w_048_2835, w_048_2837, w_048_2838, w_048_2839, w_048_2845, w_048_2851, w_048_2853, w_048_2858, w_048_2859, w_048_2860, w_048_2861, w_048_2864, w_048_2865, w_048_2869, w_048_2870, w_048_2871, w_048_2872, w_048_2874, w_048_2875, w_048_2876, w_048_2877, w_048_2879, w_048_2880, w_048_2884, w_048_2890, w_048_2891, w_048_2892, w_048_2894, w_048_2896, w_048_2899, w_048_2901, w_048_2906, w_048_2908, w_048_2909, w_048_2911, w_048_2912, w_048_2913, w_048_2915, w_048_2916, w_048_2917, w_048_2918, w_048_2919, w_048_2924, w_048_2925, w_048_2929, w_048_2932, w_048_2933, w_048_2934, w_048_2935, w_048_2939, w_048_2941, w_048_2942, w_048_2945, w_048_2946, w_048_2947, w_048_2950, w_048_2952, w_048_2955, w_048_2957, w_048_2964, w_048_2966, w_048_2967, w_048_2968, w_048_2969, w_048_2972, w_048_2975, w_048_2976, w_048_2978, w_048_2980, w_048_2981, w_048_2982, w_048_2983, w_048_2986, w_048_2987, w_048_2988, w_048_2990, w_048_2992, w_048_2994, w_048_2998, w_048_3004, w_048_3006, w_048_3011, w_048_3013, w_048_3014, w_048_3015, w_048_3016, w_048_3018, w_048_3020, w_048_3023, w_048_3024, w_048_3027, w_048_3029, w_048_3031, w_048_3039, w_048_3040, w_048_3042, w_048_3045, w_048_3049, w_048_3050, w_048_3051, w_048_3053, w_048_3055, w_048_3056, w_048_3059, w_048_3060, w_048_3061, w_048_3062, w_048_3066, w_048_3067, w_048_3073, w_048_3074, w_048_3075, w_048_3078, w_048_3082, w_048_3084, w_048_3088, w_048_3089, w_048_3093, w_048_3098, w_048_3101, w_048_3103, w_048_3104, w_048_3105, w_048_3106, w_048_3107, w_048_3112, w_048_3116, w_048_3117, w_048_3118, w_048_3119, w_048_3120, w_048_3122, w_048_3125, w_048_3127, w_048_3129, w_048_3132, w_048_3135, w_048_3136, w_048_3137, w_048_3138, w_048_3140, w_048_3141, w_048_3142, w_048_3143, w_048_3148, w_048_3152, w_048_3153, w_048_3156, w_048_3157, w_048_3158, w_048_3159, w_048_3161, w_048_3162, w_048_3163, w_048_3164, w_048_3165, w_048_3167, w_048_3171, w_048_3173, w_048_3174, w_048_3175, w_048_3176, w_048_3177, w_048_3181, w_048_3184, w_048_3185, w_048_3188, w_048_3194, w_048_3197, w_048_3198, w_048_3199, w_048_3201, w_048_3203, w_048_3204, w_048_3207, w_048_3210, w_048_3212, w_048_3216, w_048_3217, w_048_3219, w_048_3222, w_048_3223, w_048_3225, w_048_3231, w_048_3232, w_048_3236, w_048_3239, w_048_3240, w_048_3243, w_048_3244, w_048_3246, w_048_3247, w_048_3248, w_048_3249, w_048_3260, w_048_3263, w_048_3268, w_048_3269, w_048_3270, w_048_3275, w_048_3276, w_048_3277, w_048_3278, w_048_3279, w_048_3280, w_048_3281, w_048_3282, w_048_3283, w_048_3284, w_048_3287, w_048_3292, w_048_3293, w_048_3294, w_048_3295, w_048_3297, w_048_3299, w_048_3301, w_048_3302, w_048_3303, w_048_3308, w_048_3311, w_048_3312, w_048_3313, w_048_3315, w_048_3316, w_048_3317, w_048_3319, w_048_3320, w_048_3321, w_048_3323, w_048_3324, w_048_3325, w_048_3326, w_048_3329, w_048_3330, w_048_3334, w_048_3335, w_048_3336, w_048_3337, w_048_3339, w_048_3340, w_048_3342, w_048_3343, w_048_3348, w_048_3350, w_048_3351, w_048_3352, w_048_3353, w_048_3354, w_048_3355, w_048_3356, w_048_3357, w_048_3360, w_048_3361, w_048_3362, w_048_3369, w_048_3370, w_048_3373, w_048_3378, w_048_3379, w_048_3381, w_048_3382, w_048_3385, w_048_3386, w_048_3387, w_048_3388, w_048_3389, w_048_3390, w_048_3391, w_048_3392, w_048_3398, w_048_3401, w_048_3402, w_048_3403, w_048_3404, w_048_3405, w_048_3407, w_048_3408, w_048_3409, w_048_3410, w_048_3411, w_048_3414, w_048_3418, w_048_3420, w_048_3421, w_048_3422, w_048_3424, w_048_3428, w_048_3432, w_048_3435, w_048_3438, w_048_3439, w_048_3442, w_048_3443, w_048_3445, w_048_3446, w_048_3447, w_048_3448, w_048_3449, w_048_3451, w_048_3452, w_048_3453, w_048_3454, w_048_3455, w_048_3456, w_048_3457, w_048_3458, w_048_3460, w_048_3464, w_048_3465, w_048_3466, w_048_3467, w_048_3470, w_048_3472, w_048_3474, w_048_3475, w_048_3477, w_048_3478, w_048_3481, w_048_3483, w_048_3484, w_048_3485, w_048_3486, w_048_3487, w_048_3489, w_048_3491, w_048_3492, w_048_3494, w_048_3495, w_048_3496, w_048_3497, w_048_3499, w_048_3500, w_048_3503, w_048_3504, w_048_3505, w_048_3506, w_048_3507, w_048_3511, w_048_3512, w_048_3515, w_048_3516, w_048_3519, w_048_3520, w_048_3522, w_048_3523, w_048_3524, w_048_3526, w_048_3529, w_048_3533, w_048_3536, w_048_3539, w_048_3541, w_048_3542, w_048_3544, w_048_3545, w_048_3548, w_048_3549, w_048_3550, w_048_3552, w_048_3555, w_048_3556, w_048_3558, w_048_3560, w_048_3561, w_048_3563, w_048_3571, w_048_3573, w_048_3575, w_048_3577, w_048_3578, w_048_3579, w_048_3581, w_048_3584, w_048_3589, w_048_3591, w_048_3595, w_048_3596, w_048_3597, w_048_3599, w_048_3601, w_048_3602, w_048_3603, w_048_3608, w_048_3613, w_048_3614, w_048_3615, w_048_3616, w_048_3617, w_048_3618, w_048_3623, w_048_3625, w_048_3627, w_048_3628, w_048_3634, w_048_3643, w_048_3648, w_048_3650, w_048_3651, w_048_3653, w_048_3654, w_048_3656, w_048_3657, w_048_3659, w_048_3661, w_048_3665, w_048_3666, w_048_3667, w_048_3671, w_048_3672, w_048_3677, w_048_3678, w_048_3679, w_048_3680, w_048_3681, w_048_3682, w_048_3684, w_048_3685, w_048_3687, w_048_3688, w_048_3690, w_048_3692, w_048_3693, w_048_3694, w_048_3697, w_048_3698, w_048_3699, w_048_3701, w_048_3703, w_048_3710, w_048_3713, w_048_3715, w_048_3716, w_048_3717, w_048_3718, w_048_3723, w_048_3725, w_048_3726, w_048_3729, w_048_3731, w_048_3732, w_048_3734, w_048_3735, w_048_3736, w_048_3737, w_048_3738, w_048_3739, w_048_3740, w_048_3741, w_048_3746, w_048_3750, w_048_3752, w_048_3753, w_048_3756, w_048_3758, w_048_3759, w_048_3760, w_048_3761, w_048_3762, w_048_3764, w_048_3767, w_048_3768, w_048_3769, w_048_3776, w_048_3779, w_048_3781, w_048_3786, w_048_3787, w_048_3788, w_048_3789, w_048_3792, w_048_3798, w_048_3799, w_048_3800, w_048_3801, w_048_3803, w_048_3806, w_048_3807, w_048_3809, w_048_3810, w_048_3815, w_048_3817, w_048_3818, w_048_3820, w_048_3821, w_048_3825, w_048_3826, w_048_3831, w_048_3832, w_048_3833, w_048_3836, w_048_3838, w_048_3839, w_048_3840, w_048_3841, w_048_3843, w_048_3844, w_048_3845, w_048_3848, w_048_3849, w_048_3851, w_048_3852, w_048_3853, w_048_3857, w_048_3860, w_048_3861, w_048_3863, w_048_3865, w_048_3869, w_048_3874, w_048_3876, w_048_3879, w_048_3881, w_048_3883, w_048_3886, w_048_3888, w_048_3889, w_048_3891, w_048_3894, w_048_3898, w_048_3899, w_048_3901, w_048_3903, w_048_3904, w_048_3906, w_048_3907, w_048_3909, w_048_3910, w_048_3912, w_048_3914, w_048_3919, w_048_3920, w_048_3922, w_048_3923, w_048_3924, w_048_3926, w_048_3927, w_048_3930, w_048_3931, w_048_3935, w_048_3936, w_048_3939, w_048_3947, w_048_3949, w_048_3950, w_048_3955, w_048_3961, w_048_3967, w_048_3968, w_048_3969, w_048_3974, w_048_3976, w_048_3979, w_048_3980, w_048_3985, w_048_3986, w_048_3990, w_048_3991, w_048_3993, w_048_3994, w_048_4001, w_048_4002, w_048_4005, w_048_4008, w_048_4009, w_048_4010, w_048_4012, w_048_4013, w_048_4014, w_048_4018, w_048_4020, w_048_4026, w_048_4027, w_048_4028, w_048_4029, w_048_4030, w_048_4033, w_048_4034, w_048_4038, w_048_4041, w_048_4042, w_048_4043, w_048_4048, w_048_4050, w_048_4051, w_048_4053, w_048_4055, w_048_4056, w_048_4057, w_048_4058, w_048_4059, w_048_4060, w_048_4061, w_048_4066, w_048_4068, w_048_4072, w_048_4073, w_048_4074, w_048_4075, w_048_4079, w_048_4080, w_048_4081, w_048_4083, w_048_4084, w_048_4088, w_048_4091, w_048_4094, w_048_4096, w_048_4097, w_048_4098, w_048_4101, w_048_4103, w_048_4104, w_048_4105, w_048_4108, w_048_4110, w_048_4112, w_048_4113, w_048_4114, w_048_4115, w_048_4120, w_048_4123, w_048_4125, w_048_4126, w_048_4128, w_048_4130, w_048_4131, w_048_4133, w_048_4136, w_048_4141, w_048_4142, w_048_4146, w_048_4151, w_048_4154, w_048_4155, w_048_4157, w_048_4158, w_048_4160, w_048_4161, w_048_4164, w_048_4167, w_048_4168, w_048_4169, w_048_4170, w_048_4173, w_048_4175, w_048_4177, w_048_4178, w_048_4181, w_048_4183, w_048_4184, w_048_4187, w_048_4189, w_048_4192, w_048_4193, w_048_4195, w_048_4197, w_048_4199, w_048_4200, w_048_4201, w_048_4202, w_048_4203, w_048_4206, w_048_4213, w_048_4216, w_048_4218, w_048_4219, w_048_4220, w_048_4221, w_048_4227, w_048_4228, w_048_4233, w_048_4234, w_048_4235, w_048_4237, w_048_4239, w_048_4242, w_048_4243, w_048_4244, w_048_4247, w_048_4248, w_048_4249, w_048_4251, w_048_4252, w_048_4254, w_048_4255, w_048_4258, w_048_4259, w_048_4260, w_048_4261, w_048_4266, w_048_4272, w_048_4274, w_048_4275, w_048_4279, w_048_4282, w_048_4283, w_048_4284, w_048_4285, w_048_4290, w_048_4292, w_048_4293, w_048_4295, w_048_4296, w_048_4300, w_048_4303, w_048_4304, w_048_4305, w_048_4308, w_048_4311, w_048_4313, w_048_4314, w_048_4317, w_048_4319, w_048_4320, w_048_4322, w_048_4327, w_048_4329, w_048_4332, w_048_4333, w_048_4335, w_048_4338, w_048_4340, w_048_4341, w_048_4345, w_048_4346, w_048_4350, w_048_4354, w_048_4359, w_048_4360, w_048_4361, w_048_4363, w_048_4367, w_048_4368, w_048_4369, w_048_4372, w_048_4373, w_048_4374, w_048_4375, w_048_4379, w_048_4380, w_048_4382, w_048_4384, w_048_4385, w_048_4388, w_048_4390, w_048_4391, w_048_4395, w_048_4396, w_048_4399, w_048_4400, w_048_4401, w_048_4410, w_048_4413, w_048_4414, w_048_4416, w_048_4418, w_048_4420, w_048_4421, w_048_4422, w_048_4423, w_048_4424, w_048_4426, w_048_4427, w_048_4428, w_048_4431, w_048_4434, w_048_4435, w_048_4438, w_048_4440, w_048_4441, w_048_4442, w_048_4443, w_048_4444, w_048_4445, w_048_4446, w_048_4447, w_048_4448, w_048_4450, w_048_4452, w_048_4455, w_048_4456, w_048_4461, w_048_4462, w_048_4465, w_048_4468, w_048_4469, w_048_4472, w_048_4475, w_048_4476, w_048_4481, w_048_4488, w_048_4493, w_048_4495, w_048_4499, w_048_4501, w_048_4502, w_048_4503, w_048_4505, w_048_4506, w_048_4508, w_048_4510, w_048_4511, w_048_4516, w_048_4518, w_048_4519, w_048_4520, w_048_4521, w_048_4523, w_048_4525, w_048_4527, w_048_4528, w_048_4531, w_048_4535, w_048_4539, w_048_4540, w_048_4541, w_048_4542, w_048_4544, w_048_4548, w_048_4550, w_048_4551, w_048_4554, w_048_4556, w_048_4557, w_048_4558, w_048_4559, w_048_4560, w_048_4563, w_048_4565;
  wire w_049_000, w_049_001, w_049_003, w_049_004, w_049_005, w_049_006, w_049_007, w_049_008, w_049_009, w_049_011, w_049_012, w_049_015, w_049_016, w_049_018, w_049_019, w_049_020, w_049_022, w_049_023, w_049_025, w_049_026, w_049_028, w_049_029, w_049_030, w_049_031, w_049_032, w_049_033, w_049_035, w_049_036, w_049_037, w_049_038, w_049_039, w_049_040, w_049_041, w_049_042, w_049_043, w_049_046, w_049_047, w_049_048, w_049_050, w_049_051, w_049_052, w_049_053, w_049_054, w_049_056, w_049_057, w_049_058, w_049_059, w_049_060, w_049_061, w_049_062, w_049_063, w_049_065, w_049_066, w_049_067, w_049_069, w_049_071, w_049_072, w_049_073, w_049_074, w_049_075, w_049_076, w_049_078, w_049_079, w_049_080, w_049_081, w_049_082, w_049_083, w_049_086, w_049_088, w_049_089, w_049_090, w_049_092, w_049_093, w_049_094, w_049_095, w_049_096, w_049_097, w_049_098, w_049_099, w_049_100, w_049_102, w_049_103, w_049_104, w_049_105, w_049_107, w_049_108, w_049_109, w_049_111, w_049_112, w_049_119, w_049_120, w_049_121, w_049_122, w_049_123, w_049_124, w_049_125, w_049_126, w_049_127, w_049_128, w_049_129, w_049_130, w_049_132, w_049_133, w_049_136, w_049_138, w_049_139, w_049_142, w_049_145, w_049_147, w_049_148, w_049_149, w_049_150, w_049_151, w_049_152, w_049_153, w_049_155, w_049_156, w_049_157, w_049_158, w_049_159, w_049_160, w_049_163, w_049_164, w_049_165, w_049_166, w_049_170, w_049_171, w_049_172, w_049_173, w_049_174, w_049_175, w_049_176, w_049_177, w_049_179, w_049_180, w_049_181, w_049_182, w_049_183, w_049_184, w_049_188, w_049_189, w_049_190, w_049_191, w_049_192, w_049_193, w_049_194, w_049_197, w_049_199, w_049_200, w_049_201, w_049_202, w_049_204, w_049_205, w_049_207, w_049_208, w_049_209, w_049_210, w_049_211, w_049_213, w_049_214, w_049_215, w_049_216, w_049_217, w_049_219, w_049_220, w_049_221, w_049_225, w_049_226, w_049_227, w_049_228, w_049_229, w_049_231, w_049_232, w_049_233, w_049_234, w_049_235, w_049_238, w_049_239, w_049_240, w_049_241, w_049_242, w_049_243, w_049_245, w_049_247, w_049_248, w_049_250, w_049_252, w_049_253, w_049_254, w_049_255, w_049_256, w_049_258, w_049_259, w_049_260, w_049_261, w_049_262, w_049_264, w_049_265, w_049_266, w_049_267, w_049_269, w_049_270, w_049_271, w_049_273, w_049_274, w_049_277, w_049_278, w_049_279, w_049_280, w_049_281, w_049_282, w_049_283, w_049_284, w_049_285, w_049_286, w_049_287, w_049_288, w_049_289, w_049_290, w_049_293, w_049_294, w_049_295, w_049_296, w_049_297, w_049_298, w_049_299, w_049_300, w_049_301, w_049_302, w_049_303, w_049_304, w_049_305, w_049_307, w_049_308, w_049_309, w_049_310, w_049_311, w_049_312, w_049_313, w_049_314, w_049_315, w_049_316, w_049_318, w_049_319, w_049_320, w_049_322, w_049_323, w_049_324, w_049_325, w_049_327, w_049_328, w_049_329, w_049_331, w_049_333, w_049_334, w_049_335, w_049_336, w_049_337, w_049_338, w_049_339, w_049_340, w_049_341, w_049_342, w_049_343, w_049_344, w_049_345, w_049_347, w_049_348, w_049_349, w_049_350, w_049_352, w_049_354, w_049_355, w_049_356, w_049_357, w_049_359, w_049_360, w_049_361, w_049_362, w_049_363, w_049_364, w_049_366, w_049_367, w_049_368, w_049_369, w_049_370, w_049_371, w_049_372, w_049_373, w_049_374, w_049_375, w_049_376, w_049_377, w_049_378, w_049_379, w_049_380, w_049_381, w_049_382, w_049_383, w_049_384, w_049_386, w_049_387, w_049_389, w_049_390, w_049_391, w_049_392, w_049_393, w_049_394, w_049_395, w_049_396, w_049_397, w_049_401, w_049_402, w_049_403, w_049_404, w_049_405, w_049_406, w_049_409, w_049_410, w_049_411, w_049_412, w_049_414, w_049_415, w_049_416, w_049_417, w_049_418, w_049_419, w_049_420, w_049_421, w_049_422, w_049_423, w_049_424, w_049_427, w_049_430, w_049_433, w_049_434, w_049_435, w_049_436, w_049_437, w_049_439, w_049_440, w_049_441, w_049_442, w_049_443, w_049_444, w_049_446, w_049_448, w_049_449, w_049_450, w_049_451, w_049_453, w_049_454, w_049_455, w_049_456, w_049_457, w_049_458, w_049_459, w_049_460, w_049_461, w_049_463, w_049_465, w_049_466, w_049_468, w_049_469, w_049_470, w_049_471, w_049_475, w_049_476, w_049_477, w_049_478, w_049_480, w_049_481, w_049_483, w_049_484, w_049_485, w_049_488, w_049_489, w_049_492, w_049_493, w_049_495, w_049_496, w_049_498, w_049_499, w_049_500, w_049_502, w_049_503, w_049_504, w_049_505, w_049_506, w_049_507, w_049_508, w_049_509, w_049_512, w_049_513, w_049_514, w_049_515, w_049_516, w_049_518, w_049_519, w_049_520, w_049_522, w_049_523, w_049_524, w_049_525, w_049_526, w_049_528, w_049_530, w_049_531, w_049_532, w_049_533, w_049_534, w_049_535, w_049_536, w_049_537, w_049_539, w_049_541, w_049_542, w_049_543, w_049_547, w_049_549, w_049_550, w_049_551, w_049_552, w_049_553, w_049_555, w_049_556, w_049_557, w_049_558, w_049_559, w_049_560, w_049_563, w_049_564, w_049_566, w_049_567, w_049_568, w_049_569, w_049_571, w_049_572, w_049_573, w_049_574, w_049_575, w_049_576, w_049_577, w_049_578, w_049_581, w_049_582, w_049_583, w_049_584, w_049_587, w_049_588, w_049_589, w_049_591, w_049_594, w_049_595, w_049_596, w_049_598, w_049_599, w_049_600, w_049_601, w_049_603, w_049_604, w_049_605, w_049_606, w_049_608, w_049_609, w_049_610, w_049_611, w_049_612, w_049_614, w_049_615, w_049_621, w_049_622, w_049_623, w_049_624, w_049_625, w_049_626, w_049_627, w_049_629, w_049_630, w_049_631, w_049_632, w_049_634, w_049_635, w_049_636, w_049_637, w_049_638, w_049_640, w_049_641, w_049_642, w_049_643, w_049_644, w_049_645, w_049_646, w_049_647, w_049_649, w_049_650, w_049_652, w_049_654, w_049_657, w_049_658, w_049_659, w_049_660, w_049_661, w_049_662, w_049_664, w_049_665, w_049_666, w_049_668, w_049_669, w_049_670, w_049_672, w_049_673, w_049_674, w_049_675, w_049_676, w_049_678, w_049_679, w_049_681, w_049_686, w_049_689, w_049_691, w_049_693, w_049_694, w_049_695, w_049_696, w_049_697, w_049_698, w_049_700, w_049_702, w_049_703, w_049_707, w_049_708, w_049_709, w_049_715, w_049_718, w_049_719, w_049_722, w_049_723, w_049_727, w_049_729, w_049_733, w_049_734, w_049_735, w_049_737, w_049_739, w_049_745, w_049_746, w_049_748, w_049_749, w_049_750, w_049_751, w_049_752, w_049_753, w_049_754, w_049_755, w_049_757, w_049_758, w_049_766, w_049_767, w_049_768, w_049_771, w_049_772, w_049_774, w_049_775, w_049_776, w_049_778, w_049_779, w_049_783, w_049_786, w_049_787, w_049_788, w_049_789, w_049_791, w_049_793, w_049_795, w_049_798, w_049_799, w_049_800, w_049_804, w_049_805, w_049_812, w_049_814, w_049_816, w_049_818, w_049_820, w_049_822, w_049_829, w_049_830, w_049_831, w_049_835, w_049_841, w_049_842, w_049_848, w_049_849, w_049_855, w_049_856, w_049_857, w_049_859, w_049_860, w_049_864, w_049_866, w_049_873, w_049_874, w_049_876, w_049_877, w_049_883, w_049_886, w_049_890, w_049_893, w_049_894, w_049_895, w_049_898, w_049_900, w_049_901, w_049_902, w_049_905, w_049_908, w_049_910, w_049_912, w_049_917, w_049_919, w_049_922, w_049_925, w_049_928, w_049_930, w_049_931, w_049_932, w_049_933, w_049_935, w_049_939, w_049_941, w_049_942, w_049_944, w_049_945, w_049_946, w_049_947, w_049_949, w_049_952, w_049_954, w_049_955, w_049_958, w_049_960, w_049_961, w_049_963, w_049_964, w_049_967, w_049_968, w_049_971, w_049_973, w_049_977, w_049_979, w_049_980, w_049_981, w_049_984, w_049_985, w_049_987, w_049_988, w_049_989, w_049_990, w_049_991, w_049_992, w_049_995, w_049_996, w_049_999, w_049_1000, w_049_1001, w_049_1002, w_049_1003, w_049_1004, w_049_1007, w_049_1011, w_049_1012, w_049_1015, w_049_1020, w_049_1023, w_049_1024, w_049_1026, w_049_1028, w_049_1032, w_049_1037, w_049_1040, w_049_1043, w_049_1045, w_049_1047, w_049_1051, w_049_1052, w_049_1053, w_049_1058, w_049_1059, w_049_1060, w_049_1061, w_049_1064, w_049_1068, w_049_1071, w_049_1078, w_049_1079, w_049_1080, w_049_1081, w_049_1087, w_049_1090, w_049_1091, w_049_1092, w_049_1093, w_049_1097, w_049_1099, w_049_1100, w_049_1101, w_049_1103, w_049_1104, w_049_1105, w_049_1107, w_049_1108, w_049_1110, w_049_1111, w_049_1112, w_049_1113, w_049_1114, w_049_1115, w_049_1116, w_049_1117, w_049_1119, w_049_1120, w_049_1121, w_049_1122, w_049_1123, w_049_1125, w_049_1129, w_049_1130, w_049_1136, w_049_1137, w_049_1146, w_049_1149, w_049_1150, w_049_1152, w_049_1154, w_049_1155, w_049_1156, w_049_1157, w_049_1158, w_049_1159, w_049_1161, w_049_1163, w_049_1164, w_049_1165, w_049_1167, w_049_1169, w_049_1172, w_049_1175, w_049_1177, w_049_1178, w_049_1180, w_049_1182, w_049_1183, w_049_1186, w_049_1188, w_049_1191, w_049_1192, w_049_1193, w_049_1194, w_049_1195, w_049_1196, w_049_1197, w_049_1200, w_049_1203, w_049_1205, w_049_1206, w_049_1208, w_049_1210, w_049_1212, w_049_1213, w_049_1214, w_049_1216, w_049_1224, w_049_1226, w_049_1227, w_049_1228, w_049_1233, w_049_1234, w_049_1235, w_049_1244, w_049_1245, w_049_1247, w_049_1251, w_049_1252, w_049_1255, w_049_1256, w_049_1258, w_049_1259, w_049_1267, w_049_1268, w_049_1270, w_049_1273, w_049_1275, w_049_1283, w_049_1284, w_049_1290, w_049_1294, w_049_1295, w_049_1296, w_049_1298, w_049_1300, w_049_1303, w_049_1306, w_049_1307, w_049_1310, w_049_1312, w_049_1314, w_049_1316, w_049_1317, w_049_1322, w_049_1325, w_049_1326, w_049_1328, w_049_1330, w_049_1333, w_049_1334, w_049_1336, w_049_1337, w_049_1338, w_049_1339, w_049_1341, w_049_1343, w_049_1345, w_049_1349, w_049_1351, w_049_1352, w_049_1355, w_049_1356, w_049_1357, w_049_1358, w_049_1361, w_049_1363, w_049_1364, w_049_1370, w_049_1372, w_049_1375, w_049_1376, w_049_1377, w_049_1379, w_049_1380, w_049_1381, w_049_1382, w_049_1387, w_049_1388, w_049_1389, w_049_1390, w_049_1391, w_049_1393, w_049_1394, w_049_1395, w_049_1397, w_049_1401, w_049_1402, w_049_1403, w_049_1405, w_049_1406, w_049_1407, w_049_1408, w_049_1409, w_049_1411, w_049_1415, w_049_1419, w_049_1420, w_049_1422, w_049_1424, w_049_1427, w_049_1428, w_049_1432, w_049_1433, w_049_1434, w_049_1436, w_049_1437, w_049_1438, w_049_1441, w_049_1444, w_049_1449, w_049_1450, w_049_1451, w_049_1453, w_049_1454, w_049_1458, w_049_1459, w_049_1461, w_049_1462, w_049_1465, w_049_1467, w_049_1468, w_049_1469, w_049_1471, w_049_1474, w_049_1476, w_049_1477, w_049_1478, w_049_1480, w_049_1481, w_049_1486, w_049_1487, w_049_1489, w_049_1490, w_049_1492, w_049_1495, w_049_1497, w_049_1498, w_049_1503, w_049_1505, w_049_1506, w_049_1508, w_049_1509, w_049_1510, w_049_1512, w_049_1514, w_049_1515, w_049_1517, w_049_1519, w_049_1522, w_049_1524, w_049_1529, w_049_1532, w_049_1534, w_049_1535, w_049_1538, w_049_1539, w_049_1540, w_049_1542, w_049_1545, w_049_1547, w_049_1548, w_049_1550, w_049_1551, w_049_1552, w_049_1554, w_049_1557, w_049_1560, w_049_1563, w_049_1565, w_049_1569, w_049_1572, w_049_1573, w_049_1575, w_049_1577, w_049_1585, w_049_1589, w_049_1590, w_049_1591, w_049_1594, w_049_1596, w_049_1602, w_049_1603, w_049_1604, w_049_1606, w_049_1607, w_049_1608, w_049_1609, w_049_1610, w_049_1613, w_049_1615, w_049_1617, w_049_1619, w_049_1624, w_049_1625, w_049_1628, w_049_1630, w_049_1631, w_049_1635, w_049_1638, w_049_1641, w_049_1643, w_049_1645, w_049_1646, w_049_1647, w_049_1650, w_049_1651, w_049_1655, w_049_1656, w_049_1657, w_049_1659, w_049_1664, w_049_1666, w_049_1667, w_049_1668, w_049_1670, w_049_1671, w_049_1675, w_049_1677, w_049_1679, w_049_1680, w_049_1681, w_049_1684, w_049_1687, w_049_1688, w_049_1690, w_049_1691, w_049_1692, w_049_1693, w_049_1694, w_049_1695, w_049_1696, w_049_1697, w_049_1698, w_049_1702, w_049_1707, w_049_1710, w_049_1711, w_049_1712, w_049_1713, w_049_1715, w_049_1720, w_049_1721, w_049_1722, w_049_1727, w_049_1733, w_049_1734, w_049_1736, w_049_1737, w_049_1738, w_049_1739, w_049_1740, w_049_1747, w_049_1748, w_049_1749, w_049_1750, w_049_1751, w_049_1755, w_049_1758, w_049_1759, w_049_1760, w_049_1761, w_049_1762, w_049_1766, w_049_1767, w_049_1768, w_049_1770, w_049_1772, w_049_1773, w_049_1774, w_049_1775, w_049_1780, w_049_1785, w_049_1787, w_049_1790, w_049_1795, w_049_1803, w_049_1804, w_049_1805, w_049_1806, w_049_1807, w_049_1810, w_049_1811, w_049_1813, w_049_1815, w_049_1816, w_049_1819, w_049_1820, w_049_1821, w_049_1822, w_049_1823, w_049_1824, w_049_1826, w_049_1829, w_049_1831, w_049_1834, w_049_1835, w_049_1836, w_049_1837, w_049_1841, w_049_1843, w_049_1844, w_049_1845, w_049_1847, w_049_1848, w_049_1850, w_049_1852, w_049_1853, w_049_1855, w_049_1857, w_049_1858, w_049_1861, w_049_1862, w_049_1864, w_049_1866, w_049_1867, w_049_1868, w_049_1869, w_049_1873, w_049_1874, w_049_1876, w_049_1877, w_049_1879, w_049_1881, w_049_1883, w_049_1885, w_049_1887, w_049_1888, w_049_1889, w_049_1890, w_049_1891, w_049_1892, w_049_1893, w_049_1894, w_049_1895, w_049_1896, w_049_1898, w_049_1900, w_049_1901, w_049_1902, w_049_1903, w_049_1908, w_049_1910, w_049_1912, w_049_1913, w_049_1914, w_049_1916, w_049_1917, w_049_1919, w_049_1920, w_049_1922, w_049_1926, w_049_1927, w_049_1929, w_049_1930, w_049_1933, w_049_1934, w_049_1935, w_049_1937, w_049_1939, w_049_1940, w_049_1943, w_049_1944, w_049_1949, w_049_1950, w_049_1952, w_049_1955, w_049_1957, w_049_1959, w_049_1961, w_049_1962, w_049_1965, w_049_1967, w_049_1968, w_049_1972, w_049_1974, w_049_1975, w_049_1976, w_049_1978, w_049_1983, w_049_1988, w_049_1989, w_049_1990, w_049_1991, w_049_1993, w_049_1995, w_049_1996, w_049_1997, w_049_2000, w_049_2005, w_049_2006, w_049_2008, w_049_2009, w_049_2011, w_049_2012, w_049_2013, w_049_2017, w_049_2018, w_049_2020, w_049_2021, w_049_2022, w_049_2023, w_049_2024, w_049_2025, w_049_2026, w_049_2028, w_049_2032, w_049_2033, w_049_2037, w_049_2038, w_049_2039, w_049_2040, w_049_2041, w_049_2046, w_049_2047, w_049_2048, w_049_2049, w_049_2052, w_049_2053, w_049_2054, w_049_2056, w_049_2057, w_049_2060, w_049_2061, w_049_2063, w_049_2064, w_049_2065, w_049_2068, w_049_2070, w_049_2072, w_049_2073, w_049_2074, w_049_2076, w_049_2077, w_049_2078, w_049_2083, w_049_2084, w_049_2085, w_049_2086, w_049_2087, w_049_2090, w_049_2091, w_049_2093, w_049_2094, w_049_2095, w_049_2104, w_049_2106, w_049_2107, w_049_2110, w_049_2113, w_049_2114, w_049_2116, w_049_2117, w_049_2118, w_049_2120, w_049_2121, w_049_2122, w_049_2124, w_049_2126, w_049_2130, w_049_2131, w_049_2132, w_049_2135, w_049_2138, w_049_2139, w_049_2140, w_049_2141, w_049_2144, w_049_2145, w_049_2146, w_049_2149, w_049_2154, w_049_2155, w_049_2159, w_049_2161, w_049_2162, w_049_2164, w_049_2170, w_049_2171, w_049_2172, w_049_2174, w_049_2175, w_049_2178, w_049_2179, w_049_2182, w_049_2183, w_049_2185, w_049_2186, w_049_2187, w_049_2188, w_049_2191, w_049_2192, w_049_2193, w_049_2194, w_049_2195, w_049_2196, w_049_2197, w_049_2199, w_049_2201, w_049_2203, w_049_2205, w_049_2212, w_049_2213, w_049_2215, w_049_2216, w_049_2219, w_049_2220, w_049_2223, w_049_2224, w_049_2226, w_049_2227, w_049_2229, w_049_2230, w_049_2231, w_049_2232, w_049_2233, w_049_2234, w_049_2235, w_049_2237, w_049_2238, w_049_2240, w_049_2241, w_049_2242, w_049_2244, w_049_2245, w_049_2246, w_049_2248, w_049_2250, w_049_2253, w_049_2259, w_049_2260, w_049_2262, w_049_2264, w_049_2266, w_049_2268, w_049_2269, w_049_2271, w_049_2272, w_049_2275, w_049_2277, w_049_2279, w_049_2282, w_049_2283, w_049_2285, w_049_2286, w_049_2287, w_049_2288, w_049_2290, w_049_2291, w_049_2292, w_049_2293, w_049_2294, w_049_2295, w_049_2296, w_049_2298, w_049_2299, w_049_2300, w_049_2302, w_049_2303, w_049_2305, w_049_2310, w_049_2314, w_049_2315, w_049_2316, w_049_2319, w_049_2320, w_049_2321, w_049_2322, w_049_2323, w_049_2325, w_049_2331, w_049_2332, w_049_2333, w_049_2334, w_049_2335, w_049_2336, w_049_2337, w_049_2338, w_049_2340, w_049_2343, w_049_2344, w_049_2345, w_049_2346, w_049_2349, w_049_2350, w_049_2353, w_049_2354, w_049_2357, w_049_2358, w_049_2364, w_049_2370, w_049_2371, w_049_2372, w_049_2375, w_049_2376, w_049_2377, w_049_2378, w_049_2379, w_049_2382, w_049_2383, w_049_2384, w_049_2385, w_049_2386, w_049_2387, w_049_2388, w_049_2390, w_049_2393, w_049_2402, w_049_2403, w_049_2406, w_049_2407, w_049_2408, w_049_2409, w_049_2410, w_049_2411, w_049_2414, w_049_2417, w_049_2418, w_049_2420, w_049_2423, w_049_2425, w_049_2427, w_049_2428, w_049_2429, w_049_2431, w_049_2432, w_049_2438, w_049_2439, w_049_2440, w_049_2441, w_049_2447, w_049_2449, w_049_2450, w_049_2451, w_049_2452, w_049_2454, w_049_2455, w_049_2456, w_049_2457, w_049_2461, w_049_2462, w_049_2463, w_049_2464, w_049_2465, w_049_2466, w_049_2467, w_049_2468, w_049_2469, w_049_2471, w_049_2474, w_049_2478, w_049_2479, w_049_2483, w_049_2484, w_049_2486, w_049_2487, w_049_2488, w_049_2492, w_049_2498, w_049_2499, w_049_2500, w_049_2501, w_049_2506, w_049_2508, w_049_2511, w_049_2512, w_049_2513, w_049_2514, w_049_2515, w_049_2516, w_049_2517, w_049_2520, w_049_2525, w_049_2526, w_049_2527, w_049_2528, w_049_2536, w_049_2540, w_049_2542, w_049_2543, w_049_2544, w_049_2545, w_049_2548, w_049_2549, w_049_2552, w_049_2553, w_049_2556, w_049_2561, w_049_2562, w_049_2565, w_049_2566, w_049_2569, w_049_2570, w_049_2578, w_049_2580, w_049_2581, w_049_2582, w_049_2584, w_049_2585, w_049_2586, w_049_2588, w_049_2589, w_049_2590, w_049_2592, w_049_2594, w_049_2599, w_049_2601, w_049_2603, w_049_2604, w_049_2607, w_049_2608, w_049_2609, w_049_2616, w_049_2618, w_049_2621, w_049_2623, w_049_2625, w_049_2626, w_049_2628, w_049_2629, w_049_2634, w_049_2635, w_049_2639, w_049_2642, w_049_2643, w_049_2644, w_049_2646, w_049_2647, w_049_2651, w_049_2653, w_049_2654, w_049_2659, w_049_2661, w_049_2662, w_049_2664, w_049_2669, w_049_2670, w_049_2672, w_049_2677, w_049_2681, w_049_2686, w_049_2687, w_049_2688, w_049_2689, w_049_2690, w_049_2692, w_049_2693, w_049_2695, w_049_2696, w_049_2701, w_049_2702, w_049_2705, w_049_2707, w_049_2715, w_049_2716, w_049_2717, w_049_2718, w_049_2722, w_049_2723, w_049_2728, w_049_2729, w_049_2731, w_049_2732, w_049_2735, w_049_2736, w_049_2739, w_049_2742, w_049_2753, w_049_2755, w_049_2757, w_049_2759, w_049_2762, w_049_2766, w_049_2770, w_049_2771, w_049_2772, w_049_2773, w_049_2776, w_049_2777, w_049_2784, w_049_2786, w_049_2787, w_049_2788, w_049_2789, w_049_2790, w_049_2792, w_049_2793, w_049_2794, w_049_2796, w_049_2798, w_049_2799, w_049_2801, w_049_2802, w_049_2803, w_049_2804, w_049_2807, w_049_2810, w_049_2811, w_049_2812, w_049_2814, w_049_2817, w_049_2818, w_049_2819, w_049_2821, w_049_2824, w_049_2826, w_049_2827, w_049_2829, w_049_2831, w_049_2835, w_049_2836, w_049_2838, w_049_2840, w_049_2843, w_049_2845, w_049_2846, w_049_2849, w_049_2850, w_049_2852, w_049_2853, w_049_2854, w_049_2856, w_049_2858, w_049_2860, w_049_2862, w_049_2863, w_049_2865, w_049_2866, w_049_2867, w_049_2868, w_049_2871, w_049_2875, w_049_2878, w_049_2885, w_049_2887, w_049_2888, w_049_2890, w_049_2891, w_049_2893, w_049_2894, w_049_2896, w_049_2898, w_049_2899, w_049_2900, w_049_2903, w_049_2907, w_049_2910, w_049_2911, w_049_2914, w_049_2917, w_049_2919, w_049_2920, w_049_2922, w_049_2923, w_049_2927, w_049_2928, w_049_2930, w_049_2933, w_049_2935, w_049_2936, w_049_2937, w_049_2939, w_049_2942, w_049_2943, w_049_2944, w_049_2947, w_049_2950, w_049_2951, w_049_2954, w_049_2955, w_049_2957, w_049_2960, w_049_2962, w_049_2965, w_049_2967, w_049_2968, w_049_2972, w_049_2973, w_049_2974, w_049_2976, w_049_2977, w_049_2978, w_049_2980, w_049_2982, w_049_2986, w_049_2987, w_049_2988, w_049_2990, w_049_2991, w_049_2998, w_049_2999, w_049_3002, w_049_3005, w_049_3008, w_049_3010, w_049_3011, w_049_3014, w_049_3018, w_049_3021, w_049_3024, w_049_3025, w_049_3028, w_049_3031, w_049_3034, w_049_3035, w_049_3036, w_049_3040, w_049_3043, w_049_3044, w_049_3046, w_049_3051, w_049_3052, w_049_3053, w_049_3054, w_049_3060, w_049_3061, w_049_3062, w_049_3063, w_049_3064, w_049_3066, w_049_3067, w_049_3068, w_049_3073, w_049_3074, w_049_3077, w_049_3078, w_049_3079, w_049_3084, w_049_3085, w_049_3086, w_049_3089, w_049_3093, w_049_3094, w_049_3095, w_049_3096, w_049_3100, w_049_3101, w_049_3102, w_049_3103, w_049_3105, w_049_3106, w_049_3107, w_049_3109, w_049_3110, w_049_3111, w_049_3113, w_049_3115, w_049_3116, w_049_3119, w_049_3122, w_049_3123, w_049_3124, w_049_3127, w_049_3132, w_049_3133, w_049_3135, w_049_3137, w_049_3138, w_049_3141, w_049_3143, w_049_3144, w_049_3145, w_049_3147, w_049_3150, w_049_3151, w_049_3152, w_049_3153, w_049_3157, w_049_3160, w_049_3163, w_049_3164, w_049_3165, w_049_3167, w_049_3168, w_049_3170, w_049_3172, w_049_3173, w_049_3175, w_049_3176, w_049_3178, w_049_3179, w_049_3182, w_049_3183, w_049_3184, w_049_3185, w_049_3186, w_049_3189, w_049_3190, w_049_3198, w_049_3199, w_049_3200, w_049_3202, w_049_3205, w_049_3206, w_049_3207, w_049_3209, w_049_3210, w_049_3212, w_049_3213, w_049_3215, w_049_3216, w_049_3217, w_049_3219, w_049_3220, w_049_3221, w_049_3223, w_049_3225, w_049_3228, w_049_3229, w_049_3231, w_049_3234, w_049_3236, w_049_3237, w_049_3238, w_049_3239, w_049_3241, w_049_3242, w_049_3243, w_049_3247, w_049_3251, w_049_3253, w_049_3256, w_049_3258, w_049_3260, w_049_3264, w_049_3266, w_049_3268, w_049_3269, w_049_3270, w_049_3274, w_049_3275, w_049_3276, w_049_3278, w_049_3279, w_049_3280, w_049_3282, w_049_3284, w_049_3290, w_049_3291, w_049_3295, w_049_3298, w_049_3299, w_049_3302, w_049_3303, w_049_3305, w_049_3307, w_049_3308, w_049_3313, w_049_3315, w_049_3316, w_049_3319, w_049_3320, w_049_3321, w_049_3322, w_049_3323, w_049_3324, w_049_3326, w_049_3327, w_049_3330, w_049_3331, w_049_3333, w_049_3334, w_049_3335, w_049_3336, w_049_3337, w_049_3338, w_049_3339, w_049_3340, w_049_3345, w_049_3346, w_049_3348, w_049_3349, w_049_3351, w_049_3353, w_049_3356, w_049_3357, w_049_3359, w_049_3360, w_049_3361, w_049_3362, w_049_3365, w_049_3367, w_049_3368, w_049_3371, w_049_3372, w_049_3378, w_049_3379, w_049_3381, w_049_3385, w_049_3387, w_049_3388, w_049_3390, w_049_3391, w_049_3392, w_049_3393, w_049_3394, w_049_3395, w_049_3396, w_049_3401, w_049_3403, w_049_3405, w_049_3406, w_049_3408, w_049_3409, w_049_3411, w_049_3412, w_049_3414, w_049_3415, w_049_3417, w_049_3419, w_049_3421, w_049_3422, w_049_3426, w_049_3427, w_049_3429, w_049_3432, w_049_3434, w_049_3435, w_049_3436, w_049_3437, w_049_3441, w_049_3443, w_049_3444, w_049_3446, w_049_3454, w_049_3456, w_049_3457, w_049_3458, w_049_3460, w_049_3464, w_049_3465, w_049_3466, w_049_3471, w_049_3474, w_049_3475, w_049_3477, w_049_3478, w_049_3480, w_049_3481, w_049_3484, w_049_3485, w_049_3486, w_049_3487, w_049_3488, w_049_3489, w_049_3495, w_049_3499, w_049_3500, w_049_3503, w_049_3504, w_049_3508, w_049_3510, w_049_3513, w_049_3517, w_049_3518, w_049_3520, w_049_3522, w_049_3523, w_049_3525, w_049_3526, w_049_3529, w_049_3531, w_049_3532, w_049_3533, w_049_3534, w_049_3535, w_049_3537, w_049_3540, w_049_3541, w_049_3542, w_049_3543, w_049_3545, w_049_3546, w_049_3547, w_049_3548, w_049_3550, w_049_3551, w_049_3552, w_049_3553, w_049_3556, w_049_3559, w_049_3560, w_049_3561, w_049_3562, w_049_3563, w_049_3564, w_049_3566, w_049_3568, w_049_3569, w_049_3572, w_049_3575, w_049_3577, w_049_3578, w_049_3581, w_049_3583, w_049_3584, w_049_3587, w_049_3591, w_049_3592, w_049_3593, w_049_3594, w_049_3595, w_049_3600, w_049_3602, w_049_3603, w_049_3605, w_049_3606, w_049_3607, w_049_3609, w_049_3610, w_049_3612, w_049_3614, w_049_3615, w_049_3618, w_049_3620, w_049_3621, w_049_3622, w_049_3623, w_049_3624, w_049_3625, w_049_3628, w_049_3630, w_049_3633, w_049_3635, w_049_3638, w_049_3642, w_049_3643, w_049_3645, w_049_3646, w_049_3647, w_049_3649, w_049_3650, w_049_3651, w_049_3652, w_049_3656, w_049_3663, w_049_3664, w_049_3667, w_049_3668, w_049_3670, w_049_3671, w_049_3672, w_049_3674, w_049_3675, w_049_3676, w_049_3677, w_049_3678, w_049_3681, w_049_3683, w_049_3684, w_049_3685, w_049_3686, w_049_3687, w_049_3688, w_049_3689, w_049_3691, w_049_3692, w_049_3695, w_049_3698, w_049_3700, w_049_3702, w_049_3705, w_049_3706, w_049_3709, w_049_3710, w_049_3711, w_049_3718, w_049_3719, w_049_3722, w_049_3723, w_049_3725, w_049_3728, w_049_3730, w_049_3733, w_049_3735, w_049_3736, w_049_3737, w_049_3738, w_049_3742, w_049_3743, w_049_3747, w_049_3751, w_049_3752, w_049_3754, w_049_3756, w_049_3760, w_049_3761, w_049_3762, w_049_3764, w_049_3767, w_049_3771, w_049_3774, w_049_3776, w_049_3777, w_049_3778, w_049_3779, w_049_3780, w_049_3784, w_049_3785, w_049_3786, w_049_3788, w_049_3795, w_049_3796, w_049_3797, w_049_3798, w_049_3799, w_049_3800, w_049_3801, w_049_3803, w_049_3806, w_049_3808, w_049_3809, w_049_3813, w_049_3814, w_049_3815, w_049_3816, w_049_3817, w_049_3818, w_049_3822, w_049_3824, w_049_3825, w_049_3826, w_049_3829, w_049_3831, w_049_3832, w_049_3836, w_049_3838, w_049_3840, w_049_3841, w_049_3844, w_049_3845, w_049_3846, w_049_3847, w_049_3848, w_049_3849, w_049_3850, w_049_3851, w_049_3852, w_049_3853, w_049_3854, w_049_3859, w_049_3860, w_049_3861, w_049_3862, w_049_3863, w_049_3869, w_049_3871, w_049_3875, w_049_3877, w_049_3878, w_049_3879, w_049_3883, w_049_3884, w_049_3886, w_049_3887, w_049_3888, w_049_3889, w_049_3891, w_049_3895, w_049_3896, w_049_3902, w_049_3903, w_049_3905, w_049_3909, w_049_3912, w_049_3916, w_049_3917, w_049_3919, w_049_3921, w_049_3922, w_049_3928, w_049_3929, w_049_3931, w_049_3933, w_049_3936, w_049_3938, w_049_3940, w_049_3943, w_049_3944, w_049_3947, w_049_3948, w_049_3958, w_049_3959, w_049_3965, w_049_3967, w_049_3970, w_049_3972, w_049_3974, w_049_3975, w_049_3978, w_049_3979, w_049_3980, w_049_3981, w_049_3982, w_049_3983, w_049_3988, w_049_3989, w_049_3990, w_049_3991, w_049_3992, w_049_3993, w_049_3994, w_049_3996, w_049_3997, w_049_3998, w_049_4005, w_049_4006, w_049_4007, w_049_4011, w_049_4012, w_049_4013, w_049_4015, w_049_4016, w_049_4017, w_049_4018, w_049_4019, w_049_4020, w_049_4024, w_049_4025, w_049_4027, w_049_4028, w_049_4029, w_049_4031, w_049_4032, w_049_4033, w_049_4035, w_049_4037, w_049_4038, w_049_4039, w_049_4041, w_049_4043, w_049_4047, w_049_4049, w_049_4051, w_049_4052, w_049_4053, w_049_4059, w_049_4062, w_049_4063, w_049_4066, w_049_4067, w_049_4068, w_049_4073, w_049_4075, w_049_4079, w_049_4080, w_049_4082, w_049_4088, w_049_4089, w_049_4091, w_049_4092, w_049_4093, w_049_4094, w_049_4096, w_049_4097, w_049_4098, w_049_4102, w_049_4104, w_049_4106, w_049_4107, w_049_4108, w_049_4111, w_049_4112, w_049_4113, w_049_4114, w_049_4115, w_049_4118, w_049_4121, w_049_4122, w_049_4123, w_049_4126, w_049_4127, w_049_4131, w_049_4132, w_049_4133, w_049_4134, w_049_4135, w_049_4139, w_049_4140, w_049_4141, w_049_4142, w_049_4143, w_049_4148, w_049_4149, w_049_4150, w_049_4151, w_049_4153, w_049_4154, w_049_4155, w_049_4157, w_049_4158, w_049_4161, w_049_4162, w_049_4163, w_049_4166, w_049_4167, w_049_4171, w_049_4172, w_049_4174, w_049_4176, w_049_4178, w_049_4179, w_049_4187, w_049_4190, w_049_4195, w_049_4205, w_049_4206, w_049_4209, w_049_4210, w_049_4212, w_049_4216, w_049_4218, w_049_4220, w_049_4225, w_049_4226, w_049_4228, w_049_4229, w_049_4234, w_049_4235, w_049_4236, w_049_4237, w_049_4241, w_049_4242, w_049_4243, w_049_4245, w_049_4249, w_049_4252, w_049_4253, w_049_4254, w_049_4255, w_049_4257, w_049_4258, w_049_4260, w_049_4261, w_049_4262, w_049_4263, w_049_4264, w_049_4265, w_049_4266, w_049_4268, w_049_4270, w_049_4272, w_049_4273, w_049_4276, w_049_4277, w_049_4278, w_049_4281, w_049_4283, w_049_4289, w_049_4290, w_049_4292, w_049_4294, w_049_4295, w_049_4297, w_049_4303, w_049_4304, w_049_4306, w_049_4310, w_049_4313, w_049_4314, w_049_4317, w_049_4320, w_049_4321, w_049_4323, w_049_4324, w_049_4325, w_049_4326, w_049_4327, w_049_4328, w_049_4329, w_049_4330, w_049_4332;
  wire w_050_001, w_050_003, w_050_004, w_050_006, w_050_008, w_050_009, w_050_010, w_050_011, w_050_013, w_050_014, w_050_016, w_050_017, w_050_018, w_050_019, w_050_020, w_050_024, w_050_025, w_050_026, w_050_027, w_050_028, w_050_030, w_050_031, w_050_032, w_050_033, w_050_034, w_050_035, w_050_036, w_050_037, w_050_038, w_050_039, w_050_041, w_050_042, w_050_047, w_050_048, w_050_050, w_050_051, w_050_054, w_050_055, w_050_057, w_050_058, w_050_061, w_050_062, w_050_063, w_050_064, w_050_065, w_050_066, w_050_067, w_050_068, w_050_069, w_050_070, w_050_071, w_050_072, w_050_073, w_050_076, w_050_078, w_050_080, w_050_082, w_050_083, w_050_084, w_050_085, w_050_086, w_050_087, w_050_088, w_050_089, w_050_090, w_050_091, w_050_092, w_050_095, w_050_096, w_050_098, w_050_100, w_050_101, w_050_102, w_050_103, w_050_105, w_050_106, w_050_107, w_050_110, w_050_113, w_050_115, w_050_116, w_050_118, w_050_119, w_050_122, w_050_123, w_050_125, w_050_126, w_050_130, w_050_132, w_050_134, w_050_135, w_050_137, w_050_139, w_050_140, w_050_141, w_050_143, w_050_144, w_050_145, w_050_147, w_050_148, w_050_149, w_050_150, w_050_151, w_050_153, w_050_158, w_050_159, w_050_160, w_050_161, w_050_163, w_050_164, w_050_165, w_050_166, w_050_167, w_050_168, w_050_169, w_050_170, w_050_171, w_050_172, w_050_173, w_050_174, w_050_175, w_050_177, w_050_178, w_050_179, w_050_180, w_050_181, w_050_182, w_050_183, w_050_185, w_050_186, w_050_188, w_050_189, w_050_190, w_050_191, w_050_192, w_050_196, w_050_197, w_050_198, w_050_200, w_050_201, w_050_202, w_050_205, w_050_207, w_050_209, w_050_210, w_050_211, w_050_212, w_050_213, w_050_215, w_050_216, w_050_217, w_050_218, w_050_219, w_050_220, w_050_221, w_050_222, w_050_223, w_050_224, w_050_226, w_050_228, w_050_229, w_050_230, w_050_231, w_050_232, w_050_233, w_050_234, w_050_235, w_050_236, w_050_237, w_050_238, w_050_239, w_050_240, w_050_241, w_050_243, w_050_244, w_050_245, w_050_246, w_050_248, w_050_249, w_050_250, w_050_251, w_050_253, w_050_254, w_050_256, w_050_257, w_050_258, w_050_259, w_050_261, w_050_262, w_050_263, w_050_264, w_050_265, w_050_267, w_050_268, w_050_270, w_050_271, w_050_272, w_050_274, w_050_275, w_050_276, w_050_277, w_050_278, w_050_279, w_050_280, w_050_282, w_050_283, w_050_285, w_050_286, w_050_288, w_050_289, w_050_291, w_050_292, w_050_294, w_050_295, w_050_296, w_050_297, w_050_299, w_050_300, w_050_301, w_050_302, w_050_303, w_050_306, w_050_309, w_050_310, w_050_311, w_050_312, w_050_314, w_050_316, w_050_317, w_050_318, w_050_320, w_050_321, w_050_323, w_050_324, w_050_325, w_050_326, w_050_327, w_050_328, w_050_329, w_050_330, w_050_332, w_050_333, w_050_334, w_050_335, w_050_336, w_050_338, w_050_339, w_050_340, w_050_341, w_050_342, w_050_343, w_050_344, w_050_345, w_050_347, w_050_348, w_050_349, w_050_350, w_050_351, w_050_352, w_050_353, w_050_354, w_050_356, w_050_357, w_050_358, w_050_360, w_050_361, w_050_363, w_050_364, w_050_365, w_050_366, w_050_369, w_050_373, w_050_374, w_050_375, w_050_376, w_050_377, w_050_378, w_050_379, w_050_381, w_050_382, w_050_383, w_050_386, w_050_387, w_050_388, w_050_389, w_050_390, w_050_391, w_050_392, w_050_393, w_050_394, w_050_395, w_050_397, w_050_398, w_050_399, w_050_401, w_050_402, w_050_403, w_050_404, w_050_405, w_050_406, w_050_409, w_050_410, w_050_411, w_050_414, w_050_415, w_050_416, w_050_417, w_050_418, w_050_419, w_050_420, w_050_421, w_050_422, w_050_423, w_050_424, w_050_425, w_050_428, w_050_429, w_050_431, w_050_432, w_050_435, w_050_437, w_050_438, w_050_439, w_050_440, w_050_441, w_050_443, w_050_444, w_050_445, w_050_447, w_050_450, w_050_451, w_050_452, w_050_453, w_050_454, w_050_456, w_050_457, w_050_460, w_050_464, w_050_465, w_050_467, w_050_469, w_050_470, w_050_474, w_050_475, w_050_476, w_050_477, w_050_478, w_050_480, w_050_481, w_050_482, w_050_483, w_050_487, w_050_488, w_050_489, w_050_490, w_050_491, w_050_493, w_050_494, w_050_496, w_050_497, w_050_499, w_050_500, w_050_502, w_050_503, w_050_504, w_050_505, w_050_509, w_050_510, w_050_512, w_050_514, w_050_515, w_050_516, w_050_517, w_050_519, w_050_520, w_050_522, w_050_523, w_050_524, w_050_526, w_050_527, w_050_528, w_050_529, w_050_530, w_050_531, w_050_535, w_050_536, w_050_538, w_050_539, w_050_543, w_050_544, w_050_545, w_050_546, w_050_548, w_050_549, w_050_551, w_050_553, w_050_554, w_050_555, w_050_556, w_050_557, w_050_559, w_050_560, w_050_561, w_050_562, w_050_563, w_050_565, w_050_567, w_050_568, w_050_569, w_050_571, w_050_573, w_050_574, w_050_575, w_050_577, w_050_579, w_050_581, w_050_582, w_050_584, w_050_585, w_050_586, w_050_587, w_050_588, w_050_589, w_050_590, w_050_592, w_050_593, w_050_595, w_050_599, w_050_600, w_050_601, w_050_602, w_050_604, w_050_605, w_050_606, w_050_607, w_050_608, w_050_610, w_050_611, w_050_612, w_050_613, w_050_614, w_050_615, w_050_616, w_050_618, w_050_619, w_050_620, w_050_621, w_050_622, w_050_624, w_050_625, w_050_627, w_050_628, w_050_630, w_050_631, w_050_632, w_050_634, w_050_635, w_050_636, w_050_638, w_050_639, w_050_640, w_050_641, w_050_642, w_050_645, w_050_646, w_050_647, w_050_648, w_050_650, w_050_651, w_050_653, w_050_654, w_050_655, w_050_657, w_050_658, w_050_659, w_050_661, w_050_662, w_050_663, w_050_666, w_050_668, w_050_669, w_050_670, w_050_671, w_050_672, w_050_673, w_050_674, w_050_675, w_050_676, w_050_677, w_050_678, w_050_679, w_050_680, w_050_681, w_050_682, w_050_685, w_050_686, w_050_687, w_050_689, w_050_690, w_050_692, w_050_693, w_050_694, w_050_695, w_050_696, w_050_698, w_050_699, w_050_701, w_050_704, w_050_706, w_050_708, w_050_709, w_050_710, w_050_711, w_050_712, w_050_713, w_050_715, w_050_716, w_050_717, w_050_718, w_050_719, w_050_720, w_050_725, w_050_726, w_050_727, w_050_728, w_050_729, w_050_731, w_050_733, w_050_734, w_050_735, w_050_736, w_050_737, w_050_738, w_050_739, w_050_741, w_050_743, w_050_745, w_050_746, w_050_747, w_050_748, w_050_749, w_050_750, w_050_751, w_050_752, w_050_753, w_050_754, w_050_755, w_050_757, w_050_758, w_050_759, w_050_761, w_050_763, w_050_764, w_050_766, w_050_767, w_050_769, w_050_770, w_050_771, w_050_772, w_050_773, w_050_775, w_050_776, w_050_777, w_050_778, w_050_779, w_050_780, w_050_781, w_050_782, w_050_783, w_050_784, w_050_785, w_050_786, w_050_787, w_050_788, w_050_789, w_050_790, w_050_792, w_050_793, w_050_795, w_050_796, w_050_797, w_050_798, w_050_799, w_050_801, w_050_802, w_050_803, w_050_804, w_050_805, w_050_808, w_050_809, w_050_810, w_050_812, w_050_813, w_050_814, w_050_815, w_050_816, w_050_817, w_050_818, w_050_821, w_050_823, w_050_825, w_050_826, w_050_827, w_050_828, w_050_829, w_050_830, w_050_831, w_050_832, w_050_833, w_050_834, w_050_837, w_050_838, w_050_840, w_050_842, w_050_843, w_050_844, w_050_846, w_050_847, w_050_848, w_050_849, w_050_851, w_050_852, w_050_853, w_050_854, w_050_855, w_050_856, w_050_857, w_050_859, w_050_860, w_050_861, w_050_862, w_050_863, w_050_865, w_050_866, w_050_867, w_050_868, w_050_869, w_050_870, w_050_871, w_050_872, w_050_874, w_050_879, w_050_880, w_050_881, w_050_882, w_050_883, w_050_884, w_050_885, w_050_886, w_050_888, w_050_890, w_050_892, w_050_893, w_050_894, w_050_896, w_050_897, w_050_898, w_050_899, w_050_900, w_050_901, w_050_902, w_050_907, w_050_908, w_050_909, w_050_910, w_050_911, w_050_912, w_050_913, w_050_915, w_050_916, w_050_917, w_050_918, w_050_919, w_050_920, w_050_921, w_050_922, w_050_923, w_050_924, w_050_926, w_050_931, w_050_933, w_050_935, w_050_936, w_050_937, w_050_938, w_050_939, w_050_941, w_050_943, w_050_945, w_050_946, w_050_947, w_050_948, w_050_949, w_050_950, w_050_952, w_050_954, w_050_955, w_050_956, w_050_957, w_050_958, w_050_959, w_050_960, w_050_962, w_050_963, w_050_964, w_050_965, w_050_966, w_050_967, w_050_969, w_050_970, w_050_973, w_050_974, w_050_976, w_050_978, w_050_979, w_050_981, w_050_983, w_050_984, w_050_985, w_050_986, w_050_987, w_050_989, w_050_990, w_050_993, w_050_994, w_050_995, w_050_996, w_050_997, w_050_999, w_050_1001, w_050_1006, w_050_1008, w_050_1009, w_050_1010, w_050_1011, w_050_1012, w_050_1013, w_050_1015, w_050_1016, w_050_1017, w_050_1018, w_050_1019, w_050_1020, w_050_1021, w_050_1022, w_050_1023, w_050_1024, w_050_1025, w_050_1026, w_050_1027, w_050_1029, w_050_1030, w_050_1031, w_050_1032, w_050_1034, w_050_1037, w_050_1038, w_050_1039, w_050_1040, w_050_1041, w_050_1042, w_050_1044, w_050_1046, w_050_1048, w_050_1049, w_050_1050, w_050_1051, w_050_1052, w_050_1053, w_050_1054, w_050_1055, w_050_1059, w_050_1064, w_050_1066, w_050_1068, w_050_1069, w_050_1070, w_050_1072, w_050_1073, w_050_1074, w_050_1075, w_050_1076, w_050_1077, w_050_1078, w_050_1079, w_050_1080, w_050_1081, w_050_1083, w_050_1085, w_050_1086, w_050_1087, w_050_1088, w_050_1089, w_050_1090, w_050_1091, w_050_1092, w_050_1093, w_050_1094, w_050_1096, w_050_1097, w_050_1098, w_050_1100, w_050_1102, w_050_1103, w_050_1105, w_050_1106, w_050_1109, w_050_1111, w_050_1113, w_050_1115, w_050_1116, w_050_1117, w_050_1119, w_050_1120, w_050_1121, w_050_1122, w_050_1124, w_050_1125, w_050_1127, w_050_1129, w_050_1132, w_050_1133, w_050_1134, w_050_1136, w_050_1137, w_050_1138, w_050_1140, w_050_1142, w_050_1143, w_050_1144, w_050_1145, w_050_1147, w_050_1148, w_050_1150, w_050_1151, w_050_1152, w_050_1153, w_050_1154, w_050_1155, w_050_1157, w_050_1158, w_050_1159, w_050_1161, w_050_1162, w_050_1163, w_050_1164, w_050_1165, w_050_1166, w_050_1167, w_050_1168, w_050_1169, w_050_1172, w_050_1173, w_050_1174, w_050_1175, w_050_1176, w_050_1178, w_050_1179, w_050_1181, w_050_1183, w_050_1184, w_050_1185, w_050_1187, w_050_1188, w_050_1189, w_050_1192, w_050_1194, w_050_1197, w_050_1199, w_050_1201, w_050_1202, w_050_1204, w_050_1205, w_050_1206, w_050_1207, w_050_1208, w_050_1210, w_050_1211, w_050_1213, w_050_1214, w_050_1215, w_050_1216, w_050_1217, w_050_1219, w_050_1220, w_050_1221, w_050_1222, w_050_1224, w_050_1225, w_050_1226, w_050_1228, w_050_1229, w_050_1230, w_050_1231, w_050_1233, w_050_1234, w_050_1236, w_050_1237, w_050_1238, w_050_1241, w_050_1242, w_050_1243, w_050_1244, w_050_1245, w_050_1246, w_050_1248, w_050_1250, w_050_1251, w_050_1252, w_050_1255, w_050_1256, w_050_1257, w_050_1259, w_050_1261, w_050_1262, w_050_1264, w_050_1265, w_050_1266, w_050_1267, w_050_1269, w_050_1270, w_050_1271, w_050_1272, w_050_1273, w_050_1274, w_050_1275, w_050_1276, w_050_1277, w_050_1279, w_050_1280, w_050_1281, w_050_1282, w_050_1283, w_050_1284, w_050_1285, w_050_1286, w_050_1287, w_050_1288, w_050_1291, w_050_1292, w_050_1294, w_050_1295, w_050_1297, w_050_1298, w_050_1299, w_050_1300, w_050_1302, w_050_1303, w_050_1305, w_050_1306, w_050_1307, w_050_1308, w_050_1309, w_050_1310, w_050_1311, w_050_1312, w_050_1313, w_050_1314, w_050_1316, w_050_1317, w_050_1318, w_050_1319, w_050_1321, w_050_1322, w_050_1324, w_050_1325, w_050_1327, w_050_1328, w_050_1329, w_050_1330, w_050_1331, w_050_1333, w_050_1334, w_050_1335, w_050_1336, w_050_1339, w_050_1341, w_050_1342, w_050_1344, w_050_1345, w_050_1347, w_050_1349, w_050_1351, w_050_1353, w_050_1354, w_050_1358, w_050_1359, w_050_1361, w_050_1362, w_050_1363, w_050_1365, w_050_1368, w_050_1369, w_050_1370, w_050_1372, w_050_1373, w_050_1374, w_050_1375, w_050_1376, w_050_1378, w_050_1379, w_050_1380, w_050_1381, w_050_1384, w_050_1385, w_050_1387, w_050_1388, w_050_1389, w_050_1390, w_050_1392, w_050_1393, w_050_1394, w_050_1395, w_050_1396, w_050_1397, w_050_1398, w_050_1399, w_050_1400, w_050_1401, w_050_1402, w_050_1403, w_050_1404, w_050_1406, w_050_1407, w_050_1408, w_050_1409, w_050_1411, w_050_1414, w_050_1415, w_050_1416, w_050_1417, w_050_1418, w_050_1419, w_050_1420, w_050_1421, w_050_1422, w_050_1423, w_050_1424, w_050_1425, w_050_1426, w_050_1427, w_050_1428, w_050_1429, w_050_1430, w_050_1431, w_050_1432, w_050_1433, w_050_1435, w_050_1436, w_050_1437, w_050_1438, w_050_1439, w_050_1441, w_050_1442, w_050_1444, w_050_1445, w_050_1446, w_050_1447, w_050_1448, w_050_1449, w_050_1451, w_050_1453, w_050_1458, w_050_1459, w_050_1460, w_050_1461, w_050_1462, w_050_1464, w_050_1468, w_050_1470, w_050_1472, w_050_1473, w_050_1474, w_050_1475, w_050_1478, w_050_1479, w_050_1480, w_050_1481, w_050_1484, w_050_1486, w_050_1487, w_050_1491, w_050_1492, w_050_1493, w_050_1494, w_050_1497, w_050_1499, w_050_1500, w_050_1504, w_050_1505, w_050_1506, w_050_1507, w_050_1509, w_050_1510, w_050_1512, w_050_1514, w_050_1515, w_050_1516, w_050_1517, w_050_1518, w_050_1519, w_050_1521, w_050_1523, w_050_1524, w_050_1525, w_050_1526, w_050_1527, w_050_1528, w_050_1529, w_050_1531, w_050_1533, w_050_1534, w_050_1535, w_050_1536, w_050_1538, w_050_1539, w_050_1542, w_050_1543, w_050_1544, w_050_1547, w_050_1548, w_050_1549, w_050_1550, w_050_1552, w_050_1553, w_050_1554, w_050_1555, w_050_1557, w_050_1559, w_050_1560, w_050_1563, w_050_1564, w_050_1565, w_050_1569, w_050_1570, w_050_1571, w_050_1575, w_050_1576, w_050_1577, w_050_1578, w_050_1579, w_050_1581, w_050_1582, w_050_1583, w_050_1584, w_050_1585, w_050_1586, w_050_1589, w_050_1590, w_050_1591, w_050_1592, w_050_1593, w_050_1595, w_050_1598, w_050_1599, w_050_1600, w_050_1602, w_050_1603, w_050_1604, w_050_1605, w_050_1606, w_050_1607, w_050_1608, w_050_1609, w_050_1610, w_050_1613, w_050_1614, w_050_1615, w_050_1619, w_050_1621, w_050_1625, w_050_1626, w_050_1627, w_050_1629, w_050_1630, w_050_1631, w_050_1632, w_050_1633, w_050_1634, w_050_1636, w_050_1637, w_050_1638, w_050_1639, w_050_1640, w_050_1641, w_050_1643, w_050_1644, w_050_1645, w_050_1646, w_050_1648, w_050_1649, w_050_1650, w_050_1651, w_050_1652, w_050_1653, w_050_1654, w_050_1656, w_050_1657, w_050_1658, w_050_1659, w_050_1660, w_050_1661, w_050_1662, w_050_1663, w_050_1664, w_050_1665, w_050_1666, w_050_1667, w_050_1668, w_050_1669, w_050_1670, w_050_1671, w_050_1672, w_050_1674, w_050_1675, w_050_1676, w_050_1678, w_050_1679, w_050_1680, w_050_1681, w_050_1682, w_050_1683, w_050_1688, w_050_1689, w_050_1691, w_050_1692, w_050_1693, w_050_1694, w_050_1695, w_050_1697, w_050_1698, w_050_1700, w_050_1702, w_050_1705, w_050_1706, w_050_1707, w_050_1708, w_050_1709, w_050_1711, w_050_1712, w_050_1713, w_050_1716, w_050_1718, w_050_1719, w_050_1720, w_050_1721, w_050_1722, w_050_1723, w_050_1724, w_050_1725, w_050_1726, w_050_1727, w_050_1728, w_050_1729, w_050_1730, w_050_1731, w_050_1732, w_050_1733, w_050_1734, w_050_1735, w_050_1736, w_050_1737, w_050_1738, w_050_1740, w_050_1741, w_050_1742, w_050_1743, w_050_1744, w_050_1747, w_050_1748, w_050_1750, w_050_1751, w_050_1752, w_050_1753, w_050_1754, w_050_1755, w_050_1756, w_050_1757, w_050_1758, w_050_1759, w_050_1760, w_050_1761, w_050_1763, w_050_1765, w_050_1766, w_050_1770, w_050_1771, w_050_1772, w_050_1773, w_050_1774, w_050_1775, w_050_1776, w_050_1777, w_050_1780, w_050_1781, w_050_1784, w_050_1785, w_050_1787, w_050_1788, w_050_1792, w_050_1793, w_050_1794, w_050_1795, w_050_1797, w_050_1798, w_050_1799, w_050_1800, w_050_1802, w_050_1803, w_050_1804, w_050_1806, w_050_1808, w_050_1809, w_050_1811, w_050_1813, w_050_1814, w_050_1815, w_050_1816, w_050_1817, w_050_1818, w_050_1819, w_050_1820, w_050_1821, w_050_1822, w_050_1823, w_050_1824, w_050_1825, w_050_1826, w_050_1827, w_050_1828, w_050_1831, w_050_1833, w_050_1834, w_050_1835, w_050_1836, w_050_1839, w_050_1841, w_050_1842, w_050_1843, w_050_1845, w_050_1846, w_050_1851, w_050_1854, w_050_1855, w_050_1858, w_050_1860, w_050_1861, w_050_1862, w_050_1863, w_050_1864, w_050_1865, w_050_1866, w_050_1867, w_050_1868, w_050_1869, w_050_1871, w_050_1872, w_050_1873, w_050_1874, w_050_1875, w_050_1876, w_050_1878, w_050_1879, w_050_1881, w_050_1882, w_050_1883, w_050_1884, w_050_1886, w_050_1887, w_050_1888, w_050_1889, w_050_1891, w_050_1892, w_050_1893, w_050_1894, w_050_1895, w_050_1897, w_050_1899, w_050_1900, w_050_1901, w_050_1902, w_050_1903, w_050_1905, w_050_1906, w_050_1907, w_050_1908, w_050_1910, w_050_1912, w_050_1913, w_050_1914, w_050_1915, w_050_1917, w_050_1918, w_050_1919, w_050_1920, w_050_1921, w_050_1922, w_050_1923, w_050_1924, w_050_1925, w_050_1926, w_050_1927, w_050_1928, w_050_1929, w_050_1931, w_050_1932, w_050_1933, w_050_1934, w_050_1935, w_050_1936, w_050_1938, w_050_1939, w_050_1940, w_050_1941, w_050_1942, w_050_1943, w_050_1944, w_050_1946, w_050_1947, w_050_1948, w_050_1949, w_050_1952, w_050_1954, w_050_1955, w_050_1956, w_050_1957, w_050_1958, w_050_1959, w_050_1960, w_050_1963, w_050_1964, w_050_1965, w_050_1967, w_050_1968, w_050_1969, w_050_1970, w_050_1971, w_050_1972, w_050_1973, w_050_1974, w_050_1975, w_050_1977, w_050_1979, w_050_1980, w_050_1982, w_050_1983, w_050_1985, w_050_1988, w_050_1989, w_050_1990, w_050_1992, w_050_1994, w_050_1996, w_050_1997, w_050_1998, w_050_1999, w_050_2000, w_050_2001, w_050_2002, w_050_2003, w_050_2004, w_050_2005, w_050_2006, w_050_2007, w_050_2009, w_050_2010, w_050_2011, w_050_2012, w_050_2013, w_050_2014, w_050_2016, w_050_2017, w_050_2018, w_050_2019, w_050_2020, w_050_2023, w_050_2024, w_050_2025, w_050_2026, w_050_2027, w_050_2028, w_050_2030, w_050_2031, w_050_2034, w_050_2035, w_050_2036, w_050_2039, w_050_2040, w_050_2042, w_050_2044, w_050_2046, w_050_2050, w_050_2051, w_050_2052, w_050_2054, w_050_2056, w_050_2057, w_050_2059, w_050_2060, w_050_2061, w_050_2062, w_050_2063, w_050_2065, w_050_2066, w_050_2067, w_050_2068, w_050_2070, w_050_2071, w_050_2072, w_050_2073, w_050_2074, w_050_2075, w_050_2076, w_050_2077, w_050_2078, w_050_2079, w_050_2080, w_050_2082, w_050_2084, w_050_2085, w_050_2086, w_050_2087, w_050_2088, w_050_2090, w_050_2093, w_050_2094, w_050_2095, w_050_2097, w_050_2100, w_050_2102, w_050_2103, w_050_2104, w_050_2106, w_050_2107, w_050_2108, w_050_2109, w_050_2110, w_050_2111, w_050_2113, w_050_2114, w_050_2115, w_050_2118, w_050_2120, w_050_2122, w_050_2123, w_050_2124, w_050_2127, w_050_2128, w_050_2132, w_050_2134, w_050_2135, w_050_2136, w_050_2137, w_050_2140, w_050_2141, w_050_2142, w_050_2144, w_050_2145, w_050_2146, w_050_2148, w_050_2149, w_050_2151, w_050_2152, w_050_2154, w_050_2155, w_050_2156, w_050_2157, w_050_2158, w_050_2159, w_050_2160, w_050_2161, w_050_2162, w_050_2163, w_050_2165, w_050_2166, w_050_2167, w_050_2168, w_050_2169, w_050_2170, w_050_2171, w_050_2172, w_050_2173, w_050_2174, w_050_2177, w_050_2178, w_050_2179, w_050_2181, w_050_2182, w_050_2183, w_050_2184, w_050_2185, w_050_2186, w_050_2187, w_050_2189, w_050_2191, w_050_2192, w_050_2193, w_050_2195, w_050_2197, w_050_2198, w_050_2199, w_050_2201, w_050_2203, w_050_2205, w_050_2206, w_050_2207, w_050_2209, w_050_2210, w_050_2211, w_050_2212, w_050_2213, w_050_2214, w_050_2215, w_050_2216, w_050_2217, w_050_2218, w_050_2220, w_050_2221, w_050_2222, w_050_2223, w_050_2224, w_050_2225, w_050_2228, w_050_2229, w_050_2230, w_050_2232, w_050_2233, w_050_2235, w_050_2236, w_050_2239, w_050_2240, w_050_2241, w_050_2242, w_050_2245, w_050_2246, w_050_2247, w_050_2249, w_050_2250, w_050_2251, w_050_2252, w_050_2253, w_050_2254, w_050_2255, w_050_2256, w_050_2257, w_050_2258, w_050_2260, w_050_2261, w_050_2262, w_050_2263, w_050_2264, w_050_2265, w_050_2266, w_050_2267, w_050_2268, w_050_2269, w_050_2272, w_050_2274, w_050_2275, w_050_2279, w_050_2280, w_050_2282, w_050_2283, w_050_2284, w_050_2286, w_050_2287, w_050_2288, w_050_2289, w_050_2290, w_050_2292, w_050_2295, w_050_2296, w_050_2297, w_050_2298, w_050_2299, w_050_2300, w_050_2301, w_050_2303, w_050_2304, w_050_2308, w_050_2309, w_050_2310, w_050_2311, w_050_2312, w_050_2313, w_050_2314, w_050_2315, w_050_2316, w_050_2317, w_050_2318, w_050_2320, w_050_2321, w_050_2322, w_050_2323, w_050_2324, w_050_2326, w_050_2327, w_050_2328, w_050_2329, w_050_2331, w_050_2332, w_050_2333, w_050_2335, w_050_2336, w_050_2337, w_050_2338, w_050_2339, w_050_2340, w_050_2341, w_050_2342, w_050_2343, w_050_2344, w_050_2345, w_050_2346, w_050_2347, w_050_2348, w_050_2349, w_050_2350, w_050_2351, w_050_2352, w_050_2353, w_050_2354, w_050_2356, w_050_2357, w_050_2358, w_050_2362, w_050_2363, w_050_2364, w_050_2367, w_050_2369, w_050_2370, w_050_2371, w_050_2374, w_050_2375, w_050_2379, w_050_2380, w_050_2381, w_050_2384, w_050_2385, w_050_2386, w_050_2387, w_050_2388, w_050_2389, w_050_2390, w_050_2391, w_050_2393, w_050_2394, w_050_2395, w_050_2396, w_050_2398, w_050_2400, w_050_2401, w_050_2403, w_050_2405, w_050_2406, w_050_2409, w_050_2410, w_050_2412, w_050_2413, w_050_2414, w_050_2415, w_050_2416, w_050_2417, w_050_2419, w_050_2420, w_050_2421, w_050_2424, w_050_2426, w_050_2427, w_050_2429, w_050_2430, w_050_2431, w_050_2433, w_050_2434, w_050_2435, w_050_2436, w_050_2437, w_050_2438, w_050_2440, w_050_2442, w_050_2443, w_050_2444, w_050_2446, w_050_2447, w_050_2448, w_050_2450, w_050_2453, w_050_2454, w_050_2455, w_050_2456, w_050_2457, w_050_2459, w_050_2460, w_050_2464, w_050_2465, w_050_2466, w_050_2467, w_050_2468, w_050_2469, w_050_2470, w_050_2471, w_050_2472, w_050_2476, w_050_2477, w_050_2479, w_050_2480, w_050_2481, w_050_2482, w_050_2483, w_050_2487, w_050_2489, w_050_2490, w_050_2491, w_050_2492, w_050_2494, w_050_2502, w_050_2504, w_050_2506, w_050_2507, w_050_2510, w_050_2511, w_050_2512, w_050_2513, w_050_2514, w_050_2515, w_050_2516, w_050_2517, w_050_2518, w_050_2519, w_050_2520, w_050_2521, w_050_2525, w_050_2526, w_050_2527, w_050_2528, w_050_2529, w_050_2530, w_050_2531, w_050_2532, w_050_2533, w_050_2534, w_050_2535, w_050_2537;
  wire w_051_002, w_051_004, w_051_005, w_051_006, w_051_007, w_051_008, w_051_010, w_051_011, w_051_012, w_051_013, w_051_015, w_051_017, w_051_018, w_051_019, w_051_020, w_051_022, w_051_023, w_051_024, w_051_026, w_051_027, w_051_028, w_051_029, w_051_030, w_051_031, w_051_033, w_051_036, w_051_037, w_051_038, w_051_039, w_051_041, w_051_044, w_051_045, w_051_046, w_051_048, w_051_049, w_051_050, w_051_051, w_051_053, w_051_055, w_051_056, w_051_057, w_051_060, w_051_061, w_051_063, w_051_065, w_051_066, w_051_067, w_051_068, w_051_069, w_051_070, w_051_071, w_051_072, w_051_073, w_051_074, w_051_075, w_051_076, w_051_078, w_051_079, w_051_081, w_051_082, w_051_083, w_051_084, w_051_087, w_051_088, w_051_090, w_051_092, w_051_093, w_051_094, w_051_096, w_051_097, w_051_099, w_051_100, w_051_102, w_051_103, w_051_104, w_051_106, w_051_107, w_051_108, w_051_109, w_051_110, w_051_111, w_051_112, w_051_114, w_051_116, w_051_118, w_051_119, w_051_120, w_051_121, w_051_122, w_051_123, w_051_125, w_051_126, w_051_129, w_051_131, w_051_133, w_051_134, w_051_135, w_051_137, w_051_138, w_051_140, w_051_141, w_051_142, w_051_143, w_051_144, w_051_145, w_051_146, w_051_147, w_051_149, w_051_150, w_051_151, w_051_152, w_051_155, w_051_157, w_051_158, w_051_159, w_051_160, w_051_161, w_051_162, w_051_163, w_051_164, w_051_165, w_051_166, w_051_167, w_051_169, w_051_170, w_051_171, w_051_172, w_051_173, w_051_174, w_051_177, w_051_178, w_051_180, w_051_181, w_051_182, w_051_184, w_051_185, w_051_188, w_051_190, w_051_191, w_051_193, w_051_194, w_051_195, w_051_196, w_051_197, w_051_201, w_051_202, w_051_203, w_051_207, w_051_208, w_051_209, w_051_211, w_051_212, w_051_213, w_051_215, w_051_216, w_051_217, w_051_218, w_051_219, w_051_220, w_051_223, w_051_224, w_051_225, w_051_226, w_051_229, w_051_230, w_051_231, w_051_232, w_051_233, w_051_234, w_051_237, w_051_239, w_051_240, w_051_241, w_051_242, w_051_243, w_051_244, w_051_245, w_051_246, w_051_247, w_051_249, w_051_250, w_051_251, w_051_252, w_051_254, w_051_256, w_051_258, w_051_259, w_051_260, w_051_261, w_051_262, w_051_264, w_051_265, w_051_266, w_051_268, w_051_269, w_051_270, w_051_271, w_051_272, w_051_273, w_051_274, w_051_275, w_051_276, w_051_277, w_051_278, w_051_279, w_051_281, w_051_282, w_051_283, w_051_284, w_051_285, w_051_287, w_051_288, w_051_289, w_051_290, w_051_292, w_051_293, w_051_294, w_051_295, w_051_296, w_051_297, w_051_301, w_051_302, w_051_303, w_051_304, w_051_305, w_051_306, w_051_307, w_051_308, w_051_310, w_051_312, w_051_313, w_051_314, w_051_315, w_051_316, w_051_317, w_051_318, w_051_319, w_051_321, w_051_322, w_051_323, w_051_324, w_051_325, w_051_326, w_051_327, w_051_328, w_051_329, w_051_330, w_051_334, w_051_335, w_051_336, w_051_338, w_051_339, w_051_340, w_051_341, w_051_342, w_051_343, w_051_346, w_051_349, w_051_350, w_051_351, w_051_352, w_051_353, w_051_355, w_051_356, w_051_358, w_051_361, w_051_362, w_051_363, w_051_364, w_051_368, w_051_370, w_051_373, w_051_374, w_051_375, w_051_377, w_051_378, w_051_379, w_051_383, w_051_384, w_051_385, w_051_386, w_051_388, w_051_390, w_051_394, w_051_396, w_051_397, w_051_398, w_051_400, w_051_404, w_051_405, w_051_409, w_051_410, w_051_412, w_051_413, w_051_414, w_051_415, w_051_416, w_051_417, w_051_418, w_051_420, w_051_423, w_051_425, w_051_426, w_051_427, w_051_428, w_051_429, w_051_430, w_051_432, w_051_434, w_051_436, w_051_437, w_051_438, w_051_439, w_051_441, w_051_442, w_051_445, w_051_447, w_051_449, w_051_451, w_051_452, w_051_456, w_051_457, w_051_458, w_051_460, w_051_462, w_051_463, w_051_464, w_051_465, w_051_468, w_051_469, w_051_473, w_051_474, w_051_475, w_051_476, w_051_477, w_051_479, w_051_480, w_051_481, w_051_483, w_051_484, w_051_485, w_051_487, w_051_488, w_051_489, w_051_490, w_051_491, w_051_493, w_051_494, w_051_495, w_051_496, w_051_497, w_051_498, w_051_499, w_051_500, w_051_502, w_051_503, w_051_504, w_051_508, w_051_509, w_051_511, w_051_512, w_051_513, w_051_514, w_051_515, w_051_516, w_051_517, w_051_518, w_051_519, w_051_520, w_051_522, w_051_523, w_051_524, w_051_526, w_051_527, w_051_528, w_051_529, w_051_531, w_051_532, w_051_533, w_051_536, w_051_540, w_051_541, w_051_542, w_051_543, w_051_544, w_051_545, w_051_546, w_051_548, w_051_552, w_051_553, w_051_554, w_051_555, w_051_557, w_051_559, w_051_561, w_051_564, w_051_565, w_051_566, w_051_567, w_051_569, w_051_571, w_051_572, w_051_573, w_051_574, w_051_575, w_051_576, w_051_578, w_051_579, w_051_580, w_051_581, w_051_583, w_051_584, w_051_586, w_051_588, w_051_589, w_051_590, w_051_591, w_051_592, w_051_593, w_051_594, w_051_595, w_051_597, w_051_599, w_051_600, w_051_603, w_051_604, w_051_605, w_051_609, w_051_610, w_051_611, w_051_613, w_051_614, w_051_616, w_051_617, w_051_618, w_051_620, w_051_623, w_051_625, w_051_626, w_051_629, w_051_630, w_051_632, w_051_634, w_051_636, w_051_639, w_051_640, w_051_641, w_051_642, w_051_644, w_051_645, w_051_646, w_051_647, w_051_648, w_051_649, w_051_650, w_051_651, w_051_652, w_051_658, w_051_659, w_051_661, w_051_662, w_051_663, w_051_665, w_051_666, w_051_667, w_051_671, w_051_672, w_051_673, w_051_675, w_051_677, w_051_678, w_051_679, w_051_680, w_051_681, w_051_682, w_051_683, w_051_684, w_051_685, w_051_686, w_051_688, w_051_689, w_051_690, w_051_692, w_051_693, w_051_694, w_051_695, w_051_696, w_051_697, w_051_700, w_051_701, w_051_702, w_051_703, w_051_704, w_051_706, w_051_707, w_051_708, w_051_710, w_051_712, w_051_713, w_051_714, w_051_716, w_051_717, w_051_719, w_051_720, w_051_721, w_051_722, w_051_723, w_051_725, w_051_726, w_051_728, w_051_729, w_051_730, w_051_731, w_051_734, w_051_735, w_051_736, w_051_737, w_051_738, w_051_740, w_051_741, w_051_742, w_051_743, w_051_745, w_051_746, w_051_747, w_051_749, w_051_751, w_051_753, w_051_754, w_051_755, w_051_757, w_051_761, w_051_762, w_051_763, w_051_764, w_051_766, w_051_767, w_051_768, w_051_769, w_051_771, w_051_772, w_051_773, w_051_774, w_051_775, w_051_776, w_051_778, w_051_779, w_051_780, w_051_781, w_051_782, w_051_783, w_051_784, w_051_785, w_051_787, w_051_788, w_051_789, w_051_790, w_051_792, w_051_793, w_051_795, w_051_796, w_051_797, w_051_798, w_051_799, w_051_800, w_051_801, w_051_802, w_051_803, w_051_804, w_051_806, w_051_807, w_051_808, w_051_809, w_051_810, w_051_811, w_051_812, w_051_813, w_051_814, w_051_815, w_051_816, w_051_817, w_051_818, w_051_819, w_051_820, w_051_821, w_051_822, w_051_823, w_051_824, w_051_827, w_051_830, w_051_831, w_051_832, w_051_833, w_051_835, w_051_836, w_051_838, w_051_839, w_051_840, w_051_841, w_051_845, w_051_846, w_051_847, w_051_849, w_051_850, w_051_851, w_051_852, w_051_853, w_051_855, w_051_856, w_051_857, w_051_858, w_051_859, w_051_861, w_051_862, w_051_863, w_051_864, w_051_867, w_051_869, w_051_870, w_051_871, w_051_872, w_051_873, w_051_875, w_051_876, w_051_877, w_051_878, w_051_881, w_051_884, w_051_885, w_051_886, w_051_887, w_051_888, w_051_889, w_051_891, w_051_892, w_051_894, w_051_895, w_051_896, w_051_897, w_051_899, w_051_901, w_051_903, w_051_904, w_051_906, w_051_908, w_051_910, w_051_911, w_051_912, w_051_913, w_051_914, w_051_915, w_051_916, w_051_917, w_051_918, w_051_921, w_051_922, w_051_923, w_051_924, w_051_925, w_051_926, w_051_927, w_051_928, w_051_929, w_051_930, w_051_931, w_051_932, w_051_934, w_051_937, w_051_938, w_051_939, w_051_940, w_051_942, w_051_943, w_051_944, w_051_945, w_051_946, w_051_947, w_051_948, w_051_951, w_051_953, w_051_954, w_051_955, w_051_956, w_051_957, w_051_959, w_051_960, w_051_961, w_051_962, w_051_965, w_051_966, w_051_967, w_051_968, w_051_969, w_051_970, w_051_971, w_051_972, w_051_973, w_051_975, w_051_976, w_051_977, w_051_978, w_051_979, w_051_980, w_051_981, w_051_982, w_051_983, w_051_984, w_051_986, w_051_987, w_051_988, w_051_989, w_051_990, w_051_991, w_051_993, w_051_994, w_051_995, w_051_997, w_051_998, w_051_999, w_051_1000, w_051_1002, w_051_1005, w_051_1009, w_051_1010, w_051_1012, w_051_1014, w_051_1017, w_051_1019, w_051_1021, w_051_1022, w_051_1023, w_051_1024, w_051_1025, w_051_1026, w_051_1027, w_051_1029, w_051_1030, w_051_1031, w_051_1032, w_051_1034, w_051_1036, w_051_1037, w_051_1038, w_051_1039, w_051_1040, w_051_1043, w_051_1044, w_051_1045, w_051_1046, w_051_1047, w_051_1048, w_051_1049, w_051_1050, w_051_1052, w_051_1055, w_051_1056, w_051_1057, w_051_1058, w_051_1059, w_051_1061, w_051_1062, w_051_1063, w_051_1064, w_051_1068, w_051_1069, w_051_1070, w_051_1071, w_051_1072, w_051_1073, w_051_1074, w_051_1075, w_051_1079, w_051_1083, w_051_1085, w_051_1086, w_051_1088, w_051_1089, w_051_1091, w_051_1092, w_051_1093, w_051_1096, w_051_1097, w_051_1099, w_051_1100, w_051_1101, w_051_1102, w_051_1103, w_051_1108, w_051_1109, w_051_1110, w_051_1112, w_051_1113, w_051_1114, w_051_1115, w_051_1116, w_051_1117, w_051_1120, w_051_1123, w_051_1124, w_051_1125, w_051_1126, w_051_1127, w_051_1128, w_051_1130, w_051_1131, w_051_1132, w_051_1133, w_051_1134, w_051_1135, w_051_1136, w_051_1137, w_051_1138, w_051_1139, w_051_1140, w_051_1141, w_051_1142, w_051_1143, w_051_1144, w_051_1145, w_051_1146, w_051_1148, w_051_1149, w_051_1150, w_051_1151, w_051_1153, w_051_1154, w_051_1157, w_051_1158, w_051_1159, w_051_1160, w_051_1162, w_051_1163, w_051_1164, w_051_1165, w_051_1166, w_051_1169, w_051_1171, w_051_1173, w_051_1174, w_051_1175, w_051_1177, w_051_1178, w_051_1181, w_051_1182, w_051_1183, w_051_1185, w_051_1186, w_051_1188, w_051_1189, w_051_1190, w_051_1192, w_051_1193, w_051_1194, w_051_1197, w_051_1198, w_051_1199, w_051_1200, w_051_1201, w_051_1203, w_051_1204, w_051_1206, w_051_1207, w_051_1210, w_051_1211, w_051_1212, w_051_1213, w_051_1214, w_051_1218, w_051_1220, w_051_1221, w_051_1222, w_051_1223, w_051_1226, w_051_1227, w_051_1228, w_051_1229, w_051_1230, w_051_1231, w_051_1232, w_051_1233, w_051_1234, w_051_1237, w_051_1238, w_051_1239, w_051_1240, w_051_1243, w_051_1244, w_051_1245, w_051_1246, w_051_1248, w_051_1249, w_051_1250, w_051_1251, w_051_1253, w_051_1254, w_051_1255, w_051_1256, w_051_1259, w_051_1260, w_051_1261, w_051_1262, w_051_1263, w_051_1264, w_051_1265, w_051_1268, w_051_1269, w_051_1270, w_051_1271, w_051_1273, w_051_1274, w_051_1276, w_051_1277, w_051_1278, w_051_1280, w_051_1283, w_051_1284, w_051_1285, w_051_1286, w_051_1287, w_051_1288, w_051_1289, w_051_1292, w_051_1293, w_051_1294, w_051_1295, w_051_1297, w_051_1298, w_051_1299, w_051_1301, w_051_1302, w_051_1303, w_051_1305, w_051_1306, w_051_1307, w_051_1308, w_051_1309, w_051_1310, w_051_1312, w_051_1313, w_051_1316, w_051_1318, w_051_1319, w_051_1321, w_051_1322, w_051_1325, w_051_1328, w_051_1330, w_051_1331, w_051_1332, w_051_1334, w_051_1335, w_051_1336, w_051_1338, w_051_1339, w_051_1340, w_051_1341, w_051_1343, w_051_1345, w_051_1347, w_051_1348, w_051_1349, w_051_1351, w_051_1353, w_051_1355, w_051_1356, w_051_1357, w_051_1358, w_051_1359, w_051_1360, w_051_1361, w_051_1362, w_051_1363, w_051_1365, w_051_1368, w_051_1369, w_051_1373, w_051_1374, w_051_1376, w_051_1377, w_051_1379, w_051_1380, w_051_1381, w_051_1382, w_051_1383, w_051_1384, w_051_1385, w_051_1386, w_051_1387, w_051_1389, w_051_1390, w_051_1391, w_051_1392, w_051_1393, w_051_1395, w_051_1396, w_051_1399, w_051_1400, w_051_1401, w_051_1403, w_051_1407, w_051_1410, w_051_1412, w_051_1413, w_051_1414, w_051_1415, w_051_1416, w_051_1417, w_051_1419, w_051_1420, w_051_1422, w_051_1423, w_051_1424, w_051_1425, w_051_1426, w_051_1427, w_051_1428, w_051_1429, w_051_1430, w_051_1431, w_051_1432, w_051_1433, w_051_1434, w_051_1435, w_051_1436, w_051_1437, w_051_1438, w_051_1439, w_051_1440, w_051_1441, w_051_1443, w_051_1444, w_051_1445, w_051_1446, w_051_1447, w_051_1448, w_051_1450, w_051_1451, w_051_1452, w_051_1453, w_051_1455, w_051_1456, w_051_1457, w_051_1459, w_051_1461, w_051_1463, w_051_1464, w_051_1465, w_051_1467, w_051_1468, w_051_1469, w_051_1470, w_051_1471, w_051_1472, w_051_1473, w_051_1474, w_051_1475, w_051_1476, w_051_1477, w_051_1478, w_051_1479, w_051_1480, w_051_1482, w_051_1483, w_051_1484, w_051_1488, w_051_1489, w_051_1490, w_051_1491, w_051_1493, w_051_1494, w_051_1496, w_051_1497, w_051_1498, w_051_1499, w_051_1500, w_051_1501, w_051_1502, w_051_1503, w_051_1505, w_051_1508, w_051_1509, w_051_1510, w_051_1511, w_051_1512, w_051_1513, w_051_1514, w_051_1515, w_051_1516, w_051_1517, w_051_1520, w_051_1521, w_051_1522, w_051_1525, w_051_1526, w_051_1528, w_051_1529, w_051_1530, w_051_1531, w_051_1533, w_051_1535, w_051_1537, w_051_1538, w_051_1539, w_051_1540, w_051_1541, w_051_1542, w_051_1543, w_051_1544, w_051_1545, w_051_1546, w_051_1547, w_051_1548, w_051_1549, w_051_1551, w_051_1554, w_051_1555, w_051_1556, w_051_1558, w_051_1559, w_051_1562, w_051_1563, w_051_1564, w_051_1565, w_051_1567, w_051_1568, w_051_1569, w_051_1570, w_051_1571, w_051_1574, w_051_1577, w_051_1579, w_051_1581, w_051_1583, w_051_1585, w_051_1586, w_051_1587, w_051_1589, w_051_1590, w_051_1591, w_051_1592, w_051_1593, w_051_1594, w_051_1596, w_051_1597, w_051_1598, w_051_1599, w_051_1602, w_051_1603, w_051_1605, w_051_1606, w_051_1607, w_051_1608, w_051_1609, w_051_1610, w_051_1611, w_051_1612, w_051_1613, w_051_1614, w_051_1615, w_051_1616, w_051_1618, w_051_1619, w_051_1620, w_051_1621, w_051_1622, w_051_1623, w_051_1624, w_051_1625, w_051_1626, w_051_1627, w_051_1629, w_051_1631, w_051_1632, w_051_1634, w_051_1635, w_051_1636, w_051_1637, w_051_1638, w_051_1639, w_051_1640, w_051_1641, w_051_1642, w_051_1643, w_051_1644, w_051_1645, w_051_1648, w_051_1650, w_051_1652, w_051_1654, w_051_1655, w_051_1656, w_051_1657, w_051_1658, w_051_1659, w_051_1661, w_051_1662, w_051_1663, w_051_1664, w_051_1665, w_051_1666, w_051_1668, w_051_1669, w_051_1670, w_051_1675, w_051_1676, w_051_1677, w_051_1678, w_051_1679, w_051_1681, w_051_1682, w_051_1684, w_051_1685, w_051_1686, w_051_1687, w_051_1688, w_051_1689, w_051_1690, w_051_1691, w_051_1692, w_051_1694, w_051_1695, w_051_1696, w_051_1697, w_051_1698, w_051_1699, w_051_1700, w_051_1701, w_051_1702, w_051_1705, w_051_1706, w_051_1707, w_051_1708, w_051_1709, w_051_1710, w_051_1712, w_051_1714, w_051_1715, w_051_1716, w_051_1717, w_051_1718, w_051_1720, w_051_1721, w_051_1722, w_051_1723, w_051_1724, w_051_1727, w_051_1728, w_051_1730, w_051_1731, w_051_1732, w_051_1733, w_051_1734, w_051_1735, w_051_1736, w_051_1738, w_051_1742, w_051_1745, w_051_1746, w_051_1747, w_051_1749, w_051_1750, w_051_1753, w_051_1754, w_051_1757, w_051_1758, w_051_1759, w_051_1762, w_051_1764, w_051_1765, w_051_1766, w_051_1768, w_051_1769, w_051_1770, w_051_1772, w_051_1774, w_051_1775, w_051_1776, w_051_1777, w_051_1779, w_051_1780, w_051_1781, w_051_1786, w_051_1787, w_051_1789, w_051_1790, w_051_1791, w_051_1792, w_051_1793, w_051_1794, w_051_1795, w_051_1796, w_051_1797, w_051_1798, w_051_1799, w_051_1801, w_051_1802, w_051_1803, w_051_1804, w_051_1805, w_051_1806, w_051_1807, w_051_1808, w_051_1809, w_051_1810, w_051_1811, w_051_1812, w_051_1813, w_051_1814, w_051_1815, w_051_1817, w_051_1818, w_051_1819, w_051_1820, w_051_1822, w_051_1824, w_051_1825, w_051_1827, w_051_1829, w_051_1830, w_051_1831, w_051_1832, w_051_1834, w_051_1835, w_051_1836, w_051_1837, w_051_1838, w_051_1840, w_051_1843, w_051_1846, w_051_1850, w_051_1851, w_051_1852, w_051_1853, w_051_1854, w_051_1855, w_051_1856, w_051_1857, w_051_1858, w_051_1859, w_051_1860, w_051_1861, w_051_1862, w_051_1863, w_051_1864, w_051_1867, w_051_1868, w_051_1869, w_051_1870, w_051_1871, w_051_1873, w_051_1874, w_051_1876, w_051_1878, w_051_1879, w_051_1880, w_051_1881, w_051_1882, w_051_1883, w_051_1884, w_051_1885, w_051_1886, w_051_1888, w_051_1890, w_051_1891, w_051_1893, w_051_1894, w_051_1896, w_051_1897, w_051_1898, w_051_1899, w_051_1900, w_051_1901, w_051_1902, w_051_1904, w_051_1905, w_051_1906, w_051_1907, w_051_1908, w_051_1912, w_051_1913, w_051_1914, w_051_1915, w_051_1916, w_051_1918, w_051_1919, w_051_1921, w_051_1923, w_051_1925, w_051_1927, w_051_1928, w_051_1929, w_051_1931, w_051_1932, w_051_1933, w_051_1934, w_051_1936, w_051_1938, w_051_1939, w_051_1940, w_051_1942, w_051_1943, w_051_1944, w_051_1945, w_051_1946, w_051_1947, w_051_1948, w_051_1949, w_051_1950, w_051_1951, w_051_1952, w_051_1953, w_051_1954, w_051_1955, w_051_1956, w_051_1957, w_051_1958, w_051_1959, w_051_1960, w_051_1961, w_051_1964, w_051_1965, w_051_1966, w_051_1967, w_051_1969, w_051_1970, w_051_1971, w_051_1972, w_051_1973, w_051_1975, w_051_1977, w_051_1978, w_051_1979, w_051_1980, w_051_1981, w_051_1982, w_051_1985, w_051_1986, w_051_1987, w_051_1988, w_051_1992, w_051_1993, w_051_1994, w_051_1995, w_051_1996, w_051_1997, w_051_1998, w_051_1999, w_051_2000, w_051_2001, w_051_2003, w_051_2004, w_051_2005, w_051_2007, w_051_2008, w_051_2009, w_051_2010, w_051_2013, w_051_2015, w_051_2017, w_051_2018, w_051_2019, w_051_2020, w_051_2021, w_051_2022, w_051_2023, w_051_2024, w_051_2025, w_051_2029, w_051_2030, w_051_2031, w_051_2032, w_051_2034, w_051_2035, w_051_2036, w_051_2037, w_051_2038, w_051_2043, w_051_2044, w_051_2045, w_051_2046, w_051_2047, w_051_2048, w_051_2050, w_051_2053, w_051_2054, w_051_2056, w_051_2057, w_051_2058, w_051_2061, w_051_2062, w_051_2063, w_051_2065, w_051_2066, w_051_2067, w_051_2068, w_051_2069, w_051_2070, w_051_2071, w_051_2072, w_051_2073, w_051_2074, w_051_2075, w_051_2076, w_051_2077, w_051_2078, w_051_2079, w_051_2080, w_051_2081, w_051_2082, w_051_2083, w_051_2084, w_051_2086, w_051_2087, w_051_2088, w_051_2089, w_051_2091, w_051_2093, w_051_2095, w_051_2096, w_051_2097, w_051_2098, w_051_2099, w_051_2100, w_051_2101, w_051_2102, w_051_2103, w_051_2104, w_051_2106, w_051_2107, w_051_2108, w_051_2109, w_051_2110, w_051_2112, w_051_2114, w_051_2115, w_051_2116, w_051_2117, w_051_2118, w_051_2119, w_051_2120, w_051_2121, w_051_2122, w_051_2124, w_051_2125, w_051_2126, w_051_2127, w_051_2128, w_051_2129, w_051_2132, w_051_2133, w_051_2134, w_051_2135, w_051_2136, w_051_2137, w_051_2138, w_051_2140, w_051_2141, w_051_2142, w_051_2143, w_051_2144, w_051_2145, w_051_2146, w_051_2150, w_051_2151, w_051_2152, w_051_2153, w_051_2154, w_051_2155, w_051_2156, w_051_2158, w_051_2159, w_051_2163, w_051_2164, w_051_2165, w_051_2166, w_051_2168, w_051_2170, w_051_2171, w_051_2174, w_051_2175, w_051_2176, w_051_2178, w_051_2179, w_051_2180, w_051_2181, w_051_2182, w_051_2183, w_051_2184, w_051_2187, w_051_2189, w_051_2194, w_051_2195, w_051_2197, w_051_2198, w_051_2199, w_051_2200, w_051_2202, w_051_2203, w_051_2204, w_051_2206, w_051_2208, w_051_2210, w_051_2211, w_051_2212, w_051_2213, w_051_2214, w_051_2216, w_051_2217, w_051_2219, w_051_2220, w_051_2221, w_051_2222, w_051_2223, w_051_2224, w_051_2226, w_051_2227, w_051_2228, w_051_2229, w_051_2231, w_051_2232, w_051_2234, w_051_2235, w_051_2236, w_051_2237, w_051_2238, w_051_2239, w_051_2240, w_051_2241, w_051_2242, w_051_2243, w_051_2245, w_051_2246, w_051_2247, w_051_2249, w_051_2252, w_051_2254, w_051_2255, w_051_2256, w_051_2257, w_051_2258, w_051_2259, w_051_2260, w_051_2261, w_051_2262, w_051_2263, w_051_2264, w_051_2265, w_051_2266, w_051_2267, w_051_2268, w_051_2270, w_051_2271, w_051_2272, w_051_2276, w_051_2279, w_051_2282, w_051_2283, w_051_2284, w_051_2285, w_051_2286, w_051_2287, w_051_2288, w_051_2291, w_051_2292, w_051_2293, w_051_2295, w_051_2296, w_051_2298, w_051_2299, w_051_2301, w_051_2302, w_051_2303, w_051_2304, w_051_2305, w_051_2306, w_051_2307, w_051_2308, w_051_2309, w_051_2310, w_051_2311, w_051_2312, w_051_2313, w_051_2314, w_051_2315, w_051_2321, w_051_2325, w_051_2327, w_051_2328, w_051_2332, w_051_2333, w_051_2334, w_051_2336, w_051_2337, w_051_2340, w_051_2343, w_051_2344, w_051_2346, w_051_2347, w_051_2348, w_051_2349, w_051_2350, w_051_2352, w_051_2355, w_051_2357, w_051_2365, w_051_2366, w_051_2368, w_051_2369, w_051_2375, w_051_2377, w_051_2379, w_051_2384, w_051_2385, w_051_2386, w_051_2387, w_051_2388, w_051_2392, w_051_2393, w_051_2394, w_051_2396, w_051_2399, w_051_2400, w_051_2401, w_051_2402, w_051_2405, w_051_2406, w_051_2411, w_051_2414, w_051_2416, w_051_2418, w_051_2420, w_051_2421, w_051_2422, w_051_2423, w_051_2424, w_051_2425, w_051_2426, w_051_2428, w_051_2429, w_051_2430, w_051_2431, w_051_2432, w_051_2433, w_051_2436, w_051_2439, w_051_2440, w_051_2441, w_051_2443, w_051_2445, w_051_2449, w_051_2451, w_051_2452, w_051_2460, w_051_2466, w_051_2467, w_051_2469, w_051_2475, w_051_2478, w_051_2480, w_051_2481, w_051_2482, w_051_2484, w_051_2488, w_051_2489, w_051_2491, w_051_2494, w_051_2497, w_051_2498, w_051_2499, w_051_2501, w_051_2503, w_051_2508, w_051_2514, w_051_2515, w_051_2516, w_051_2522, w_051_2523, w_051_2527, w_051_2531, w_051_2532, w_051_2535, w_051_2540, w_051_2548, w_051_2549, w_051_2552, w_051_2554, w_051_2555, w_051_2556, w_051_2557, w_051_2559, w_051_2566, w_051_2575, w_051_2580, w_051_2581, w_051_2583, w_051_2585, w_051_2586, w_051_2587, w_051_2590, w_051_2591, w_051_2592, w_051_2593, w_051_2595, w_051_2598, w_051_2599, w_051_2601, w_051_2602, w_051_2606, w_051_2608, w_051_2610, w_051_2611, w_051_2613, w_051_2614, w_051_2616, w_051_2618, w_051_2619, w_051_2629, w_051_2631, w_051_2632, w_051_2635, w_051_2637, w_051_2642, w_051_2647, w_051_2649, w_051_2650, w_051_2651, w_051_2652, w_051_2653, w_051_2654, w_051_2655, w_051_2657, w_051_2659, w_051_2665, w_051_2666, w_051_2667, w_051_2668, w_051_2669, w_051_2671, w_051_2672, w_051_2673, w_051_2674, w_051_2675, w_051_2676, w_051_2678, w_051_2682, w_051_2683, w_051_2684, w_051_2686, w_051_2687, w_051_2688, w_051_2689, w_051_2691, w_051_2693, w_051_2694, w_051_2695, w_051_2696, w_051_2698, w_051_2700, w_051_2701, w_051_2702, w_051_2703, w_051_2704, w_051_2705, w_051_2706, w_051_2707, w_051_2711, w_051_2712, w_051_2713, w_051_2714, w_051_2715, w_051_2716, w_051_2717, w_051_2718, w_051_2720;
  wire w_052_002, w_052_003, w_052_005, w_052_006, w_052_007, w_052_008, w_052_009, w_052_011, w_052_012, w_052_013, w_052_014, w_052_015, w_052_016, w_052_017, w_052_020, w_052_021, w_052_022, w_052_023, w_052_024, w_052_025, w_052_026, w_052_027, w_052_028, w_052_029, w_052_030, w_052_031, w_052_032, w_052_033, w_052_034, w_052_035, w_052_036, w_052_037, w_052_038, w_052_040, w_052_041, w_052_042, w_052_044, w_052_045, w_052_046, w_052_047, w_052_049, w_052_051, w_052_052, w_052_053, w_052_055, w_052_056, w_052_058, w_052_059, w_052_060, w_052_063, w_052_064, w_052_065, w_052_066, w_052_067, w_052_069, w_052_071, w_052_072, w_052_073, w_052_074, w_052_075, w_052_077, w_052_078, w_052_079, w_052_082, w_052_083, w_052_090, w_052_093, w_052_096, w_052_100, w_052_101, w_052_104, w_052_105, w_052_106, w_052_107, w_052_108, w_052_110, w_052_111, w_052_112, w_052_115, w_052_116, w_052_120, w_052_122, w_052_125, w_052_126, w_052_127, w_052_128, w_052_129, w_052_130, w_052_132, w_052_140, w_052_143, w_052_146, w_052_147, w_052_148, w_052_149, w_052_150, w_052_151, w_052_153, w_052_155, w_052_161, w_052_171, w_052_172, w_052_173, w_052_174, w_052_179, w_052_180, w_052_182, w_052_189, w_052_190, w_052_196, w_052_199, w_052_200, w_052_201, w_052_202, w_052_207, w_052_209, w_052_210, w_052_211, w_052_212, w_052_213, w_052_216, w_052_218, w_052_219, w_052_223, w_052_227, w_052_228, w_052_230, w_052_233, w_052_234, w_052_235, w_052_236, w_052_237, w_052_238, w_052_239, w_052_240, w_052_241, w_052_243, w_052_244, w_052_247, w_052_248, w_052_250, w_052_251, w_052_252, w_052_255, w_052_257, w_052_259, w_052_261, w_052_263, w_052_264, w_052_265, w_052_267, w_052_268, w_052_269, w_052_271, w_052_272, w_052_275, w_052_277, w_052_278, w_052_279, w_052_281, w_052_284, w_052_285, w_052_288, w_052_291, w_052_292, w_052_294, w_052_303, w_052_306, w_052_307, w_052_308, w_052_310, w_052_313, w_052_316, w_052_317, w_052_320, w_052_321, w_052_323, w_052_324, w_052_325, w_052_326, w_052_327, w_052_330, w_052_331, w_052_335, w_052_337, w_052_338, w_052_339, w_052_340, w_052_341, w_052_343, w_052_345, w_052_346, w_052_347, w_052_348, w_052_350, w_052_354, w_052_356, w_052_358, w_052_362, w_052_365, w_052_366, w_052_367, w_052_370, w_052_371, w_052_378, w_052_379, w_052_380, w_052_382, w_052_383, w_052_384, w_052_385, w_052_386, w_052_389, w_052_390, w_052_391, w_052_392, w_052_393, w_052_394, w_052_395, w_052_396, w_052_400, w_052_401, w_052_405, w_052_407, w_052_408, w_052_412, w_052_414, w_052_418, w_052_420, w_052_421, w_052_423, w_052_426, w_052_433, w_052_434, w_052_435, w_052_436, w_052_443, w_052_445, w_052_446, w_052_447, w_052_449, w_052_450, w_052_453, w_052_454, w_052_457, w_052_465, w_052_467, w_052_469, w_052_470, w_052_475, w_052_481, w_052_482, w_052_484, w_052_485, w_052_486, w_052_487, w_052_489, w_052_491, w_052_493, w_052_495, w_052_498, w_052_502, w_052_506, w_052_509, w_052_515, w_052_516, w_052_517, w_052_519, w_052_521, w_052_524, w_052_529, w_052_530, w_052_533, w_052_534, w_052_535, w_052_536, w_052_541, w_052_542, w_052_543, w_052_546, w_052_547, w_052_551, w_052_553, w_052_556, w_052_557, w_052_572, w_052_579, w_052_580, w_052_581, w_052_582, w_052_583, w_052_585, w_052_587, w_052_589, w_052_590, w_052_592, w_052_593, w_052_594, w_052_595, w_052_596, w_052_599, w_052_600, w_052_601, w_052_602, w_052_604, w_052_605, w_052_606, w_052_609, w_052_610, w_052_614, w_052_619, w_052_621, w_052_623, w_052_626, w_052_627, w_052_628, w_052_629, w_052_631, w_052_632, w_052_633, w_052_634, w_052_637, w_052_639, w_052_641, w_052_643, w_052_647, w_052_649, w_052_652, w_052_653, w_052_662, w_052_664, w_052_665, w_052_666, w_052_668, w_052_670, w_052_671, w_052_674, w_052_675, w_052_680, w_052_687, w_052_688, w_052_690, w_052_691, w_052_692, w_052_694, w_052_695, w_052_696, w_052_697, w_052_699, w_052_701, w_052_702, w_052_704, w_052_707, w_052_708, w_052_710, w_052_713, w_052_715, w_052_716, w_052_719, w_052_720, w_052_721, w_052_722, w_052_725, w_052_726, w_052_727, w_052_731, w_052_732, w_052_736, w_052_737, w_052_738, w_052_739, w_052_742, w_052_743, w_052_747, w_052_749, w_052_753, w_052_754, w_052_755, w_052_760, w_052_766, w_052_767, w_052_771, w_052_773, w_052_774, w_052_776, w_052_779, w_052_780, w_052_782, w_052_783, w_052_786, w_052_787, w_052_789, w_052_795, w_052_801, w_052_802, w_052_805, w_052_806, w_052_809, w_052_811, w_052_812, w_052_813, w_052_815, w_052_820, w_052_822, w_052_825, w_052_827, w_052_828, w_052_832, w_052_833, w_052_836, w_052_839, w_052_841, w_052_842, w_052_844, w_052_846, w_052_848, w_052_850, w_052_853, w_052_854, w_052_859, w_052_860, w_052_862, w_052_870, w_052_872, w_052_875, w_052_876, w_052_877, w_052_881, w_052_883, w_052_886, w_052_888, w_052_890, w_052_891, w_052_892, w_052_894, w_052_895, w_052_898, w_052_900, w_052_906, w_052_909, w_052_911, w_052_912, w_052_914, w_052_917, w_052_919, w_052_921, w_052_923, w_052_924, w_052_925, w_052_926, w_052_927, w_052_928, w_052_929, w_052_930, w_052_933, w_052_935, w_052_939, w_052_942, w_052_944, w_052_947, w_052_949, w_052_952, w_052_957, w_052_963, w_052_964, w_052_965, w_052_968, w_052_974, w_052_977, w_052_978, w_052_988, w_052_989, w_052_993, w_052_994, w_052_995, w_052_996, w_052_998, w_052_1000, w_052_1001, w_052_1002, w_052_1005, w_052_1006, w_052_1008, w_052_1011, w_052_1012, w_052_1013, w_052_1014, w_052_1015, w_052_1017, w_052_1018, w_052_1019, w_052_1020, w_052_1021, w_052_1023, w_052_1024, w_052_1027, w_052_1028, w_052_1029, w_052_1031, w_052_1034, w_052_1035, w_052_1036, w_052_1044, w_052_1048, w_052_1050, w_052_1052, w_052_1054, w_052_1057, w_052_1062, w_052_1064, w_052_1066, w_052_1067, w_052_1068, w_052_1070, w_052_1072, w_052_1073, w_052_1074, w_052_1076, w_052_1082, w_052_1083, w_052_1084, w_052_1085, w_052_1086, w_052_1090, w_052_1091, w_052_1093, w_052_1094, w_052_1095, w_052_1096, w_052_1100, w_052_1101, w_052_1105, w_052_1106, w_052_1108, w_052_1110, w_052_1112, w_052_1116, w_052_1118, w_052_1122, w_052_1123, w_052_1125, w_052_1127, w_052_1131, w_052_1132, w_052_1134, w_052_1135, w_052_1136, w_052_1137, w_052_1139, w_052_1145, w_052_1149, w_052_1150, w_052_1152, w_052_1154, w_052_1156, w_052_1166, w_052_1169, w_052_1171, w_052_1173, w_052_1174, w_052_1178, w_052_1180, w_052_1185, w_052_1186, w_052_1188, w_052_1190, w_052_1194, w_052_1195, w_052_1201, w_052_1207, w_052_1209, w_052_1210, w_052_1211, w_052_1215, w_052_1217, w_052_1220, w_052_1223, w_052_1224, w_052_1228, w_052_1231, w_052_1232, w_052_1234, w_052_1238, w_052_1245, w_052_1247, w_052_1250, w_052_1253, w_052_1254, w_052_1258, w_052_1266, w_052_1269, w_052_1271, w_052_1272, w_052_1274, w_052_1275, w_052_1276, w_052_1277, w_052_1281, w_052_1285, w_052_1287, w_052_1288, w_052_1290, w_052_1292, w_052_1294, w_052_1297, w_052_1298, w_052_1299, w_052_1300, w_052_1302, w_052_1303, w_052_1304, w_052_1305, w_052_1310, w_052_1314, w_052_1317, w_052_1318, w_052_1319, w_052_1320, w_052_1321, w_052_1329, w_052_1330, w_052_1331, w_052_1333, w_052_1339, w_052_1340, w_052_1343, w_052_1344, w_052_1345, w_052_1347, w_052_1349, w_052_1355, w_052_1356, w_052_1358, w_052_1361, w_052_1362, w_052_1363, w_052_1364, w_052_1366, w_052_1368, w_052_1369, w_052_1371, w_052_1373, w_052_1374, w_052_1375, w_052_1376, w_052_1378, w_052_1379, w_052_1380, w_052_1384, w_052_1387, w_052_1389, w_052_1391, w_052_1393, w_052_1396, w_052_1402, w_052_1403, w_052_1404, w_052_1405, w_052_1408, w_052_1410, w_052_1411, w_052_1416, w_052_1418, w_052_1424, w_052_1425, w_052_1426, w_052_1427, w_052_1429, w_052_1430, w_052_1431, w_052_1434, w_052_1436, w_052_1441, w_052_1442, w_052_1443, w_052_1444, w_052_1449, w_052_1459, w_052_1462, w_052_1463, w_052_1464, w_052_1465, w_052_1467, w_052_1469, w_052_1470, w_052_1471, w_052_1473, w_052_1474, w_052_1476, w_052_1477, w_052_1478, w_052_1482, w_052_1483, w_052_1484, w_052_1485, w_052_1486, w_052_1489, w_052_1490, w_052_1494, w_052_1495, w_052_1496, w_052_1499, w_052_1500, w_052_1501, w_052_1503, w_052_1504, w_052_1505, w_052_1506, w_052_1507, w_052_1509, w_052_1510, w_052_1512, w_052_1519, w_052_1525, w_052_1527, w_052_1528, w_052_1529, w_052_1534, w_052_1536, w_052_1542, w_052_1543, w_052_1547, w_052_1548, w_052_1553, w_052_1555, w_052_1559, w_052_1561, w_052_1568, w_052_1572, w_052_1574, w_052_1575, w_052_1577, w_052_1580, w_052_1582, w_052_1583, w_052_1588, w_052_1591, w_052_1597, w_052_1599, w_052_1603, w_052_1605, w_052_1606, w_052_1608, w_052_1612, w_052_1613, w_052_1614, w_052_1615, w_052_1618, w_052_1619, w_052_1620, w_052_1621, w_052_1623, w_052_1624, w_052_1625, w_052_1630, w_052_1631, w_052_1633, w_052_1634, w_052_1637, w_052_1638, w_052_1640, w_052_1641, w_052_1643, w_052_1647, w_052_1648, w_052_1651, w_052_1657, w_052_1658, w_052_1659, w_052_1662, w_052_1668, w_052_1669, w_052_1673, w_052_1676, w_052_1677, w_052_1681, w_052_1683, w_052_1684, w_052_1685, w_052_1686, w_052_1687, w_052_1688, w_052_1689, w_052_1691, w_052_1692, w_052_1694, w_052_1696, w_052_1700, w_052_1701, w_052_1703, w_052_1708, w_052_1709, w_052_1712, w_052_1716, w_052_1718, w_052_1721, w_052_1724, w_052_1725, w_052_1726, w_052_1727, w_052_1728, w_052_1729, w_052_1731, w_052_1735, w_052_1737, w_052_1738, w_052_1739, w_052_1743, w_052_1745, w_052_1753, w_052_1756, w_052_1757, w_052_1759, w_052_1762, w_052_1770, w_052_1772, w_052_1774, w_052_1775, w_052_1778, w_052_1779, w_052_1780, w_052_1781, w_052_1784, w_052_1787, w_052_1790, w_052_1792, w_052_1793, w_052_1795, w_052_1797, w_052_1798, w_052_1801, w_052_1802, w_052_1803, w_052_1804, w_052_1805, w_052_1806, w_052_1807, w_052_1808, w_052_1809, w_052_1810, w_052_1811, w_052_1812, w_052_1816, w_052_1820, w_052_1821, w_052_1822, w_052_1823, w_052_1824, w_052_1825, w_052_1826, w_052_1828, w_052_1829, w_052_1834, w_052_1838, w_052_1840, w_052_1842, w_052_1843, w_052_1846, w_052_1854, w_052_1859, w_052_1861, w_052_1862, w_052_1863, w_052_1865, w_052_1870, w_052_1871, w_052_1872, w_052_1873, w_052_1876, w_052_1878, w_052_1880, w_052_1882, w_052_1883, w_052_1884, w_052_1886, w_052_1888, w_052_1890, w_052_1896, w_052_1898, w_052_1903, w_052_1904, w_052_1907, w_052_1910, w_052_1911, w_052_1913, w_052_1918, w_052_1922, w_052_1924, w_052_1926, w_052_1932, w_052_1934, w_052_1935, w_052_1937, w_052_1939, w_052_1942, w_052_1943, w_052_1944, w_052_1947, w_052_1948, w_052_1951, w_052_1954, w_052_1955, w_052_1956, w_052_1957, w_052_1960, w_052_1962, w_052_1963, w_052_1965, w_052_1967, w_052_1968, w_052_1971, w_052_1972, w_052_1975, w_052_1976, w_052_1978, w_052_1979, w_052_1986, w_052_1995, w_052_1996, w_052_2000, w_052_2009, w_052_2011, w_052_2015, w_052_2022, w_052_2025, w_052_2026, w_052_2028, w_052_2030, w_052_2031, w_052_2033, w_052_2035, w_052_2038, w_052_2041, w_052_2042, w_052_2048, w_052_2049, w_052_2050, w_052_2053, w_052_2055, w_052_2060, w_052_2061, w_052_2062, w_052_2066, w_052_2069, w_052_2075, w_052_2079, w_052_2083, w_052_2084, w_052_2085, w_052_2089, w_052_2090, w_052_2091, w_052_2093, w_052_2094, w_052_2095, w_052_2097, w_052_2099, w_052_2100, w_052_2103, w_052_2104, w_052_2105, w_052_2106, w_052_2108, w_052_2110, w_052_2113, w_052_2116, w_052_2119, w_052_2126, w_052_2127, w_052_2128, w_052_2130, w_052_2133, w_052_2136, w_052_2137, w_052_2138, w_052_2140, w_052_2141, w_052_2142, w_052_2151, w_052_2153, w_052_2157, w_052_2159, w_052_2160, w_052_2161, w_052_2162, w_052_2163, w_052_2165, w_052_2166, w_052_2167, w_052_2172, w_052_2173, w_052_2177, w_052_2188, w_052_2190, w_052_2191, w_052_2192, w_052_2194, w_052_2197, w_052_2200, w_052_2204, w_052_2205, w_052_2206, w_052_2207, w_052_2209, w_052_2213, w_052_2214, w_052_2215, w_052_2216, w_052_2220, w_052_2222, w_052_2224, w_052_2228, w_052_2229, w_052_2233, w_052_2234, w_052_2235, w_052_2239, w_052_2242, w_052_2245, w_052_2248, w_052_2250, w_052_2251, w_052_2252, w_052_2253, w_052_2257, w_052_2263, w_052_2264, w_052_2265, w_052_2267, w_052_2271, w_052_2272, w_052_2273, w_052_2277, w_052_2278, w_052_2281, w_052_2286, w_052_2287, w_052_2289, w_052_2293, w_052_2297, w_052_2303, w_052_2305, w_052_2306, w_052_2309, w_052_2312, w_052_2313, w_052_2317, w_052_2319, w_052_2321, w_052_2324, w_052_2325, w_052_2326, w_052_2327, w_052_2329, w_052_2332, w_052_2338, w_052_2340, w_052_2342, w_052_2343, w_052_2345, w_052_2346, w_052_2347, w_052_2350, w_052_2351, w_052_2353, w_052_2356, w_052_2358, w_052_2361, w_052_2365, w_052_2366, w_052_2368, w_052_2369, w_052_2370, w_052_2374, w_052_2378, w_052_2381, w_052_2382, w_052_2385, w_052_2389, w_052_2391, w_052_2394, w_052_2396, w_052_2397, w_052_2398, w_052_2400, w_052_2401, w_052_2402, w_052_2403, w_052_2405, w_052_2406, w_052_2407, w_052_2408, w_052_2409, w_052_2410, w_052_2412, w_052_2419, w_052_2423, w_052_2425, w_052_2426, w_052_2427, w_052_2430, w_052_2431, w_052_2432, w_052_2433, w_052_2434, w_052_2436, w_052_2437, w_052_2439, w_052_2440, w_052_2441, w_052_2442, w_052_2444, w_052_2447, w_052_2451, w_052_2454, w_052_2459, w_052_2461, w_052_2463, w_052_2466, w_052_2468, w_052_2474, w_052_2478, w_052_2481, w_052_2483, w_052_2484, w_052_2485, w_052_2486, w_052_2490, w_052_2493, w_052_2494, w_052_2496, w_052_2498, w_052_2501, w_052_2502, w_052_2509, w_052_2511, w_052_2512, w_052_2513, w_052_2514, w_052_2516, w_052_2517, w_052_2518, w_052_2519, w_052_2521, w_052_2523, w_052_2529, w_052_2531, w_052_2533, w_052_2535, w_052_2539, w_052_2540, w_052_2541, w_052_2545, w_052_2547, w_052_2549, w_052_2550, w_052_2551, w_052_2552, w_052_2553, w_052_2554, w_052_2555, w_052_2557, w_052_2558, w_052_2561, w_052_2563, w_052_2565, w_052_2569, w_052_2574, w_052_2576, w_052_2578, w_052_2579, w_052_2581, w_052_2586, w_052_2588, w_052_2589, w_052_2595, w_052_2597, w_052_2598, w_052_2613, w_052_2614, w_052_2618, w_052_2623, w_052_2626, w_052_2627, w_052_2628, w_052_2629, w_052_2630, w_052_2632, w_052_2633, w_052_2635, w_052_2636, w_052_2638, w_052_2641, w_052_2644, w_052_2645, w_052_2648, w_052_2649, w_052_2650, w_052_2651, w_052_2652, w_052_2654, w_052_2656, w_052_2662, w_052_2664, w_052_2667, w_052_2668, w_052_2669, w_052_2670, w_052_2671, w_052_2672, w_052_2674, w_052_2675, w_052_2677, w_052_2678, w_052_2679, w_052_2680, w_052_2681, w_052_2683, w_052_2687, w_052_2688, w_052_2689, w_052_2691, w_052_2692, w_052_2695, w_052_2698, w_052_2700, w_052_2702, w_052_2705, w_052_2708, w_052_2712, w_052_2714, w_052_2720, w_052_2723, w_052_2727, w_052_2729, w_052_2732, w_052_2733, w_052_2734, w_052_2738, w_052_2741, w_052_2745, w_052_2747, w_052_2749, w_052_2750, w_052_2754, w_052_2755, w_052_2757, w_052_2758, w_052_2761, w_052_2762, w_052_2764, w_052_2765, w_052_2769, w_052_2770, w_052_2775, w_052_2776, w_052_2777, w_052_2779, w_052_2780, w_052_2781, w_052_2785, w_052_2788, w_052_2789, w_052_2790, w_052_2792, w_052_2793, w_052_2796, w_052_2797, w_052_2799, w_052_2800, w_052_2806, w_052_2808, w_052_2810, w_052_2812, w_052_2814, w_052_2816, w_052_2819, w_052_2820, w_052_2821, w_052_2826, w_052_2827, w_052_2831, w_052_2833, w_052_2836, w_052_2840, w_052_2842, w_052_2848, w_052_2849, w_052_2850, w_052_2853, w_052_2858, w_052_2859, w_052_2860, w_052_2863, w_052_2865, w_052_2866, w_052_2867, w_052_2868, w_052_2869, w_052_2870, w_052_2871, w_052_2872, w_052_2874, w_052_2878, w_052_2880, w_052_2881, w_052_2882, w_052_2883, w_052_2885, w_052_2886, w_052_2887, w_052_2888, w_052_2889, w_052_2890, w_052_2891, w_052_2892, w_052_2893, w_052_2894, w_052_2895, w_052_2898, w_052_2900, w_052_2901, w_052_2902, w_052_2903, w_052_2904, w_052_2905, w_052_2908, w_052_2912, w_052_2913, w_052_2914, w_052_2915, w_052_2916, w_052_2918, w_052_2919, w_052_2920, w_052_2922, w_052_2923, w_052_2924, w_052_2925, w_052_2927, w_052_2930, w_052_2933, w_052_2934, w_052_2935, w_052_2936, w_052_2937, w_052_2939, w_052_2940, w_052_2942, w_052_2943, w_052_2945, w_052_2946, w_052_2947, w_052_2948, w_052_2949, w_052_2953, w_052_2955, w_052_2957, w_052_2958, w_052_2959, w_052_2960, w_052_2961, w_052_2962, w_052_2963, w_052_2965, w_052_2968, w_052_2969, w_052_2971, w_052_2972, w_052_2976, w_052_2979, w_052_2980, w_052_2983, w_052_2985, w_052_2987, w_052_2988, w_052_2993, w_052_2994, w_052_2998, w_052_3002, w_052_3003, w_052_3005, w_052_3006, w_052_3008, w_052_3009, w_052_3010, w_052_3011, w_052_3016, w_052_3019, w_052_3021, w_052_3022, w_052_3023, w_052_3025, w_052_3026, w_052_3027, w_052_3028, w_052_3029, w_052_3031, w_052_3032, w_052_3033, w_052_3036, w_052_3037, w_052_3038, w_052_3039, w_052_3043, w_052_3045, w_052_3048, w_052_3049, w_052_3052, w_052_3053, w_052_3056, w_052_3057, w_052_3059, w_052_3060, w_052_3063, w_052_3064, w_052_3067, w_052_3068, w_052_3069, w_052_3070, w_052_3072, w_052_3073, w_052_3074, w_052_3077, w_052_3079, w_052_3080, w_052_3081, w_052_3082, w_052_3083, w_052_3084, w_052_3085, w_052_3086, w_052_3089, w_052_3090, w_052_3091, w_052_3095, w_052_3099, w_052_3100, w_052_3102, w_052_3104, w_052_3106, w_052_3107, w_052_3108, w_052_3112, w_052_3115, w_052_3116, w_052_3117, w_052_3121, w_052_3122, w_052_3124, w_052_3125, w_052_3128, w_052_3129, w_052_3132, w_052_3134, w_052_3135, w_052_3136, w_052_3137, w_052_3140, w_052_3142, w_052_3145, w_052_3146, w_052_3147, w_052_3149, w_052_3150, w_052_3154, w_052_3157, w_052_3158, w_052_3160, w_052_3161, w_052_3162, w_052_3164, w_052_3165, w_052_3166, w_052_3169, w_052_3174, w_052_3180, w_052_3185, w_052_3186, w_052_3187, w_052_3189, w_052_3190, w_052_3191, w_052_3193, w_052_3194, w_052_3195, w_052_3197, w_052_3206, w_052_3209, w_052_3210, w_052_3211, w_052_3213, w_052_3214, w_052_3215, w_052_3216, w_052_3221, w_052_3224, w_052_3225, w_052_3228, w_052_3229, w_052_3230, w_052_3232, w_052_3234, w_052_3236, w_052_3237, w_052_3238, w_052_3242, w_052_3243, w_052_3245, w_052_3247, w_052_3248, w_052_3250, w_052_3258, w_052_3262, w_052_3264, w_052_3266, w_052_3268, w_052_3269, w_052_3270, w_052_3273, w_052_3275, w_052_3281, w_052_3283, w_052_3287, w_052_3291, w_052_3292, w_052_3297, w_052_3298, w_052_3299, w_052_3300, w_052_3301, w_052_3302, w_052_3304, w_052_3308, w_052_3309, w_052_3310, w_052_3311, w_052_3314, w_052_3315, w_052_3316, w_052_3318, w_052_3320, w_052_3329, w_052_3330, w_052_3331, w_052_3332, w_052_3333, w_052_3335, w_052_3336, w_052_3337, w_052_3339, w_052_3340, w_052_3342, w_052_3344, w_052_3348, w_052_3352, w_052_3355, w_052_3356, w_052_3357, w_052_3358, w_052_3359, w_052_3360, w_052_3363, w_052_3364, w_052_3368, w_052_3369, w_052_3372, w_052_3376, w_052_3377, w_052_3381, w_052_3383, w_052_3389, w_052_3390, w_052_3391, w_052_3394, w_052_3395, w_052_3396, w_052_3401, w_052_3403, w_052_3411, w_052_3414, w_052_3415, w_052_3416, w_052_3418, w_052_3419, w_052_3420, w_052_3421, w_052_3425, w_052_3427, w_052_3429, w_052_3430, w_052_3431, w_052_3433, w_052_3435, w_052_3436, w_052_3437, w_052_3438, w_052_3441, w_052_3446, w_052_3449, w_052_3451, w_052_3455, w_052_3456, w_052_3457, w_052_3458, w_052_3460, w_052_3461, w_052_3463, w_052_3464, w_052_3469, w_052_3470, w_052_3473, w_052_3474, w_052_3477, w_052_3479, w_052_3485, w_052_3486, w_052_3487, w_052_3489, w_052_3490, w_052_3494, w_052_3495, w_052_3499, w_052_3500, w_052_3501, w_052_3505, w_052_3509, w_052_3517, w_052_3518, w_052_3520, w_052_3522, w_052_3524, w_052_3526, w_052_3529, w_052_3533, w_052_3534, w_052_3536, w_052_3537, w_052_3538, w_052_3541, w_052_3551, w_052_3552, w_052_3558, w_052_3559, w_052_3560, w_052_3561, w_052_3562, w_052_3567, w_052_3570, w_052_3571, w_052_3572, w_052_3573, w_052_3577, w_052_3580, w_052_3581, w_052_3582, w_052_3583, w_052_3589, w_052_3590, w_052_3591, w_052_3596, w_052_3597, w_052_3598, w_052_3602, w_052_3603, w_052_3609, w_052_3611, w_052_3618, w_052_3620, w_052_3622, w_052_3624, w_052_3626, w_052_3627, w_052_3628, w_052_3633, w_052_3634, w_052_3636, w_052_3638, w_052_3639, w_052_3642, w_052_3643, w_052_3647, w_052_3650, w_052_3652, w_052_3653, w_052_3655, w_052_3656, w_052_3658, w_052_3660, w_052_3662, w_052_3663, w_052_3668, w_052_3672, w_052_3673, w_052_3675, w_052_3677, w_052_3683, w_052_3684, w_052_3685, w_052_3686, w_052_3688, w_052_3689, w_052_3692, w_052_3693, w_052_3694, w_052_3696, w_052_3700, w_052_3701, w_052_3702, w_052_3704, w_052_3705, w_052_3708, w_052_3710, w_052_3711, w_052_3713, w_052_3715, w_052_3717, w_052_3720, w_052_3722, w_052_3724, w_052_3726, w_052_3729, w_052_3734, w_052_3735, w_052_3736, w_052_3738, w_052_3739, w_052_3747, w_052_3748, w_052_3749, w_052_3750, w_052_3758, w_052_3759, w_052_3760, w_052_3761, w_052_3762, w_052_3763, w_052_3764, w_052_3765, w_052_3767, w_052_3771, w_052_3772, w_052_3775, w_052_3776, w_052_3777, w_052_3783, w_052_3785, w_052_3786, w_052_3788, w_052_3790, w_052_3791, w_052_3792, w_052_3794, w_052_3795, w_052_3796, w_052_3797, w_052_3803, w_052_3804, w_052_3805, w_052_3811, w_052_3819, w_052_3820, w_052_3821, w_052_3822, w_052_3826, w_052_3827, w_052_3828, w_052_3829, w_052_3831, w_052_3833, w_052_3834, w_052_3836, w_052_3837, w_052_3838, w_052_3840, w_052_3842, w_052_3844, w_052_3849, w_052_3850, w_052_3851, w_052_3852, w_052_3855, w_052_3857, w_052_3862, w_052_3863, w_052_3864, w_052_3866, w_052_3868, w_052_3872, w_052_3873, w_052_3878, w_052_3882, w_052_3883, w_052_3884, w_052_3886, w_052_3887, w_052_3888, w_052_3891, w_052_3892, w_052_3896, w_052_3898, w_052_3899, w_052_3900, w_052_3903, w_052_3904, w_052_3907, w_052_3912, w_052_3914, w_052_3915, w_052_3917, w_052_3918, w_052_3922, w_052_3923, w_052_3924, w_052_3925, w_052_3926, w_052_3928, w_052_3934, w_052_3935, w_052_3938, w_052_3941, w_052_3943, w_052_3945, w_052_3946, w_052_3950, w_052_3953, w_052_3956, w_052_3958, w_052_3960, w_052_3964, w_052_3965, w_052_3969, w_052_3970, w_052_3972, w_052_3974, w_052_3976, w_052_3977, w_052_3978, w_052_3980, w_052_3982, w_052_3985, w_052_3987, w_052_3988, w_052_3990, w_052_3992, w_052_3993, w_052_3997, w_052_3998, w_052_3999, w_052_4000, w_052_4005, w_052_4008, w_052_4010, w_052_4012, w_052_4014, w_052_4016, w_052_4017, w_052_4018, w_052_4021, w_052_4022, w_052_4023, w_052_4024, w_052_4025, w_052_4026, w_052_4029, w_052_4031, w_052_4033, w_052_4035, w_052_4036, w_052_4038, w_052_4039, w_052_4042, w_052_4043, w_052_4044, w_052_4045, w_052_4046, w_052_4051, w_052_4054, w_052_4055, w_052_4058, w_052_4065, w_052_4067, w_052_4069, w_052_4070, w_052_4071, w_052_4073, w_052_4077, w_052_4078, w_052_4080, w_052_4082, w_052_4083, w_052_4084, w_052_4086, w_052_4088, w_052_4091, w_052_4092, w_052_4095, w_052_4102, w_052_4103, w_052_4107, w_052_4108, w_052_4114, w_052_4116, w_052_4119, w_052_4120, w_052_4124, w_052_4128, w_052_4130, w_052_4132, w_052_4134, w_052_4136, w_052_4138, w_052_4140, w_052_4142, w_052_4144, w_052_4147, w_052_4148, w_052_4149, w_052_4150, w_052_4152, w_052_4153, w_052_4156, w_052_4159, w_052_4163, w_052_4164, w_052_4165, w_052_4167, w_052_4175, w_052_4182, w_052_4183, w_052_4184, w_052_4186, w_052_4187, w_052_4188, w_052_4189, w_052_4190, w_052_4191, w_052_4192, w_052_4193, w_052_4194, w_052_4197, w_052_4198, w_052_4199, w_052_4202, w_052_4204, w_052_4206, w_052_4208, w_052_4211, w_052_4212, w_052_4215, w_052_4216, w_052_4218, w_052_4221, w_052_4223, w_052_4225, w_052_4229, w_052_4232, w_052_4234, w_052_4235, w_052_4236, w_052_4243, w_052_4246, w_052_4248, w_052_4249, w_052_4254, w_052_4257, w_052_4260, w_052_4261, w_052_4262, w_052_4268, w_052_4270, w_052_4271, w_052_4273, w_052_4274, w_052_4278, w_052_4279, w_052_4280, w_052_4281, w_052_4282, w_052_4284, w_052_4288, w_052_4290, w_052_4291, w_052_4292, w_052_4293, w_052_4296, w_052_4297, w_052_4298, w_052_4302, w_052_4303, w_052_4305, w_052_4306, w_052_4309, w_052_4310, w_052_4311, w_052_4312, w_052_4314, w_052_4318, w_052_4319, w_052_4320, w_052_4321, w_052_4326, w_052_4328, w_052_4329, w_052_4330, w_052_4334, w_052_4335, w_052_4336, w_052_4337, w_052_4338, w_052_4339, w_052_4342, w_052_4343, w_052_4344, w_052_4346, w_052_4347, w_052_4352, w_052_4354, w_052_4357, w_052_4360, w_052_4361, w_052_4364, w_052_4365, w_052_4366, w_052_4368, w_052_4369, w_052_4370, w_052_4372, w_052_4382, w_052_4386, w_052_4392, w_052_4393, w_052_4397, w_052_4398, w_052_4399, w_052_4400, w_052_4405, w_052_4406, w_052_4407, w_052_4408, w_052_4409, w_052_4412, w_052_4414, w_052_4415, w_052_4417, w_052_4418, w_052_4420, w_052_4421, w_052_4422, w_052_4425, w_052_4428, w_052_4430, w_052_4431, w_052_4432, w_052_4433, w_052_4434, w_052_4438, w_052_4441, w_052_4443, w_052_4445, w_052_4447, w_052_4452, w_052_4458, w_052_4464, w_052_4465, w_052_4468, w_052_4469, w_052_4471, w_052_4472, w_052_4473, w_052_4474, w_052_4477, w_052_4478, w_052_4479, w_052_4480, w_052_4481, w_052_4483, w_052_4484, w_052_4485, w_052_4487, w_052_4489, w_052_4490, w_052_4492, w_052_4494, w_052_4495, w_052_4498, w_052_4499, w_052_4500, w_052_4501, w_052_4506, w_052_4510, w_052_4512, w_052_4514, w_052_4515, w_052_4520, w_052_4522, w_052_4524, w_052_4525, w_052_4530, w_052_4531, w_052_4532, w_052_4535, w_052_4540, w_052_4542, w_052_4543, w_052_4545, w_052_4546, w_052_4548, w_052_4556, w_052_4560, w_052_4561, w_052_4562, w_052_4566, w_052_4569, w_052_4570, w_052_4571, w_052_4574, w_052_4576, w_052_4578, w_052_4579, w_052_4582, w_052_4583, w_052_4585, w_052_4586, w_052_4587, w_052_4590, w_052_4591, w_052_4598, w_052_4600, w_052_4603, w_052_4604, w_052_4608, w_052_4612, w_052_4613, w_052_4614, w_052_4615, w_052_4618, w_052_4621, w_052_4623, w_052_4624, w_052_4625, w_052_4630, w_052_4632, w_052_4637, w_052_4639, w_052_4640, w_052_4641, w_052_4642, w_052_4643, w_052_4644, w_052_4645, w_052_4646, w_052_4647, w_052_4650, w_052_4651, w_052_4654, w_052_4655, w_052_4656, w_052_4657, w_052_4658, w_052_4659, w_052_4660, w_052_4661, w_052_4662, w_052_4663, w_052_4664, w_052_4666, w_052_4669, w_052_4671, w_052_4677, w_052_4678, w_052_4679, w_052_4688, w_052_4690, w_052_4691, w_052_4692, w_052_4695, w_052_4696, w_052_4701, w_052_4702, w_052_4703, w_052_4707, w_052_4709, w_052_4710, w_052_4712, w_052_4713, w_052_4715, w_052_4717, w_052_4720, w_052_4723, w_052_4724, w_052_4726, w_052_4727, w_052_4729, w_052_4734, w_052_4736, w_052_4737, w_052_4739, w_052_4743, w_052_4744, w_052_4746, w_052_4747, w_052_4748, w_052_4749, w_052_4751, w_052_4753, w_052_4754, w_052_4755, w_052_4758, w_052_4759, w_052_4763, w_052_4765, w_052_4766, w_052_4768, w_052_4769, w_052_4770, w_052_4774, w_052_4779, w_052_4782, w_052_4783, w_052_4784, w_052_4787, w_052_4788, w_052_4789, w_052_4793, w_052_4798, w_052_4801, w_052_4802, w_052_4805, w_052_4810, w_052_4816, w_052_4817, w_052_4821, w_052_4822, w_052_4825, w_052_4826, w_052_4827, w_052_4828, w_052_4837, w_052_4839, w_052_4841, w_052_4843, w_052_4846, w_052_4848, w_052_4849, w_052_4851, w_052_4854, w_052_4855, w_052_4856, w_052_4857, w_052_4859, w_052_4863, w_052_4864, w_052_4866, w_052_4867, w_052_4868, w_052_4869, w_052_4872, w_052_4877, w_052_4880, w_052_4882, w_052_4884, w_052_4885, w_052_4887, w_052_4888, w_052_4890, w_052_4891, w_052_4892, w_052_4895, w_052_4900, w_052_4903, w_052_4904, w_052_4906, w_052_4907, w_052_4909, w_052_4910, w_052_4911, w_052_4912, w_052_4913, w_052_4919, w_052_4920, w_052_4922, w_052_4923, w_052_4924, w_052_4925, w_052_4926, w_052_4927, w_052_4928, w_052_4930, w_052_4932, w_052_4933, w_052_4934, w_052_4935, w_052_4936, w_052_4937, w_052_4938, w_052_4939, w_052_4940, w_052_4942;
  wire w_053_000, w_053_001, w_053_002, w_053_003, w_053_004, w_053_005, w_053_006, w_053_007, w_053_008, w_053_009, w_053_011, w_053_012, w_053_013, w_053_014, w_053_017, w_053_018, w_053_019, w_053_020, w_053_021, w_053_022, w_053_023, w_053_024, w_053_025, w_053_026, w_053_027, w_053_028, w_053_029, w_053_031, w_053_032, w_053_033, w_053_035, w_053_036, w_053_037, w_053_038, w_053_039, w_053_041, w_053_042, w_053_043, w_053_044, w_053_045, w_053_046, w_053_047, w_053_049, w_053_050, w_053_051, w_053_053, w_053_054, w_053_055, w_053_056, w_053_057, w_053_059, w_053_060, w_053_061, w_053_062, w_053_063, w_053_064, w_053_065, w_053_066, w_053_068, w_053_069, w_053_070, w_053_071, w_053_072, w_053_073, w_053_074, w_053_075, w_053_076, w_053_077, w_053_078, w_053_079, w_053_080, w_053_081, w_053_082, w_053_083, w_053_084, w_053_085, w_053_086, w_053_087, w_053_088, w_053_089, w_053_090, w_053_091, w_053_092, w_053_093, w_053_094, w_053_095, w_053_096, w_053_097, w_053_098, w_053_099, w_053_102, w_053_103, w_053_104, w_053_105, w_053_106, w_053_107, w_053_108, w_053_109, w_053_110, w_053_111, w_053_113, w_053_114, w_053_115, w_053_117, w_053_119, w_053_120, w_053_121, w_053_122, w_053_123, w_053_124, w_053_125, w_053_126, w_053_127, w_053_128, w_053_130, w_053_131, w_053_132, w_053_133, w_053_134, w_053_135, w_053_136, w_053_138, w_053_139, w_053_140, w_053_141, w_053_142, w_053_143, w_053_144, w_053_145, w_053_146, w_053_148, w_053_149, w_053_151, w_053_152, w_053_154, w_053_155, w_053_156, w_053_158, w_053_159, w_053_160, w_053_161, w_053_162, w_053_163, w_053_164, w_053_165, w_053_167, w_053_169, w_053_170, w_053_172, w_053_173, w_053_174, w_053_175, w_053_176, w_053_177, w_053_179, w_053_180, w_053_181, w_053_182, w_053_183, w_053_184, w_053_185, w_053_186, w_053_187, w_053_188, w_053_189, w_053_190, w_053_191, w_053_192, w_053_193, w_053_194, w_053_195, w_053_196, w_053_197, w_053_198, w_053_199, w_053_200, w_053_201, w_053_202, w_053_203, w_053_204, w_053_207, w_053_208, w_053_210, w_053_211, w_053_212, w_053_213, w_053_214, w_053_215, w_053_216, w_053_217, w_053_218, w_053_219, w_053_220, w_053_222, w_053_223, w_053_224, w_053_225, w_053_226, w_053_227, w_053_228, w_053_229, w_053_231, w_053_232, w_053_233, w_053_234, w_053_235, w_053_236, w_053_237, w_053_238, w_053_239, w_053_240, w_053_241, w_053_242, w_053_243, w_053_245, w_053_247, w_053_248, w_053_249, w_053_250, w_053_251, w_053_252, w_053_253, w_053_254, w_053_256, w_053_257, w_053_258, w_053_259, w_053_260, w_053_261, w_053_262, w_053_263, w_053_264, w_053_265, w_053_266, w_053_267, w_053_269, w_053_271, w_053_272, w_053_274, w_053_276, w_053_277, w_053_278, w_053_279, w_053_280, w_053_281, w_053_282, w_053_283, w_053_284, w_053_286, w_053_288, w_053_289, w_053_290, w_053_291, w_053_292, w_053_293, w_053_295, w_053_296, w_053_297, w_053_298, w_053_299, w_053_300, w_053_301, w_053_302, w_053_304, w_053_305, w_053_308, w_053_309, w_053_310, w_053_311, w_053_312, w_053_313, w_053_314, w_053_315, w_053_316, w_053_317, w_053_318, w_053_320, w_053_321, w_053_322, w_053_326, w_053_327, w_053_328, w_053_331, w_053_332, w_053_333, w_053_334, w_053_335, w_053_336, w_053_337, w_053_338, w_053_339, w_053_340, w_053_341, w_053_342, w_053_344, w_053_345, w_053_346, w_053_347, w_053_349, w_053_350, w_053_351, w_053_352, w_053_353, w_053_354, w_053_355, w_053_356, w_053_357, w_053_359, w_053_361, w_053_362, w_053_363, w_053_364, w_053_366, w_053_367, w_053_368, w_053_369, w_053_370, w_053_371, w_053_372, w_053_373, w_053_375, w_053_376, w_053_377, w_053_378, w_053_379, w_053_380, w_053_381, w_053_382, w_053_383, w_053_384, w_053_385, w_053_386, w_053_387, w_053_388, w_053_389, w_053_390, w_053_391, w_053_392, w_053_393, w_053_394, w_053_395, w_053_396, w_053_397, w_053_399, w_053_400, w_053_401, w_053_402, w_053_403, w_053_404, w_053_405, w_053_406, w_053_408, w_053_409, w_053_410, w_053_411, w_053_412, w_053_413, w_053_414, w_053_415, w_053_416, w_053_417, w_053_418, w_053_419, w_053_422, w_053_423, w_053_426, w_053_427, w_053_429, w_053_430, w_053_431, w_053_432, w_053_433, w_053_434, w_053_435, w_053_436, w_053_437, w_053_438, w_053_439, w_053_440, w_053_441, w_053_442, w_053_443, w_053_444, w_053_445, w_053_446, w_053_447, w_053_449, w_053_450, w_053_451, w_053_452, w_053_453, w_053_454, w_053_455, w_053_456, w_053_457, w_053_458, w_053_460, w_053_461, w_053_462, w_053_463, w_053_464, w_053_465, w_053_466, w_053_467, w_053_468, w_053_469, w_053_470, w_053_471, w_053_472, w_053_473, w_053_474, w_053_475, w_053_476, w_053_477, w_053_478, w_053_479, w_053_480, w_053_481, w_053_482, w_053_483, w_053_484, w_053_485, w_053_486, w_053_487, w_053_488, w_053_489, w_053_490, w_053_491, w_053_492, w_053_493, w_053_494, w_053_495, w_053_496, w_053_497, w_053_498, w_053_500, w_053_501, w_053_502, w_053_503, w_053_504, w_053_505, w_053_506, w_053_507, w_053_508, w_053_509, w_053_510, w_053_512, w_053_513, w_053_514, w_053_515, w_053_516, w_053_517, w_053_518, w_053_519, w_053_524, w_053_526, w_053_527, w_053_528, w_053_529, w_053_531, w_053_532, w_053_533, w_053_534, w_053_535, w_053_536, w_053_537, w_053_538, w_053_539, w_053_541, w_053_543, w_053_544, w_053_545, w_053_546, w_053_547, w_053_549, w_053_551, w_053_552, w_053_553, w_053_554, w_053_555, w_053_556, w_053_557, w_053_558, w_053_560, w_053_561, w_053_562, w_053_564, w_053_565, w_053_566, w_053_567, w_053_568, w_053_569, w_053_570, w_053_571, w_053_572, w_053_573, w_053_574, w_053_575, w_053_576, w_053_577, w_053_578, w_053_579, w_053_580, w_053_581, w_053_582, w_053_583, w_053_584, w_053_585, w_053_586, w_053_588, w_053_589, w_053_590, w_053_591, w_053_592, w_053_593, w_053_594, w_053_595, w_053_596, w_053_597, w_053_598, w_053_599, w_053_600, w_053_601, w_053_602, w_053_603, w_053_604, w_053_605, w_053_606, w_053_607, w_053_608, w_053_609, w_053_610, w_053_611, w_053_613, w_053_614, w_053_615, w_053_616, w_053_617, w_053_619, w_053_620, w_053_621, w_053_623, w_053_624, w_053_625, w_053_626, w_053_627, w_053_628, w_053_629, w_053_631, w_053_632, w_053_633, w_053_634, w_053_635, w_053_636, w_053_638, w_053_640, w_053_641, w_053_643, w_053_644, w_053_645, w_053_646, w_053_650, w_053_653, w_053_654, w_053_655, w_053_656, w_053_657, w_053_658, w_053_659, w_053_660, w_053_661, w_053_662, w_053_663, w_053_664, w_053_665, w_053_667, w_053_668, w_053_669, w_053_670, w_053_671, w_053_672, w_053_673, w_053_676, w_053_678, w_053_680, w_053_681, w_053_683, w_053_684, w_053_685, w_053_686, w_053_687, w_053_688, w_053_689, w_053_691, w_053_692, w_053_693, w_053_694, w_053_695, w_053_696, w_053_697, w_053_698, w_053_699, w_053_700, w_053_701, w_053_702, w_053_703, w_053_704, w_053_705, w_053_708, w_053_709, w_053_710, w_053_713, w_053_714, w_053_715, w_053_716, w_053_717, w_053_718, w_053_719, w_053_720, w_053_721, w_053_722, w_053_723, w_053_724, w_053_726, w_053_727, w_053_729, w_053_730, w_053_731, w_053_732, w_053_733, w_053_735, w_053_736, w_053_737, w_053_739, w_053_740, w_053_741, w_053_742, w_053_743, w_053_744, w_053_745, w_053_746, w_053_747, w_053_750, w_053_751, w_053_752, w_053_753, w_053_754, w_053_756, w_053_757, w_053_758, w_053_759, w_053_760, w_053_762, w_053_763, w_053_764, w_053_765, w_053_766, w_053_767, w_053_769, w_053_770, w_053_772, w_053_773, w_053_774, w_053_775, w_053_776, w_053_777, w_053_778, w_053_779, w_053_780, w_053_782, w_053_783, w_053_784, w_053_785, w_053_786, w_053_787, w_053_788, w_053_789, w_053_790, w_053_791, w_053_792, w_053_793, w_053_795, w_053_796, w_053_798, w_053_799, w_053_800, w_053_801, w_053_802, w_053_803, w_053_805, w_053_806, w_053_807, w_053_808, w_053_809, w_053_810, w_053_812, w_053_813, w_053_816, w_053_819, w_053_820, w_053_821, w_053_822, w_053_823, w_053_824, w_053_825, w_053_826, w_053_827, w_053_830, w_053_832, w_053_833, w_053_834, w_053_835, w_053_836, w_053_837, w_053_838, w_053_840, w_053_841, w_053_842, w_053_843, w_053_844, w_053_845, w_053_848, w_053_849, w_053_850, w_053_851, w_053_852, w_053_853, w_053_854, w_053_855, w_053_856, w_053_857, w_053_858, w_053_859, w_053_861, w_053_862, w_053_863, w_053_864, w_053_865, w_053_866, w_053_867, w_053_868, w_053_871, w_053_872, w_053_873, w_053_874, w_053_875, w_053_876, w_053_877, w_053_878, w_053_879, w_053_880, w_053_881, w_053_882, w_053_883, w_053_884, w_053_885, w_053_886, w_053_888, w_053_889, w_053_891, w_053_892, w_053_893, w_053_895, w_053_896, w_053_897, w_053_898, w_053_901, w_053_902, w_053_903, w_053_904, w_053_905, w_053_906, w_053_907, w_053_908, w_053_909, w_053_910, w_053_911, w_053_912, w_053_913, w_053_914, w_053_915, w_053_916, w_053_918, w_053_919, w_053_920, w_053_921, w_053_922, w_053_923, w_053_924, w_053_925, w_053_928, w_053_930, w_053_931, w_053_932, w_053_933, w_053_934, w_053_935, w_053_938, w_053_940, w_053_941, w_053_943, w_053_944, w_053_945, w_053_946, w_053_947, w_053_948, w_053_950, w_053_951, w_053_952, w_053_953, w_053_954, w_053_955, w_053_957, w_053_958, w_053_960, w_053_961, w_053_962, w_053_963, w_053_964, w_053_966, w_053_967, w_053_968, w_053_969, w_053_970, w_053_971, w_053_972, w_053_973, w_053_975, w_053_976, w_053_977, w_053_978, w_053_979, w_053_982, w_053_983, w_053_984, w_053_985, w_053_987, w_053_988, w_053_989, w_053_990, w_053_991, w_053_992, w_053_993, w_053_994, w_053_995, w_053_996, w_053_1000, w_053_1001, w_053_1002, w_053_1003, w_053_1005, w_053_1007, w_053_1008, w_053_1009, w_053_1010, w_053_1011, w_053_1012, w_053_1013, w_053_1014, w_053_1015, w_053_1016, w_053_1017, w_053_1018, w_053_1019, w_053_1020, w_053_1022, w_053_1023, w_053_1024, w_053_1026, w_053_1028, w_053_1029, w_053_1031, w_053_1032, w_053_1033, w_053_1034, w_053_1036, w_053_1037, w_053_1039, w_053_1040, w_053_1041, w_053_1042, w_053_1043, w_053_1044, w_053_1045, w_053_1046, w_053_1047, w_053_1048, w_053_1049, w_053_1050, w_053_1051, w_053_1052, w_053_1053, w_053_1054, w_053_1055, w_053_1056, w_053_1057, w_053_1058, w_053_1059, w_053_1062, w_053_1063, w_053_1065, w_053_1067, w_053_1069, w_053_1070, w_053_1071, w_053_1072, w_053_1073, w_053_1079, w_053_1080, w_053_1082, w_053_1083, w_053_1084, w_053_1085, w_053_1086, w_053_1087, w_053_1089, w_053_1090, w_053_1091, w_053_1092, w_053_1094, w_053_1095, w_053_1096, w_053_1098, w_053_1099, w_053_1101, w_053_1102, w_053_1103, w_053_1104, w_053_1105, w_053_1106, w_053_1107, w_053_1113, w_053_1115, w_053_1117, w_053_1118, w_053_1120, w_053_1122, w_053_1125, w_053_1126, w_053_1127, w_053_1128, w_053_1129, w_053_1131, w_053_1132, w_053_1133, w_053_1134, w_053_1135, w_053_1136, w_053_1137, w_053_1139, w_053_1140, w_053_1141, w_053_1143, w_053_1145, w_053_1149, w_053_1150, w_053_1151, w_053_1155, w_053_1156, w_053_1157, w_053_1158, w_053_1161, w_053_1162, w_053_1163, w_053_1164, w_053_1165, w_053_1168, w_053_1171, w_053_1176, w_053_1177, w_053_1178, w_053_1179, w_053_1180, w_053_1181, w_053_1183, w_053_1184, w_053_1185, w_053_1187, w_053_1188, w_053_1190, w_053_1191, w_053_1193, w_053_1194, w_053_1195, w_053_1196, w_053_1197, w_053_1198, w_053_1199, w_053_1200, w_053_1202, w_053_1203, w_053_1204, w_053_1205, w_053_1207, w_053_1213, w_053_1215, w_053_1216, w_053_1217, w_053_1218, w_053_1220, w_053_1221, w_053_1222, w_053_1223, w_053_1224, w_053_1225, w_053_1227, w_053_1228, w_053_1229, w_053_1231, w_053_1232, w_053_1233, w_053_1234, w_053_1235, w_053_1236, w_053_1238, w_053_1240, w_053_1241, w_053_1242, w_053_1243, w_053_1244, w_053_1245, w_053_1246, w_053_1248, w_053_1251, w_053_1252, w_053_1253, w_053_1254, w_053_1255, w_053_1257, w_053_1258, w_053_1259, w_053_1260, w_053_1261, w_053_1264, w_053_1266, w_053_1267, w_053_1270, w_053_1271, w_053_1273, w_053_1274, w_053_1275, w_053_1277, w_053_1278, w_053_1280, w_053_1282, w_053_1283, w_053_1284, w_053_1286, w_053_1287, w_053_1288, w_053_1289, w_053_1291, w_053_1292, w_053_1294, w_053_1295, w_053_1296, w_053_1297, w_053_1298, w_053_1299, w_053_1301, w_053_1302, w_053_1304, w_053_1306, w_053_1307, w_053_1309, w_053_1310, w_053_1311, w_053_1313, w_053_1314, w_053_1315, w_053_1317, w_053_1320, w_053_1321, w_053_1322, w_053_1323, w_053_1324, w_053_1325, w_053_1326, w_053_1328, w_053_1330, w_053_1332, w_053_1333, w_053_1334, w_053_1335, w_053_1337, w_053_1340, w_053_1341, w_053_1342, w_053_1343, w_053_1344, w_053_1346, w_053_1347, w_053_1348, w_053_1350, w_053_1351, w_053_1352, w_053_1353, w_053_1354, w_053_1356, w_053_1360, w_053_1362, w_053_1364, w_053_1366, w_053_1368, w_053_1369, w_053_1370, w_053_1371, w_053_1372, w_053_1373, w_053_1374, w_053_1378, w_053_1379, w_053_1383, w_053_1384, w_053_1385, w_053_1386, w_053_1391, w_053_1392, w_053_1394, w_053_1395, w_053_1398, w_053_1401, w_053_1402, w_053_1403, w_053_1404, w_053_1405, w_053_1406, w_053_1407, w_053_1410, w_053_1411, w_053_1412, w_053_1413, w_053_1414, w_053_1415, w_053_1416, w_053_1418, w_053_1419, w_053_1420, w_053_1421, w_053_1423, w_053_1426, w_053_1427, w_053_1428, w_053_1429, w_053_1431, w_053_1432, w_053_1433, w_053_1436, w_053_1438, w_053_1439, w_053_1440, w_053_1441, w_053_1442, w_053_1443, w_053_1444, w_053_1446, w_053_1447, w_053_1448, w_053_1449, w_053_1451, w_053_1452, w_053_1453, w_053_1455, w_053_1459, w_053_1460, w_053_1464, w_053_1465, w_053_1467, w_053_1468, w_053_1470, w_053_1471, w_053_1472, w_053_1473, w_053_1474, w_053_1475, w_053_1476, w_053_1483, w_053_1485, w_053_1486, w_053_1488, w_053_1489, w_053_1490, w_053_1491, w_053_1493, w_053_1494, w_053_1495, w_053_1496, w_053_1497, w_053_1499, w_053_1500, w_053_1501, w_053_1502, w_053_1503, w_053_1504, w_053_1506, w_053_1507, w_053_1508, w_053_1509, w_053_1510, w_053_1512, w_053_1513, w_053_1515, w_053_1516, w_053_1518, w_053_1519, w_053_1521, w_053_1522, w_053_1524, w_053_1527, w_053_1528, w_053_1529, w_053_1531, w_053_1532, w_053_1533, w_053_1534, w_053_1535, w_053_1536, w_053_1537, w_053_1538, w_053_1540, w_053_1542, w_053_1547, w_053_1548, w_053_1552, w_053_1553, w_053_1554, w_053_1557, w_053_1558, w_053_1561, w_053_1562, w_053_1563, w_053_1564, w_053_1565, w_053_1568, w_053_1569, w_053_1570, w_053_1571, w_053_1572, w_053_1573, w_053_1576, w_053_1577, w_053_1578, w_053_1579, w_053_1581, w_053_1582, w_053_1583, w_053_1584, w_053_1585, w_053_1586, w_053_1589, w_053_1590, w_053_1591, w_053_1592, w_053_1593, w_053_1594, w_053_1595, w_053_1597, w_053_1598, w_053_1599, w_053_1600, w_053_1601, w_053_1603, w_053_1604, w_053_1605, w_053_1606, w_053_1607, w_053_1609, w_053_1612, w_053_1613, w_053_1615, w_053_1619, w_053_1620, w_053_1621, w_053_1623, w_053_1624, w_053_1625, w_053_1629, w_053_1630, w_053_1632, w_053_1634, w_053_1635, w_053_1636, w_053_1638, w_053_1640, w_053_1642, w_053_1644, w_053_1645, w_053_1647, w_053_1648, w_053_1649, w_053_1650, w_053_1651, w_053_1652, w_053_1653, w_053_1654, w_053_1655, w_053_1656, w_053_1657, w_053_1658, w_053_1659, w_053_1661, w_053_1662, w_053_1663, w_053_1664, w_053_1665, w_053_1666, w_053_1667, w_053_1668, w_053_1669, w_053_1670, w_053_1671, w_053_1672, w_053_1673, w_053_1674, w_053_1675, w_053_1678, w_053_1679, w_053_1680, w_053_1681, w_053_1682, w_053_1683, w_053_1684, w_053_1685, w_053_1686, w_053_1687, w_053_1688, w_053_1690, w_053_1691, w_053_1692, w_053_1695, w_053_1697, w_053_1698, w_053_1699, w_053_1700, w_053_1701, w_053_1702, w_053_1703, w_053_1708, w_053_1709, w_053_1710, w_053_1714, w_053_1715, w_053_1717, w_053_1718, w_053_1719, w_053_1722, w_053_1725, w_053_1726, w_053_1727, w_053_1728, w_053_1729, w_053_1730, w_053_1735, w_053_1736, w_053_1737, w_053_1740, w_053_1741, w_053_1742, w_053_1745, w_053_1746, w_053_1747, w_053_1748, w_053_1749, w_053_1750, w_053_1751, w_053_1752, w_053_1753, w_053_1754, w_053_1755, w_053_1757, w_053_1758, w_053_1760, w_053_1761, w_053_1762, w_053_1763, w_053_1764, w_053_1765, w_053_1767, w_053_1768, w_053_1770, w_053_1772, w_053_1773, w_053_1774, w_053_1775, w_053_1776, w_053_1777, w_053_1778, w_053_1779, w_053_1780, w_053_1781, w_053_1783, w_053_1785, w_053_1786, w_053_1787, w_053_1788, w_053_1790, w_053_1792, w_053_1793, w_053_1794, w_053_1795, w_053_1797, w_053_1798, w_053_1799, w_053_1800, w_053_1801, w_053_1803, w_053_1805, w_053_1806, w_053_1808, w_053_1809, w_053_1810, w_053_1811, w_053_1812, w_053_1813, w_053_1814, w_053_1815, w_053_1816, w_053_1820, w_053_1821, w_053_1822, w_053_1825, w_053_1826, w_053_1828, w_053_1829, w_053_1832, w_053_1833, w_053_1834, w_053_1835, w_053_1836, w_053_1839, w_053_1840, w_053_1842, w_053_1846, w_053_1847, w_053_1849, w_053_1850, w_053_1851, w_053_1854, w_053_1855, w_053_1857, w_053_1860, w_053_1862, w_053_1863, w_053_1864, w_053_1865, w_053_1867, w_053_1868, w_053_1869, w_053_1871, w_053_1872, w_053_1874, w_053_1875, w_053_1876, w_053_1877, w_053_1878, w_053_1880, w_053_1881, w_053_1882, w_053_1883, w_053_1884, w_053_1885, w_053_1886, w_053_1887, w_053_1890, w_053_1891, w_053_1892, w_053_1895, w_053_1896, w_053_1899, w_053_1900, w_053_1901, w_053_1902, w_053_1903, w_053_1904, w_053_1905, w_053_1907, w_053_1908, w_053_1909, w_053_1910, w_053_1911, w_053_1914, w_053_1915, w_053_1916, w_053_1917, w_053_1919, w_053_1921, w_053_1923, w_053_1924, w_053_1928, w_053_1931, w_053_1932, w_053_1933, w_053_1935, w_053_1936, w_053_1938, w_053_1939, w_053_1943, w_053_1944, w_053_1945, w_053_1946, w_053_1947, w_053_1950, w_053_1951, w_053_1952, w_053_1954, w_053_1956, w_053_1957, w_053_1959, w_053_1960, w_053_1962;
  wire w_054_000, w_054_003, w_054_004, w_054_006, w_054_008, w_054_009, w_054_011, w_054_012, w_054_013, w_054_014, w_054_015, w_054_017, w_054_018, w_054_019, w_054_020, w_054_021, w_054_022, w_054_023, w_054_024, w_054_025, w_054_026, w_054_027, w_054_028, w_054_029, w_054_030, w_054_031, w_054_032, w_054_033, w_054_035, w_054_037, w_054_038, w_054_039, w_054_040, w_054_041, w_054_042, w_054_043, w_054_045, w_054_046, w_054_047, w_054_049, w_054_050, w_054_051, w_054_052, w_054_053, w_054_055, w_054_056, w_054_057, w_054_058, w_054_059, w_054_060, w_054_061, w_054_062, w_054_064, w_054_065, w_054_067, w_054_068, w_054_069, w_054_071, w_054_073, w_054_078, w_054_081, w_054_082, w_054_083, w_054_084, w_054_086, w_054_088, w_054_089, w_054_091, w_054_095, w_054_097, w_054_101, w_054_102, w_054_103, w_054_107, w_054_108, w_054_110, w_054_111, w_054_114, w_054_117, w_054_118, w_054_121, w_054_124, w_054_125, w_054_126, w_054_127, w_054_129, w_054_130, w_054_131, w_054_133, w_054_134, w_054_135, w_054_137, w_054_139, w_054_146, w_054_149, w_054_150, w_054_151, w_054_152, w_054_156, w_054_157, w_054_160, w_054_164, w_054_165, w_054_167, w_054_170, w_054_171, w_054_172, w_054_178, w_054_179, w_054_180, w_054_181, w_054_184, w_054_187, w_054_192, w_054_196, w_054_197, w_054_199, w_054_203, w_054_204, w_054_207, w_054_213, w_054_215, w_054_218, w_054_219, w_054_221, w_054_222, w_054_223, w_054_224, w_054_229, w_054_234, w_054_235, w_054_238, w_054_239, w_054_241, w_054_244, w_054_245, w_054_247, w_054_248, w_054_250, w_054_251, w_054_252, w_054_253, w_054_255, w_054_256, w_054_258, w_054_260, w_054_262, w_054_264, w_054_266, w_054_267, w_054_271, w_054_281, w_054_282, w_054_286, w_054_289, w_054_290, w_054_291, w_054_293, w_054_294, w_054_295, w_054_296, w_054_297, w_054_298, w_054_300, w_054_301, w_054_302, w_054_304, w_054_305, w_054_307, w_054_308, w_054_312, w_054_314, w_054_315, w_054_316, w_054_321, w_054_322, w_054_323, w_054_326, w_054_327, w_054_328, w_054_329, w_054_332, w_054_333, w_054_336, w_054_345, w_054_347, w_054_348, w_054_354, w_054_356, w_054_360, w_054_365, w_054_366, w_054_369, w_054_371, w_054_373, w_054_376, w_054_378, w_054_379, w_054_380, w_054_382, w_054_386, w_054_387, w_054_389, w_054_396, w_054_398, w_054_399, w_054_400, w_054_401, w_054_402, w_054_403, w_054_406, w_054_407, w_054_409, w_054_410, w_054_412, w_054_416, w_054_417, w_054_418, w_054_419, w_054_421, w_054_431, w_054_434, w_054_437, w_054_442, w_054_446, w_054_449, w_054_450, w_054_451, w_054_452, w_054_453, w_054_456, w_054_457, w_054_458, w_054_460, w_054_463, w_054_466, w_054_468, w_054_471, w_054_473, w_054_476, w_054_481, w_054_482, w_054_485, w_054_486, w_054_487, w_054_488, w_054_489, w_054_493, w_054_495, w_054_497, w_054_499, w_054_500, w_054_504, w_054_506, w_054_510, w_054_513, w_054_514, w_054_518, w_054_519, w_054_520, w_054_524, w_054_528, w_054_533, w_054_536, w_054_537, w_054_541, w_054_543, w_054_544, w_054_547, w_054_550, w_054_553, w_054_554, w_054_555, w_054_557, w_054_560, w_054_561, w_054_562, w_054_564, w_054_566, w_054_574, w_054_577, w_054_581, w_054_583, w_054_584, w_054_587, w_054_593, w_054_594, w_054_595, w_054_596, w_054_598, w_054_601, w_054_602, w_054_603, w_054_604, w_054_605, w_054_610, w_054_613, w_054_614, w_054_615, w_054_617, w_054_618, w_054_619, w_054_621, w_054_624, w_054_625, w_054_629, w_054_630, w_054_631, w_054_636, w_054_646, w_054_648, w_054_650, w_054_652, w_054_655, w_054_657, w_054_660, w_054_661, w_054_662, w_054_663, w_054_665, w_054_666, w_054_667, w_054_671, w_054_673, w_054_678, w_054_679, w_054_683, w_054_684, w_054_692, w_054_697, w_054_698, w_054_699, w_054_701, w_054_703, w_054_705, w_054_707, w_054_713, w_054_714, w_054_723, w_054_725, w_054_727, w_054_729, w_054_730, w_054_732, w_054_734, w_054_735, w_054_737, w_054_739, w_054_742, w_054_744, w_054_746, w_054_751, w_054_752, w_054_754, w_054_756, w_054_760, w_054_761, w_054_764, w_054_765, w_054_768, w_054_769, w_054_770, w_054_771, w_054_772, w_054_774, w_054_775, w_054_776, w_054_778, w_054_781, w_054_782, w_054_783, w_054_784, w_054_785, w_054_786, w_054_787, w_054_789, w_054_794, w_054_795, w_054_796, w_054_798, w_054_799, w_054_802, w_054_805, w_054_808, w_054_813, w_054_816, w_054_823, w_054_825, w_054_826, w_054_832, w_054_834, w_054_839, w_054_843, w_054_848, w_054_849, w_054_852, w_054_853, w_054_856, w_054_858, w_054_859, w_054_860, w_054_862, w_054_864, w_054_865, w_054_866, w_054_867, w_054_869, w_054_872, w_054_873, w_054_874, w_054_876, w_054_879, w_054_880, w_054_882, w_054_886, w_054_888, w_054_890, w_054_896, w_054_897, w_054_898, w_054_899, w_054_901, w_054_905, w_054_906, w_054_913, w_054_917, w_054_921, w_054_923, w_054_924, w_054_927, w_054_929, w_054_930, w_054_935, w_054_936, w_054_938, w_054_939, w_054_940, w_054_943, w_054_946, w_054_950, w_054_957, w_054_961, w_054_962, w_054_963, w_054_966, w_054_968, w_054_970, w_054_974, w_054_976, w_054_978, w_054_982, w_054_983, w_054_984, w_054_987, w_054_992, w_054_997, w_054_998, w_054_999, w_054_1002, w_054_1004, w_054_1006, w_054_1009, w_054_1013, w_054_1015, w_054_1018, w_054_1019, w_054_1020, w_054_1024, w_054_1025, w_054_1026, w_054_1027, w_054_1028, w_054_1029, w_054_1030, w_054_1031, w_054_1032, w_054_1036, w_054_1038, w_054_1039, w_054_1041, w_054_1043, w_054_1044, w_054_1045, w_054_1046, w_054_1047, w_054_1048, w_054_1049, w_054_1051, w_054_1053, w_054_1059, w_054_1062, w_054_1070, w_054_1076, w_054_1078, w_054_1079, w_054_1080, w_054_1081, w_054_1082, w_054_1083, w_054_1085, w_054_1087, w_054_1091, w_054_1093, w_054_1094, w_054_1096, w_054_1097, w_054_1100, w_054_1104, w_054_1110, w_054_1114, w_054_1115, w_054_1119, w_054_1122, w_054_1123, w_054_1124, w_054_1129, w_054_1131, w_054_1132, w_054_1135, w_054_1137, w_054_1141, w_054_1143, w_054_1144, w_054_1145, w_054_1151, w_054_1152, w_054_1155, w_054_1157, w_054_1158, w_054_1160, w_054_1161, w_054_1162, w_054_1163, w_054_1166, w_054_1169, w_054_1171, w_054_1173, w_054_1179, w_054_1180, w_054_1182, w_054_1184, w_054_1185, w_054_1188, w_054_1189, w_054_1191, w_054_1192, w_054_1193, w_054_1194, w_054_1195, w_054_1198, w_054_1199, w_054_1205, w_054_1207, w_054_1210, w_054_1211, w_054_1213, w_054_1217, w_054_1220, w_054_1224, w_054_1225, w_054_1235, w_054_1236, w_054_1238, w_054_1239, w_054_1242, w_054_1243, w_054_1244, w_054_1245, w_054_1246, w_054_1247, w_054_1248, w_054_1249, w_054_1250, w_054_1251, w_054_1255, w_054_1256, w_054_1257, w_054_1258, w_054_1259, w_054_1261, w_054_1264, w_054_1268, w_054_1272, w_054_1273, w_054_1275, w_054_1282, w_054_1284, w_054_1286, w_054_1287, w_054_1289, w_054_1294, w_054_1295, w_054_1296, w_054_1297, w_054_1298, w_054_1299, w_054_1301, w_054_1302, w_054_1308, w_054_1310, w_054_1311, w_054_1312, w_054_1314, w_054_1318, w_054_1319, w_054_1320, w_054_1322, w_054_1327, w_054_1329, w_054_1333, w_054_1334, w_054_1335, w_054_1336, w_054_1337, w_054_1344, w_054_1348, w_054_1349, w_054_1350, w_054_1351, w_054_1354, w_054_1355, w_054_1357, w_054_1361, w_054_1363, w_054_1364, w_054_1365, w_054_1367, w_054_1369, w_054_1371, w_054_1373, w_054_1378, w_054_1379, w_054_1380, w_054_1382, w_054_1386, w_054_1388, w_054_1392, w_054_1393, w_054_1394, w_054_1400, w_054_1401, w_054_1402, w_054_1403, w_054_1405, w_054_1408, w_054_1415, w_054_1417, w_054_1418, w_054_1420, w_054_1422, w_054_1423, w_054_1424, w_054_1426, w_054_1427, w_054_1428, w_054_1430, w_054_1434, w_054_1435, w_054_1437, w_054_1442, w_054_1443, w_054_1447, w_054_1448, w_054_1450, w_054_1451, w_054_1452, w_054_1460, w_054_1461, w_054_1462, w_054_1463, w_054_1466, w_054_1468, w_054_1469, w_054_1471, w_054_1472, w_054_1474, w_054_1477, w_054_1480, w_054_1481, w_054_1482, w_054_1484, w_054_1485, w_054_1486, w_054_1492, w_054_1494, w_054_1495, w_054_1496, w_054_1497, w_054_1499, w_054_1501, w_054_1502, w_054_1505, w_054_1511, w_054_1514, w_054_1515, w_054_1516, w_054_1517, w_054_1518, w_054_1520, w_054_1521, w_054_1525, w_054_1526, w_054_1528, w_054_1530, w_054_1534, w_054_1535, w_054_1541, w_054_1544, w_054_1545, w_054_1546, w_054_1547, w_054_1550, w_054_1551, w_054_1552, w_054_1555, w_054_1556, w_054_1557, w_054_1559, w_054_1561, w_054_1562, w_054_1563, w_054_1564, w_054_1565, w_054_1567, w_054_1568, w_054_1574, w_054_1576, w_054_1582, w_054_1583, w_054_1584, w_054_1585, w_054_1586, w_054_1587, w_054_1592, w_054_1597, w_054_1605, w_054_1609, w_054_1611, w_054_1612, w_054_1613, w_054_1616, w_054_1619, w_054_1620, w_054_1627, w_054_1630, w_054_1632, w_054_1634, w_054_1638, w_054_1641, w_054_1646, w_054_1648, w_054_1649, w_054_1650, w_054_1653, w_054_1654, w_054_1655, w_054_1658, w_054_1662, w_054_1663, w_054_1665, w_054_1666, w_054_1669, w_054_1670, w_054_1674, w_054_1675, w_054_1676, w_054_1677, w_054_1679, w_054_1680, w_054_1681, w_054_1682, w_054_1686, w_054_1687, w_054_1688, w_054_1690, w_054_1695, w_054_1696, w_054_1697, w_054_1701, w_054_1710, w_054_1711, w_054_1713, w_054_1714, w_054_1716, w_054_1717, w_054_1720, w_054_1721, w_054_1723, w_054_1724, w_054_1725, w_054_1727, w_054_1731, w_054_1732, w_054_1733, w_054_1735, w_054_1736, w_054_1739, w_054_1740, w_054_1746, w_054_1747, w_054_1749, w_054_1750, w_054_1751, w_054_1752, w_054_1753, w_054_1754, w_054_1757, w_054_1761, w_054_1763, w_054_1778, w_054_1779, w_054_1781, w_054_1782, w_054_1783, w_054_1784, w_054_1787, w_054_1788, w_054_1791, w_054_1792, w_054_1798, w_054_1800, w_054_1804, w_054_1805, w_054_1806, w_054_1807, w_054_1808, w_054_1811, w_054_1814, w_054_1816, w_054_1818, w_054_1823, w_054_1825, w_054_1830, w_054_1832, w_054_1833, w_054_1834, w_054_1838, w_054_1841, w_054_1843, w_054_1844, w_054_1845, w_054_1846, w_054_1849, w_054_1852, w_054_1853, w_054_1854, w_054_1856, w_054_1857, w_054_1858, w_054_1859, w_054_1860, w_054_1863, w_054_1864, w_054_1867, w_054_1868, w_054_1873, w_054_1875, w_054_1878, w_054_1881, w_054_1884, w_054_1886, w_054_1887, w_054_1892, w_054_1893, w_054_1897, w_054_1898, w_054_1899, w_054_1900, w_054_1904, w_054_1905, w_054_1906, w_054_1907, w_054_1908, w_054_1911, w_054_1915, w_054_1922, w_054_1923, w_054_1925, w_054_1929, w_054_1930, w_054_1931, w_054_1932, w_054_1935, w_054_1937, w_054_1944, w_054_1945, w_054_1946, w_054_1947, w_054_1949, w_054_1955, w_054_1958, w_054_1963, w_054_1965, w_054_1967, w_054_1969, w_054_1971, w_054_1972, w_054_1977, w_054_1982, w_054_1984, w_054_1987, w_054_1989, w_054_1992, w_054_1994, w_054_1996, w_054_1997, w_054_2000, w_054_2004, w_054_2007, w_054_2008, w_054_2009, w_054_2013, w_054_2019, w_054_2022, w_054_2023, w_054_2024, w_054_2025, w_054_2031, w_054_2032, w_054_2033, w_054_2035, w_054_2036, w_054_2037, w_054_2038, w_054_2039, w_054_2040, w_054_2043, w_054_2044, w_054_2047, w_054_2048, w_054_2049, w_054_2051, w_054_2055, w_054_2058, w_054_2059, w_054_2060, w_054_2061, w_054_2062, w_054_2063, w_054_2074, w_054_2075, w_054_2076, w_054_2077, w_054_2080, w_054_2081, w_054_2083, w_054_2086, w_054_2087, w_054_2088, w_054_2097, w_054_2098, w_054_2099, w_054_2102, w_054_2105, w_054_2106, w_054_2108, w_054_2109, w_054_2110, w_054_2114, w_054_2115, w_054_2116, w_054_2117, w_054_2124, w_054_2125, w_054_2126, w_054_2128, w_054_2129, w_054_2134, w_054_2138, w_054_2142, w_054_2147, w_054_2148, w_054_2149, w_054_2150, w_054_2151, w_054_2155, w_054_2157, w_054_2163, w_054_2164, w_054_2166, w_054_2168, w_054_2169, w_054_2171, w_054_2172, w_054_2173, w_054_2174, w_054_2178, w_054_2179, w_054_2181, w_054_2184, w_054_2188, w_054_2189, w_054_2191, w_054_2192, w_054_2194, w_054_2195, w_054_2196, w_054_2197, w_054_2198, w_054_2200, w_054_2201, w_054_2202, w_054_2203, w_054_2208, w_054_2209, w_054_2210, w_054_2211, w_054_2212, w_054_2214, w_054_2215, w_054_2216, w_054_2218, w_054_2219, w_054_2222, w_054_2223, w_054_2224, w_054_2228, w_054_2229, w_054_2233, w_054_2235, w_054_2238, w_054_2240, w_054_2242, w_054_2244, w_054_2246, w_054_2250, w_054_2254, w_054_2255, w_054_2256, w_054_2259, w_054_2261, w_054_2263, w_054_2264, w_054_2268, w_054_2270, w_054_2271, w_054_2275, w_054_2276, w_054_2279, w_054_2284, w_054_2285, w_054_2286, w_054_2290, w_054_2292, w_054_2293, w_054_2299, w_054_2303, w_054_2309, w_054_2311, w_054_2313, w_054_2315, w_054_2317, w_054_2318, w_054_2319, w_054_2320, w_054_2324, w_054_2327, w_054_2328, w_054_2329, w_054_2331, w_054_2335, w_054_2338, w_054_2339, w_054_2343, w_054_2346, w_054_2347, w_054_2349, w_054_2350, w_054_2355, w_054_2356, w_054_2358, w_054_2359, w_054_2362, w_054_2363, w_054_2364, w_054_2365, w_054_2368, w_054_2369, w_054_2370, w_054_2373, w_054_2374, w_054_2375, w_054_2380, w_054_2382, w_054_2385, w_054_2388, w_054_2393, w_054_2394, w_054_2395, w_054_2398, w_054_2399, w_054_2400, w_054_2402, w_054_2404, w_054_2405, w_054_2406, w_054_2410, w_054_2411, w_054_2412, w_054_2415, w_054_2417, w_054_2420, w_054_2421, w_054_2425, w_054_2426, w_054_2431, w_054_2434, w_054_2436, w_054_2439, w_054_2440, w_054_2442, w_054_2443, w_054_2452, w_054_2453, w_054_2456, w_054_2457, w_054_2460, w_054_2463, w_054_2464, w_054_2466, w_054_2468, w_054_2470, w_054_2472, w_054_2474, w_054_2476, w_054_2477, w_054_2480, w_054_2481, w_054_2485, w_054_2489, w_054_2490, w_054_2492, w_054_2501, w_054_2502, w_054_2503, w_054_2506, w_054_2507, w_054_2508, w_054_2509, w_054_2511, w_054_2516, w_054_2519, w_054_2522, w_054_2523, w_054_2525, w_054_2527, w_054_2528, w_054_2530, w_054_2533, w_054_2534, w_054_2536, w_054_2539, w_054_2540, w_054_2543, w_054_2544, w_054_2545, w_054_2546, w_054_2549, w_054_2550, w_054_2551, w_054_2552, w_054_2553, w_054_2554, w_054_2557, w_054_2558, w_054_2559, w_054_2562, w_054_2564, w_054_2566, w_054_2567, w_054_2569, w_054_2570, w_054_2572, w_054_2576, w_054_2577, w_054_2579, w_054_2583, w_054_2584, w_054_2586, w_054_2589, w_054_2591, w_054_2599, w_054_2604, w_054_2607, w_054_2608, w_054_2611, w_054_2612, w_054_2614, w_054_2616, w_054_2618, w_054_2620, w_054_2623, w_054_2625, w_054_2628, w_054_2631, w_054_2633, w_054_2634, w_054_2635, w_054_2637, w_054_2638, w_054_2639, w_054_2640, w_054_2641, w_054_2642, w_054_2645, w_054_2654, w_054_2656, w_054_2659, w_054_2661, w_054_2663, w_054_2667, w_054_2668, w_054_2669, w_054_2670, w_054_2673, w_054_2677, w_054_2679, w_054_2680, w_054_2682, w_054_2685, w_054_2687, w_054_2689, w_054_2692, w_054_2698, w_054_2702, w_054_2703, w_054_2704, w_054_2705, w_054_2706, w_054_2707, w_054_2708, w_054_2709, w_054_2710, w_054_2711, w_054_2712, w_054_2713, w_054_2714, w_054_2716, w_054_2717, w_054_2721, w_054_2722, w_054_2724, w_054_2725, w_054_2727, w_054_2730, w_054_2731, w_054_2732, w_054_2734, w_054_2736, w_054_2737, w_054_2739, w_054_2741, w_054_2742, w_054_2743, w_054_2744, w_054_2745, w_054_2746, w_054_2749, w_054_2750, w_054_2751, w_054_2753, w_054_2755, w_054_2756, w_054_2757, w_054_2758, w_054_2767, w_054_2771, w_054_2773, w_054_2777, w_054_2778, w_054_2784, w_054_2794, w_054_2796, w_054_2798, w_054_2799, w_054_2801, w_054_2802, w_054_2805, w_054_2806, w_054_2808, w_054_2809, w_054_2810, w_054_2811, w_054_2812, w_054_2816, w_054_2818, w_054_2820, w_054_2821, w_054_2823, w_054_2826, w_054_2830, w_054_2835, w_054_2837, w_054_2838, w_054_2845, w_054_2848, w_054_2849, w_054_2850, w_054_2854, w_054_2855, w_054_2858, w_054_2859, w_054_2862, w_054_2864, w_054_2865, w_054_2868, w_054_2869, w_054_2871, w_054_2872, w_054_2873, w_054_2875, w_054_2876, w_054_2880, w_054_2882, w_054_2884, w_054_2888, w_054_2890, w_054_2891, w_054_2892, w_054_2893, w_054_2894, w_054_2897, w_054_2899, w_054_2900, w_054_2901, w_054_2902, w_054_2903, w_054_2904, w_054_2905, w_054_2906, w_054_2910, w_054_2912, w_054_2913, w_054_2916, w_054_2917, w_054_2919, w_054_2923, w_054_2924, w_054_2925, w_054_2929, w_054_2930, w_054_2932, w_054_2933, w_054_2934, w_054_2935, w_054_2936, w_054_2939, w_054_2940, w_054_2942, w_054_2946, w_054_2947, w_054_2948, w_054_2951, w_054_2952, w_054_2953, w_054_2954, w_054_2957, w_054_2959, w_054_2960, w_054_2963, w_054_2964, w_054_2966, w_054_2969, w_054_2970, w_054_2971, w_054_2974, w_054_2977, w_054_2978, w_054_2980, w_054_2992, w_054_2994, w_054_2997, w_054_2998, w_054_2999, w_054_3000, w_054_3001, w_054_3002, w_054_3007, w_054_3008, w_054_3009, w_054_3013, w_054_3014, w_054_3016, w_054_3019, w_054_3020, w_054_3022, w_054_3023, w_054_3025, w_054_3030, w_054_3031, w_054_3033, w_054_3038, w_054_3040, w_054_3041, w_054_3044, w_054_3052, w_054_3053, w_054_3054, w_054_3056, w_054_3061, w_054_3065, w_054_3067, w_054_3068, w_054_3069, w_054_3070, w_054_3076, w_054_3077, w_054_3082, w_054_3084, w_054_3085, w_054_3090, w_054_3092, w_054_3094, w_054_3097, w_054_3098, w_054_3100, w_054_3101, w_054_3104, w_054_3105, w_054_3106, w_054_3114, w_054_3117, w_054_3118, w_054_3121, w_054_3122, w_054_3123, w_054_3125, w_054_3127, w_054_3128, w_054_3129, w_054_3132, w_054_3136, w_054_3138, w_054_3139, w_054_3140, w_054_3142, w_054_3147, w_054_3149, w_054_3150, w_054_3153, w_054_3154, w_054_3156, w_054_3159, w_054_3161, w_054_3165, w_054_3168, w_054_3170, w_054_3172, w_054_3173, w_054_3174, w_054_3177, w_054_3180, w_054_3182, w_054_3185, w_054_3187, w_054_3188, w_054_3192, w_054_3193, w_054_3195, w_054_3196, w_054_3200, w_054_3203, w_054_3209, w_054_3210, w_054_3212, w_054_3218, w_054_3219, w_054_3221, w_054_3223, w_054_3224, w_054_3226, w_054_3227, w_054_3229, w_054_3230, w_054_3231, w_054_3232, w_054_3235, w_054_3237, w_054_3239, w_054_3242, w_054_3243, w_054_3245, w_054_3247, w_054_3248, w_054_3250, w_054_3253, w_054_3254, w_054_3256, w_054_3258, w_054_3261, w_054_3262, w_054_3263, w_054_3264, w_054_3268, w_054_3269, w_054_3270, w_054_3272, w_054_3275, w_054_3276, w_054_3277, w_054_3278, w_054_3281, w_054_3286, w_054_3290, w_054_3291, w_054_3292, w_054_3293, w_054_3294, w_054_3295, w_054_3297, w_054_3298, w_054_3301, w_054_3304, w_054_3305, w_054_3308, w_054_3314, w_054_3316, w_054_3319, w_054_3321, w_054_3322, w_054_3324, w_054_3326, w_054_3327, w_054_3328, w_054_3330, w_054_3332, w_054_3338, w_054_3339, w_054_3340, w_054_3344, w_054_3349, w_054_3351, w_054_3354, w_054_3356, w_054_3357, w_054_3358, w_054_3359, w_054_3361, w_054_3363, w_054_3369, w_054_3370, w_054_3372, w_054_3374, w_054_3375, w_054_3377, w_054_3378, w_054_3379, w_054_3380, w_054_3382, w_054_3388, w_054_3390, w_054_3392, w_054_3396, w_054_3399, w_054_3400, w_054_3402, w_054_3403, w_054_3404, w_054_3405, w_054_3409, w_054_3410, w_054_3411, w_054_3413, w_054_3419, w_054_3427, w_054_3430, w_054_3432, w_054_3436, w_054_3438, w_054_3439, w_054_3441, w_054_3442, w_054_3445, w_054_3446, w_054_3447, w_054_3449, w_054_3452, w_054_3455, w_054_3456, w_054_3457, w_054_3458, w_054_3461, w_054_3462, w_054_3465, w_054_3471, w_054_3476, w_054_3479, w_054_3482, w_054_3483, w_054_3487, w_054_3488, w_054_3490, w_054_3491, w_054_3492, w_054_3493, w_054_3494, w_054_3495, w_054_3496, w_054_3501, w_054_3506, w_054_3507, w_054_3509, w_054_3510, w_054_3511, w_054_3513, w_054_3520, w_054_3521, w_054_3525, w_054_3526, w_054_3527, w_054_3529, w_054_3532, w_054_3533, w_054_3536, w_054_3537, w_054_3538, w_054_3543, w_054_3544, w_054_3545, w_054_3548, w_054_3552, w_054_3554, w_054_3560, w_054_3561, w_054_3566, w_054_3567, w_054_3569, w_054_3572, w_054_3577, w_054_3580, w_054_3581, w_054_3583, w_054_3585, w_054_3586, w_054_3592, w_054_3593, w_054_3597, w_054_3598, w_054_3599, w_054_3600, w_054_3601, w_054_3603, w_054_3604, w_054_3605, w_054_3608, w_054_3609, w_054_3610, w_054_3611, w_054_3612, w_054_3615, w_054_3617, w_054_3619, w_054_3621, w_054_3622, w_054_3624, w_054_3630, w_054_3632, w_054_3634, w_054_3635, w_054_3636, w_054_3637, w_054_3643, w_054_3645, w_054_3646, w_054_3649, w_054_3651, w_054_3653, w_054_3655, w_054_3656, w_054_3659, w_054_3662, w_054_3663, w_054_3668, w_054_3669, w_054_3670, w_054_3671, w_054_3672, w_054_3675, w_054_3682, w_054_3683, w_054_3687, w_054_3688, w_054_3689, w_054_3690, w_054_3694, w_054_3696, w_054_3697, w_054_3698, w_054_3699, w_054_3704, w_054_3706, w_054_3707, w_054_3709, w_054_3710, w_054_3713, w_054_3714, w_054_3716, w_054_3717, w_054_3718, w_054_3719, w_054_3722, w_054_3725, w_054_3730, w_054_3732, w_054_3735, w_054_3738, w_054_3739, w_054_3741, w_054_3742, w_054_3743, w_054_3746, w_054_3747, w_054_3748, w_054_3749, w_054_3750, w_054_3751, w_054_3753, w_054_3754, w_054_3755, w_054_3758, w_054_3760, w_054_3762, w_054_3763, w_054_3766, w_054_3768, w_054_3770, w_054_3771, w_054_3772, w_054_3773, w_054_3777, w_054_3786, w_054_3787, w_054_3790, w_054_3792, w_054_3794, w_054_3795, w_054_3796, w_054_3798, w_054_3799, w_054_3801, w_054_3802, w_054_3804, w_054_3805, w_054_3807, w_054_3809, w_054_3813, w_054_3814, w_054_3817, w_054_3818, w_054_3819, w_054_3823, w_054_3827, w_054_3829, w_054_3831, w_054_3832, w_054_3833, w_054_3834, w_054_3835, w_054_3840, w_054_3843, w_054_3845, w_054_3848, w_054_3849, w_054_3851, w_054_3852, w_054_3856, w_054_3857, w_054_3859, w_054_3862, w_054_3863, w_054_3864, w_054_3866, w_054_3868, w_054_3870, w_054_3871, w_054_3872, w_054_3873, w_054_3874, w_054_3878, w_054_3879, w_054_3883, w_054_3885, w_054_3886, w_054_3887, w_054_3890, w_054_3893, w_054_3894, w_054_3897, w_054_3898, w_054_3902, w_054_3905, w_054_3906, w_054_3910, w_054_3911, w_054_3914, w_054_3918, w_054_3919, w_054_3920, w_054_3923, w_054_3925, w_054_3928, w_054_3933, w_054_3939, w_054_3940, w_054_3945, w_054_3946, w_054_3947, w_054_3948, w_054_3949, w_054_3951, w_054_3955, w_054_3957, w_054_3958, w_054_3963, w_054_3964, w_054_3966, w_054_3972, w_054_3977, w_054_3978, w_054_3979, w_054_3980, w_054_3986, w_054_3990, w_054_3993, w_054_3996, w_054_3997, w_054_4006, w_054_4009, w_054_4010, w_054_4013, w_054_4014, w_054_4016, w_054_4018, w_054_4022, w_054_4026, w_054_4028, w_054_4036, w_054_4038, w_054_4039, w_054_4040, w_054_4041, w_054_4043, w_054_4048, w_054_4050, w_054_4051, w_054_4053, w_054_4054, w_054_4056, w_054_4057, w_054_4058, w_054_4059, w_054_4060, w_054_4064, w_054_4065, w_054_4074, w_054_4077, w_054_4080, w_054_4083, w_054_4084, w_054_4085, w_054_4089, w_054_4092, w_054_4093, w_054_4094, w_054_4098, w_054_4099, w_054_4103, w_054_4105, w_054_4111, w_054_4113, w_054_4115, w_054_4116, w_054_4118, w_054_4120, w_054_4122, w_054_4125, w_054_4127, w_054_4128, w_054_4130, w_054_4133, w_054_4134, w_054_4136, w_054_4138, w_054_4139, w_054_4143, w_054_4146, w_054_4148, w_054_4151, w_054_4152, w_054_4153, w_054_4155, w_054_4158, w_054_4159, w_054_4160, w_054_4161, w_054_4162, w_054_4164, w_054_4165, w_054_4166, w_054_4167, w_054_4170, w_054_4171, w_054_4172, w_054_4174, w_054_4175, w_054_4176, w_054_4177, w_054_4183, w_054_4184, w_054_4186, w_054_4187, w_054_4192, w_054_4195, w_054_4196, w_054_4199, w_054_4200, w_054_4203, w_054_4204, w_054_4206, w_054_4208, w_054_4209, w_054_4210, w_054_4211, w_054_4212, w_054_4214, w_054_4216, w_054_4218, w_054_4219, w_054_4220, w_054_4221, w_054_4223, w_054_4224, w_054_4225, w_054_4229, w_054_4230, w_054_4231, w_054_4233, w_054_4237, w_054_4239, w_054_4243, w_054_4246, w_054_4248, w_054_4250, w_054_4251, w_054_4253, w_054_4254, w_054_4258, w_054_4259, w_054_4260, w_054_4261, w_054_4263, w_054_4265, w_054_4270, w_054_4271, w_054_4272, w_054_4274, w_054_4277, w_054_4285, w_054_4286, w_054_4287, w_054_4288, w_054_4289, w_054_4291, w_054_4294, w_054_4296, w_054_4297, w_054_4298, w_054_4303, w_054_4306, w_054_4308, w_054_4311, w_054_4312, w_054_4316, w_054_4321, w_054_4322, w_054_4325, w_054_4327, w_054_4328, w_054_4329, w_054_4332, w_054_4333, w_054_4334, w_054_4336, w_054_4338, w_054_4342, w_054_4343, w_054_4349, w_054_4353, w_054_4354, w_054_4357, w_054_4360, w_054_4362, w_054_4365, w_054_4368, w_054_4369, w_054_4370, w_054_4380, w_054_4381, w_054_4382, w_054_4391, w_054_4394, w_054_4397, w_054_4398, w_054_4399, w_054_4401, w_054_4403, w_054_4404, w_054_4408, w_054_4409, w_054_4415, w_054_4418, w_054_4419, w_054_4421, w_054_4422, w_054_4424, w_054_4427, w_054_4429, w_054_4433, w_054_4434, w_054_4435, w_054_4436, w_054_4438, w_054_4439, w_054_4440, w_054_4442, w_054_4444, w_054_4445, w_054_4448, w_054_4449, w_054_4451, w_054_4452, w_054_4454, w_054_4455, w_054_4459, w_054_4460, w_054_4461, w_054_4464, w_054_4468, w_054_4473, w_054_4474, w_054_4476, w_054_4479, w_054_4482, w_054_4484, w_054_4485, w_054_4489, w_054_4490, w_054_4494, w_054_4500, w_054_4504, w_054_4506, w_054_4508, w_054_4509, w_054_4512, w_054_4513, w_054_4514, w_054_4515, w_054_4516, w_054_4517, w_054_4519, w_054_4520, w_054_4521, w_054_4525, w_054_4526, w_054_4529, w_054_4531, w_054_4538, w_054_4542, w_054_4544, w_054_4546, w_054_4548, w_054_4550, w_054_4551, w_054_4553, w_054_4555, w_054_4557, w_054_4558, w_054_4559, w_054_4562, w_054_4564, w_054_4565, w_054_4566, w_054_4569, w_054_4570, w_054_4573, w_054_4574, w_054_4575, w_054_4579, w_054_4581, w_054_4582, w_054_4583, w_054_4584, w_054_4589, w_054_4592, w_054_4593, w_054_4594, w_054_4596, w_054_4597, w_054_4599, w_054_4600, w_054_4603, w_054_4606, w_054_4612, w_054_4615, w_054_4617, w_054_4619, w_054_4622, w_054_4624, w_054_4626, w_054_4628, w_054_4629, w_054_4631, w_054_4636, w_054_4637, w_054_4638, w_054_4639, w_054_4644, w_054_4645, w_054_4648, w_054_4649, w_054_4651, w_054_4654, w_054_4656, w_054_4657, w_054_4659, w_054_4660, w_054_4662, w_054_4663, w_054_4664, w_054_4666, w_054_4668, w_054_4672, w_054_4673, w_054_4675, w_054_4676, w_054_4677, w_054_4678, w_054_4679, w_054_4681, w_054_4687, w_054_4688, w_054_4689, w_054_4691, w_054_4693, w_054_4698, w_054_4701, w_054_4705, w_054_4707, w_054_4710, w_054_4711, w_054_4712, w_054_4718, w_054_4722, w_054_4723, w_054_4725, w_054_4726, w_054_4727, w_054_4728, w_054_4736, w_054_4739, w_054_4740, w_054_4741, w_054_4742, w_054_4744, w_054_4745, w_054_4746, w_054_4749, w_054_4753, w_054_4758, w_054_4760, w_054_4764, w_054_4766, w_054_4772, w_054_4774, w_054_4777, w_054_4778, w_054_4779, w_054_4784, w_054_4788, w_054_4791, w_054_4796, w_054_4800, w_054_4802, w_054_4804, w_054_4805, w_054_4806, w_054_4807, w_054_4813, w_054_4814, w_054_4815, w_054_4816, w_054_4817, w_054_4819, w_054_4820, w_054_4822, w_054_4823, w_054_4824, w_054_4825, w_054_4826, w_054_4833, w_054_4838, w_054_4839, w_054_4840, w_054_4846, w_054_4849, w_054_4850, w_054_4853, w_054_4854, w_054_4855, w_054_4856, w_054_4857, w_054_4859, w_054_4860, w_054_4864, w_054_4865, w_054_4867, w_054_4870, w_054_4871, w_054_4873, w_054_4875, w_054_4876, w_054_4877, w_054_4878, w_054_4879, w_054_4882, w_054_4885, w_054_4886, w_054_4887, w_054_4888, w_054_4891, w_054_4892, w_054_4895, w_054_4899, w_054_4900, w_054_4906, w_054_4908, w_054_4909, w_054_4911, w_054_4912, w_054_4913, w_054_4915, w_054_4917, w_054_4919, w_054_4921, w_054_4923, w_054_4925;
  wire w_055_001, w_055_002, w_055_004, w_055_005, w_055_006, w_055_008, w_055_011, w_055_012, w_055_013, w_055_014, w_055_015, w_055_016, w_055_017, w_055_018, w_055_020, w_055_021, w_055_022, w_055_024, w_055_025, w_055_027, w_055_028, w_055_029, w_055_030, w_055_031, w_055_033, w_055_034, w_055_035, w_055_036, w_055_037, w_055_040, w_055_042, w_055_043, w_055_045, w_055_048, w_055_050, w_055_051, w_055_052, w_055_053, w_055_054, w_055_055, w_055_057, w_055_058, w_055_059, w_055_060, w_055_061, w_055_062, w_055_064, w_055_065, w_055_066, w_055_067, w_055_072, w_055_073, w_055_076, w_055_078, w_055_079, w_055_080, w_055_084, w_055_085, w_055_086, w_055_088, w_055_091, w_055_092, w_055_094, w_055_095, w_055_096, w_055_097, w_055_099, w_055_101, w_055_102, w_055_104, w_055_105, w_055_106, w_055_107, w_055_108, w_055_109, w_055_110, w_055_111, w_055_112, w_055_115, w_055_117, w_055_118, w_055_120, w_055_123, w_055_124, w_055_125, w_055_126, w_055_127, w_055_128, w_055_132, w_055_133, w_055_134, w_055_135, w_055_136, w_055_139, w_055_140, w_055_142, w_055_145, w_055_146, w_055_147, w_055_148, w_055_149, w_055_151, w_055_152, w_055_153, w_055_154, w_055_155, w_055_156, w_055_160, w_055_161, w_055_162, w_055_163, w_055_164, w_055_165, w_055_166, w_055_168, w_055_169, w_055_171, w_055_172, w_055_174, w_055_175, w_055_178, w_055_180, w_055_181, w_055_182, w_055_183, w_055_184, w_055_185, w_055_186, w_055_187, w_055_188, w_055_190, w_055_195, w_055_196, w_055_197, w_055_199, w_055_200, w_055_201, w_055_202, w_055_204, w_055_206, w_055_209, w_055_210, w_055_211, w_055_212, w_055_213, w_055_214, w_055_215, w_055_216, w_055_217, w_055_218, w_055_219, w_055_220, w_055_222, w_055_223, w_055_224, w_055_225, w_055_228, w_055_229, w_055_230, w_055_231, w_055_232, w_055_235, w_055_236, w_055_237, w_055_239, w_055_241, w_055_243, w_055_244, w_055_245, w_055_246, w_055_247, w_055_248, w_055_250, w_055_252, w_055_253, w_055_254, w_055_255, w_055_257, w_055_258, w_055_259, w_055_260, w_055_261, w_055_263, w_055_265, w_055_266, w_055_267, w_055_271, w_055_273, w_055_275, w_055_276, w_055_277, w_055_278, w_055_279, w_055_280, w_055_281, w_055_285, w_055_287, w_055_289, w_055_290, w_055_291, w_055_292, w_055_293, w_055_295, w_055_296, w_055_297, w_055_298, w_055_299, w_055_302, w_055_303, w_055_304, w_055_305, w_055_306, w_055_308, w_055_310, w_055_311, w_055_312, w_055_313, w_055_314, w_055_315, w_055_316, w_055_317, w_055_318, w_055_321, w_055_322, w_055_323, w_055_325, w_055_326, w_055_327, w_055_328, w_055_330, w_055_332, w_055_333, w_055_334, w_055_336, w_055_337, w_055_338, w_055_339, w_055_340, w_055_341, w_055_343, w_055_345, w_055_346, w_055_350, w_055_352, w_055_353, w_055_356, w_055_357, w_055_359, w_055_360, w_055_363, w_055_364, w_055_366, w_055_369, w_055_370, w_055_371, w_055_372, w_055_374, w_055_376, w_055_377, w_055_378, w_055_380, w_055_383, w_055_385, w_055_386, w_055_390, w_055_393, w_055_394, w_055_395, w_055_396, w_055_397, w_055_398, w_055_399, w_055_400, w_055_401, w_055_402, w_055_404, w_055_405, w_055_411, w_055_414, w_055_415, w_055_416, w_055_417, w_055_419, w_055_420, w_055_422, w_055_423, w_055_424, w_055_425, w_055_427, w_055_428, w_055_431, w_055_432, w_055_433, w_055_434, w_055_435, w_055_438, w_055_439, w_055_440, w_055_441, w_055_442, w_055_443, w_055_445, w_055_446, w_055_447, w_055_448, w_055_449, w_055_451, w_055_452, w_055_454, w_055_455, w_055_460, w_055_461, w_055_462, w_055_463, w_055_467, w_055_468, w_055_469, w_055_470, w_055_472, w_055_473, w_055_474, w_055_475, w_055_476, w_055_477, w_055_478, w_055_479, w_055_480, w_055_481, w_055_482, w_055_484, w_055_486, w_055_487, w_055_488, w_055_489, w_055_490, w_055_491, w_055_492, w_055_493, w_055_494, w_055_495, w_055_496, w_055_498, w_055_499, w_055_501, w_055_502, w_055_503, w_055_504, w_055_505, w_055_506, w_055_507, w_055_508, w_055_509, w_055_510, w_055_511, w_055_513, w_055_516, w_055_517, w_055_518, w_055_519, w_055_520, w_055_521, w_055_523, w_055_524, w_055_525, w_055_527, w_055_528, w_055_530, w_055_531, w_055_532, w_055_533, w_055_534, w_055_535, w_055_537, w_055_539, w_055_540, w_055_541, w_055_542, w_055_544, w_055_545, w_055_546, w_055_547, w_055_548, w_055_549, w_055_550, w_055_551, w_055_552, w_055_553, w_055_554, w_055_556, w_055_558, w_055_559, w_055_560, w_055_561, w_055_564, w_055_566, w_055_567, w_055_568, w_055_569, w_055_570, w_055_571, w_055_573, w_055_574, w_055_575, w_055_576, w_055_577, w_055_578, w_055_579, w_055_582, w_055_584, w_055_586, w_055_587, w_055_588, w_055_592, w_055_593, w_055_594, w_055_595, w_055_596, w_055_597, w_055_598, w_055_599, w_055_600, w_055_601, w_055_602, w_055_603, w_055_604, w_055_606, w_055_607, w_055_608, w_055_611, w_055_612, w_055_613, w_055_614, w_055_615, w_055_616, w_055_617, w_055_619, w_055_620, w_055_621, w_055_622, w_055_623, w_055_624, w_055_625, w_055_626, w_055_629, w_055_633, w_055_634, w_055_637, w_055_638, w_055_640, w_055_642, w_055_643, w_055_644, w_055_646, w_055_648, w_055_649, w_055_651, w_055_652, w_055_653, w_055_655, w_055_656, w_055_658, w_055_660, w_055_661, w_055_662, w_055_663, w_055_664, w_055_665, w_055_666, w_055_667, w_055_670, w_055_671, w_055_672, w_055_674, w_055_676, w_055_678, w_055_679, w_055_681, w_055_682, w_055_687, w_055_688, w_055_689, w_055_690, w_055_691, w_055_692, w_055_694, w_055_695, w_055_697, w_055_698, w_055_700, w_055_703, w_055_704, w_055_705, w_055_706, w_055_709, w_055_713, w_055_714, w_055_715, w_055_717, w_055_719, w_055_720, w_055_721, w_055_723, w_055_724, w_055_725, w_055_726, w_055_727, w_055_728, w_055_729, w_055_730, w_055_731, w_055_732, w_055_733, w_055_735, w_055_738, w_055_741, w_055_742, w_055_745, w_055_748, w_055_750, w_055_752, w_055_753, w_055_756, w_055_757, w_055_758, w_055_759, w_055_760, w_055_762, w_055_763, w_055_765, w_055_766, w_055_767, w_055_768, w_055_770, w_055_772, w_055_773, w_055_774, w_055_781, w_055_782, w_055_783, w_055_784, w_055_787, w_055_788, w_055_790, w_055_791, w_055_793, w_055_796, w_055_797, w_055_799, w_055_800, w_055_802, w_055_804, w_055_806, w_055_807, w_055_808, w_055_809, w_055_810, w_055_811, w_055_812, w_055_813, w_055_814, w_055_816, w_055_820, w_055_821, w_055_824, w_055_826, w_055_829, w_055_830, w_055_832, w_055_833, w_055_834, w_055_835, w_055_836, w_055_837, w_055_838, w_055_839, w_055_840, w_055_842, w_055_843, w_055_844, w_055_845, w_055_846, w_055_848, w_055_849, w_055_851, w_055_852, w_055_853, w_055_856, w_055_857, w_055_859, w_055_860, w_055_862, w_055_863, w_055_864, w_055_865, w_055_867, w_055_869, w_055_870, w_055_872, w_055_873, w_055_875, w_055_876, w_055_878, w_055_879, w_055_880, w_055_881, w_055_882, w_055_883, w_055_884, w_055_886, w_055_888, w_055_894, w_055_895, w_055_897, w_055_901, w_055_902, w_055_903, w_055_905, w_055_906, w_055_908, w_055_909, w_055_910, w_055_912, w_055_913, w_055_915, w_055_916, w_055_917, w_055_918, w_055_921, w_055_922, w_055_923, w_055_924, w_055_925, w_055_927, w_055_928, w_055_930, w_055_935, w_055_937, w_055_938, w_055_942, w_055_943, w_055_945, w_055_946, w_055_948, w_055_950, w_055_952, w_055_955, w_055_959, w_055_961, w_055_963, w_055_967, w_055_970, w_055_971, w_055_972, w_055_979, w_055_980, w_055_988, w_055_989, w_055_990, w_055_993, w_055_994, w_055_996, w_055_998, w_055_999, w_055_1001, w_055_1002, w_055_1005, w_055_1006, w_055_1007, w_055_1009, w_055_1010, w_055_1012, w_055_1017, w_055_1018, w_055_1020, w_055_1022, w_055_1023, w_055_1024, w_055_1025, w_055_1027, w_055_1028, w_055_1032, w_055_1033, w_055_1036, w_055_1040, w_055_1043, w_055_1044, w_055_1045, w_055_1046, w_055_1047, w_055_1051, w_055_1054, w_055_1055, w_055_1057, w_055_1058, w_055_1060, w_055_1064, w_055_1065, w_055_1067, w_055_1069, w_055_1071, w_055_1073, w_055_1075, w_055_1080, w_055_1081, w_055_1082, w_055_1083, w_055_1084, w_055_1085, w_055_1087, w_055_1094, w_055_1095, w_055_1096, w_055_1100, w_055_1102, w_055_1108, w_055_1109, w_055_1111, w_055_1113, w_055_1117, w_055_1119, w_055_1121, w_055_1122, w_055_1123, w_055_1125, w_055_1126, w_055_1129, w_055_1132, w_055_1138, w_055_1140, w_055_1141, w_055_1146, w_055_1147, w_055_1148, w_055_1152, w_055_1153, w_055_1155, w_055_1157, w_055_1160, w_055_1163, w_055_1164, w_055_1165, w_055_1172, w_055_1173, w_055_1175, w_055_1178, w_055_1180, w_055_1181, w_055_1182, w_055_1186, w_055_1188, w_055_1189, w_055_1190, w_055_1195, w_055_1197, w_055_1202, w_055_1203, w_055_1205, w_055_1209, w_055_1211, w_055_1212, w_055_1213, w_055_1214, w_055_1215, w_055_1219, w_055_1222, w_055_1223, w_055_1225, w_055_1226, w_055_1229, w_055_1230, w_055_1232, w_055_1234, w_055_1238, w_055_1241, w_055_1242, w_055_1244, w_055_1249, w_055_1251, w_055_1256, w_055_1258, w_055_1260, w_055_1261, w_055_1262, w_055_1263, w_055_1266, w_055_1268, w_055_1269, w_055_1271, w_055_1272, w_055_1274, w_055_1275, w_055_1278, w_055_1279, w_055_1281, w_055_1282, w_055_1285, w_055_1287, w_055_1289, w_055_1290, w_055_1291, w_055_1293, w_055_1294, w_055_1296, w_055_1297, w_055_1298, w_055_1300, w_055_1301, w_055_1302, w_055_1305, w_055_1306, w_055_1307, w_055_1309, w_055_1311, w_055_1313, w_055_1314, w_055_1317, w_055_1318, w_055_1319, w_055_1322, w_055_1323, w_055_1326, w_055_1328, w_055_1330, w_055_1332, w_055_1335, w_055_1338, w_055_1339, w_055_1340, w_055_1343, w_055_1344, w_055_1346, w_055_1349, w_055_1350, w_055_1356, w_055_1358, w_055_1359, w_055_1360, w_055_1361, w_055_1363, w_055_1364, w_055_1367, w_055_1369, w_055_1370, w_055_1371, w_055_1375, w_055_1376, w_055_1378, w_055_1380, w_055_1384, w_055_1386, w_055_1392, w_055_1393, w_055_1394, w_055_1396, w_055_1397, w_055_1399, w_055_1404, w_055_1405, w_055_1412, w_055_1414, w_055_1415, w_055_1416, w_055_1417, w_055_1419, w_055_1425, w_055_1426, w_055_1427, w_055_1429, w_055_1430, w_055_1431, w_055_1432, w_055_1433, w_055_1435, w_055_1437, w_055_1441, w_055_1443, w_055_1444, w_055_1446, w_055_1447, w_055_1448, w_055_1449, w_055_1451, w_055_1452, w_055_1456, w_055_1457, w_055_1458, w_055_1460, w_055_1461, w_055_1464, w_055_1468, w_055_1472, w_055_1474, w_055_1476, w_055_1477, w_055_1478, w_055_1479, w_055_1480, w_055_1481, w_055_1485, w_055_1486, w_055_1488, w_055_1492, w_055_1493, w_055_1494, w_055_1497, w_055_1498, w_055_1501, w_055_1504, w_055_1505, w_055_1507, w_055_1508, w_055_1509, w_055_1510, w_055_1512, w_055_1515, w_055_1517, w_055_1518, w_055_1520, w_055_1525, w_055_1530, w_055_1532, w_055_1541, w_055_1545, w_055_1548, w_055_1550, w_055_1552, w_055_1557, w_055_1560, w_055_1562, w_055_1563, w_055_1564, w_055_1565, w_055_1567, w_055_1568, w_055_1570, w_055_1572, w_055_1573, w_055_1575, w_055_1578, w_055_1579, w_055_1581, w_055_1582, w_055_1583, w_055_1584, w_055_1585, w_055_1586, w_055_1587, w_055_1589, w_055_1591, w_055_1592, w_055_1595, w_055_1596, w_055_1597, w_055_1598, w_055_1603, w_055_1605, w_055_1609, w_055_1614, w_055_1615, w_055_1617, w_055_1618, w_055_1619, w_055_1622, w_055_1623, w_055_1624, w_055_1625, w_055_1626, w_055_1627, w_055_1631, w_055_1632, w_055_1633, w_055_1634, w_055_1636, w_055_1637, w_055_1638, w_055_1639, w_055_1640, w_055_1642, w_055_1648, w_055_1649, w_055_1650, w_055_1653, w_055_1658, w_055_1661, w_055_1665, w_055_1667, w_055_1668, w_055_1670, w_055_1675, w_055_1676, w_055_1680, w_055_1683, w_055_1685, w_055_1687, w_055_1689, w_055_1690, w_055_1692, w_055_1694, w_055_1695, w_055_1696, w_055_1697, w_055_1701, w_055_1703, w_055_1705, w_055_1707, w_055_1712, w_055_1714, w_055_1719, w_055_1720, w_055_1721, w_055_1722, w_055_1723, w_055_1725, w_055_1726, w_055_1729, w_055_1731, w_055_1734, w_055_1736, w_055_1740, w_055_1741, w_055_1747, w_055_1748, w_055_1749, w_055_1751, w_055_1754, w_055_1755, w_055_1759, w_055_1760, w_055_1762, w_055_1763, w_055_1764, w_055_1768, w_055_1769, w_055_1770, w_055_1771, w_055_1773, w_055_1774, w_055_1777, w_055_1778, w_055_1780, w_055_1781, w_055_1787, w_055_1789, w_055_1793, w_055_1799, w_055_1800, w_055_1801, w_055_1805, w_055_1806, w_055_1817, w_055_1818, w_055_1821, w_055_1832, w_055_1833, w_055_1834, w_055_1836, w_055_1837, w_055_1838, w_055_1839, w_055_1840, w_055_1841, w_055_1842, w_055_1844, w_055_1845, w_055_1850, w_055_1851, w_055_1854, w_055_1856, w_055_1861, w_055_1862, w_055_1865, w_055_1872, w_055_1873, w_055_1874, w_055_1879, w_055_1880, w_055_1881, w_055_1882, w_055_1883, w_055_1885, w_055_1886, w_055_1888, w_055_1893, w_055_1896, w_055_1897, w_055_1899, w_055_1900, w_055_1901, w_055_1903, w_055_1905, w_055_1906, w_055_1908, w_055_1913, w_055_1915, w_055_1918, w_055_1921, w_055_1923, w_055_1924, w_055_1925, w_055_1926, w_055_1928, w_055_1929, w_055_1930, w_055_1934, w_055_1943, w_055_1952, w_055_1953, w_055_1956, w_055_1957, w_055_1959, w_055_1962, w_055_1964, w_055_1968, w_055_1969, w_055_1970, w_055_1973, w_055_1975, w_055_1976, w_055_1984, w_055_1989, w_055_1991, w_055_1992, w_055_1999, w_055_2001, w_055_2002, w_055_2004, w_055_2009, w_055_2011, w_055_2013, w_055_2015, w_055_2021, w_055_2022, w_055_2025, w_055_2028, w_055_2029, w_055_2031, w_055_2033, w_055_2035, w_055_2038, w_055_2043, w_055_2045, w_055_2048, w_055_2049, w_055_2053, w_055_2054, w_055_2055, w_055_2057, w_055_2058, w_055_2059, w_055_2061, w_055_2063, w_055_2064, w_055_2068, w_055_2069, w_055_2070, w_055_2071, w_055_2072, w_055_2074, w_055_2076, w_055_2081, w_055_2083, w_055_2085, w_055_2087, w_055_2089, w_055_2092, w_055_2096, w_055_2097, w_055_2099, w_055_2100, w_055_2104, w_055_2106, w_055_2107, w_055_2110, w_055_2111, w_055_2112, w_055_2115, w_055_2116, w_055_2119, w_055_2124, w_055_2125, w_055_2128, w_055_2130, w_055_2133, w_055_2135, w_055_2136, w_055_2137, w_055_2139, w_055_2142, w_055_2143, w_055_2144, w_055_2146, w_055_2152, w_055_2153, w_055_2154, w_055_2156, w_055_2157, w_055_2158, w_055_2168, w_055_2175, w_055_2176, w_055_2177, w_055_2186, w_055_2188, w_055_2190, w_055_2191, w_055_2192, w_055_2194, w_055_2196, w_055_2197, w_055_2198, w_055_2202, w_055_2203, w_055_2207, w_055_2208, w_055_2209, w_055_2212, w_055_2213, w_055_2214, w_055_2215, w_055_2217, w_055_2220, w_055_2223, w_055_2224, w_055_2225, w_055_2226, w_055_2229, w_055_2230, w_055_2236, w_055_2238, w_055_2241, w_055_2246, w_055_2251, w_055_2262, w_055_2266, w_055_2267, w_055_2270, w_055_2272, w_055_2273, w_055_2274, w_055_2276, w_055_2277, w_055_2280, w_055_2281, w_055_2284, w_055_2286, w_055_2288, w_055_2291, w_055_2296, w_055_2297, w_055_2302, w_055_2304, w_055_2307, w_055_2309, w_055_2310, w_055_2312, w_055_2314, w_055_2315, w_055_2317, w_055_2318, w_055_2319, w_055_2320, w_055_2324, w_055_2327, w_055_2329, w_055_2331, w_055_2333, w_055_2336, w_055_2342, w_055_2343, w_055_2344, w_055_2346, w_055_2352, w_055_2353, w_055_2354, w_055_2356, w_055_2358, w_055_2360, w_055_2362, w_055_2363, w_055_2365, w_055_2366, w_055_2367, w_055_2370, w_055_2373, w_055_2375, w_055_2376, w_055_2378, w_055_2382, w_055_2384, w_055_2385, w_055_2388, w_055_2389, w_055_2394, w_055_2395, w_055_2397, w_055_2398, w_055_2401, w_055_2406, w_055_2407, w_055_2410, w_055_2411, w_055_2413, w_055_2414, w_055_2415, w_055_2416, w_055_2417, w_055_2420, w_055_2422, w_055_2424, w_055_2427, w_055_2433, w_055_2434, w_055_2435, w_055_2436, w_055_2438, w_055_2442, w_055_2443, w_055_2444, w_055_2447, w_055_2448, w_055_2451, w_055_2455, w_055_2458, w_055_2459, w_055_2465, w_055_2467, w_055_2469, w_055_2470, w_055_2472, w_055_2474, w_055_2478, w_055_2480, w_055_2481, w_055_2482, w_055_2484, w_055_2485, w_055_2487, w_055_2489, w_055_2492, w_055_2494, w_055_2495, w_055_2496, w_055_2501, w_055_2502, w_055_2506, w_055_2509, w_055_2512, w_055_2513, w_055_2514, w_055_2517, w_055_2523, w_055_2525, w_055_2526, w_055_2529, w_055_2530, w_055_2533, w_055_2535, w_055_2539, w_055_2540, w_055_2541, w_055_2546, w_055_2552, w_055_2553, w_055_2554, w_055_2556, w_055_2558, w_055_2559, w_055_2563, w_055_2567, w_055_2569, w_055_2572, w_055_2574, w_055_2575, w_055_2576, w_055_2577, w_055_2578, w_055_2580, w_055_2581, w_055_2584, w_055_2585, w_055_2588, w_055_2590, w_055_2595, w_055_2597, w_055_2599, w_055_2601, w_055_2605, w_055_2606, w_055_2608, w_055_2609, w_055_2615, w_055_2617, w_055_2622, w_055_2624, w_055_2630, w_055_2631, w_055_2633, w_055_2635, w_055_2636, w_055_2637, w_055_2645, w_055_2646, w_055_2650, w_055_2651, w_055_2654, w_055_2655, w_055_2656, w_055_2657, w_055_2667, w_055_2669, w_055_2672, w_055_2674, w_055_2675, w_055_2681, w_055_2682, w_055_2688, w_055_2695, w_055_2697, w_055_2702, w_055_2704, w_055_2708, w_055_2709, w_055_2710, w_055_2712, w_055_2713, w_055_2715, w_055_2716, w_055_2721, w_055_2728, w_055_2730, w_055_2731, w_055_2733, w_055_2735, w_055_2737, w_055_2739, w_055_2744, w_055_2746, w_055_2751, w_055_2752, w_055_2758, w_055_2759, w_055_2761, w_055_2763, w_055_2764, w_055_2765, w_055_2772, w_055_2774, w_055_2776, w_055_2778, w_055_2781, w_055_2784, w_055_2787, w_055_2788, w_055_2790, w_055_2791, w_055_2793, w_055_2794, w_055_2798, w_055_2801, w_055_2802, w_055_2803, w_055_2804, w_055_2805, w_055_2806, w_055_2807, w_055_2809, w_055_2810, w_055_2811, w_055_2814, w_055_2815, w_055_2821, w_055_2823, w_055_2826, w_055_2830, w_055_2831, w_055_2832, w_055_2834, w_055_2838, w_055_2844, w_055_2849, w_055_2852, w_055_2853, w_055_2856, w_055_2861, w_055_2862, w_055_2863, w_055_2864, w_055_2865, w_055_2871, w_055_2872, w_055_2877, w_055_2878, w_055_2879, w_055_2881, w_055_2882, w_055_2885, w_055_2886, w_055_2894, w_055_2896, w_055_2897, w_055_2899, w_055_2900, w_055_2903, w_055_2905, w_055_2906, w_055_2907, w_055_2909, w_055_2912, w_055_2915, w_055_2916, w_055_2918, w_055_2920, w_055_2921, w_055_2923, w_055_2926, w_055_2927, w_055_2929, w_055_2932, w_055_2933, w_055_2939, w_055_2942, w_055_2943, w_055_2944, w_055_2949, w_055_2950, w_055_2951, w_055_2953, w_055_2956, w_055_2958, w_055_2959, w_055_2960, w_055_2964, w_055_2966, w_055_2967, w_055_2968, w_055_2970, w_055_2975, w_055_2978, w_055_2980, w_055_2986, w_055_2989, w_055_2992, w_055_2993, w_055_2994, w_055_2996, w_055_3000, w_055_3002, w_055_3003, w_055_3008, w_055_3011, w_055_3019, w_055_3022, w_055_3023, w_055_3024, w_055_3027, w_055_3034, w_055_3037, w_055_3038, w_055_3043, w_055_3047, w_055_3049, w_055_3050, w_055_3052, w_055_3058, w_055_3061, w_055_3062, w_055_3069, w_055_3072, w_055_3074, w_055_3076, w_055_3077, w_055_3079, w_055_3081, w_055_3084, w_055_3088, w_055_3089, w_055_3093, w_055_3094, w_055_3096, w_055_3097, w_055_3101, w_055_3102, w_055_3103, w_055_3105, w_055_3106, w_055_3112, w_055_3113, w_055_3116, w_055_3117, w_055_3118, w_055_3121, w_055_3122, w_055_3124, w_055_3127, w_055_3130, w_055_3131, w_055_3134, w_055_3137, w_055_3138, w_055_3144, w_055_3149, w_055_3154, w_055_3155, w_055_3158, w_055_3159, w_055_3160, w_055_3161, w_055_3162, w_055_3165, w_055_3174, w_055_3181, w_055_3183, w_055_3185, w_055_3191, w_055_3194, w_055_3196, w_055_3203, w_055_3206, w_055_3207, w_055_3208, w_055_3209, w_055_3210, w_055_3212, w_055_3213, w_055_3214, w_055_3219, w_055_3221, w_055_3223, w_055_3225, w_055_3227, w_055_3228, w_055_3230, w_055_3231, w_055_3238, w_055_3239, w_055_3242, w_055_3243, w_055_3244, w_055_3245, w_055_3247, w_055_3248, w_055_3250, w_055_3255, w_055_3259, w_055_3261, w_055_3262, w_055_3266, w_055_3267, w_055_3269, w_055_3272, w_055_3276, w_055_3280, w_055_3283, w_055_3284, w_055_3285, w_055_3286, w_055_3288, w_055_3292, w_055_3293, w_055_3295, w_055_3299, w_055_3302, w_055_3303, w_055_3305, w_055_3309, w_055_3311, w_055_3316, w_055_3318, w_055_3319, w_055_3322, w_055_3324, w_055_3325, w_055_3332, w_055_3333, w_055_3335, w_055_3337, w_055_3339, w_055_3340, w_055_3343, w_055_3346, w_055_3347, w_055_3349, w_055_3352, w_055_3354, w_055_3355, w_055_3356, w_055_3357, w_055_3358, w_055_3360, w_055_3362, w_055_3363, w_055_3364, w_055_3366, w_055_3368, w_055_3369, w_055_3376, w_055_3385, w_055_3387, w_055_3389, w_055_3391, w_055_3393, w_055_3394, w_055_3395, w_055_3399, w_055_3401, w_055_3404, w_055_3405, w_055_3408, w_055_3409, w_055_3410, w_055_3412, w_055_3413, w_055_3415, w_055_3417, w_055_3418, w_055_3419, w_055_3422, w_055_3423, w_055_3426, w_055_3427, w_055_3428, w_055_3430, w_055_3433, w_055_3435, w_055_3437, w_055_3438, w_055_3439, w_055_3440, w_055_3445, w_055_3446, w_055_3448, w_055_3450, w_055_3451, w_055_3452, w_055_3454, w_055_3456, w_055_3457, w_055_3458, w_055_3459, w_055_3461, w_055_3463, w_055_3464, w_055_3466, w_055_3467, w_055_3470, w_055_3471, w_055_3475, w_055_3476, w_055_3478, w_055_3479, w_055_3480, w_055_3482, w_055_3484, w_055_3485, w_055_3486, w_055_3487, w_055_3488, w_055_3489, w_055_3497, w_055_3498, w_055_3501, w_055_3502, w_055_3504, w_055_3508, w_055_3509, w_055_3515, w_055_3517, w_055_3520, w_055_3521, w_055_3522, w_055_3523, w_055_3525, w_055_3529, w_055_3530, w_055_3534, w_055_3536, w_055_3541, w_055_3544, w_055_3545, w_055_3551, w_055_3552, w_055_3554, w_055_3555, w_055_3558, w_055_3560, w_055_3563, w_055_3566, w_055_3571, w_055_3572, w_055_3573, w_055_3581, w_055_3583, w_055_3584, w_055_3588, w_055_3593, w_055_3594, w_055_3596, w_055_3598, w_055_3599, w_055_3600, w_055_3602, w_055_3603, w_055_3611, w_055_3614, w_055_3619, w_055_3621, w_055_3624, w_055_3626, w_055_3631, w_055_3634, w_055_3635, w_055_3636, w_055_3641, w_055_3649, w_055_3657, w_055_3659, w_055_3660, w_055_3663, w_055_3665, w_055_3669, w_055_3670, w_055_3671, w_055_3675, w_055_3677, w_055_3679, w_055_3682, w_055_3684, w_055_3685, w_055_3689, w_055_3690, w_055_3694, w_055_3700, w_055_3701, w_055_3704, w_055_3707, w_055_3710, w_055_3711, w_055_3717, w_055_3718, w_055_3720, w_055_3722, w_055_3724, w_055_3725, w_055_3726, w_055_3727, w_055_3729, w_055_3730, w_055_3732, w_055_3733, w_055_3734, w_055_3735, w_055_3739, w_055_3741, w_055_3746, w_055_3748, w_055_3749, w_055_3754, w_055_3760, w_055_3768, w_055_3769, w_055_3775, w_055_3776, w_055_3778, w_055_3779, w_055_3784, w_055_3785, w_055_3786, w_055_3787, w_055_3788, w_055_3790, w_055_3791, w_055_3792, w_055_3793, w_055_3795, w_055_3798, w_055_3799, w_055_3800, w_055_3801, w_055_3806, w_055_3807, w_055_3809, w_055_3810, w_055_3811, w_055_3812, w_055_3813, w_055_3814, w_055_3818, w_055_3819, w_055_3826, w_055_3827, w_055_3832, w_055_3835, w_055_3837, w_055_3839, w_055_3840, w_055_3845, w_055_3847, w_055_3848, w_055_3851, w_055_3855, w_055_3860, w_055_3863, w_055_3865, w_055_3866, w_055_3868, w_055_3873, w_055_3874, w_055_3875, w_055_3879, w_055_3880, w_055_3884, w_055_3886, w_055_3892, w_055_3893, w_055_3894, w_055_3896, w_055_3897, w_055_3898, w_055_3899, w_055_3900, w_055_3901, w_055_3902, w_055_3903, w_055_3904, w_055_3905, w_055_3906, w_055_3910, w_055_3913, w_055_3918, w_055_3920, w_055_3921, w_055_3922, w_055_3924, w_055_3926, w_055_3928, w_055_3929, w_055_3936, w_055_3938, w_055_3939, w_055_3940, w_055_3943, w_055_3946, w_055_3947, w_055_3948, w_055_3949, w_055_3951, w_055_3952, w_055_3954, w_055_3955, w_055_3956, w_055_3959, w_055_3960, w_055_3963, w_055_3964, w_055_3966, w_055_3972, w_055_3973, w_055_3976, w_055_3977, w_055_3978, w_055_3982, w_055_3983, w_055_3984, w_055_3986, w_055_3989, w_055_3991, w_055_3993, w_055_3994, w_055_3996, w_055_3997, w_055_3998, w_055_3999, w_055_4000, w_055_4005, w_055_4007, w_055_4008, w_055_4009, w_055_4010, w_055_4011, w_055_4012, w_055_4017, w_055_4018, w_055_4021, w_055_4022, w_055_4023, w_055_4026, w_055_4028, w_055_4035, w_055_4038, w_055_4040, w_055_4042, w_055_4044, w_055_4046, w_055_4051, w_055_4056, w_055_4057, w_055_4059, w_055_4060, w_055_4061, w_055_4062, w_055_4065, w_055_4067, w_055_4068, w_055_4075, w_055_4078, w_055_4080;
  wire w_056_000, w_056_001, w_056_002, w_056_003, w_056_004, w_056_006, w_056_008, w_056_011, w_056_012, w_056_013, w_056_014, w_056_015, w_056_016, w_056_018, w_056_019, w_056_020, w_056_021, w_056_023, w_056_025, w_056_027, w_056_029, w_056_031, w_056_032, w_056_033, w_056_034, w_056_035, w_056_036, w_056_037, w_056_038, w_056_039, w_056_041, w_056_042, w_056_046, w_056_047, w_056_049, w_056_050, w_056_051, w_056_053, w_056_054, w_056_056, w_056_060, w_056_061, w_056_062, w_056_063, w_056_066, w_056_070, w_056_072, w_056_073, w_056_074, w_056_075, w_056_076, w_056_077, w_056_078, w_056_079, w_056_080, w_056_082, w_056_085, w_056_086, w_056_087, w_056_088, w_056_090, w_056_091, w_056_093, w_056_094, w_056_095, w_056_096, w_056_097, w_056_098, w_056_099, w_056_100, w_056_101, w_056_104, w_056_105, w_056_106, w_056_107, w_056_108, w_056_109, w_056_110, w_056_111, w_056_113, w_056_116, w_056_118, w_056_119, w_056_120, w_056_121, w_056_123, w_056_124, w_056_126, w_056_127, w_056_128, w_056_129, w_056_130, w_056_134, w_056_135, w_056_136, w_056_137, w_056_138, w_056_139, w_056_142, w_056_143, w_056_145, w_056_146, w_056_147, w_056_148, w_056_149, w_056_150, w_056_152, w_056_153, w_056_157, w_056_159, w_056_162, w_056_163, w_056_164, w_056_166, w_056_168, w_056_170, w_056_171, w_056_173, w_056_174, w_056_175, w_056_176, w_056_178, w_056_179, w_056_181, w_056_182, w_056_184, w_056_185, w_056_187, w_056_188, w_056_189, w_056_191, w_056_192, w_056_193, w_056_194, w_056_196, w_056_197, w_056_200, w_056_201, w_056_202, w_056_203, w_056_205, w_056_206, w_056_207, w_056_208, w_056_209, w_056_210, w_056_212, w_056_213, w_056_215, w_056_218, w_056_222, w_056_225, w_056_226, w_056_228, w_056_229, w_056_231, w_056_233, w_056_235, w_056_236, w_056_239, w_056_240, w_056_241, w_056_242, w_056_243, w_056_244, w_056_245, w_056_246, w_056_247, w_056_249, w_056_251, w_056_252, w_056_254, w_056_257, w_056_258, w_056_260, w_056_261, w_056_262, w_056_263, w_056_265, w_056_266, w_056_267, w_056_268, w_056_269, w_056_270, w_056_271, w_056_272, w_056_273, w_056_274, w_056_275, w_056_277, w_056_279, w_056_280, w_056_282, w_056_284, w_056_285, w_056_286, w_056_290, w_056_291, w_056_292, w_056_293, w_056_294, w_056_295, w_056_297, w_056_298, w_056_299, w_056_300, w_056_301, w_056_302, w_056_303, w_056_304, w_056_305, w_056_306, w_056_308, w_056_309, w_056_314, w_056_318, w_056_319, w_056_320, w_056_322, w_056_324, w_056_326, w_056_327, w_056_328, w_056_329, w_056_331, w_056_332, w_056_333, w_056_334, w_056_335, w_056_336, w_056_337, w_056_338, w_056_339, w_056_340, w_056_341, w_056_342, w_056_344, w_056_347, w_056_348, w_056_349, w_056_350, w_056_353, w_056_354, w_056_355, w_056_356, w_056_357, w_056_359, w_056_360, w_056_361, w_056_364, w_056_365, w_056_367, w_056_368, w_056_371, w_056_373, w_056_374, w_056_376, w_056_377, w_056_379, w_056_380, w_056_381, w_056_385, w_056_386, w_056_389, w_056_391, w_056_394, w_056_395, w_056_396, w_056_398, w_056_399, w_056_403, w_056_404, w_056_405, w_056_406, w_056_408, w_056_409, w_056_410, w_056_412, w_056_414, w_056_416, w_056_417, w_056_418, w_056_419, w_056_420, w_056_421, w_056_422, w_056_424, w_056_425, w_056_428, w_056_431, w_056_433, w_056_434, w_056_435, w_056_437, w_056_438, w_056_439, w_056_441, w_056_442, w_056_443, w_056_445, w_056_446, w_056_447, w_056_448, w_056_449, w_056_450, w_056_451, w_056_452, w_056_454, w_056_455, w_056_457, w_056_459, w_056_460, w_056_461, w_056_462, w_056_463, w_056_465, w_056_468, w_056_469, w_056_470, w_056_471, w_056_472, w_056_473, w_056_474, w_056_475, w_056_477, w_056_478, w_056_479, w_056_480, w_056_483, w_056_484, w_056_487, w_056_488, w_056_489, w_056_490, w_056_491, w_056_493, w_056_494, w_056_495, w_056_496, w_056_497, w_056_498, w_056_499, w_056_501, w_056_503, w_056_504, w_056_505, w_056_506, w_056_507, w_056_510, w_056_514, w_056_515, w_056_516, w_056_519, w_056_520, w_056_522, w_056_523, w_056_524, w_056_526, w_056_527, w_056_528, w_056_529, w_056_530, w_056_531, w_056_533, w_056_535, w_056_537, w_056_538, w_056_540, w_056_541, w_056_543, w_056_544, w_056_545, w_056_547, w_056_548, w_056_549, w_056_551, w_056_552, w_056_553, w_056_555, w_056_557, w_056_558, w_056_559, w_056_560, w_056_561, w_056_562, w_056_563, w_056_564, w_056_566, w_056_569, w_056_571, w_056_573, w_056_574, w_056_575, w_056_576, w_056_578, w_056_580, w_056_582, w_056_583, w_056_584, w_056_585, w_056_586, w_056_587, w_056_588, w_056_589, w_056_590, w_056_592, w_056_593, w_056_594, w_056_596, w_056_600, w_056_601, w_056_602, w_056_603, w_056_604, w_056_605, w_056_606, w_056_608, w_056_609, w_056_610, w_056_611, w_056_612, w_056_613, w_056_614, w_056_616, w_056_620, w_056_621, w_056_622, w_056_623, w_056_624, w_056_625, w_056_628, w_056_629, w_056_630, w_056_631, w_056_633, w_056_635, w_056_636, w_056_637, w_056_639, w_056_640, w_056_641, w_056_642, w_056_643, w_056_644, w_056_645, w_056_646, w_056_648, w_056_649, w_056_653, w_056_654, w_056_655, w_056_656, w_056_658, w_056_660, w_056_661, w_056_662, w_056_664, w_056_665, w_056_666, w_056_667, w_056_668, w_056_670, w_056_671, w_056_672, w_056_675, w_056_676, w_056_677, w_056_680, w_056_682, w_056_684, w_056_686, w_056_687, w_056_688, w_056_690, w_056_691, w_056_692, w_056_693, w_056_697, w_056_698, w_056_699, w_056_700, w_056_701, w_056_703, w_056_704, w_056_705, w_056_708, w_056_710, w_056_711, w_056_713, w_056_714, w_056_715, w_056_716, w_056_718, w_056_719, w_056_720, w_056_722, w_056_727, w_056_728, w_056_729, w_056_731, w_056_733, w_056_735, w_056_737, w_056_738, w_056_739, w_056_741, w_056_742, w_056_743, w_056_745, w_056_746, w_056_747, w_056_749, w_056_750, w_056_753, w_056_754, w_056_755, w_056_756, w_056_757, w_056_758, w_056_759, w_056_760, w_056_761, w_056_764, w_056_765, w_056_766, w_056_767, w_056_768, w_056_769, w_056_770, w_056_773, w_056_776, w_056_777, w_056_778, w_056_779, w_056_780, w_056_781, w_056_782, w_056_783, w_056_784, w_056_785, w_056_786, w_056_787, w_056_788, w_056_789, w_056_790, w_056_791, w_056_793, w_056_795, w_056_797, w_056_798, w_056_799, w_056_801, w_056_803, w_056_806, w_056_809, w_056_811, w_056_812, w_056_814, w_056_816, w_056_818, w_056_823, w_056_824, w_056_825, w_056_826, w_056_827, w_056_828, w_056_830, w_056_831, w_056_832, w_056_833, w_056_835, w_056_836, w_056_837, w_056_838, w_056_839, w_056_841, w_056_842, w_056_843, w_056_846, w_056_847, w_056_848, w_056_849, w_056_853, w_056_854, w_056_855, w_056_857, w_056_859, w_056_860, w_056_861, w_056_863, w_056_864, w_056_870, w_056_871, w_056_873, w_056_874, w_056_875, w_056_876, w_056_878, w_056_879, w_056_880, w_056_881, w_056_884, w_056_885, w_056_888, w_056_890, w_056_892, w_056_895, w_056_897, w_056_898, w_056_899, w_056_900, w_056_901, w_056_904, w_056_905, w_056_907, w_056_908, w_056_910, w_056_911, w_056_913, w_056_914, w_056_915, w_056_917, w_056_918, w_056_919, w_056_920, w_056_921, w_056_923, w_056_924, w_056_925, w_056_926, w_056_927, w_056_928, w_056_929, w_056_931, w_056_932, w_056_935, w_056_937, w_056_938, w_056_940, w_056_941, w_056_942, w_056_944, w_056_945, w_056_946, w_056_947, w_056_948, w_056_949, w_056_950, w_056_952, w_056_953, w_056_954, w_056_955, w_056_956, w_056_959, w_056_960, w_056_962, w_056_963, w_056_966, w_056_967, w_056_968, w_056_969, w_056_971, w_056_972, w_056_974, w_056_975, w_056_976, w_056_977, w_056_979, w_056_980, w_056_981, w_056_982, w_056_983, w_056_984, w_056_985, w_056_986, w_056_987, w_056_988, w_056_990, w_056_991, w_056_992, w_056_993, w_056_994, w_056_995, w_056_996, w_056_997, w_056_998, w_056_999, w_056_1001, w_056_1004, w_056_1005, w_056_1006, w_056_1007, w_056_1008, w_056_1010, w_056_1011, w_056_1012, w_056_1014, w_056_1015, w_056_1016, w_056_1017, w_056_1019, w_056_1023, w_056_1024, w_056_1026, w_056_1027, w_056_1028, w_056_1031, w_056_1032, w_056_1033, w_056_1035, w_056_1036, w_056_1037, w_056_1038, w_056_1039, w_056_1040, w_056_1041, w_056_1042, w_056_1043, w_056_1045, w_056_1046, w_056_1047, w_056_1049, w_056_1051, w_056_1052, w_056_1053, w_056_1054, w_056_1055, w_056_1057, w_056_1058, w_056_1060, w_056_1061, w_056_1062, w_056_1063, w_056_1064, w_056_1066, w_056_1067, w_056_1068, w_056_1069, w_056_1070, w_056_1072, w_056_1074, w_056_1075, w_056_1076, w_056_1077, w_056_1078, w_056_1079, w_056_1082, w_056_1083, w_056_1084, w_056_1085, w_056_1086, w_056_1090, w_056_1091, w_056_1093, w_056_1094, w_056_1095, w_056_1097, w_056_1098, w_056_1100, w_056_1101, w_056_1102, w_056_1103, w_056_1104, w_056_1106, w_056_1108, w_056_1109, w_056_1111, w_056_1112, w_056_1113, w_056_1114, w_056_1115, w_056_1116, w_056_1117, w_056_1119, w_056_1120, w_056_1121, w_056_1123, w_056_1124, w_056_1125, w_056_1127, w_056_1129, w_056_1132, w_056_1133, w_056_1134, w_056_1135, w_056_1137, w_056_1140, w_056_1142, w_056_1143, w_056_1144, w_056_1145, w_056_1146, w_056_1147, w_056_1150, w_056_1152, w_056_1155, w_056_1157, w_056_1158, w_056_1160, w_056_1162, w_056_1164, w_056_1165, w_056_1166, w_056_1167, w_056_1170, w_056_1171, w_056_1172, w_056_1173, w_056_1174, w_056_1176, w_056_1180, w_056_1181, w_056_1182, w_056_1184, w_056_1186, w_056_1188, w_056_1189, w_056_1191, w_056_1195, w_056_1196, w_056_1198, w_056_1199, w_056_1201, w_056_1202, w_056_1204, w_056_1206, w_056_1208, w_056_1209, w_056_1210, w_056_1211, w_056_1212, w_056_1214, w_056_1215, w_056_1217, w_056_1219, w_056_1220, w_056_1221, w_056_1222, w_056_1224, w_056_1226, w_056_1232, w_056_1234, w_056_1235, w_056_1236, w_056_1237, w_056_1239, w_056_1241, w_056_1242, w_056_1243, w_056_1245, w_056_1246, w_056_1247, w_056_1248, w_056_1249, w_056_1250, w_056_1253, w_056_1254, w_056_1255, w_056_1258, w_056_1259, w_056_1262, w_056_1263, w_056_1264, w_056_1266, w_056_1267, w_056_1268, w_056_1269, w_056_1270, w_056_1271, w_056_1272, w_056_1273, w_056_1274, w_056_1276, w_056_1278, w_056_1279, w_056_1281, w_056_1282, w_056_1283, w_056_1284, w_056_1286, w_056_1288, w_056_1290, w_056_1293, w_056_1295, w_056_1297, w_056_1298, w_056_1299, w_056_1300, w_056_1301, w_056_1302, w_056_1304, w_056_1305, w_056_1306, w_056_1308, w_056_1310, w_056_1311, w_056_1312, w_056_1313, w_056_1314, w_056_1315, w_056_1316, w_056_1318, w_056_1319, w_056_1321, w_056_1322, w_056_1324, w_056_1326, w_056_1327, w_056_1329, w_056_1330, w_056_1331, w_056_1332, w_056_1333, w_056_1335, w_056_1337, w_056_1338, w_056_1339, w_056_1342, w_056_1343, w_056_1344, w_056_1346, w_056_1348, w_056_1349, w_056_1353, w_056_1354, w_056_1355, w_056_1356, w_056_1357, w_056_1360, w_056_1362, w_056_1363, w_056_1365, w_056_1368, w_056_1369, w_056_1370, w_056_1371, w_056_1373, w_056_1374, w_056_1375, w_056_1376, w_056_1378, w_056_1379, w_056_1380, w_056_1382, w_056_1383, w_056_1384, w_056_1387, w_056_1388, w_056_1389, w_056_1390, w_056_1392, w_056_1394, w_056_1396, w_056_1397, w_056_1398, w_056_1399, w_056_1400, w_056_1402, w_056_1405, w_056_1406, w_056_1407, w_056_1408, w_056_1409, w_056_1410, w_056_1411, w_056_1412, w_056_1413, w_056_1414, w_056_1415, w_056_1416, w_056_1419, w_056_1420, w_056_1422, w_056_1423, w_056_1424, w_056_1425, w_056_1426, w_056_1427, w_056_1430, w_056_1431, w_056_1433, w_056_1434, w_056_1435, w_056_1437, w_056_1438, w_056_1439, w_056_1440, w_056_1443, w_056_1444, w_056_1446, w_056_1448, w_056_1451, w_056_1452, w_056_1454, w_056_1456, w_056_1457, w_056_1458, w_056_1460, w_056_1461, w_056_1462, w_056_1463, w_056_1465, w_056_1466, w_056_1467, w_056_1469, w_056_1470, w_056_1471, w_056_1472, w_056_1473, w_056_1474, w_056_1476, w_056_1477, w_056_1478, w_056_1479, w_056_1480, w_056_1482, w_056_1484, w_056_1485, w_056_1486, w_056_1487, w_056_1488, w_056_1489, w_056_1490, w_056_1491, w_056_1492, w_056_1493, w_056_1494, w_056_1497, w_056_1501, w_056_1502, w_056_1503, w_056_1505, w_056_1507, w_056_1508, w_056_1509, w_056_1510, w_056_1511, w_056_1512, w_056_1514, w_056_1516, w_056_1517, w_056_1518, w_056_1522, w_056_1523, w_056_1524, w_056_1525, w_056_1526, w_056_1527, w_056_1528, w_056_1529, w_056_1531, w_056_1532, w_056_1533, w_056_1534, w_056_1535, w_056_1539, w_056_1540, w_056_1541, w_056_1543, w_056_1544, w_056_1547, w_056_1548, w_056_1549, w_056_1550, w_056_1553, w_056_1554, w_056_1556, w_056_1559, w_056_1562, w_056_1564, w_056_1565, w_056_1566, w_056_1568, w_056_1569, w_056_1570, w_056_1571, w_056_1575, w_056_1577, w_056_1580, w_056_1581, w_056_1584, w_056_1585, w_056_1586, w_056_1591, w_056_1595, w_056_1596, w_056_1597, w_056_1599, w_056_1600, w_056_1601, w_056_1602, w_056_1603, w_056_1605, w_056_1606, w_056_1607, w_056_1608, w_056_1609, w_056_1610, w_056_1611, w_056_1612, w_056_1613, w_056_1615, w_056_1617, w_056_1618, w_056_1619, w_056_1620, w_056_1621, w_056_1622, w_056_1623, w_056_1624, w_056_1626, w_056_1627, w_056_1628, w_056_1629, w_056_1632, w_056_1634, w_056_1635, w_056_1636, w_056_1638, w_056_1639, w_056_1642, w_056_1643, w_056_1645, w_056_1646, w_056_1647, w_056_1648, w_056_1649, w_056_1651, w_056_1652, w_056_1654, w_056_1656, w_056_1657, w_056_1658, w_056_1660, w_056_1663, w_056_1665, w_056_1667, w_056_1669, w_056_1670, w_056_1671, w_056_1672, w_056_1673, w_056_1674, w_056_1675, w_056_1676, w_056_1677, w_056_1681, w_056_1682, w_056_1683, w_056_1684, w_056_1685, w_056_1686, w_056_1687, w_056_1688, w_056_1689, w_056_1691, w_056_1692, w_056_1693, w_056_1694, w_056_1695, w_056_1697, w_056_1698, w_056_1699, w_056_1701, w_056_1702, w_056_1703, w_056_1705, w_056_1707, w_056_1708, w_056_1710, w_056_1711, w_056_1712, w_056_1713, w_056_1714, w_056_1716, w_056_1717, w_056_1718, w_056_1719, w_056_1720, w_056_1722, w_056_1724, w_056_1725, w_056_1726, w_056_1727, w_056_1728, w_056_1730, w_056_1731, w_056_1732, w_056_1735, w_056_1736, w_056_1737, w_056_1739, w_056_1740, w_056_1741, w_056_1744, w_056_1746, w_056_1747, w_056_1748, w_056_1749, w_056_1750, w_056_1753, w_056_1754, w_056_1755, w_056_1756, w_056_1757, w_056_1758, w_056_1759, w_056_1760, w_056_1761, w_056_1763, w_056_1764, w_056_1766, w_056_1767, w_056_1769, w_056_1771, w_056_1772, w_056_1773, w_056_1775, w_056_1777, w_056_1778, w_056_1779, w_056_1780, w_056_1783, w_056_1784, w_056_1785, w_056_1786, w_056_1787, w_056_1788, w_056_1789, w_056_1791, w_056_1793, w_056_1794, w_056_1795, w_056_1796, w_056_1797, w_056_1798, w_056_1799, w_056_1800, w_056_1801, w_056_1803, w_056_1805, w_056_1808, w_056_1811, w_056_1812, w_056_1813, w_056_1814, w_056_1815, w_056_1816, w_056_1818, w_056_1819, w_056_1822, w_056_1823, w_056_1826, w_056_1828, w_056_1829, w_056_1830, w_056_1833, w_056_1835, w_056_1837, w_056_1838, w_056_1839, w_056_1840, w_056_1842, w_056_1843, w_056_1849, w_056_1850, w_056_1851, w_056_1852, w_056_1853, w_056_1856, w_056_1858, w_056_1862, w_056_1863, w_056_1864, w_056_1865, w_056_1867, w_056_1868, w_056_1869, w_056_1870, w_056_1871, w_056_1873, w_056_1874, w_056_1875, w_056_1876, w_056_1879, w_056_1882, w_056_1885, w_056_1887, w_056_1888, w_056_1890, w_056_1891, w_056_1894, w_056_1895, w_056_1896, w_056_1897, w_056_1899, w_056_1900, w_056_1901, w_056_1902, w_056_1905, w_056_1906, w_056_1907, w_056_1908, w_056_1911, w_056_1912, w_056_1913, w_056_1916, w_056_1918, w_056_1920, w_056_1921, w_056_1923, w_056_1924, w_056_1925, w_056_1926, w_056_1927, w_056_1929, w_056_1930, w_056_1931, w_056_1932, w_056_1934, w_056_1935, w_056_1936, w_056_1938, w_056_1939, w_056_1940, w_056_1941, w_056_1943, w_056_1944, w_056_1945, w_056_1947, w_056_1948, w_056_1950, w_056_1951, w_056_1953, w_056_1954, w_056_1955, w_056_1956, w_056_1957, w_056_1958, w_056_1959, w_056_1960, w_056_1962, w_056_1964, w_056_1966, w_056_1967, w_056_1968, w_056_1969, w_056_1970, w_056_1973, w_056_1974, w_056_1976, w_056_1977, w_056_1978, w_056_1979, w_056_1980, w_056_1981, w_056_1982, w_056_1984, w_056_1985, w_056_1987, w_056_1988, w_056_1991, w_056_1992, w_056_1994, w_056_1995, w_056_1997, w_056_1998, w_056_1999, w_056_2000, w_056_2002, w_056_2004, w_056_2006, w_056_2007, w_056_2008, w_056_2009, w_056_2011, w_056_2012, w_056_2014, w_056_2015, w_056_2016, w_056_2017, w_056_2018, w_056_2020, w_056_2023, w_056_2024, w_056_2027, w_056_2028, w_056_2029, w_056_2031, w_056_2032, w_056_2033, w_056_2035, w_056_2036, w_056_2038, w_056_2040, w_056_2041, w_056_2043, w_056_2044, w_056_2045, w_056_2046, w_056_2047, w_056_2049, w_056_2051, w_056_2052, w_056_2053, w_056_2054, w_056_2055, w_056_2056, w_056_2058, w_056_2059, w_056_2060, w_056_2061, w_056_2062, w_056_2064, w_056_2065, w_056_2066, w_056_2067, w_056_2068, w_056_2069, w_056_2070, w_056_2071, w_056_2072, w_056_2075, w_056_2076, w_056_2078, w_056_2079, w_056_2081, w_056_2082, w_056_2083, w_056_2085, w_056_2087, w_056_2088, w_056_2089, w_056_2090, w_056_2091, w_056_2092, w_056_2094, w_056_2098, w_056_2099, w_056_2100, w_056_2101, w_056_2102, w_056_2103, w_056_2105, w_056_2106, w_056_2107, w_056_2110, w_056_2112, w_056_2113, w_056_2114, w_056_2115, w_056_2116, w_056_2117, w_056_2118, w_056_2120, w_056_2121, w_056_2122, w_056_2124, w_056_2125, w_056_2127, w_056_2128, w_056_2129, w_056_2130, w_056_2134, w_056_2135, w_056_2136, w_056_2137, w_056_2138, w_056_2139, w_056_2141, w_056_2142, w_056_2143, w_056_2144, w_056_2147, w_056_2148, w_056_2149, w_056_2150, w_056_2152, w_056_2154, w_056_2155, w_056_2156, w_056_2157, w_056_2158, w_056_2159, w_056_2160, w_056_2161, w_056_2164, w_056_2167, w_056_2168, w_056_2170, w_056_2172, w_056_2173, w_056_2174, w_056_2175, w_056_2180, w_056_2182, w_056_2184, w_056_2185, w_056_2186, w_056_2188, w_056_2191, w_056_2193, w_056_2195, w_056_2196, w_056_2199, w_056_2201, w_056_2202, w_056_2203, w_056_2204, w_056_2206, w_056_2207, w_056_2209, w_056_2212, w_056_2213, w_056_2214, w_056_2219, w_056_2220, w_056_2221, w_056_2222, w_056_2223, w_056_2224, w_056_2228, w_056_2229, w_056_2230, w_056_2231, w_056_2232, w_056_2233, w_056_2234, w_056_2236, w_056_2237, w_056_2238, w_056_2239, w_056_2240, w_056_2241, w_056_2242, w_056_2244, w_056_2246, w_056_2247, w_056_2249, w_056_2251, w_056_2253, w_056_2255, w_056_2257, w_056_2258, w_056_2259, w_056_2260, w_056_2263, w_056_2266, w_056_2267, w_056_2268, w_056_2272, w_056_2274, w_056_2277, w_056_2278, w_056_2279, w_056_2280, w_056_2282, w_056_2284, w_056_2286, w_056_2287, w_056_2288, w_056_2291, w_056_2292, w_056_2293, w_056_2295, w_056_2296, w_056_2298, w_056_2300, w_056_2302, w_056_2303, w_056_2309, w_056_2310, w_056_2311, w_056_2315, w_056_2317, w_056_2321, w_056_2325, w_056_2327, w_056_2328, w_056_2329, w_056_2330, w_056_2331, w_056_2333, w_056_2337, w_056_2339, w_056_2343, w_056_2348, w_056_2349, w_056_2353, w_056_2357, w_056_2358, w_056_2360, w_056_2365, w_056_2374, w_056_2376, w_056_2379, w_056_2381, w_056_2382, w_056_2386, w_056_2387, w_056_2388, w_056_2389, w_056_2390, w_056_2393, w_056_2395, w_056_2399, w_056_2401, w_056_2402, w_056_2403, w_056_2406, w_056_2407, w_056_2409, w_056_2412, w_056_2415, w_056_2419, w_056_2423, w_056_2424, w_056_2425, w_056_2428, w_056_2429, w_056_2430, w_056_2431, w_056_2432, w_056_2437, w_056_2438, w_056_2440, w_056_2447, w_056_2448, w_056_2450, w_056_2451, w_056_2452, w_056_2453, w_056_2459, w_056_2460, w_056_2461, w_056_2462, w_056_2463, w_056_2464, w_056_2465, w_056_2466, w_056_2467, w_056_2472, w_056_2474, w_056_2475, w_056_2478, w_056_2480, w_056_2484, w_056_2486, w_056_2489, w_056_2490, w_056_2497, w_056_2499, w_056_2500, w_056_2502, w_056_2504, w_056_2505, w_056_2506, w_056_2510, w_056_2511, w_056_2513, w_056_2517, w_056_2518, w_056_2520, w_056_2523, w_056_2526, w_056_2530, w_056_2531, w_056_2532, w_056_2534, w_056_2535, w_056_2536, w_056_2540, w_056_2542, w_056_2544, w_056_2546, w_056_2548, w_056_2551, w_056_2553, w_056_2556, w_056_2561, w_056_2562, w_056_2563, w_056_2564, w_056_2565, w_056_2572, w_056_2574, w_056_2575, w_056_2576, w_056_2577, w_056_2578, w_056_2581, w_056_2591, w_056_2592, w_056_2595, w_056_2596, w_056_2602, w_056_2605, w_056_2607, w_056_2608, w_056_2610, w_056_2612, w_056_2614, w_056_2617, w_056_2618, w_056_2619, w_056_2620, w_056_2621, w_056_2622, w_056_2626, w_056_2627, w_056_2629, w_056_2632, w_056_2634, w_056_2635, w_056_2637, w_056_2639, w_056_2640, w_056_2641, w_056_2642, w_056_2644, w_056_2647, w_056_2648, w_056_2649, w_056_2650, w_056_2651, w_056_2652, w_056_2657, w_056_2658, w_056_2659, w_056_2664, w_056_2665, w_056_2670, w_056_2671, w_056_2673, w_056_2674, w_056_2676, w_056_2678, w_056_2679, w_056_2681, w_056_2683, w_056_2685, w_056_2686, w_056_2687, w_056_2688, w_056_2689, w_056_2690, w_056_2691, w_056_2697, w_056_2701, w_056_2704, w_056_2705, w_056_2706, w_056_2707, w_056_2708, w_056_2709, w_056_2713, w_056_2714, w_056_2715, w_056_2716, w_056_2717, w_056_2718, w_056_2719, w_056_2720, w_056_2721, w_056_2722, w_056_2723, w_056_2725;
  wire w_057_000, w_057_001, w_057_002, w_057_003, w_057_004, w_057_006, w_057_007, w_057_008, w_057_009, w_057_010, w_057_011, w_057_012, w_057_013, w_057_015, w_057_016, w_057_017, w_057_018, w_057_019, w_057_020, w_057_021, w_057_022, w_057_023, w_057_024, w_057_025, w_057_027, w_057_028, w_057_029, w_057_030, w_057_031, w_057_032, w_057_033, w_057_034, w_057_035, w_057_036, w_057_037, w_057_038, w_057_039, w_057_040, w_057_041, w_057_042, w_057_043, w_057_044, w_057_045, w_057_046, w_057_047, w_057_048, w_057_049, w_057_050, w_057_051, w_057_052, w_057_053, w_057_054, w_057_055, w_057_056, w_057_057, w_057_058, w_057_059, w_057_060, w_057_061, w_057_062, w_057_063, w_057_064, w_057_065, w_057_066, w_057_067, w_057_069, w_057_070, w_057_071, w_057_072, w_057_074, w_057_076, w_057_077, w_057_078, w_057_079, w_057_080, w_057_081, w_057_082, w_057_083, w_057_084, w_057_085, w_057_086, w_057_087, w_057_088, w_057_089, w_057_090, w_057_091, w_057_092, w_057_093, w_057_094, w_057_095, w_057_096, w_057_097, w_057_098, w_057_099, w_057_100, w_057_101, w_057_102, w_057_103, w_057_104, w_057_105, w_057_106, w_057_107, w_057_108, w_057_109, w_057_110, w_057_111, w_057_112, w_057_114, w_057_115, w_057_116, w_057_117, w_057_118, w_057_119, w_057_120, w_057_121, w_057_122, w_057_123, w_057_124, w_057_125, w_057_126, w_057_127, w_057_128, w_057_129, w_057_130, w_057_131, w_057_132, w_057_133, w_057_134, w_057_135, w_057_136, w_057_137, w_057_138, w_057_139, w_057_140, w_057_141, w_057_142, w_057_143, w_057_144, w_057_145, w_057_146, w_057_147, w_057_148, w_057_149, w_057_150, w_057_151, w_057_152, w_057_153, w_057_154, w_057_155, w_057_156, w_057_157, w_057_158, w_057_159, w_057_160, w_057_161, w_057_162, w_057_163, w_057_164, w_057_165, w_057_166, w_057_167, w_057_168, w_057_169, w_057_170, w_057_172, w_057_173, w_057_174, w_057_175, w_057_176, w_057_177, w_057_178, w_057_179, w_057_180, w_057_181, w_057_182, w_057_183, w_057_184, w_057_185, w_057_186, w_057_187, w_057_188, w_057_189, w_057_190, w_057_191, w_057_192, w_057_193, w_057_194, w_057_195, w_057_196, w_057_197, w_057_198, w_057_199, w_057_200, w_057_201, w_057_202, w_057_203, w_057_204, w_057_205, w_057_206, w_057_207, w_057_208, w_057_209, w_057_210, w_057_211, w_057_212, w_057_213, w_057_214, w_057_215, w_057_216, w_057_217, w_057_218, w_057_219, w_057_220, w_057_221, w_057_222, w_057_224, w_057_225, w_057_226, w_057_227, w_057_228, w_057_229, w_057_230, w_057_231, w_057_232, w_057_233, w_057_234, w_057_235, w_057_236, w_057_237, w_057_238, w_057_240, w_057_241, w_057_242, w_057_243, w_057_244, w_057_245, w_057_246, w_057_247, w_057_248, w_057_249, w_057_250, w_057_251, w_057_252, w_057_253, w_057_254, w_057_255, w_057_256, w_057_257, w_057_258, w_057_259, w_057_260, w_057_261, w_057_262, w_057_263, w_057_264, w_057_265, w_057_266, w_057_267, w_057_268, w_057_269, w_057_270, w_057_271, w_057_272, w_057_273, w_057_274, w_057_275, w_057_276, w_057_277, w_057_278, w_057_279, w_057_280, w_057_281, w_057_282, w_057_283, w_057_284, w_057_285, w_057_286, w_057_287, w_057_288, w_057_289, w_057_290, w_057_291, w_057_292, w_057_293, w_057_294, w_057_295, w_057_296, w_057_297, w_057_298, w_057_299, w_057_300, w_057_301, w_057_302, w_057_303, w_057_304, w_057_305, w_057_306, w_057_307, w_057_308, w_057_309, w_057_310, w_057_311, w_057_312, w_057_313, w_057_314, w_057_315, w_057_316, w_057_317, w_057_318, w_057_319, w_057_320, w_057_321, w_057_322, w_057_324, w_057_326, w_057_327, w_057_328, w_057_329, w_057_330, w_057_331, w_057_332, w_057_333, w_057_334, w_057_335, w_057_336, w_057_337, w_057_338, w_057_339, w_057_340, w_057_341, w_057_342, w_057_343, w_057_344, w_057_345, w_057_346, w_057_347, w_057_348, w_057_349, w_057_350, w_057_351, w_057_352, w_057_353, w_057_354, w_057_355, w_057_356, w_057_357, w_057_358, w_057_359, w_057_360, w_057_361, w_057_362, w_057_363, w_057_364, w_057_365, w_057_366, w_057_367, w_057_369, w_057_370, w_057_371, w_057_372, w_057_373, w_057_374, w_057_375, w_057_376, w_057_377, w_057_378, w_057_379, w_057_380, w_057_381, w_057_382, w_057_383, w_057_384, w_057_385, w_057_386, w_057_387, w_057_388, w_057_389, w_057_390, w_057_391, w_057_393, w_057_395, w_057_396, w_057_397, w_057_398, w_057_399, w_057_400, w_057_401, w_057_402, w_057_403, w_057_404, w_057_405, w_057_407, w_057_408, w_057_409, w_057_410, w_057_411, w_057_412, w_057_413, w_057_414, w_057_415, w_057_416, w_057_417, w_057_418, w_057_419, w_057_420, w_057_421, w_057_422, w_057_424, w_057_425, w_057_426, w_057_427, w_057_428, w_057_429, w_057_430, w_057_431, w_057_432, w_057_433, w_057_434, w_057_435, w_057_436, w_057_437, w_057_438, w_057_439, w_057_440, w_057_441, w_057_442, w_057_443, w_057_445, w_057_446, w_057_447, w_057_448, w_057_449, w_057_450, w_057_451, w_057_453, w_057_454, w_057_455, w_057_456, w_057_457, w_057_458, w_057_459, w_057_460, w_057_461, w_057_462, w_057_463, w_057_464, w_057_465, w_057_466, w_057_467, w_057_468, w_057_469, w_057_470, w_057_471, w_057_472, w_057_473, w_057_474, w_057_475, w_057_476, w_057_477, w_057_478, w_057_479, w_057_481, w_057_483, w_057_484, w_057_485, w_057_486, w_057_487, w_057_488, w_057_489, w_057_490, w_057_491, w_057_492, w_057_493, w_057_494, w_057_495, w_057_496, w_057_497, w_057_498, w_057_499, w_057_500, w_057_501, w_057_502, w_057_503, w_057_504, w_057_506, w_057_507, w_057_508, w_057_509, w_057_510, w_057_511, w_057_512, w_057_513, w_057_514, w_057_515, w_057_516, w_057_518, w_057_519, w_057_520, w_057_521, w_057_522, w_057_523, w_057_524, w_057_525, w_057_526, w_057_527, w_057_528, w_057_529, w_057_530, w_057_531, w_057_532, w_057_533, w_057_534, w_057_535, w_057_536, w_057_537, w_057_538, w_057_539, w_057_540, w_057_541, w_057_542, w_057_543, w_057_544, w_057_545, w_057_546, w_057_547, w_057_548, w_057_549, w_057_550, w_057_551, w_057_552, w_057_553, w_057_554, w_057_555, w_057_556, w_057_557, w_057_558, w_057_559, w_057_560, w_057_562, w_057_563, w_057_564, w_057_565, w_057_566, w_057_567, w_057_568, w_057_569, w_057_570, w_057_571, w_057_572, w_057_573, w_057_574, w_057_575, w_057_576, w_057_577, w_057_578, w_057_579, w_057_580, w_057_581, w_057_582, w_057_583, w_057_584, w_057_585, w_057_586, w_057_587, w_057_588, w_057_589, w_057_590, w_057_591, w_057_592, w_057_593, w_057_594, w_057_595, w_057_596, w_057_598, w_057_599, w_057_600, w_057_601, w_057_602, w_057_603, w_057_604, w_057_605, w_057_606, w_057_607, w_057_608, w_057_609, w_057_610, w_057_611, w_057_612, w_057_613, w_057_614, w_057_615, w_057_616, w_057_617, w_057_618, w_057_619, w_057_620, w_057_621, w_057_622, w_057_623, w_057_624, w_057_625, w_057_626, w_057_627, w_057_628, w_057_629, w_057_630, w_057_631, w_057_632, w_057_633, w_057_634, w_057_635, w_057_636, w_057_637, w_057_638, w_057_639, w_057_640, w_057_641, w_057_642, w_057_643, w_057_644, w_057_645, w_057_646, w_057_647, w_057_649, w_057_650, w_057_651, w_057_652, w_057_653, w_057_654, w_057_655, w_057_656, w_057_657, w_057_658, w_057_659, w_057_660, w_057_661, w_057_662, w_057_663, w_057_664, w_057_665, w_057_667, w_057_668, w_057_669, w_057_670, w_057_671, w_057_672, w_057_673, w_057_674, w_057_675, w_057_676, w_057_677, w_057_678, w_057_679, w_057_680, w_057_681, w_057_682, w_057_683, w_057_684, w_057_685, w_057_686, w_057_687, w_057_688, w_057_689, w_057_690, w_057_691, w_057_692, w_057_693, w_057_694, w_057_695, w_057_696, w_057_697, w_057_698, w_057_699, w_057_700, w_057_701, w_057_702, w_057_703, w_057_704, w_057_705, w_057_706, w_057_707, w_057_708, w_057_709, w_057_710, w_057_711, w_057_712, w_057_713, w_057_714, w_057_715, w_057_716, w_057_718, w_057_719, w_057_720, w_057_721, w_057_722, w_057_723, w_057_724, w_057_725, w_057_726, w_057_727, w_057_728, w_057_729, w_057_730, w_057_731, w_057_732, w_057_733, w_057_734, w_057_735, w_057_736, w_057_737, w_057_738, w_057_739, w_057_740, w_057_741, w_057_742, w_057_743, w_057_744, w_057_745, w_057_746, w_057_747, w_057_748, w_057_749, w_057_750, w_057_751, w_057_752, w_057_753, w_057_754, w_057_755, w_057_756, w_057_757, w_057_758, w_057_759, w_057_760, w_057_761, w_057_762, w_057_763, w_057_764, w_057_765, w_057_766, w_057_767, w_057_768, w_057_770, w_057_771, w_057_772, w_057_773, w_057_775, w_057_776, w_057_777, w_057_779, w_057_780, w_057_781, w_057_782, w_057_783, w_057_784, w_057_785, w_057_786, w_057_787, w_057_788, w_057_789, w_057_790, w_057_791, w_057_792, w_057_793, w_057_794, w_057_795, w_057_796, w_057_797, w_057_798, w_057_799, w_057_800, w_057_801, w_057_802, w_057_803, w_057_804, w_057_805, w_057_806, w_057_807, w_057_808, w_057_809, w_057_810, w_057_811, w_057_812, w_057_813, w_057_814, w_057_815, w_057_816, w_057_817, w_057_818, w_057_819, w_057_820, w_057_821, w_057_822, w_057_823, w_057_824, w_057_825, w_057_826, w_057_827, w_057_828, w_057_829, w_057_830, w_057_831, w_057_832, w_057_833, w_057_834;
  wire w_058_001, w_058_002, w_058_003, w_058_005, w_058_006, w_058_008, w_058_009, w_058_010, w_058_012, w_058_013, w_058_014, w_058_015, w_058_017, w_058_020, w_058_022, w_058_023, w_058_024, w_058_028, w_058_031, w_058_032, w_058_035, w_058_036, w_058_040, w_058_041, w_058_042, w_058_044, w_058_045, w_058_046, w_058_047, w_058_048, w_058_049, w_058_050, w_058_051, w_058_052, w_058_053, w_058_055, w_058_056, w_058_057, w_058_059, w_058_060, w_058_061, w_058_065, w_058_066, w_058_068, w_058_069, w_058_070, w_058_071, w_058_072, w_058_073, w_058_074, w_058_079, w_058_080, w_058_081, w_058_082, w_058_083, w_058_085, w_058_087, w_058_088, w_058_090, w_058_091, w_058_092, w_058_093, w_058_094, w_058_095, w_058_096, w_058_097, w_058_098, w_058_099, w_058_101, w_058_102, w_058_103, w_058_104, w_058_105, w_058_106, w_058_107, w_058_108, w_058_111, w_058_113, w_058_115, w_058_117, w_058_118, w_058_119, w_058_121, w_058_123, w_058_126, w_058_128, w_058_129, w_058_131, w_058_132, w_058_133, w_058_134, w_058_136, w_058_140, w_058_143, w_058_144, w_058_145, w_058_146, w_058_147, w_058_150, w_058_151, w_058_152, w_058_154, w_058_155, w_058_156, w_058_157, w_058_158, w_058_160, w_058_162, w_058_164, w_058_166, w_058_169, w_058_172, w_058_173, w_058_175, w_058_176, w_058_177, w_058_179, w_058_181, w_058_182, w_058_183, w_058_184, w_058_186, w_058_189, w_058_190, w_058_192, w_058_195, w_058_196, w_058_197, w_058_199, w_058_201, w_058_202, w_058_203, w_058_204, w_058_205, w_058_206, w_058_208, w_058_209, w_058_210, w_058_212, w_058_216, w_058_217, w_058_219, w_058_220, w_058_224, w_058_225, w_058_226, w_058_227, w_058_228, w_058_229, w_058_230, w_058_232, w_058_236, w_058_237, w_058_238, w_058_239, w_058_240, w_058_242, w_058_243, w_058_244, w_058_245, w_058_246, w_058_250, w_058_253, w_058_254, w_058_255, w_058_256, w_058_257, w_058_259, w_058_261, w_058_262, w_058_263, w_058_264, w_058_266, w_058_267, w_058_268, w_058_269, w_058_271, w_058_274, w_058_275, w_058_276, w_058_278, w_058_279, w_058_282, w_058_284, w_058_285, w_058_286, w_058_288, w_058_289, w_058_290, w_058_292, w_058_295, w_058_296, w_058_297, w_058_298, w_058_300, w_058_304, w_058_306, w_058_307, w_058_308, w_058_309, w_058_310, w_058_311, w_058_312, w_058_314, w_058_315, w_058_316, w_058_317, w_058_319, w_058_320, w_058_321, w_058_322, w_058_323, w_058_324, w_058_325, w_058_326, w_058_327, w_058_331, w_058_332, w_058_336, w_058_337, w_058_338, w_058_339, w_058_340, w_058_344, w_058_345, w_058_346, w_058_348, w_058_349, w_058_350, w_058_351, w_058_353, w_058_355, w_058_357, w_058_358, w_058_359, w_058_360, w_058_361, w_058_365, w_058_367, w_058_369, w_058_370, w_058_371, w_058_372, w_058_373, w_058_374, w_058_376, w_058_377, w_058_379, w_058_380, w_058_381, w_058_384, w_058_385, w_058_386, w_058_387, w_058_388, w_058_389, w_058_390, w_058_392, w_058_394, w_058_396, w_058_397, w_058_398, w_058_399, w_058_401, w_058_402, w_058_403, w_058_404, w_058_405, w_058_407, w_058_408, w_058_410, w_058_417, w_058_419, w_058_420, w_058_421, w_058_422, w_058_423, w_058_424, w_058_425, w_058_426, w_058_427, w_058_428, w_058_430, w_058_431, w_058_433, w_058_434, w_058_435, w_058_436, w_058_438, w_058_439, w_058_440, w_058_441, w_058_442, w_058_443, w_058_444, w_058_446, w_058_447, w_058_448, w_058_449, w_058_451, w_058_452, w_058_453, w_058_455, w_058_458, w_058_459, w_058_460, w_058_461, w_058_462, w_058_463, w_058_465, w_058_466, w_058_467, w_058_469, w_058_470, w_058_471, w_058_474, w_058_476, w_058_477, w_058_478, w_058_480, w_058_482, w_058_483, w_058_484, w_058_487, w_058_489, w_058_490, w_058_491, w_058_492, w_058_493, w_058_494, w_058_496, w_058_498, w_058_499, w_058_500, w_058_502, w_058_503, w_058_504, w_058_506, w_058_508, w_058_509, w_058_510, w_058_511, w_058_512, w_058_513, w_058_517, w_058_518, w_058_519, w_058_520, w_058_521, w_058_522, w_058_526, w_058_527, w_058_529, w_058_530, w_058_531, w_058_532, w_058_534, w_058_535, w_058_536, w_058_537, w_058_538, w_058_539, w_058_540, w_058_542, w_058_547, w_058_548, w_058_549, w_058_550, w_058_551, w_058_552, w_058_555, w_058_556, w_058_557, w_058_558, w_058_559, w_058_560, w_058_561, w_058_562, w_058_563, w_058_565, w_058_568, w_058_570, w_058_571, w_058_572, w_058_573, w_058_574, w_058_575, w_058_576, w_058_578, w_058_581, w_058_583, w_058_584, w_058_585, w_058_586, w_058_587, w_058_588, w_058_589, w_058_591, w_058_594, w_058_596, w_058_597, w_058_598, w_058_601, w_058_603, w_058_604, w_058_605, w_058_608, w_058_609, w_058_610, w_058_611, w_058_612, w_058_613, w_058_614, w_058_616, w_058_617, w_058_619, w_058_620, w_058_623, w_058_624, w_058_625, w_058_626, w_058_628, w_058_631, w_058_632, w_058_633, w_058_636, w_058_637, w_058_639, w_058_640, w_058_641, w_058_642, w_058_643, w_058_644, w_058_645, w_058_647, w_058_648, w_058_649, w_058_650, w_058_651, w_058_652, w_058_653, w_058_657, w_058_658, w_058_659, w_058_660, w_058_662, w_058_663, w_058_664, w_058_665, w_058_668, w_058_669, w_058_670, w_058_671, w_058_673, w_058_674, w_058_676, w_058_678, w_058_679, w_058_681, w_058_683, w_058_685, w_058_688, w_058_690, w_058_693, w_058_694, w_058_695, w_058_696, w_058_697, w_058_699, w_058_705, w_058_707, w_058_710, w_058_711, w_058_712, w_058_714, w_058_715, w_058_716, w_058_717, w_058_718, w_058_721, w_058_722, w_058_723, w_058_724, w_058_726, w_058_728, w_058_730, w_058_731, w_058_732, w_058_734, w_058_735, w_058_736, w_058_737, w_058_738, w_058_740, w_058_741, w_058_744, w_058_746, w_058_747, w_058_749, w_058_750, w_058_751, w_058_753, w_058_755, w_058_756, w_058_760, w_058_761, w_058_762, w_058_763, w_058_764, w_058_765, w_058_766, w_058_771, w_058_772, w_058_774, w_058_778, w_058_780, w_058_781, w_058_783, w_058_785, w_058_786, w_058_787, w_058_789, w_058_790, w_058_791, w_058_792, w_058_793, w_058_794, w_058_795, w_058_796, w_058_797, w_058_798, w_058_799, w_058_800, w_058_801, w_058_802, w_058_803, w_058_804, w_058_806, w_058_808, w_058_810, w_058_811, w_058_812, w_058_814, w_058_816, w_058_817, w_058_819, w_058_820, w_058_821, w_058_822, w_058_823, w_058_824, w_058_825, w_058_826, w_058_827, w_058_829, w_058_831, w_058_832, w_058_834, w_058_835, w_058_837, w_058_838, w_058_839, w_058_840, w_058_842, w_058_843, w_058_844, w_058_845, w_058_848, w_058_849, w_058_850, w_058_857, w_058_858, w_058_860, w_058_861, w_058_862, w_058_863, w_058_864, w_058_865, w_058_866, w_058_867, w_058_868, w_058_870, w_058_871, w_058_872, w_058_873, w_058_874, w_058_875, w_058_876, w_058_877, w_058_879, w_058_880, w_058_881, w_058_884, w_058_886, w_058_887, w_058_889, w_058_890, w_058_891, w_058_892, w_058_893, w_058_894, w_058_895, w_058_896, w_058_897, w_058_898, w_058_899, w_058_900, w_058_901, w_058_902, w_058_903, w_058_905, w_058_907, w_058_908, w_058_909, w_058_910, w_058_911, w_058_912, w_058_913, w_058_915, w_058_916, w_058_917, w_058_918, w_058_922, w_058_925, w_058_926, w_058_928, w_058_930, w_058_931, w_058_934, w_058_936, w_058_937, w_058_939, w_058_941, w_058_942, w_058_943, w_058_944, w_058_945, w_058_946, w_058_947, w_058_948, w_058_950, w_058_953, w_058_954, w_058_955, w_058_957, w_058_958, w_058_960, w_058_963, w_058_966, w_058_967, w_058_968, w_058_969, w_058_971, w_058_974, w_058_975, w_058_977, w_058_979, w_058_980, w_058_981, w_058_982, w_058_984, w_058_985, w_058_990, w_058_993, w_058_994, w_058_995, w_058_996, w_058_997, w_058_998, w_058_999, w_058_1000, w_058_1001, w_058_1002, w_058_1003, w_058_1004, w_058_1005, w_058_1006, w_058_1008, w_058_1009, w_058_1010, w_058_1011, w_058_1012, w_058_1013, w_058_1015, w_058_1016, w_058_1017, w_058_1019, w_058_1020, w_058_1021, w_058_1022, w_058_1026, w_058_1027, w_058_1028, w_058_1031, w_058_1032, w_058_1033, w_058_1034, w_058_1036, w_058_1039, w_058_1041, w_058_1045, w_058_1046, w_058_1048, w_058_1052, w_058_1053, w_058_1054, w_058_1055, w_058_1057, w_058_1058, w_058_1059, w_058_1061, w_058_1062, w_058_1063, w_058_1064, w_058_1067, w_058_1070, w_058_1072, w_058_1073, w_058_1075, w_058_1076, w_058_1077, w_058_1078, w_058_1079, w_058_1082, w_058_1083, w_058_1084, w_058_1085, w_058_1087, w_058_1089, w_058_1090, w_058_1091, w_058_1094, w_058_1095, w_058_1096, w_058_1102, w_058_1103, w_058_1105, w_058_1107, w_058_1110, w_058_1111, w_058_1112, w_058_1113, w_058_1115, w_058_1116, w_058_1117, w_058_1118, w_058_1119, w_058_1120, w_058_1121, w_058_1123, w_058_1124, w_058_1125, w_058_1126, w_058_1128, w_058_1130, w_058_1131, w_058_1132, w_058_1133, w_058_1135, w_058_1136, w_058_1137, w_058_1138, w_058_1141, w_058_1142, w_058_1143, w_058_1145, w_058_1146, w_058_1148, w_058_1149, w_058_1150, w_058_1152, w_058_1153, w_058_1154, w_058_1155, w_058_1157, w_058_1158, w_058_1159, w_058_1163, w_058_1165, w_058_1166, w_058_1167, w_058_1168, w_058_1170, w_058_1171, w_058_1172, w_058_1173, w_058_1174, w_058_1178, w_058_1180, w_058_1182, w_058_1184, w_058_1185, w_058_1186, w_058_1187, w_058_1188, w_058_1190, w_058_1192, w_058_1193, w_058_1197, w_058_1198, w_058_1199, w_058_1200, w_058_1201, w_058_1202, w_058_1203, w_058_1204, w_058_1205, w_058_1208, w_058_1209, w_058_1211, w_058_1212, w_058_1213, w_058_1214, w_058_1216, w_058_1217, w_058_1218, w_058_1220, w_058_1221, w_058_1222, w_058_1223, w_058_1224, w_058_1225, w_058_1228, w_058_1231, w_058_1234, w_058_1235, w_058_1237, w_058_1238, w_058_1241, w_058_1242, w_058_1243, w_058_1244, w_058_1245, w_058_1246, w_058_1247, w_058_1249, w_058_1250, w_058_1251, w_058_1252, w_058_1254, w_058_1255, w_058_1258, w_058_1261, w_058_1262, w_058_1263, w_058_1264, w_058_1265, w_058_1266, w_058_1267, w_058_1270, w_058_1271, w_058_1272, w_058_1273, w_058_1274, w_058_1276, w_058_1277, w_058_1279, w_058_1280, w_058_1281, w_058_1283, w_058_1285, w_058_1287, w_058_1288, w_058_1289, w_058_1291, w_058_1292, w_058_1294, w_058_1296, w_058_1297, w_058_1298, w_058_1299, w_058_1303, w_058_1307, w_058_1308, w_058_1310, w_058_1312, w_058_1314, w_058_1315, w_058_1316, w_058_1319, w_058_1321, w_058_1323, w_058_1324, w_058_1326, w_058_1328, w_058_1329, w_058_1330, w_058_1331, w_058_1332, w_058_1333, w_058_1334, w_058_1335, w_058_1336, w_058_1337, w_058_1339, w_058_1342, w_058_1343, w_058_1344, w_058_1346, w_058_1347, w_058_1348, w_058_1349, w_058_1350, w_058_1351, w_058_1353, w_058_1354, w_058_1355, w_058_1357, w_058_1358, w_058_1359, w_058_1360, w_058_1364, w_058_1368, w_058_1369, w_058_1370, w_058_1371, w_058_1372, w_058_1375, w_058_1377, w_058_1378, w_058_1379, w_058_1380, w_058_1384, w_058_1385, w_058_1386, w_058_1388, w_058_1389, w_058_1391, w_058_1395, w_058_1396, w_058_1397, w_058_1398, w_058_1400, w_058_1401, w_058_1405, w_058_1406, w_058_1407, w_058_1408, w_058_1409, w_058_1410, w_058_1413, w_058_1415, w_058_1416, w_058_1417, w_058_1418, w_058_1419, w_058_1420, w_058_1421, w_058_1422, w_058_1424, w_058_1425, w_058_1426, w_058_1427, w_058_1432, w_058_1433, w_058_1434, w_058_1437, w_058_1440, w_058_1442, w_058_1443, w_058_1444, w_058_1445, w_058_1446, w_058_1447, w_058_1448, w_058_1450, w_058_1452, w_058_1453, w_058_1454, w_058_1456, w_058_1458, w_058_1459, w_058_1460, w_058_1461, w_058_1463, w_058_1465, w_058_1466, w_058_1467, w_058_1468, w_058_1469, w_058_1470, w_058_1471, w_058_1472, w_058_1473, w_058_1475, w_058_1476, w_058_1477, w_058_1478, w_058_1480, w_058_1482, w_058_1484, w_058_1485, w_058_1486, w_058_1489, w_058_1490, w_058_1491, w_058_1492, w_058_1493, w_058_1494, w_058_1495, w_058_1496, w_058_1497, w_058_1498, w_058_1500, w_058_1501, w_058_1503, w_058_1504, w_058_1506, w_058_1507, w_058_1508, w_058_1509, w_058_1513, w_058_1515, w_058_1516, w_058_1517, w_058_1518, w_058_1520, w_058_1521, w_058_1525, w_058_1526, w_058_1528, w_058_1529, w_058_1531, w_058_1532, w_058_1533, w_058_1534, w_058_1538, w_058_1539, w_058_1540, w_058_1541, w_058_1542, w_058_1543, w_058_1544, w_058_1545, w_058_1546, w_058_1549, w_058_1550, w_058_1551, w_058_1553, w_058_1555, w_058_1556, w_058_1557, w_058_1558, w_058_1559, w_058_1561, w_058_1562, w_058_1563, w_058_1565, w_058_1566, w_058_1567, w_058_1568, w_058_1569, w_058_1570, w_058_1571, w_058_1574, w_058_1576, w_058_1579, w_058_1580, w_058_1581, w_058_1582, w_058_1583, w_058_1584, w_058_1587, w_058_1588, w_058_1590, w_058_1595, w_058_1596, w_058_1597, w_058_1598, w_058_1600, w_058_1601, w_058_1604, w_058_1605, w_058_1608, w_058_1609, w_058_1613, w_058_1614, w_058_1617, w_058_1620, w_058_1621, w_058_1622, w_058_1623, w_058_1624, w_058_1625, w_058_1626, w_058_1628, w_058_1630, w_058_1631, w_058_1632, w_058_1634, w_058_1635, w_058_1636, w_058_1637, w_058_1638, w_058_1640, w_058_1641, w_058_1643, w_058_1644, w_058_1645, w_058_1646, w_058_1648, w_058_1649, w_058_1650, w_058_1651, w_058_1653, w_058_1658, w_058_1661, w_058_1662, w_058_1669, w_058_1676, w_058_1678, w_058_1679, w_058_1681, w_058_1683, w_058_1685, w_058_1687, w_058_1690, w_058_1691, w_058_1693, w_058_1696, w_058_1699, w_058_1701, w_058_1702, w_058_1703, w_058_1708, w_058_1710, w_058_1712, w_058_1714, w_058_1717, w_058_1719, w_058_1720, w_058_1721, w_058_1722, w_058_1726, w_058_1727, w_058_1731, w_058_1732, w_058_1734, w_058_1743, w_058_1744, w_058_1745, w_058_1751, w_058_1753, w_058_1754, w_058_1756, w_058_1757, w_058_1758, w_058_1760, w_058_1761, w_058_1762, w_058_1763, w_058_1767, w_058_1774, w_058_1775, w_058_1776, w_058_1777, w_058_1778, w_058_1787, w_058_1789, w_058_1794, w_058_1795, w_058_1798, w_058_1801, w_058_1805, w_058_1811, w_058_1814, w_058_1817, w_058_1818, w_058_1819, w_058_1820, w_058_1822, w_058_1827, w_058_1828, w_058_1831, w_058_1835, w_058_1836, w_058_1838, w_058_1842, w_058_1843, w_058_1846, w_058_1848, w_058_1854, w_058_1855, w_058_1856, w_058_1858, w_058_1860, w_058_1861, w_058_1862, w_058_1864, w_058_1867, w_058_1868, w_058_1869, w_058_1871, w_058_1872, w_058_1874, w_058_1878, w_058_1881, w_058_1883, w_058_1884, w_058_1885, w_058_1888, w_058_1889, w_058_1895, w_058_1896, w_058_1901, w_058_1902, w_058_1903, w_058_1907, w_058_1909, w_058_1910, w_058_1911, w_058_1912, w_058_1914, w_058_1917, w_058_1921, w_058_1922, w_058_1925, w_058_1926, w_058_1929, w_058_1932, w_058_1935, w_058_1936, w_058_1939, w_058_1940, w_058_1944, w_058_1945, w_058_1947, w_058_1948, w_058_1950, w_058_1951, w_058_1955, w_058_1959, w_058_1963, w_058_1966, w_058_1967, w_058_1968, w_058_1974, w_058_1975, w_058_1978, w_058_1981, w_058_1984, w_058_1985, w_058_1986, w_058_1987, w_058_1989, w_058_1994, w_058_1995, w_058_1996, w_058_1999, w_058_2001, w_058_2003, w_058_2004, w_058_2005, w_058_2013, w_058_2016, w_058_2019, w_058_2020, w_058_2025, w_058_2028, w_058_2031, w_058_2035, w_058_2040, w_058_2042, w_058_2044, w_058_2047, w_058_2053, w_058_2055, w_058_2056, w_058_2059, w_058_2063, w_058_2065, w_058_2068, w_058_2069, w_058_2073, w_058_2074, w_058_2075, w_058_2078, w_058_2080, w_058_2082, w_058_2083, w_058_2086, w_058_2088, w_058_2093, w_058_2097, w_058_2098, w_058_2100, w_058_2103, w_058_2106, w_058_2113, w_058_2115, w_058_2117, w_058_2123, w_058_2124, w_058_2125, w_058_2126, w_058_2127, w_058_2128, w_058_2130, w_058_2131, w_058_2134, w_058_2135, w_058_2138, w_058_2140, w_058_2143, w_058_2144, w_058_2146, w_058_2147, w_058_2148, w_058_2150, w_058_2151, w_058_2152, w_058_2154, w_058_2155, w_058_2157, w_058_2158, w_058_2159, w_058_2160, w_058_2161, w_058_2162, w_058_2165, w_058_2170, w_058_2172, w_058_2173, w_058_2174, w_058_2175, w_058_2176, w_058_2181, w_058_2183, w_058_2186, w_058_2189, w_058_2190, w_058_2193, w_058_2194, w_058_2199, w_058_2203, w_058_2205, w_058_2208, w_058_2209, w_058_2210, w_058_2212, w_058_2214, w_058_2216, w_058_2217, w_058_2218, w_058_2221, w_058_2222, w_058_2223, w_058_2224, w_058_2225, w_058_2228, w_058_2229, w_058_2230, w_058_2235, w_058_2236, w_058_2237, w_058_2239, w_058_2240, w_058_2241, w_058_2243, w_058_2244, w_058_2245, w_058_2249, w_058_2250, w_058_2251, w_058_2263, w_058_2264, w_058_2265, w_058_2267, w_058_2269, w_058_2272, w_058_2276, w_058_2278, w_058_2279, w_058_2280, w_058_2284, w_058_2285, w_058_2287, w_058_2289, w_058_2293, w_058_2299, w_058_2300, w_058_2305, w_058_2307, w_058_2308, w_058_2310, w_058_2311, w_058_2314, w_058_2317, w_058_2318, w_058_2319, w_058_2320, w_058_2322, w_058_2323, w_058_2325, w_058_2327, w_058_2329, w_058_2330, w_058_2333, w_058_2338, w_058_2341, w_058_2344, w_058_2349, w_058_2352, w_058_2354, w_058_2355, w_058_2358, w_058_2361, w_058_2362, w_058_2369, w_058_2371, w_058_2372, w_058_2374, w_058_2376, w_058_2380, w_058_2382, w_058_2383, w_058_2385, w_058_2388, w_058_2389, w_058_2390, w_058_2391, w_058_2398, w_058_2399, w_058_2400, w_058_2401, w_058_2402, w_058_2403, w_058_2407, w_058_2408, w_058_2411, w_058_2412, w_058_2414, w_058_2415, w_058_2419, w_058_2420, w_058_2425, w_058_2426, w_058_2427, w_058_2428, w_058_2429, w_058_2439, w_058_2440, w_058_2441, w_058_2443, w_058_2444, w_058_2450, w_058_2452, w_058_2454, w_058_2455, w_058_2461, w_058_2465, w_058_2469, w_058_2471, w_058_2474, w_058_2488, w_058_2489, w_058_2493, w_058_2499, w_058_2502, w_058_2503, w_058_2508, w_058_2509, w_058_2514, w_058_2515, w_058_2517, w_058_2519, w_058_2520, w_058_2523, w_058_2526, w_058_2527, w_058_2528, w_058_2534, w_058_2537, w_058_2539, w_058_2543, w_058_2545, w_058_2547, w_058_2548, w_058_2549, w_058_2550, w_058_2551, w_058_2553, w_058_2554, w_058_2556, w_058_2560, w_058_2565, w_058_2569, w_058_2571, w_058_2572, w_058_2573, w_058_2574, w_058_2575, w_058_2578, w_058_2580, w_058_2586, w_058_2588, w_058_2592, w_058_2595, w_058_2596, w_058_2599, w_058_2600, w_058_2601, w_058_2603, w_058_2605, w_058_2613, w_058_2615, w_058_2616, w_058_2617, w_058_2630, w_058_2631, w_058_2632, w_058_2635, w_058_2639, w_058_2640, w_058_2641, w_058_2642, w_058_2643, w_058_2645, w_058_2646, w_058_2647, w_058_2649, w_058_2652, w_058_2656, w_058_2668, w_058_2669, w_058_2670, w_058_2672, w_058_2677, w_058_2678, w_058_2680, w_058_2683, w_058_2685, w_058_2687, w_058_2690, w_058_2693, w_058_2697, w_058_2701, w_058_2702, w_058_2703, w_058_2704, w_058_2707, w_058_2708, w_058_2709, w_058_2710, w_058_2712, w_058_2714, w_058_2717, w_058_2718, w_058_2719, w_058_2720, w_058_2721, w_058_2727, w_058_2729, w_058_2731, w_058_2732, w_058_2734, w_058_2735, w_058_2736, w_058_2737, w_058_2741, w_058_2746, w_058_2750, w_058_2752, w_058_2754, w_058_2756, w_058_2757, w_058_2760, w_058_2762, w_058_2763, w_058_2766, w_058_2768, w_058_2771, w_058_2775, w_058_2779, w_058_2784, w_058_2786, w_058_2787, w_058_2788, w_058_2789, w_058_2790, w_058_2792, w_058_2793, w_058_2796, w_058_2798, w_058_2802, w_058_2803, w_058_2805, w_058_2806, w_058_2813, w_058_2815, w_058_2818, w_058_2819, w_058_2820, w_058_2821, w_058_2823, w_058_2824, w_058_2827, w_058_2828, w_058_2829, w_058_2831, w_058_2837, w_058_2843, w_058_2844, w_058_2848, w_058_2849, w_058_2850, w_058_2852, w_058_2856, w_058_2858, w_058_2859, w_058_2862, w_058_2863, w_058_2864, w_058_2867, w_058_2869, w_058_2871, w_058_2875, w_058_2876, w_058_2878, w_058_2879, w_058_2882, w_058_2883, w_058_2884, w_058_2885, w_058_2886, w_058_2890, w_058_2893, w_058_2894, w_058_2895, w_058_2899, w_058_2904, w_058_2907, w_058_2909, w_058_2910, w_058_2915, w_058_2918, w_058_2920, w_058_2921, w_058_2925, w_058_2926, w_058_2927, w_058_2928, w_058_2933, w_058_2936, w_058_2939, w_058_2940, w_058_2942, w_058_2946, w_058_2947, w_058_2952, w_058_2957, w_058_2962, w_058_2964, w_058_2965, w_058_2966, w_058_2969, w_058_2971, w_058_2976, w_058_2980, w_058_2982, w_058_2983, w_058_2984, w_058_2987, w_058_2991, w_058_2993, w_058_2995, w_058_2996, w_058_2997, w_058_2999, w_058_3000, w_058_3002, w_058_3003, w_058_3005, w_058_3006, w_058_3007, w_058_3008, w_058_3015, w_058_3017, w_058_3018, w_058_3020, w_058_3026, w_058_3027, w_058_3031, w_058_3035, w_058_3036, w_058_3038, w_058_3041, w_058_3044, w_058_3045, w_058_3048, w_058_3051, w_058_3052, w_058_3054, w_058_3055, w_058_3056, w_058_3057, w_058_3058, w_058_3070, w_058_3071, w_058_3072, w_058_3073, w_058_3074, w_058_3076, w_058_3078, w_058_3080, w_058_3081, w_058_3082, w_058_3087, w_058_3088, w_058_3089, w_058_3095, w_058_3096, w_058_3097, w_058_3098, w_058_3100, w_058_3101, w_058_3102, w_058_3106, w_058_3107, w_058_3109, w_058_3110, w_058_3112, w_058_3119, w_058_3120, w_058_3121, w_058_3122, w_058_3125, w_058_3126, w_058_3130, w_058_3133, w_058_3135, w_058_3137, w_058_3138, w_058_3139, w_058_3141, w_058_3144, w_058_3146, w_058_3147, w_058_3148, w_058_3150, w_058_3151, w_058_3152, w_058_3153, w_058_3154, w_058_3156, w_058_3163, w_058_3164, w_058_3167, w_058_3168, w_058_3169, w_058_3175, w_058_3179, w_058_3183, w_058_3185, w_058_3186, w_058_3187, w_058_3188, w_058_3191, w_058_3193, w_058_3195, w_058_3196, w_058_3198, w_058_3199, w_058_3200, w_058_3204, w_058_3206, w_058_3210, w_058_3214, w_058_3215, w_058_3216, w_058_3217, w_058_3218, w_058_3222, w_058_3223, w_058_3225, w_058_3228, w_058_3229, w_058_3232, w_058_3233, w_058_3235, w_058_3237, w_058_3239, w_058_3240, w_058_3241, w_058_3243, w_058_3245, w_058_3246, w_058_3253, w_058_3258, w_058_3261, w_058_3263, w_058_3265, w_058_3266, w_058_3269, w_058_3275, w_058_3276, w_058_3277, w_058_3281, w_058_3283, w_058_3285, w_058_3286, w_058_3289, w_058_3291, w_058_3292, w_058_3293, w_058_3295, w_058_3296, w_058_3297, w_058_3298, w_058_3299, w_058_3301, w_058_3305, w_058_3306, w_058_3309, w_058_3310, w_058_3312, w_058_3317, w_058_3318, w_058_3321, w_058_3322, w_058_3328, w_058_3329, w_058_3331, w_058_3333, w_058_3336, w_058_3338, w_058_3339, w_058_3344, w_058_3345, w_058_3346, w_058_3348;
  wire w_059_000, w_059_002, w_059_003, w_059_004, w_059_005, w_059_006, w_059_008, w_059_009, w_059_010, w_059_011, w_059_012, w_059_014, w_059_015, w_059_016, w_059_017, w_059_018, w_059_020, w_059_021, w_059_023, w_059_024, w_059_025, w_059_026, w_059_027, w_059_028, w_059_029, w_059_030, w_059_031, w_059_032, w_059_033, w_059_035, w_059_037, w_059_038, w_059_039, w_059_040, w_059_042, w_059_045, w_059_046, w_059_049, w_059_050, w_059_052, w_059_053, w_059_054, w_059_055, w_059_056, w_059_057, w_059_058, w_059_060, w_059_061, w_059_062, w_059_063, w_059_065, w_059_066, w_059_067, w_059_068, w_059_069, w_059_070, w_059_071, w_059_072, w_059_073, w_059_074, w_059_075, w_059_076, w_059_077, w_059_079, w_059_080, w_059_081, w_059_082, w_059_083, w_059_084, w_059_085, w_059_087, w_059_090, w_059_092, w_059_093, w_059_094, w_059_095, w_059_096, w_059_097, w_059_099, w_059_100, w_059_101, w_059_102, w_059_103, w_059_104, w_059_105, w_059_106, w_059_107, w_059_108, w_059_109, w_059_110, w_059_111, w_059_114, w_059_115, w_059_116, w_059_117, w_059_118, w_059_119, w_059_120, w_059_121, w_059_122, w_059_124, w_059_125, w_059_126, w_059_128, w_059_130, w_059_131, w_059_132, w_059_134, w_059_135, w_059_136, w_059_137, w_059_138, w_059_139, w_059_141, w_059_142, w_059_143, w_059_144, w_059_145, w_059_146, w_059_147, w_059_149, w_059_151, w_059_152, w_059_154, w_059_155, w_059_156, w_059_157, w_059_158, w_059_160, w_059_162, w_059_163, w_059_164, w_059_166, w_059_167, w_059_168, w_059_169, w_059_170, w_059_172, w_059_173, w_059_174, w_059_175, w_059_177, w_059_179, w_059_181, w_059_183, w_059_184, w_059_185, w_059_186, w_059_187, w_059_189, w_059_190, w_059_191, w_059_192, w_059_193, w_059_194, w_059_196, w_059_197, w_059_198, w_059_199, w_059_200, w_059_202, w_059_204, w_059_205, w_059_206, w_059_209, w_059_210, w_059_211, w_059_212, w_059_214, w_059_215, w_059_216, w_059_217, w_059_218, w_059_219, w_059_220, w_059_221, w_059_222, w_059_223, w_059_224, w_059_225, w_059_226, w_059_227, w_059_228, w_059_229, w_059_230, w_059_231, w_059_232, w_059_233, w_059_234, w_059_235, w_059_236, w_059_237, w_059_239, w_059_240, w_059_241, w_059_242, w_059_245, w_059_246, w_059_248, w_059_249, w_059_250, w_059_252, w_059_253, w_059_254, w_059_255, w_059_256, w_059_258, w_059_260, w_059_261, w_059_263, w_059_264, w_059_266, w_059_267, w_059_268, w_059_269, w_059_270, w_059_271, w_059_272, w_059_273, w_059_274, w_059_275, w_059_276, w_059_277, w_059_278, w_059_279, w_059_280, w_059_281, w_059_282, w_059_284, w_059_285, w_059_286, w_059_288, w_059_289, w_059_290, w_059_292, w_059_293, w_059_294, w_059_295, w_059_296, w_059_297, w_059_298, w_059_299, w_059_300, w_059_301, w_059_302, w_059_304, w_059_305, w_059_306, w_059_308, w_059_310, w_059_311, w_059_312, w_059_313, w_059_314, w_059_315, w_059_316, w_059_317, w_059_318, w_059_320, w_059_321, w_059_323, w_059_324, w_059_325, w_059_326, w_059_327, w_059_328, w_059_329, w_059_330, w_059_331, w_059_333, w_059_334, w_059_335, w_059_336, w_059_337, w_059_338, w_059_339, w_059_340, w_059_341, w_059_342, w_059_344, w_059_345, w_059_346, w_059_347, w_059_348, w_059_349, w_059_350, w_059_351, w_059_352, w_059_354, w_059_355, w_059_356, w_059_357, w_059_358, w_059_359, w_059_360, w_059_361, w_059_362, w_059_364, w_059_365, w_059_366, w_059_367, w_059_368, w_059_371, w_059_372, w_059_373, w_059_375, w_059_376, w_059_378, w_059_379, w_059_381, w_059_382, w_059_383, w_059_385, w_059_387, w_059_388, w_059_389, w_059_391, w_059_393, w_059_394, w_059_395, w_059_396, w_059_397, w_059_398, w_059_399, w_059_400, w_059_401, w_059_402, w_059_403, w_059_404, w_059_405, w_059_407, w_059_408, w_059_409, w_059_412, w_059_413, w_059_414, w_059_416, w_059_417, w_059_418, w_059_420, w_059_422, w_059_423, w_059_424, w_059_425, w_059_426, w_059_427, w_059_428, w_059_429, w_059_430, w_059_431, w_059_432, w_059_433, w_059_434, w_059_436, w_059_438, w_059_439, w_059_440, w_059_441, w_059_442, w_059_443, w_059_444, w_059_445, w_059_446, w_059_447, w_059_448, w_059_450, w_059_451, w_059_453, w_059_455, w_059_457, w_059_459, w_059_460, w_059_461, w_059_464, w_059_465, w_059_466, w_059_467, w_059_468, w_059_469, w_059_471, w_059_472, w_059_473, w_059_474, w_059_475, w_059_476, w_059_477, w_059_478, w_059_479, w_059_480, w_059_482, w_059_483, w_059_484, w_059_485, w_059_486, w_059_487, w_059_488, w_059_489, w_059_490, w_059_492, w_059_493, w_059_494, w_059_495, w_059_496, w_059_498, w_059_499, w_059_500, w_059_501, w_059_502, w_059_503, w_059_505, w_059_506, w_059_507, w_059_508, w_059_509, w_059_510, w_059_511, w_059_514, w_059_515, w_059_516, w_059_517, w_059_519, w_059_521, w_059_523, w_059_524, w_059_525, w_059_526, w_059_527, w_059_528, w_059_529, w_059_530, w_059_531, w_059_532, w_059_533, w_059_539, w_059_540, w_059_541, w_059_542, w_059_543, w_059_544, w_059_545, w_059_546, w_059_547, w_059_549, w_059_550, w_059_551, w_059_553, w_059_554, w_059_555, w_059_556, w_059_557, w_059_558, w_059_559, w_059_560, w_059_561, w_059_562, w_059_563, w_059_564, w_059_565, w_059_566, w_059_567, w_059_568, w_059_569, w_059_570, w_059_571, w_059_572, w_059_573, w_059_575, w_059_577, w_059_578, w_059_579, w_059_580, w_059_581, w_059_582, w_059_583, w_059_584, w_059_585, w_059_586, w_059_587, w_059_588, w_059_589, w_059_591, w_059_592, w_059_593, w_059_595, w_059_596, w_059_597, w_059_598, w_059_599, w_059_600, w_059_601, w_059_602, w_059_603, w_059_604, w_059_605, w_059_606, w_059_611, w_059_612, w_059_613, w_059_614, w_059_616, w_059_617, w_059_618, w_059_619, w_059_620, w_059_621, w_059_622, w_059_623, w_059_624, w_059_625, w_059_626, w_059_627, w_059_628, w_059_629, w_059_630, w_059_631, w_059_632, w_059_633, w_059_634, w_059_635, w_059_637, w_059_640, w_059_641, w_059_642, w_059_643, w_059_644, w_059_646, w_059_647, w_059_648, w_059_649, w_059_650, w_059_651, w_059_652, w_059_654, w_059_655, w_059_656, w_059_657, w_059_658, w_059_659, w_059_660, w_059_661, w_059_662, w_059_663, w_059_665, w_059_666, w_059_667, w_059_668, w_059_670, w_059_671, w_059_672, w_059_673, w_059_674, w_059_676, w_059_677, w_059_678, w_059_679, w_059_680, w_059_681, w_059_682, w_059_683, w_059_684, w_059_685, w_059_686, w_059_687, w_059_688, w_059_689, w_059_690, w_059_693, w_059_694, w_059_695, w_059_696, w_059_697, w_059_699, w_059_700, w_059_701, w_059_702, w_059_703, w_059_704, w_059_705, w_059_706, w_059_707, w_059_708, w_059_709, w_059_710, w_059_711, w_059_712, w_059_713, w_059_714, w_059_715, w_059_716, w_059_718, w_059_719, w_059_720, w_059_721, w_059_722, w_059_723, w_059_724, w_059_725, w_059_728, w_059_729, w_059_730, w_059_731, w_059_732, w_059_733, w_059_734, w_059_735, w_059_737, w_059_739, w_059_740, w_059_742, w_059_743, w_059_744, w_059_746, w_059_747, w_059_749, w_059_750, w_059_751, w_059_752, w_059_753, w_059_754, w_059_755, w_059_757, w_059_759, w_059_760, w_059_761, w_059_762, w_059_763, w_059_764, w_059_766, w_059_767, w_059_768, w_059_769, w_059_770, w_059_771, w_059_772, w_059_773, w_059_774, w_059_775, w_059_776, w_059_777, w_059_778, w_059_779, w_059_780, w_059_781, w_059_782, w_059_783, w_059_784, w_059_787, w_059_788, w_059_789, w_059_790, w_059_791, w_059_793, w_059_797, w_059_798, w_059_799, w_059_800, w_059_801, w_059_802, w_059_804, w_059_805, w_059_806, w_059_807, w_059_808, w_059_809, w_059_811, w_059_813, w_059_814, w_059_815, w_059_816, w_059_817, w_059_818, w_059_819, w_059_820, w_059_821, w_059_822, w_059_823, w_059_824, w_059_825, w_059_826, w_059_828, w_059_829, w_059_830, w_059_831, w_059_832, w_059_833, w_059_834, w_059_836, w_059_838, w_059_839, w_059_840, w_059_841, w_059_842, w_059_843, w_059_844, w_059_845, w_059_846, w_059_847, w_059_848, w_059_849, w_059_850, w_059_851, w_059_855, w_059_856, w_059_857, w_059_859, w_059_860, w_059_861, w_059_863, w_059_864, w_059_865, w_059_866, w_059_867, w_059_868, w_059_869, w_059_870, w_059_871, w_059_872, w_059_873, w_059_874, w_059_875, w_059_876, w_059_878, w_059_879, w_059_880, w_059_881, w_059_883, w_059_884, w_059_885, w_059_886, w_059_887, w_059_888, w_059_889, w_059_891, w_059_892, w_059_893, w_059_894, w_059_895, w_059_896, w_059_897, w_059_899, w_059_900, w_059_902, w_059_903, w_059_904, w_059_905, w_059_906, w_059_907, w_059_909, w_059_910, w_059_911, w_059_913, w_059_914, w_059_915, w_059_916, w_059_918, w_059_919, w_059_920, w_059_921, w_059_922, w_059_924, w_059_926, w_059_928, w_059_929, w_059_930, w_059_931, w_059_932, w_059_933, w_059_934, w_059_936, w_059_937, w_059_938, w_059_939, w_059_940, w_059_941, w_059_942, w_059_943, w_059_945, w_059_946, w_059_947, w_059_948, w_059_949, w_059_950, w_059_952, w_059_953, w_059_955, w_059_956, w_059_957, w_059_958, w_059_959, w_059_962, w_059_963, w_059_964, w_059_965, w_059_966, w_059_968, w_059_969, w_059_970, w_059_971, w_059_972, w_059_974, w_059_975, w_059_976, w_059_977, w_059_979, w_059_982, w_059_983, w_059_985, w_059_986, w_059_987, w_059_989, w_059_990, w_059_991, w_059_992, w_059_995, w_059_996, w_059_998, w_059_999, w_059_1000, w_059_1001, w_059_1002, w_059_1003, w_059_1005, w_059_1006, w_059_1007, w_059_1008, w_059_1010, w_059_1012, w_059_1013, w_059_1014, w_059_1015, w_059_1016, w_059_1017, w_059_1018, w_059_1019, w_059_1020, w_059_1022, w_059_1023, w_059_1026, w_059_1028, w_059_1029, w_059_1030, w_059_1031, w_059_1032, w_059_1033, w_059_1034, w_059_1035, w_059_1037, w_059_1039, w_059_1040, w_059_1041, w_059_1042, w_059_1043, w_059_1044, w_059_1045, w_059_1046, w_059_1048, w_059_1049, w_059_1050, w_059_1051, w_059_1053, w_059_1055, w_059_1056, w_059_1057, w_059_1058, w_059_1060, w_059_1061, w_059_1062, w_059_1063, w_059_1064, w_059_1065, w_059_1066, w_059_1067, w_059_1069, w_059_1073, w_059_1074, w_059_1075, w_059_1077, w_059_1078, w_059_1079, w_059_1080, w_059_1082, w_059_1083, w_059_1084, w_059_1085, w_059_1086, w_059_1087, w_059_1088, w_059_1089, w_059_1090, w_059_1091, w_059_1093, w_059_1094, w_059_1095, w_059_1096, w_059_1097, w_059_1098, w_059_1100, w_059_1101, w_059_1102, w_059_1103, w_059_1104, w_059_1106, w_059_1107, w_059_1108, w_059_1109, w_059_1110, w_059_1111, w_059_1112, w_059_1113, w_059_1114, w_059_1115, w_059_1117, w_059_1118, w_059_1119, w_059_1120, w_059_1121, w_059_1122, w_059_1123, w_059_1124, w_059_1125, w_059_1127, w_059_1128, w_059_1129, w_059_1130, w_059_1131, w_059_1132, w_059_1133, w_059_1135, w_059_1136, w_059_1137, w_059_1139, w_059_1140, w_059_1142, w_059_1143, w_059_1144, w_059_1145, w_059_1146, w_059_1147, w_059_1148, w_059_1149, w_059_1150, w_059_1152, w_059_1153, w_059_1154, w_059_1155, w_059_1156, w_059_1157, w_059_1158, w_059_1159, w_059_1161, w_059_1162, w_059_1163, w_059_1166, w_059_1170, w_059_1171, w_059_1172, w_059_1173, w_059_1174, w_059_1175, w_059_1176, w_059_1177, w_059_1178, w_059_1179, w_059_1180, w_059_1182, w_059_1183, w_059_1184, w_059_1186, w_059_1187, w_059_1188, w_059_1190, w_059_1191, w_059_1192, w_059_1193, w_059_1195, w_059_1196, w_059_1197, w_059_1198, w_059_1199, w_059_1200, w_059_1201, w_059_1203, w_059_1204, w_059_1205, w_059_1208, w_059_1209, w_059_1210, w_059_1211, w_059_1213, w_059_1214, w_059_1215, w_059_1216, w_059_1218, w_059_1219, w_059_1221, w_059_1222, w_059_1223, w_059_1224, w_059_1225, w_059_1229, w_059_1230, w_059_1231, w_059_1233, w_059_1234, w_059_1236, w_059_1237, w_059_1239, w_059_1240, w_059_1241, w_059_1242, w_059_1244, w_059_1246, w_059_1247, w_059_1248, w_059_1249, w_059_1250, w_059_1252, w_059_1253, w_059_1254, w_059_1255, w_059_1256, w_059_1257, w_059_1259, w_059_1260, w_059_1261, w_059_1262, w_059_1263, w_059_1264, w_059_1265, w_059_1266, w_059_1267, w_059_1268, w_059_1269, w_059_1270, w_059_1271, w_059_1272, w_059_1273, w_059_1274, w_059_1275, w_059_1277, w_059_1278, w_059_1280, w_059_1281, w_059_1282, w_059_1283, w_059_1284, w_059_1285, w_059_1286, w_059_1288, w_059_1289, w_059_1290, w_059_1291, w_059_1292, w_059_1293, w_059_1296, w_059_1297, w_059_1298, w_059_1300, w_059_1302, w_059_1303, w_059_1304, w_059_1305, w_059_1306, w_059_1307, w_059_1308, w_059_1309, w_059_1310, w_059_1311, w_059_1313, w_059_1314, w_059_1315, w_059_1316, w_059_1317, w_059_1318, w_059_1319, w_059_1320, w_059_1321, w_059_1322, w_059_1323, w_059_1324, w_059_1326, w_059_1327, w_059_1328, w_059_1330, w_059_1331, w_059_1333, w_059_1334, w_059_1335, w_059_1336, w_059_1337, w_059_1338, w_059_1339, w_059_1341, w_059_1342, w_059_1343, w_059_1344, w_059_1345, w_059_1346, w_059_1347, w_059_1348, w_059_1349, w_059_1350, w_059_1351, w_059_1352, w_059_1353, w_059_1354, w_059_1355, w_059_1357, w_059_1358, w_059_1360, w_059_1362, w_059_1363, w_059_1364, w_059_1365, w_059_1367, w_059_1370, w_059_1371, w_059_1372, w_059_1373, w_059_1375, w_059_1376, w_059_1377, w_059_1378, w_059_1379, w_059_1380, w_059_1381, w_059_1382, w_059_1384, w_059_1385, w_059_1386, w_059_1387, w_059_1389, w_059_1390, w_059_1391, w_059_1392, w_059_1393, w_059_1394, w_059_1395, w_059_1396, w_059_1397, w_059_1399, w_059_1400, w_059_1401, w_059_1402, w_059_1403, w_059_1404, w_059_1405, w_059_1406, w_059_1407, w_059_1408, w_059_1409, w_059_1411, w_059_1413, w_059_1414, w_059_1415, w_059_1416, w_059_1417, w_059_1418, w_059_1419, w_059_1420, w_059_1421, w_059_1422, w_059_1424, w_059_1426, w_059_1427, w_059_1428, w_059_1429, w_059_1430, w_059_1432, w_059_1433, w_059_1435, w_059_1436, w_059_1438, w_059_1440, w_059_1442, w_059_1443, w_059_1444, w_059_1445, w_059_1446, w_059_1449, w_059_1451, w_059_1452, w_059_1453, w_059_1454, w_059_1455, w_059_1456, w_059_1457, w_059_1458, w_059_1459, w_059_1462, w_059_1463, w_059_1468, w_059_1469, w_059_1470, w_059_1471, w_059_1472, w_059_1473, w_059_1474, w_059_1475, w_059_1476, w_059_1478, w_059_1481, w_059_1482, w_059_1483, w_059_1485, w_059_1486, w_059_1487, w_059_1488, w_059_1489, w_059_1490, w_059_1491, w_059_1493, w_059_1494, w_059_1496, w_059_1497, w_059_1499, w_059_1500, w_059_1502, w_059_1503, w_059_1504, w_059_1505, w_059_1506, w_059_1507, w_059_1508, w_059_1509, w_059_1510, w_059_1511, w_059_1514, w_059_1515, w_059_1516, w_059_1517, w_059_1518, w_059_1519, w_059_1522, w_059_1523, w_059_1524, w_059_1525, w_059_1528, w_059_1529, w_059_1530, w_059_1531, w_059_1532, w_059_1533, w_059_1536, w_059_1537, w_059_1539, w_059_1540, w_059_1541, w_059_1542, w_059_1544, w_059_1546, w_059_1548, w_059_1550, w_059_1551, w_059_1552, w_059_1553, w_059_1556, w_059_1557, w_059_1558, w_059_1559, w_059_1561, w_059_1562, w_059_1564, w_059_1565, w_059_1566, w_059_1567, w_059_1569, w_059_1572, w_059_1573, w_059_1574, w_059_1576, w_059_1577, w_059_1579, w_059_1580, w_059_1582, w_059_1583, w_059_1584, w_059_1586, w_059_1587, w_059_1588, w_059_1589, w_059_1590, w_059_1592, w_059_1595, w_059_1598, w_059_1599, w_059_1600, w_059_1601, w_059_1602, w_059_1604, w_059_1608, w_059_1609, w_059_1610, w_059_1611, w_059_1613, w_059_1615, w_059_1618, w_059_1619, w_059_1622, w_059_1624, w_059_1626, w_059_1628, w_059_1629, w_059_1630, w_059_1631, w_059_1632, w_059_1634, w_059_1636, w_059_1638, w_059_1640, w_059_1641, w_059_1642, w_059_1644, w_059_1646, w_059_1648, w_059_1649, w_059_1651, w_059_1652, w_059_1653, w_059_1657, w_059_1658, w_059_1660, w_059_1664, w_059_1665, w_059_1666, w_059_1667, w_059_1669, w_059_1672, w_059_1674, w_059_1675, w_059_1676, w_059_1678, w_059_1679, w_059_1680, w_059_1683, w_059_1684, w_059_1685, w_059_1688, w_059_1689, w_059_1690, w_059_1691, w_059_1692, w_059_1694, w_059_1695, w_059_1696, w_059_1697, w_059_1698, w_059_1700, w_059_1701, w_059_1703, w_059_1706, w_059_1711, w_059_1713, w_059_1716, w_059_1717, w_059_1718, w_059_1719, w_059_1720, w_059_1722, w_059_1723, w_059_1724, w_059_1725, w_059_1726, w_059_1729, w_059_1730, w_059_1732, w_059_1733, w_059_1735, w_059_1736, w_059_1737, w_059_1738, w_059_1739, w_059_1740, w_059_1741, w_059_1743, w_059_1745, w_059_1746, w_059_1747, w_059_1748, w_059_1749, w_059_1750, w_059_1751, w_059_1752, w_059_1753;
  wire w_060_000, w_060_003, w_060_004, w_060_005, w_060_007, w_060_008, w_060_010, w_060_011, w_060_013, w_060_014, w_060_015, w_060_016, w_060_017, w_060_019, w_060_020, w_060_021, w_060_022, w_060_023, w_060_024, w_060_025, w_060_026, w_060_027, w_060_029, w_060_031, w_060_032, w_060_033, w_060_035, w_060_037, w_060_038, w_060_039, w_060_041, w_060_042, w_060_043, w_060_044, w_060_045, w_060_046, w_060_047, w_060_048, w_060_049, w_060_051, w_060_052, w_060_053, w_060_055, w_060_057, w_060_059, w_060_060, w_060_061, w_060_063, w_060_064, w_060_065, w_060_066, w_060_067, w_060_068, w_060_069, w_060_070, w_060_072, w_060_073, w_060_074, w_060_076, w_060_077, w_060_078, w_060_079, w_060_080, w_060_082, w_060_083, w_060_084, w_060_085, w_060_087, w_060_088, w_060_089, w_060_090, w_060_091, w_060_092, w_060_095, w_060_097, w_060_098, w_060_099, w_060_101, w_060_102, w_060_103, w_060_104, w_060_105, w_060_108, w_060_109, w_060_110, w_060_111, w_060_112, w_060_113, w_060_114, w_060_116, w_060_117, w_060_118, w_060_119, w_060_120, w_060_122, w_060_123, w_060_124, w_060_126, w_060_128, w_060_130, w_060_131, w_060_132, w_060_133, w_060_134, w_060_135, w_060_137, w_060_138, w_060_139, w_060_140, w_060_141, w_060_142, w_060_143, w_060_144, w_060_146, w_060_147, w_060_148, w_060_149, w_060_150, w_060_151, w_060_152, w_060_153, w_060_154, w_060_156, w_060_157, w_060_160, w_060_161, w_060_162, w_060_163, w_060_164, w_060_165, w_060_166, w_060_168, w_060_169, w_060_170, w_060_171, w_060_172, w_060_173, w_060_174, w_060_175, w_060_177, w_060_179, w_060_181, w_060_182, w_060_183, w_060_184, w_060_185, w_060_186, w_060_188, w_060_189, w_060_190, w_060_191, w_060_192, w_060_193, w_060_195, w_060_196, w_060_197, w_060_198, w_060_199, w_060_200, w_060_201, w_060_202, w_060_203, w_060_204, w_060_205, w_060_207, w_060_208, w_060_209, w_060_210, w_060_211, w_060_212, w_060_213, w_060_214, w_060_215, w_060_216, w_060_217, w_060_218, w_060_219, w_060_220, w_060_221, w_060_222, w_060_223, w_060_224, w_060_225, w_060_228, w_060_229, w_060_230, w_060_232, w_060_233, w_060_234, w_060_236, w_060_237, w_060_238, w_060_239, w_060_241, w_060_243, w_060_245, w_060_246, w_060_247, w_060_248, w_060_249, w_060_250, w_060_251, w_060_252, w_060_253, w_060_254, w_060_255, w_060_256, w_060_258, w_060_259, w_060_261, w_060_264, w_060_265, w_060_266, w_060_267, w_060_268, w_060_270, w_060_271, w_060_272, w_060_273, w_060_275, w_060_276, w_060_277, w_060_279, w_060_281, w_060_282, w_060_283, w_060_284, w_060_285, w_060_286, w_060_287, w_060_288, w_060_289, w_060_290, w_060_291, w_060_295, w_060_296, w_060_297, w_060_298, w_060_300, w_060_301, w_060_302, w_060_303, w_060_305, w_060_306, w_060_307, w_060_308, w_060_309, w_060_312, w_060_313, w_060_314, w_060_315, w_060_316, w_060_318, w_060_319, w_060_320, w_060_321, w_060_322, w_060_323, w_060_324, w_060_325, w_060_326, w_060_328, w_060_329, w_060_330, w_060_331, w_060_333, w_060_334, w_060_335, w_060_336, w_060_337, w_060_338, w_060_339, w_060_340, w_060_341, w_060_342, w_060_345, w_060_346, w_060_347, w_060_348, w_060_349, w_060_350, w_060_351, w_060_353, w_060_354, w_060_356, w_060_357, w_060_358, w_060_359, w_060_360, w_060_362, w_060_364, w_060_365, w_060_366, w_060_367, w_060_369, w_060_370, w_060_371, w_060_372, w_060_373, w_060_376, w_060_378, w_060_379, w_060_381, w_060_382, w_060_383, w_060_385, w_060_386, w_060_389, w_060_390, w_060_391, w_060_392, w_060_393, w_060_394, w_060_395, w_060_396, w_060_397, w_060_398, w_060_399, w_060_400, w_060_402, w_060_403, w_060_404, w_060_405, w_060_406, w_060_407, w_060_408, w_060_409, w_060_410, w_060_411, w_060_413, w_060_414, w_060_415, w_060_416, w_060_417, w_060_418, w_060_419, w_060_422, w_060_423, w_060_424, w_060_425, w_060_426, w_060_427, w_060_429, w_060_430, w_060_431, w_060_433, w_060_434, w_060_435, w_060_436, w_060_437, w_060_438, w_060_439, w_060_440, w_060_441, w_060_443, w_060_444, w_060_445, w_060_446, w_060_447, w_060_448, w_060_449, w_060_450, w_060_451, w_060_453, w_060_456, w_060_457, w_060_458, w_060_459, w_060_460, w_060_462, w_060_464, w_060_466, w_060_467, w_060_468, w_060_470, w_060_471, w_060_472, w_060_473, w_060_475, w_060_476, w_060_477, w_060_478, w_060_481, w_060_482, w_060_483, w_060_484, w_060_485, w_060_486, w_060_488, w_060_490, w_060_491, w_060_492, w_060_493, w_060_494, w_060_496, w_060_497, w_060_498, w_060_499, w_060_500, w_060_501, w_060_502, w_060_503, w_060_505, w_060_510, w_060_511, w_060_512, w_060_513, w_060_514, w_060_515, w_060_516, w_060_517, w_060_518, w_060_519, w_060_520, w_060_521, w_060_522, w_060_523, w_060_524, w_060_525, w_060_526, w_060_528, w_060_529, w_060_530, w_060_531, w_060_532, w_060_533, w_060_534, w_060_535, w_060_537, w_060_539, w_060_540, w_060_541, w_060_542, w_060_543, w_060_544, w_060_545, w_060_546, w_060_547, w_060_548, w_060_550, w_060_551, w_060_553, w_060_554, w_060_555, w_060_556, w_060_557, w_060_559, w_060_560, w_060_562, w_060_563, w_060_564, w_060_565, w_060_566, w_060_567, w_060_568, w_060_569, w_060_570, w_060_571, w_060_572, w_060_573, w_060_576, w_060_577, w_060_578, w_060_579, w_060_580, w_060_581, w_060_582, w_060_583, w_060_584, w_060_585, w_060_586, w_060_587, w_060_588, w_060_589, w_060_591, w_060_592, w_060_593, w_060_595, w_060_596, w_060_597, w_060_598, w_060_599, w_060_600, w_060_602, w_060_603, w_060_604, w_060_607, w_060_608, w_060_609, w_060_610, w_060_611, w_060_612, w_060_614, w_060_615, w_060_616, w_060_618, w_060_619, w_060_621, w_060_622, w_060_623, w_060_625, w_060_628, w_060_629, w_060_630, w_060_631, w_060_632, w_060_633, w_060_634, w_060_635, w_060_636, w_060_637, w_060_638, w_060_639, w_060_640, w_060_642, w_060_644, w_060_646, w_060_648, w_060_649, w_060_650, w_060_651, w_060_652, w_060_653, w_060_654, w_060_655, w_060_656, w_060_657, w_060_658, w_060_659, w_060_660, w_060_662, w_060_665, w_060_666, w_060_667, w_060_668, w_060_669, w_060_671, w_060_673, w_060_674, w_060_675, w_060_676, w_060_677, w_060_678, w_060_679, w_060_680, w_060_683, w_060_684, w_060_685, w_060_686, w_060_687, w_060_689, w_060_690, w_060_691, w_060_693, w_060_694, w_060_695, w_060_697, w_060_698, w_060_699, w_060_700, w_060_701, w_060_702, w_060_703, w_060_704, w_060_705, w_060_707, w_060_708, w_060_709, w_060_710, w_060_711, w_060_713, w_060_714, w_060_715, w_060_716, w_060_719, w_060_720, w_060_721, w_060_722, w_060_723, w_060_724, w_060_725, w_060_727, w_060_728, w_060_729, w_060_731, w_060_734, w_060_736, w_060_737, w_060_739, w_060_740, w_060_741, w_060_743, w_060_744, w_060_745, w_060_746, w_060_747, w_060_748, w_060_749, w_060_750, w_060_752, w_060_753, w_060_754, w_060_755, w_060_758, w_060_759, w_060_760, w_060_761, w_060_762, w_060_763, w_060_764, w_060_765, w_060_766, w_060_767, w_060_768, w_060_769, w_060_770, w_060_771, w_060_772, w_060_773, w_060_775, w_060_777, w_060_778, w_060_779, w_060_780, w_060_781, w_060_782, w_060_783, w_060_784, w_060_785, w_060_786, w_060_787, w_060_789, w_060_790, w_060_791, w_060_792, w_060_793, w_060_794, w_060_795, w_060_796, w_060_797, w_060_798, w_060_799, w_060_800, w_060_801, w_060_802, w_060_803, w_060_804, w_060_805, w_060_806, w_060_807, w_060_808, w_060_809, w_060_810, w_060_811, w_060_812, w_060_813, w_060_815, w_060_817, w_060_818, w_060_819, w_060_821, w_060_822, w_060_823, w_060_824, w_060_825, w_060_827, w_060_828, w_060_829, w_060_830, w_060_831, w_060_832, w_060_833, w_060_834, w_060_835, w_060_836, w_060_840, w_060_842, w_060_845, w_060_847, w_060_848, w_060_849, w_060_850, w_060_851, w_060_852, w_060_853, w_060_854, w_060_855, w_060_857, w_060_858, w_060_859, w_060_860, w_060_861, w_060_862, w_060_863, w_060_864, w_060_865, w_060_866, w_060_867, w_060_870, w_060_871, w_060_872, w_060_873, w_060_874, w_060_876, w_060_877, w_060_878, w_060_879, w_060_880, w_060_881, w_060_883, w_060_885, w_060_887, w_060_888, w_060_890, w_060_891, w_060_892, w_060_893, w_060_894, w_060_895, w_060_896, w_060_897, w_060_898, w_060_899, w_060_900, w_060_901, w_060_903, w_060_905, w_060_906, w_060_907, w_060_909, w_060_910, w_060_912, w_060_913, w_060_914, w_060_915, w_060_916, w_060_917, w_060_918, w_060_919, w_060_920, w_060_921, w_060_922, w_060_923, w_060_924, w_060_927, w_060_930, w_060_931, w_060_932, w_060_933, w_060_934, w_060_935, w_060_937, w_060_938, w_060_939, w_060_940, w_060_941, w_060_942, w_060_944, w_060_945, w_060_946, w_060_947, w_060_949, w_060_950, w_060_951, w_060_952, w_060_953, w_060_954, w_060_955, w_060_956, w_060_957, w_060_958, w_060_960, w_060_961, w_060_962, w_060_963, w_060_964, w_060_965, w_060_966, w_060_967, w_060_968, w_060_969, w_060_970, w_060_971, w_060_972, w_060_973, w_060_974, w_060_975, w_060_976, w_060_978, w_060_979, w_060_980, w_060_981, w_060_982, w_060_984, w_060_986, w_060_987, w_060_988, w_060_990, w_060_991, w_060_992, w_060_994, w_060_995, w_060_997, w_060_998, w_060_999, w_060_1000, w_060_1001, w_060_1002, w_060_1003, w_060_1005, w_060_1008, w_060_1009, w_060_1010, w_060_1011, w_060_1012, w_060_1013, w_060_1014, w_060_1015, w_060_1016, w_060_1017, w_060_1018, w_060_1019, w_060_1020, w_060_1022, w_060_1023, w_060_1024, w_060_1025, w_060_1026, w_060_1027, w_060_1028, w_060_1030, w_060_1031, w_060_1032, w_060_1033, w_060_1034, w_060_1035, w_060_1036, w_060_1038, w_060_1040, w_060_1042, w_060_1043, w_060_1044, w_060_1045, w_060_1046, w_060_1047, w_060_1048, w_060_1049, w_060_1050, w_060_1053, w_060_1054, w_060_1055, w_060_1056, w_060_1057, w_060_1059, w_060_1060, w_060_1061, w_060_1063, w_060_1064, w_060_1065, w_060_1067, w_060_1069, w_060_1070, w_060_1071, w_060_1073, w_060_1074, w_060_1075, w_060_1076, w_060_1077, w_060_1078, w_060_1079, w_060_1080, w_060_1081, w_060_1082, w_060_1083, w_060_1084, w_060_1086, w_060_1087, w_060_1088, w_060_1089, w_060_1090, w_060_1091, w_060_1092, w_060_1093, w_060_1094, w_060_1096, w_060_1097, w_060_1098, w_060_1099, w_060_1101, w_060_1102, w_060_1103, w_060_1105, w_060_1107, w_060_1108, w_060_1109, w_060_1110, w_060_1114, w_060_1115, w_060_1116, w_060_1117, w_060_1118, w_060_1119, w_060_1120, w_060_1122, w_060_1123, w_060_1124, w_060_1126, w_060_1127, w_060_1128, w_060_1129, w_060_1130, w_060_1131, w_060_1132, w_060_1133, w_060_1134, w_060_1135, w_060_1136, w_060_1140, w_060_1143, w_060_1144, w_060_1145, w_060_1146, w_060_1149, w_060_1150, w_060_1151, w_060_1154, w_060_1155, w_060_1157, w_060_1159, w_060_1160, w_060_1161, w_060_1163, w_060_1165, w_060_1167, w_060_1168, w_060_1169, w_060_1173, w_060_1174, w_060_1175, w_060_1176, w_060_1177, w_060_1180, w_060_1181, w_060_1184, w_060_1185, w_060_1186, w_060_1189, w_060_1191, w_060_1192, w_060_1193, w_060_1194, w_060_1195, w_060_1196, w_060_1197, w_060_1198, w_060_1200, w_060_1203, w_060_1206, w_060_1208, w_060_1210, w_060_1211, w_060_1212, w_060_1213, w_060_1214, w_060_1216, w_060_1217, w_060_1218, w_060_1219, w_060_1221, w_060_1222, w_060_1223, w_060_1225, w_060_1226, w_060_1227, w_060_1230, w_060_1232, w_060_1233, w_060_1234, w_060_1235, w_060_1236, w_060_1238, w_060_1239, w_060_1240, w_060_1242, w_060_1244, w_060_1245, w_060_1246, w_060_1247, w_060_1248, w_060_1249, w_060_1250, w_060_1251, w_060_1252, w_060_1254, w_060_1255, w_060_1256, w_060_1257, w_060_1259, w_060_1261, w_060_1262, w_060_1264, w_060_1265, w_060_1266, w_060_1270, w_060_1271, w_060_1273, w_060_1274, w_060_1276, w_060_1278, w_060_1279, w_060_1280, w_060_1281, w_060_1283, w_060_1284, w_060_1285, w_060_1286, w_060_1287, w_060_1292, w_060_1293, w_060_1296, w_060_1299, w_060_1300, w_060_1301, w_060_1302, w_060_1303, w_060_1305, w_060_1306, w_060_1308, w_060_1309, w_060_1310, w_060_1311, w_060_1313, w_060_1314, w_060_1315, w_060_1318, w_060_1319, w_060_1320, w_060_1322, w_060_1323, w_060_1324, w_060_1327, w_060_1330, w_060_1333, w_060_1334, w_060_1335, w_060_1336, w_060_1337, w_060_1338, w_060_1340, w_060_1341, w_060_1342, w_060_1343, w_060_1344, w_060_1345, w_060_1346, w_060_1348, w_060_1349, w_060_1350, w_060_1351, w_060_1352, w_060_1353, w_060_1356, w_060_1359, w_060_1361, w_060_1362, w_060_1363, w_060_1364, w_060_1365, w_060_1367, w_060_1370, w_060_1371, w_060_1372, w_060_1373, w_060_1374, w_060_1375, w_060_1377, w_060_1380, w_060_1381, w_060_1382, w_060_1383, w_060_1384, w_060_1385, w_060_1386, w_060_1388, w_060_1390, w_060_1391, w_060_1392, w_060_1394, w_060_1398, w_060_1399, w_060_1400, w_060_1401, w_060_1402, w_060_1403, w_060_1406, w_060_1408, w_060_1409, w_060_1413, w_060_1415, w_060_1416, w_060_1417, w_060_1418, w_060_1419, w_060_1421, w_060_1424, w_060_1426, w_060_1428, w_060_1429, w_060_1430, w_060_1432, w_060_1433, w_060_1434, w_060_1436, w_060_1437, w_060_1438, w_060_1441, w_060_1442, w_060_1445, w_060_1446, w_060_1450, w_060_1451, w_060_1452, w_060_1454, w_060_1455, w_060_1456, w_060_1457, w_060_1459, w_060_1462, w_060_1463, w_060_1464, w_060_1465, w_060_1466, w_060_1467, w_060_1468, w_060_1469, w_060_1471, w_060_1472, w_060_1473, w_060_1475, w_060_1477, w_060_1478, w_060_1479, w_060_1480, w_060_1482, w_060_1484, w_060_1488, w_060_1490, w_060_1491, w_060_1492, w_060_1493, w_060_1495, w_060_1496, w_060_1497, w_060_1498, w_060_1499, w_060_1500, w_060_1502, w_060_1503, w_060_1505, w_060_1506, w_060_1509, w_060_1510, w_060_1512, w_060_1515, w_060_1516, w_060_1517, w_060_1518, w_060_1519, w_060_1520, w_060_1523, w_060_1524, w_060_1526, w_060_1528, w_060_1532, w_060_1534, w_060_1535, w_060_1537, w_060_1538, w_060_1539, w_060_1543, w_060_1544, w_060_1545, w_060_1546, w_060_1547, w_060_1548, w_060_1549, w_060_1550, w_060_1552, w_060_1555, w_060_1556, w_060_1558, w_060_1561, w_060_1562, w_060_1564, w_060_1565, w_060_1567, w_060_1568, w_060_1569, w_060_1570, w_060_1572, w_060_1574, w_060_1575, w_060_1577, w_060_1578, w_060_1579, w_060_1580, w_060_1581, w_060_1582, w_060_1584, w_060_1586, w_060_1587, w_060_1589, w_060_1590, w_060_1592, w_060_1593, w_060_1595, w_060_1596, w_060_1597, w_060_1599, w_060_1600, w_060_1604, w_060_1606, w_060_1607, w_060_1609, w_060_1610, w_060_1611, w_060_1614, w_060_1615, w_060_1616, w_060_1617, w_060_1618, w_060_1619, w_060_1620, w_060_1621, w_060_1622, w_060_1623, w_060_1624, w_060_1627, w_060_1629, w_060_1630, w_060_1631, w_060_1633, w_060_1634, w_060_1635, w_060_1637, w_060_1638, w_060_1640, w_060_1642, w_060_1644, w_060_1645, w_060_1647, w_060_1649, w_060_1650, w_060_1652, w_060_1653, w_060_1658, w_060_1659, w_060_1661, w_060_1663, w_060_1664, w_060_1667, w_060_1669, w_060_1671, w_060_1672, w_060_1675, w_060_1677, w_060_1678, w_060_1679, w_060_1680, w_060_1681, w_060_1682, w_060_1683, w_060_1684, w_060_1685, w_060_1686, w_060_1688, w_060_1689, w_060_1690, w_060_1691, w_060_1693, w_060_1697, w_060_1699, w_060_1700, w_060_1701, w_060_1702, w_060_1703, w_060_1704, w_060_1705, w_060_1706, w_060_1708, w_060_1709, w_060_1710, w_060_1711, w_060_1713, w_060_1714, w_060_1717, w_060_1718, w_060_1719, w_060_1720, w_060_1722, w_060_1723, w_060_1724, w_060_1727, w_060_1730, w_060_1732, w_060_1734, w_060_1735, w_060_1738, w_060_1739, w_060_1742, w_060_1743, w_060_1744, w_060_1747, w_060_1750, w_060_1752, w_060_1753, w_060_1755, w_060_1756, w_060_1758, w_060_1759, w_060_1761, w_060_1764, w_060_1765, w_060_1766, w_060_1767, w_060_1768, w_060_1770, w_060_1773, w_060_1775, w_060_1777, w_060_1778, w_060_1779, w_060_1781, w_060_1782, w_060_1783, w_060_1784, w_060_1786, w_060_1792, w_060_1794, w_060_1795, w_060_1796, w_060_1799, w_060_1801, w_060_1802, w_060_1805, w_060_1806, w_060_1808, w_060_1809, w_060_1811, w_060_1813, w_060_1814, w_060_1815, w_060_1816, w_060_1817, w_060_1818, w_060_1819, w_060_1821, w_060_1822, w_060_1823, w_060_1824, w_060_1828, w_060_1829, w_060_1831, w_060_1833, w_060_1834, w_060_1835, w_060_1836, w_060_1839, w_060_1841, w_060_1842, w_060_1845, w_060_1846, w_060_1847, w_060_1848, w_060_1849, w_060_1850, w_060_1851, w_060_1852, w_060_1853, w_060_1858, w_060_1859, w_060_1860, w_060_1861, w_060_1862, w_060_1863, w_060_1865, w_060_1867, w_060_1870, w_060_1872, w_060_1874, w_060_1875, w_060_1876, w_060_1877, w_060_1878, w_060_1879, w_060_1880, w_060_1881, w_060_1882, w_060_1883, w_060_1886, w_060_1887, w_060_1889, w_060_1890, w_060_1891, w_060_1893, w_060_1894, w_060_1895, w_060_1896, w_060_1897, w_060_1898, w_060_1899, w_060_1900, w_060_1901, w_060_1903, w_060_1905, w_060_1906, w_060_1907, w_060_1908, w_060_1910, w_060_1911, w_060_1912, w_060_1915, w_060_1918, w_060_1919, w_060_1921, w_060_1922, w_060_1923, w_060_1924, w_060_1926, w_060_1927, w_060_1928, w_060_1930, w_060_1931, w_060_1932, w_060_1933, w_060_1937, w_060_1940, w_060_1941, w_060_1945, w_060_1946, w_060_1947, w_060_1948, w_060_1949;
  wire w_061_002, w_061_003, w_061_004, w_061_005, w_061_007, w_061_008, w_061_010, w_061_011, w_061_012, w_061_014, w_061_015, w_061_017, w_061_019, w_061_020, w_061_022, w_061_023, w_061_024, w_061_025, w_061_029, w_061_030, w_061_032, w_061_033, w_061_034, w_061_035, w_061_036, w_061_037, w_061_038, w_061_039, w_061_041, w_061_042, w_061_045, w_061_046, w_061_049, w_061_050, w_061_053, w_061_054, w_061_055, w_061_057, w_061_059, w_061_060, w_061_061, w_061_062, w_061_063, w_061_064, w_061_065, w_061_066, w_061_067, w_061_069, w_061_071, w_061_072, w_061_073, w_061_074, w_061_075, w_061_076, w_061_078, w_061_079, w_061_081, w_061_082, w_061_083, w_061_085, w_061_086, w_061_088, w_061_090, w_061_091, w_061_092, w_061_094, w_061_096, w_061_097, w_061_098, w_061_099, w_061_100, w_061_101, w_061_103, w_061_104, w_061_106, w_061_107, w_061_108, w_061_110, w_061_111, w_061_112, w_061_113, w_061_114, w_061_116, w_061_118, w_061_119, w_061_122, w_061_123, w_061_124, w_061_125, w_061_126, w_061_127, w_061_128, w_061_129, w_061_130, w_061_131, w_061_132, w_061_133, w_061_134, w_061_135, w_061_136, w_061_138, w_061_141, w_061_142, w_061_144, w_061_145, w_061_147, w_061_148, w_061_149, w_061_150, w_061_151, w_061_152, w_061_153, w_061_154, w_061_156, w_061_158, w_061_159, w_061_160, w_061_161, w_061_162, w_061_163, w_061_164, w_061_165, w_061_166, w_061_167, w_061_168, w_061_169, w_061_171, w_061_172, w_061_173, w_061_174, w_061_175, w_061_176, w_061_177, w_061_178, w_061_180, w_061_181, w_061_182, w_061_187, w_061_188, w_061_189, w_061_190, w_061_193, w_061_194, w_061_195, w_061_197, w_061_198, w_061_200, w_061_202, w_061_203, w_061_205, w_061_206, w_061_207, w_061_208, w_061_210, w_061_211, w_061_212, w_061_214, w_061_215, w_061_216, w_061_217, w_061_218, w_061_219, w_061_221, w_061_222, w_061_223, w_061_224, w_061_226, w_061_227, w_061_228, w_061_229, w_061_230, w_061_231, w_061_232, w_061_233, w_061_234, w_061_236, w_061_239, w_061_240, w_061_241, w_061_242, w_061_243, w_061_244, w_061_245, w_061_246, w_061_248, w_061_249, w_061_250, w_061_251, w_061_252, w_061_253, w_061_255, w_061_256, w_061_257, w_061_258, w_061_259, w_061_261, w_061_262, w_061_263, w_061_265, w_061_266, w_061_267, w_061_270, w_061_271, w_061_272, w_061_273, w_061_275, w_061_277, w_061_281, w_061_282, w_061_284, w_061_285, w_061_287, w_061_289, w_061_292, w_061_293, w_061_294, w_061_295, w_061_296, w_061_297, w_061_299, w_061_300, w_061_302, w_061_304, w_061_305, w_061_306, w_061_307, w_061_308, w_061_309, w_061_310, w_061_312, w_061_313, w_061_314, w_061_315, w_061_316, w_061_317, w_061_318, w_061_319, w_061_320, w_061_321, w_061_322, w_061_323, w_061_324, w_061_325, w_061_326, w_061_329, w_061_330, w_061_331, w_061_332, w_061_333, w_061_334, w_061_335, w_061_336, w_061_338, w_061_339, w_061_340, w_061_341, w_061_342, w_061_343, w_061_344, w_061_345, w_061_346, w_061_352, w_061_353, w_061_354, w_061_355, w_061_356, w_061_357, w_061_359, w_061_360, w_061_361, w_061_362, w_061_365, w_061_366, w_061_367, w_061_368, w_061_370, w_061_371, w_061_372, w_061_373, w_061_375, w_061_376, w_061_377, w_061_379, w_061_380, w_061_381, w_061_382, w_061_385, w_061_388, w_061_389, w_061_391, w_061_393, w_061_394, w_061_395, w_061_396, w_061_398, w_061_399, w_061_400, w_061_401, w_061_402, w_061_404, w_061_405, w_061_406, w_061_407, w_061_409, w_061_410, w_061_412, w_061_413, w_061_414, w_061_415, w_061_416, w_061_418, w_061_420, w_061_421, w_061_423, w_061_425, w_061_426, w_061_427, w_061_428, w_061_429, w_061_432, w_061_435, w_061_436, w_061_438, w_061_439, w_061_440, w_061_442, w_061_443, w_061_444, w_061_445, w_061_446, w_061_448, w_061_451, w_061_452, w_061_456, w_061_457, w_061_460, w_061_461, w_061_462, w_061_463, w_061_464, w_061_465, w_061_468, w_061_469, w_061_470, w_061_471, w_061_473, w_061_474, w_061_475, w_061_476, w_061_478, w_061_480, w_061_481, w_061_482, w_061_483, w_061_484, w_061_486, w_061_487, w_061_491, w_061_492, w_061_493, w_061_495, w_061_497, w_061_498, w_061_499, w_061_500, w_061_501, w_061_502, w_061_503, w_061_504, w_061_505, w_061_506, w_061_507, w_061_508, w_061_509, w_061_510, w_061_513, w_061_514, w_061_515, w_061_516, w_061_517, w_061_518, w_061_521, w_061_522, w_061_524, w_061_527, w_061_528, w_061_529, w_061_531, w_061_532, w_061_537, w_061_538, w_061_539, w_061_546, w_061_547, w_061_548, w_061_549, w_061_550, w_061_551, w_061_552, w_061_553, w_061_554, w_061_555, w_061_556, w_061_559, w_061_561, w_061_563, w_061_564, w_061_565, w_061_566, w_061_567, w_061_569, w_061_574, w_061_576, w_061_579, w_061_581, w_061_583, w_061_585, w_061_586, w_061_587, w_061_588, w_061_589, w_061_594, w_061_595, w_061_596, w_061_598, w_061_599, w_061_600, w_061_601, w_061_602, w_061_605, w_061_607, w_061_609, w_061_611, w_061_613, w_061_615, w_061_618, w_061_619, w_061_620, w_061_621, w_061_624, w_061_625, w_061_627, w_061_630, w_061_631, w_061_633, w_061_635, w_061_636, w_061_637, w_061_638, w_061_639, w_061_641, w_061_642, w_061_643, w_061_644, w_061_646, w_061_647, w_061_651, w_061_652, w_061_654, w_061_655, w_061_656, w_061_657, w_061_659, w_061_660, w_061_663, w_061_664, w_061_665, w_061_666, w_061_667, w_061_669, w_061_671, w_061_672, w_061_673, w_061_674, w_061_675, w_061_677, w_061_679, w_061_680, w_061_683, w_061_685, w_061_687, w_061_688, w_061_689, w_061_690, w_061_692, w_061_693, w_061_694, w_061_695, w_061_698, w_061_700, w_061_701, w_061_705, w_061_706, w_061_708, w_061_711, w_061_716, w_061_717, w_061_719, w_061_721, w_061_722, w_061_724, w_061_725, w_061_726, w_061_727, w_061_728, w_061_730, w_061_732, w_061_733, w_061_734, w_061_736, w_061_737, w_061_739, w_061_740, w_061_741, w_061_742, w_061_744, w_061_745, w_061_746, w_061_747, w_061_748, w_061_749, w_061_754, w_061_755, w_061_756, w_061_759, w_061_760, w_061_762, w_061_763, w_061_764, w_061_765, w_061_766, w_061_767, w_061_768, w_061_769, w_061_770, w_061_771, w_061_772, w_061_773, w_061_774, w_061_775, w_061_776, w_061_777, w_061_779, w_061_781, w_061_784, w_061_789, w_061_792, w_061_793, w_061_794, w_061_798, w_061_799, w_061_801, w_061_802, w_061_803, w_061_804, w_061_805, w_061_806, w_061_808, w_061_810, w_061_811, w_061_813, w_061_814, w_061_815, w_061_816, w_061_817, w_061_818, w_061_821, w_061_822, w_061_823, w_061_824, w_061_825, w_061_826, w_061_827, w_061_828, w_061_830, w_061_831, w_061_833, w_061_834, w_061_835, w_061_839, w_061_840, w_061_841, w_061_843, w_061_844, w_061_845, w_061_846, w_061_847, w_061_849, w_061_850, w_061_852, w_061_854, w_061_855, w_061_857, w_061_858, w_061_861, w_061_862, w_061_863, w_061_864, w_061_865, w_061_866, w_061_867, w_061_869, w_061_870, w_061_872, w_061_873, w_061_874, w_061_875, w_061_876, w_061_877, w_061_879, w_061_881, w_061_883, w_061_884, w_061_885, w_061_886, w_061_887, w_061_888, w_061_892, w_061_893, w_061_895, w_061_897, w_061_898, w_061_901, w_061_902, w_061_904, w_061_905, w_061_906, w_061_909, w_061_910, w_061_913, w_061_914, w_061_915, w_061_917, w_061_921, w_061_922, w_061_923, w_061_924, w_061_932, w_061_934, w_061_936, w_061_937, w_061_938, w_061_940, w_061_942, w_061_943, w_061_945, w_061_946, w_061_947, w_061_948, w_061_949, w_061_950, w_061_951, w_061_953, w_061_954, w_061_955, w_061_956, w_061_957, w_061_960, w_061_961, w_061_962, w_061_963, w_061_964, w_061_966, w_061_967, w_061_969, w_061_970, w_061_971, w_061_972, w_061_973, w_061_974, w_061_975, w_061_976, w_061_977, w_061_978, w_061_979, w_061_980, w_061_981, w_061_983, w_061_985, w_061_988, w_061_989, w_061_991, w_061_992, w_061_995, w_061_996, w_061_997, w_061_998, w_061_999, w_061_1000, w_061_1001, w_061_1003, w_061_1004, w_061_1006, w_061_1007, w_061_1009, w_061_1010, w_061_1011, w_061_1012, w_061_1014, w_061_1016, w_061_1019, w_061_1022, w_061_1025, w_061_1026, w_061_1028, w_061_1029, w_061_1030, w_061_1035, w_061_1038, w_061_1039, w_061_1040, w_061_1041, w_061_1042, w_061_1044, w_061_1046, w_061_1048, w_061_1050, w_061_1051, w_061_1053, w_061_1054, w_061_1057, w_061_1059, w_061_1061, w_061_1062, w_061_1063, w_061_1064, w_061_1065, w_061_1067, w_061_1068, w_061_1069, w_061_1070, w_061_1071, w_061_1072, w_061_1073, w_061_1074, w_061_1075, w_061_1077, w_061_1078, w_061_1079, w_061_1080, w_061_1081, w_061_1082, w_061_1083, w_061_1084, w_061_1085, w_061_1086, w_061_1087, w_061_1092, w_061_1095, w_061_1096, w_061_1097, w_061_1098, w_061_1099, w_061_1101, w_061_1105, w_061_1106, w_061_1107, w_061_1108, w_061_1109, w_061_1110, w_061_1111, w_061_1112, w_061_1116, w_061_1117, w_061_1118, w_061_1121, w_061_1124, w_061_1125, w_061_1126, w_061_1128, w_061_1130, w_061_1131, w_061_1134, w_061_1135, w_061_1137, w_061_1140, w_061_1141, w_061_1142, w_061_1143, w_061_1144, w_061_1146, w_061_1148, w_061_1150, w_061_1151, w_061_1152, w_061_1153, w_061_1155, w_061_1157, w_061_1158, w_061_1159, w_061_1162, w_061_1163, w_061_1167, w_061_1171, w_061_1172, w_061_1173, w_061_1174, w_061_1175, w_061_1179, w_061_1180, w_061_1181, w_061_1182, w_061_1184, w_061_1186, w_061_1187, w_061_1188, w_061_1190, w_061_1191, w_061_1192, w_061_1193, w_061_1194, w_061_1198, w_061_1199, w_061_1200, w_061_1203, w_061_1204, w_061_1205, w_061_1206, w_061_1207, w_061_1212, w_061_1213, w_061_1214, w_061_1215, w_061_1216, w_061_1217, w_061_1218, w_061_1219, w_061_1224, w_061_1226, w_061_1227, w_061_1228, w_061_1232, w_061_1233, w_061_1234, w_061_1235, w_061_1236, w_061_1239, w_061_1240, w_061_1241, w_061_1244, w_061_1245, w_061_1246, w_061_1247, w_061_1248, w_061_1249, w_061_1251, w_061_1255, w_061_1256, w_061_1258, w_061_1259, w_061_1260, w_061_1261, w_061_1265, w_061_1266, w_061_1268, w_061_1270, w_061_1274, w_061_1275, w_061_1276, w_061_1277, w_061_1279, w_061_1280, w_061_1282, w_061_1287, w_061_1288, w_061_1289, w_061_1291, w_061_1292, w_061_1293, w_061_1294, w_061_1295, w_061_1296, w_061_1298, w_061_1300, w_061_1301, w_061_1302, w_061_1304, w_061_1305, w_061_1307, w_061_1308, w_061_1310, w_061_1311, w_061_1315, w_061_1319, w_061_1322, w_061_1324, w_061_1325, w_061_1326, w_061_1327, w_061_1328, w_061_1330, w_061_1331, w_061_1332, w_061_1333, w_061_1334, w_061_1335, w_061_1337, w_061_1338, w_061_1339, w_061_1340, w_061_1341, w_061_1347, w_061_1348, w_061_1349, w_061_1350, w_061_1353, w_061_1355, w_061_1356, w_061_1358, w_061_1359, w_061_1360, w_061_1361, w_061_1362, w_061_1364, w_061_1368, w_061_1369, w_061_1370, w_061_1372, w_061_1373, w_061_1374, w_061_1376, w_061_1377, w_061_1379, w_061_1380, w_061_1381, w_061_1382, w_061_1383, w_061_1384, w_061_1385, w_061_1387, w_061_1388, w_061_1390, w_061_1391, w_061_1392, w_061_1394, w_061_1395, w_061_1396, w_061_1397, w_061_1398, w_061_1399, w_061_1400, w_061_1403, w_061_1404, w_061_1405, w_061_1406, w_061_1409, w_061_1410, w_061_1411, w_061_1413, w_061_1414, w_061_1417, w_061_1418, w_061_1420, w_061_1421, w_061_1424, w_061_1428, w_061_1429, w_061_1434, w_061_1436, w_061_1437, w_061_1439, w_061_1441, w_061_1442, w_061_1443, w_061_1446, w_061_1447, w_061_1449, w_061_1450, w_061_1451, w_061_1455, w_061_1460, w_061_1461, w_061_1463, w_061_1466, w_061_1467, w_061_1468, w_061_1471, w_061_1472, w_061_1473, w_061_1474, w_061_1475, w_061_1477, w_061_1478, w_061_1480, w_061_1481, w_061_1482, w_061_1483, w_061_1485, w_061_1487, w_061_1488, w_061_1489, w_061_1490, w_061_1492, w_061_1493, w_061_1494, w_061_1495, w_061_1496, w_061_1497, w_061_1498, w_061_1499, w_061_1502, w_061_1503, w_061_1504, w_061_1505, w_061_1508, w_061_1510, w_061_1515, w_061_1516, w_061_1518, w_061_1520, w_061_1521, w_061_1523, w_061_1524, w_061_1525, w_061_1526, w_061_1527, w_061_1528, w_061_1529, w_061_1530, w_061_1533, w_061_1534, w_061_1536, w_061_1537, w_061_1538, w_061_1542, w_061_1544, w_061_1546, w_061_1550, w_061_1551, w_061_1552, w_061_1554, w_061_1555, w_061_1556, w_061_1557, w_061_1558, w_061_1559, w_061_1560, w_061_1562, w_061_1563, w_061_1565, w_061_1566, w_061_1567, w_061_1568, w_061_1571, w_061_1572, w_061_1573, w_061_1574, w_061_1577, w_061_1580, w_061_1581, w_061_1582, w_061_1583, w_061_1586, w_061_1587, w_061_1590, w_061_1591, w_061_1593, w_061_1594, w_061_1595, w_061_1596, w_061_1599, w_061_1601, w_061_1602, w_061_1603, w_061_1604, w_061_1605, w_061_1606, w_061_1607, w_061_1609, w_061_1611, w_061_1614, w_061_1615, w_061_1616, w_061_1617, w_061_1620, w_061_1622, w_061_1623, w_061_1625, w_061_1627, w_061_1628, w_061_1631, w_061_1633, w_061_1636, w_061_1638, w_061_1639, w_061_1642, w_061_1644, w_061_1647, w_061_1648, w_061_1649, w_061_1650, w_061_1654, w_061_1655, w_061_1656, w_061_1659, w_061_1661, w_061_1663, w_061_1664, w_061_1666, w_061_1668, w_061_1669, w_061_1671, w_061_1675, w_061_1680, w_061_1682, w_061_1684, w_061_1685, w_061_1686, w_061_1687, w_061_1688, w_061_1691, w_061_1692, w_061_1693, w_061_1694, w_061_1699, w_061_1700, w_061_1701, w_061_1703, w_061_1704, w_061_1706, w_061_1707, w_061_1709, w_061_1710, w_061_1711, w_061_1712, w_061_1713, w_061_1714, w_061_1715, w_061_1716, w_061_1717, w_061_1719, w_061_1720, w_061_1721, w_061_1722, w_061_1725, w_061_1726, w_061_1727, w_061_1728, w_061_1729, w_061_1730, w_061_1732, w_061_1733, w_061_1734, w_061_1735, w_061_1736, w_061_1737, w_061_1738, w_061_1739, w_061_1740, w_061_1741, w_061_1742, w_061_1743, w_061_1744, w_061_1747, w_061_1748, w_061_1749, w_061_1750, w_061_1751, w_061_1753, w_061_1755, w_061_1756, w_061_1761, w_061_1763, w_061_1765, w_061_1766, w_061_1767, w_061_1768, w_061_1769, w_061_1770, w_061_1773, w_061_1774, w_061_1775, w_061_1776, w_061_1777, w_061_1778, w_061_1779, w_061_1780, w_061_1781, w_061_1782, w_061_1785, w_061_1786, w_061_1787, w_061_1788, w_061_1789, w_061_1793, w_061_1795, w_061_1796, w_061_1797, w_061_1798, w_061_1799, w_061_1800, w_061_1803, w_061_1805, w_061_1806, w_061_1807, w_061_1809, w_061_1810, w_061_1812, w_061_1813, w_061_1814, w_061_1815, w_061_1816, w_061_1817, w_061_1820, w_061_1823, w_061_1824, w_061_1825, w_061_1827, w_061_1828, w_061_1831, w_061_1832, w_061_1833, w_061_1834, w_061_1835, w_061_1836, w_061_1838, w_061_1840, w_061_1841, w_061_1842, w_061_1843, w_061_1848, w_061_1851, w_061_1852, w_061_1854, w_061_1855, w_061_1856, w_061_1858, w_061_1859, w_061_1861, w_061_1864, w_061_1866, w_061_1867, w_061_1868, w_061_1869, w_061_1870, w_061_1871, w_061_1872, w_061_1874, w_061_1876, w_061_1877, w_061_1878, w_061_1879, w_061_1881, w_061_1885, w_061_1886, w_061_1887, w_061_1888, w_061_1891, w_061_1894, w_061_1896, w_061_1897, w_061_1899, w_061_1900, w_061_1901, w_061_1903, w_061_1904, w_061_1905, w_061_1906, w_061_1907, w_061_1908, w_061_1910, w_061_1911, w_061_1914, w_061_1916, w_061_1917, w_061_1918, w_061_1919, w_061_1921, w_061_1922, w_061_1924, w_061_1926, w_061_1927, w_061_1928, w_061_1929, w_061_1930, w_061_1931, w_061_1933, w_061_1934, w_061_1935, w_061_1936, w_061_1938, w_061_1940, w_061_1941, w_061_1942, w_061_1943, w_061_1944, w_061_1946, w_061_1949, w_061_1952, w_061_1953, w_061_1957, w_061_1960, w_061_1962, w_061_1964, w_061_1965, w_061_1967, w_061_1968, w_061_1969, w_061_1971, w_061_1972, w_061_1973, w_061_1974, w_061_1976, w_061_1977, w_061_1978, w_061_1980, w_061_1981, w_061_1982, w_061_1983, w_061_1986, w_061_1987, w_061_1990, w_061_1991, w_061_1992, w_061_1993, w_061_1994, w_061_1996, w_061_1997, w_061_1998, w_061_1999, w_061_2000, w_061_2002, w_061_2004, w_061_2005, w_061_2006, w_061_2007, w_061_2008, w_061_2010, w_061_2011, w_061_2012, w_061_2014, w_061_2017, w_061_2019, w_061_2023, w_061_2024, w_061_2025, w_061_2029, w_061_2031, w_061_2032, w_061_2033, w_061_2037, w_061_2040, w_061_2041, w_061_2042, w_061_2044, w_061_2045, w_061_2046, w_061_2048, w_061_2051, w_061_2053, w_061_2054, w_061_2056, w_061_2057, w_061_2059, w_061_2061, w_061_2062, w_061_2065, w_061_2067, w_061_2070, w_061_2071, w_061_2073, w_061_2075, w_061_2076, w_061_2077, w_061_2078, w_061_2079, w_061_2080, w_061_2083, w_061_2084, w_061_2085, w_061_2088, w_061_2091, w_061_2092, w_061_2093, w_061_2096, w_061_2098, w_061_2099, w_061_2101, w_061_2104, w_061_2105, w_061_2107, w_061_2110, w_061_2111, w_061_2112, w_061_2113, w_061_2114, w_061_2115, w_061_2116, w_061_2118, w_061_2120, w_061_2121, w_061_2122, w_061_2123, w_061_2124, w_061_2125, w_061_2126, w_061_2127, w_061_2130, w_061_2131, w_061_2133, w_061_2134, w_061_2135, w_061_2136, w_061_2140, w_061_2145, w_061_2146, w_061_2147, w_061_2148, w_061_2149, w_061_2150, w_061_2152, w_061_2155, w_061_2156, w_061_2158, w_061_2162, w_061_2163, w_061_2164, w_061_2165, w_061_2166, w_061_2167, w_061_2168, w_061_2169, w_061_2170, w_061_2171, w_061_2172, w_061_2173, w_061_2174, w_061_2176, w_061_2177, w_061_2179, w_061_2181, w_061_2182, w_061_2183, w_061_2184, w_061_2185, w_061_2187, w_061_2188, w_061_2189, w_061_2190, w_061_2193, w_061_2194, w_061_2195, w_061_2197, w_061_2198, w_061_2199, w_061_2200, w_061_2201, w_061_2202, w_061_2203, w_061_2205, w_061_2207, w_061_2208, w_061_2210, w_061_2211, w_061_2214, w_061_2215, w_061_2219, w_061_2220, w_061_2226, w_061_2227, w_061_2228, w_061_2229, w_061_2230, w_061_2231, w_061_2232, w_061_2233, w_061_2238, w_061_2239, w_061_2240, w_061_2243, w_061_2244, w_061_2246, w_061_2247, w_061_2248, w_061_2249, w_061_2250, w_061_2252, w_061_2253, w_061_2255, w_061_2261, w_061_2262, w_061_2264, w_061_2265, w_061_2266, w_061_2267, w_061_2269, w_061_2271, w_061_2272, w_061_2273, w_061_2274, w_061_2275, w_061_2277, w_061_2278, w_061_2281, w_061_2284, w_061_2285, w_061_2287, w_061_2289, w_061_2290, w_061_2291, w_061_2293, w_061_2294, w_061_2295, w_061_2296, w_061_2298, w_061_2299, w_061_2301, w_061_2302, w_061_2303, w_061_2304, w_061_2306, w_061_2307, w_061_2309, w_061_2310, w_061_2311, w_061_2312, w_061_2314, w_061_2315, w_061_2316, w_061_2317, w_061_2320;
  wire w_062_000, w_062_001, w_062_002, w_062_003, w_062_004, w_062_005, w_062_006, w_062_007, w_062_008, w_062_009, w_062_010, w_062_011, w_062_012, w_062_013, w_062_014, w_062_015, w_062_016, w_062_017, w_062_018, w_062_019, w_062_020, w_062_021, w_062_022, w_062_023, w_062_024, w_062_025, w_062_026, w_062_027, w_062_028, w_062_029, w_062_030, w_062_031, w_062_032, w_062_033, w_062_034, w_062_035, w_062_036, w_062_037, w_062_038, w_062_039, w_062_040, w_062_041, w_062_042, w_062_043, w_062_044, w_062_045, w_062_046, w_062_047, w_062_048, w_062_049, w_062_050, w_062_051, w_062_052, w_062_053, w_062_054, w_062_055, w_062_056, w_062_057, w_062_058, w_062_059, w_062_060, w_062_061, w_062_062, w_062_063, w_062_064, w_062_065, w_062_066, w_062_067, w_062_068, w_062_069, w_062_070, w_062_071, w_062_072, w_062_073, w_062_074, w_062_075, w_062_076, w_062_077, w_062_078, w_062_079, w_062_080, w_062_081, w_062_082, w_062_083, w_062_084, w_062_085, w_062_086, w_062_087, w_062_088, w_062_089, w_062_090, w_062_091, w_062_092, w_062_093, w_062_094, w_062_095, w_062_096, w_062_097, w_062_098, w_062_099, w_062_100, w_062_101, w_062_102, w_062_103, w_062_104, w_062_105, w_062_106, w_062_107, w_062_108, w_062_109, w_062_110, w_062_111, w_062_112, w_062_113, w_062_114, w_062_115, w_062_116, w_062_117, w_062_118, w_062_119, w_062_120, w_062_121, w_062_122, w_062_123, w_062_124, w_062_125, w_062_126, w_062_127, w_062_128, w_062_129, w_062_130, w_062_131, w_062_132, w_062_133, w_062_134, w_062_135, w_062_136, w_062_137, w_062_138, w_062_139, w_062_140, w_062_141, w_062_142, w_062_143, w_062_144, w_062_145, w_062_146, w_062_147, w_062_148, w_062_149, w_062_150, w_062_151, w_062_152, w_062_153, w_062_154, w_062_155, w_062_156, w_062_157, w_062_158, w_062_159, w_062_160, w_062_161, w_062_162, w_062_163, w_062_164, w_062_165, w_062_166, w_062_167, w_062_168, w_062_169, w_062_170, w_062_171, w_062_172, w_062_173, w_062_174, w_062_175, w_062_176, w_062_177, w_062_178, w_062_179, w_062_180, w_062_181, w_062_182, w_062_183, w_062_184, w_062_185, w_062_186, w_062_187, w_062_188, w_062_189, w_062_190, w_062_191, w_062_192, w_062_193, w_062_194, w_062_195, w_062_196, w_062_197, w_062_198, w_062_199, w_062_200, w_062_201, w_062_202, w_062_203, w_062_204, w_062_205, w_062_206, w_062_207, w_062_208, w_062_209, w_062_210, w_062_211, w_062_212, w_062_213, w_062_214, w_062_215, w_062_216, w_062_217, w_062_218, w_062_219, w_062_220, w_062_221, w_062_222, w_062_223, w_062_224, w_062_225, w_062_226, w_062_227, w_062_228, w_062_229, w_062_230, w_062_231, w_062_232, w_062_233, w_062_234, w_062_235, w_062_236, w_062_237, w_062_238, w_062_239, w_062_240, w_062_241, w_062_242, w_062_243, w_062_244, w_062_245, w_062_246, w_062_247, w_062_248, w_062_249, w_062_250, w_062_251, w_062_252, w_062_253, w_062_254, w_062_255, w_062_256, w_062_257, w_062_258, w_062_259, w_062_260, w_062_261, w_062_262, w_062_263, w_062_264, w_062_265, w_062_266, w_062_267, w_062_268, w_062_269, w_062_270, w_062_271, w_062_272, w_062_273, w_062_274, w_062_275, w_062_276, w_062_277, w_062_278, w_062_279, w_062_280, w_062_281, w_062_282, w_062_283, w_062_284, w_062_285, w_062_286, w_062_287, w_062_288, w_062_289, w_062_290, w_062_291, w_062_292, w_062_293, w_062_294, w_062_295, w_062_296, w_062_297, w_062_298, w_062_299, w_062_300, w_062_301, w_062_302, w_062_303, w_062_304, w_062_305, w_062_306, w_062_307, w_062_308, w_062_309, w_062_310, w_062_311, w_062_312, w_062_313, w_062_314, w_062_315, w_062_316, w_062_317, w_062_318, w_062_319, w_062_320, w_062_321, w_062_322, w_062_323, w_062_324, w_062_325, w_062_326, w_062_327, w_062_328, w_062_329, w_062_330, w_062_331, w_062_332, w_062_333, w_062_334, w_062_335, w_062_336, w_062_337, w_062_338, w_062_339, w_062_340, w_062_341, w_062_342, w_062_343, w_062_344, w_062_345, w_062_346, w_062_347, w_062_348, w_062_349, w_062_350, w_062_351, w_062_352, w_062_353, w_062_354, w_062_355, w_062_356, w_062_357, w_062_358, w_062_359, w_062_360, w_062_361, w_062_362, w_062_363, w_062_364, w_062_365, w_062_366, w_062_367, w_062_368, w_062_369, w_062_370, w_062_371, w_062_372, w_062_373, w_062_374, w_062_375, w_062_376, w_062_377, w_062_378, w_062_379, w_062_380, w_062_381, w_062_382, w_062_383, w_062_384, w_062_385, w_062_386, w_062_387, w_062_388, w_062_389, w_062_390, w_062_391, w_062_392, w_062_393, w_062_394, w_062_395, w_062_396, w_062_397, w_062_398, w_062_399, w_062_400, w_062_401, w_062_402, w_062_403, w_062_404, w_062_405, w_062_406, w_062_407, w_062_408, w_062_409, w_062_410, w_062_411, w_062_412, w_062_413, w_062_414, w_062_415, w_062_416, w_062_417, w_062_418, w_062_419, w_062_420, w_062_421, w_062_422, w_062_423, w_062_424, w_062_425, w_062_426, w_062_427, w_062_428, w_062_429, w_062_430, w_062_431, w_062_432, w_062_433, w_062_434, w_062_435, w_062_436, w_062_437, w_062_438, w_062_439, w_062_440, w_062_441, w_062_442, w_062_443, w_062_444, w_062_445, w_062_446, w_062_447, w_062_448, w_062_449, w_062_450, w_062_451, w_062_452, w_062_453, w_062_454, w_062_455, w_062_456, w_062_457, w_062_458, w_062_459, w_062_460, w_062_461, w_062_462, w_062_463, w_062_464, w_062_465, w_062_466, w_062_467, w_062_468, w_062_469, w_062_470, w_062_471, w_062_472, w_062_473, w_062_474, w_062_475, w_062_476, w_062_477, w_062_478, w_062_479, w_062_480, w_062_481, w_062_482, w_062_483, w_062_484, w_062_485, w_062_486, w_062_487, w_062_488, w_062_489, w_062_490, w_062_491, w_062_492, w_062_493, w_062_494, w_062_495, w_062_496, w_062_497, w_062_498, w_062_499, w_062_500, w_062_501, w_062_502, w_062_503, w_062_504, w_062_505, w_062_506;
  wire w_063_000, w_063_002, w_063_004, w_063_005, w_063_006, w_063_007, w_063_009, w_063_010, w_063_011, w_063_012, w_063_013, w_063_016, w_063_017, w_063_019, w_063_022, w_063_024, w_063_026, w_063_029, w_063_030, w_063_031, w_063_032, w_063_034, w_063_035, w_063_036, w_063_037, w_063_038, w_063_040, w_063_042, w_063_043, w_063_044, w_063_045, w_063_046, w_063_047, w_063_050, w_063_051, w_063_052, w_063_053, w_063_054, w_063_055, w_063_056, w_063_058, w_063_059, w_063_060, w_063_061, w_063_062, w_063_063, w_063_064, w_063_065, w_063_067, w_063_068, w_063_070, w_063_071, w_063_074, w_063_077, w_063_078, w_063_079, w_063_080, w_063_082, w_063_083, w_063_084, w_063_085, w_063_086, w_063_087, w_063_090, w_063_091, w_063_092, w_063_093, w_063_094, w_063_095, w_063_096, w_063_098, w_063_100, w_063_101, w_063_102, w_063_103, w_063_105, w_063_106, w_063_108, w_063_109, w_063_111, w_063_112, w_063_113, w_063_114, w_063_115, w_063_117, w_063_118, w_063_119, w_063_121, w_063_123, w_063_124, w_063_125, w_063_126, w_063_127, w_063_128, w_063_129, w_063_130, w_063_131, w_063_132, w_063_134, w_063_135, w_063_140, w_063_141, w_063_142, w_063_143, w_063_145, w_063_147, w_063_148, w_063_149, w_063_150, w_063_151, w_063_152, w_063_153, w_063_154, w_063_155, w_063_156, w_063_157, w_063_161, w_063_164, w_063_167, w_063_169, w_063_170, w_063_171, w_063_173, w_063_174, w_063_176, w_063_177, w_063_178, w_063_179, w_063_180, w_063_181, w_063_182, w_063_184, w_063_187, w_063_188, w_063_192, w_063_193, w_063_194, w_063_195, w_063_196, w_063_198, w_063_200, w_063_202, w_063_204, w_063_206, w_063_207, w_063_208, w_063_211, w_063_212, w_063_214, w_063_223, w_063_226, w_063_227, w_063_229, w_063_232, w_063_233, w_063_234, w_063_235, w_063_236, w_063_239, w_063_241, w_063_242, w_063_243, w_063_245, w_063_246, w_063_249, w_063_250, w_063_251, w_063_252, w_063_253, w_063_255, w_063_256, w_063_258, w_063_260, w_063_261, w_063_262, w_063_263, w_063_266, w_063_267, w_063_268, w_063_269, w_063_272, w_063_273, w_063_275, w_063_277, w_063_278, w_063_279, w_063_281, w_063_282, w_063_283, w_063_284, w_063_285, w_063_286, w_063_290, w_063_291, w_063_293, w_063_294, w_063_296, w_063_297, w_063_299, w_063_301, w_063_302, w_063_304, w_063_305, w_063_306, w_063_308, w_063_310, w_063_311, w_063_313, w_063_314, w_063_315, w_063_317, w_063_318, w_063_319, w_063_321, w_063_322, w_063_323, w_063_324, w_063_326, w_063_331, w_063_332, w_063_334, w_063_335, w_063_336, w_063_337, w_063_338, w_063_339, w_063_340, w_063_341, w_063_342, w_063_343, w_063_345, w_063_347, w_063_349, w_063_350, w_063_351, w_063_352, w_063_354, w_063_355, w_063_356, w_063_357, w_063_359, w_063_361, w_063_364, w_063_365, w_063_366, w_063_368, w_063_369, w_063_371, w_063_373, w_063_374, w_063_375, w_063_376, w_063_377, w_063_379, w_063_380, w_063_381, w_063_383, w_063_384, w_063_385, w_063_386, w_063_387, w_063_388, w_063_389, w_063_395, w_063_396, w_063_397, w_063_400, w_063_401, w_063_403, w_063_404, w_063_408, w_063_409, w_063_410, w_063_411, w_063_413, w_063_415, w_063_417, w_063_418, w_063_419, w_063_420, w_063_423, w_063_424, w_063_425, w_063_427, w_063_430, w_063_432, w_063_433, w_063_434, w_063_436, w_063_437, w_063_439, w_063_441, w_063_442, w_063_443, w_063_447, w_063_449, w_063_450, w_063_451, w_063_454, w_063_455, w_063_457, w_063_458, w_063_461, w_063_463, w_063_464, w_063_465, w_063_468, w_063_469, w_063_473, w_063_474, w_063_479, w_063_481, w_063_482, w_063_484, w_063_485, w_063_486, w_063_488, w_063_489, w_063_491, w_063_492, w_063_493, w_063_494, w_063_497, w_063_500, w_063_503, w_063_504, w_063_507, w_063_508, w_063_509, w_063_510, w_063_513, w_063_518, w_063_519, w_063_520, w_063_521, w_063_522, w_063_523, w_063_525, w_063_526, w_063_527, w_063_529, w_063_530, w_063_531, w_063_532, w_063_533, w_063_534, w_063_535, w_063_536, w_063_538, w_063_539, w_063_540, w_063_541, w_063_542, w_063_545, w_063_547, w_063_548, w_063_549, w_063_554, w_063_555, w_063_558, w_063_559, w_063_560, w_063_561, w_063_562, w_063_564, w_063_565, w_063_566, w_063_567, w_063_568, w_063_569, w_063_572, w_063_574, w_063_576, w_063_577, w_063_578, w_063_579, w_063_580, w_063_581, w_063_582, w_063_583, w_063_584, w_063_586, w_063_587, w_063_590, w_063_592, w_063_593, w_063_595, w_063_596, w_063_597, w_063_598, w_063_599, w_063_600, w_063_601, w_063_603, w_063_604, w_063_605, w_063_606, w_063_607, w_063_608, w_063_609, w_063_610, w_063_612, w_063_613, w_063_614, w_063_616, w_063_617, w_063_618, w_063_619, w_063_620, w_063_622, w_063_623, w_063_624, w_063_625, w_063_626, w_063_627, w_063_629, w_063_630, w_063_631, w_063_632, w_063_633, w_063_634, w_063_635, w_063_637, w_063_638, w_063_640, w_063_641, w_063_642, w_063_643, w_063_644, w_063_647, w_063_649, w_063_650, w_063_653, w_063_654, w_063_656, w_063_657, w_063_658, w_063_659, w_063_660, w_063_661, w_063_664, w_063_665, w_063_666, w_063_667, w_063_668, w_063_669, w_063_671, w_063_674, w_063_675, w_063_676, w_063_679, w_063_680, w_063_681, w_063_685, w_063_686, w_063_687, w_063_688, w_063_690, w_063_691, w_063_692, w_063_693, w_063_694, w_063_695, w_063_696, w_063_697, w_063_698, w_063_699, w_063_700, w_063_703, w_063_704, w_063_705, w_063_706, w_063_707, w_063_708, w_063_709, w_063_710, w_063_713, w_063_714, w_063_715, w_063_717, w_063_719, w_063_721, w_063_723, w_063_725, w_063_727, w_063_728, w_063_729, w_063_731, w_063_733, w_063_734, w_063_737, w_063_738, w_063_740, w_063_741, w_063_742, w_063_745, w_063_746, w_063_751, w_063_752, w_063_753, w_063_755, w_063_756, w_063_757, w_063_758, w_063_759, w_063_761, w_063_763, w_063_764, w_063_765, w_063_766, w_063_768, w_063_769, w_063_770, w_063_772, w_063_773, w_063_775, w_063_776, w_063_777, w_063_780, w_063_782, w_063_783, w_063_784, w_063_787, w_063_788, w_063_789, w_063_791, w_063_792, w_063_793, w_063_794, w_063_795, w_063_797, w_063_798, w_063_800, w_063_801, w_063_802, w_063_805, w_063_806, w_063_807, w_063_808, w_063_809, w_063_810, w_063_811, w_063_812, w_063_813, w_063_814, w_063_815, w_063_816, w_063_817, w_063_819, w_063_821, w_063_823, w_063_825, w_063_827, w_063_830, w_063_832, w_063_834, w_063_836, w_063_837, w_063_838, w_063_840, w_063_841, w_063_843, w_063_844, w_063_846, w_063_847, w_063_848, w_063_849, w_063_851, w_063_852, w_063_855, w_063_856, w_063_857, w_063_859, w_063_861, w_063_862, w_063_863, w_063_864, w_063_868, w_063_869, w_063_870, w_063_871, w_063_873, w_063_874, w_063_875, w_063_877, w_063_878, w_063_879, w_063_880, w_063_881, w_063_882, w_063_883, w_063_884, w_063_886, w_063_887, w_063_888, w_063_889, w_063_890, w_063_891, w_063_892, w_063_893, w_063_894, w_063_895, w_063_897, w_063_898, w_063_899, w_063_900, w_063_902, w_063_903, w_063_904, w_063_906, w_063_907, w_063_908, w_063_909, w_063_910, w_063_911, w_063_913, w_063_916, w_063_919, w_063_920, w_063_921, w_063_922, w_063_923, w_063_926, w_063_928, w_063_930, w_063_931, w_063_933, w_063_936, w_063_937, w_063_942, w_063_943, w_063_944, w_063_946, w_063_947, w_063_948, w_063_949, w_063_953, w_063_954, w_063_957, w_063_958, w_063_959, w_063_960, w_063_961, w_063_962, w_063_965, w_063_966, w_063_967, w_063_969, w_063_970, w_063_973, w_063_974, w_063_975, w_063_977, w_063_978, w_063_979, w_063_982, w_063_983, w_063_984, w_063_985, w_063_986, w_063_987, w_063_988, w_063_994, w_063_995, w_063_996, w_063_999, w_063_1000, w_063_1004, w_063_1005, w_063_1007, w_063_1008, w_063_1010, w_063_1011, w_063_1015, w_063_1016, w_063_1019, w_063_1021, w_063_1022, w_063_1024, w_063_1025, w_063_1027, w_063_1030, w_063_1031, w_063_1033, w_063_1034, w_063_1035, w_063_1036, w_063_1037, w_063_1038, w_063_1040, w_063_1041, w_063_1042, w_063_1043, w_063_1044, w_063_1045, w_063_1047, w_063_1048, w_063_1050, w_063_1051, w_063_1052, w_063_1053, w_063_1057, w_063_1060, w_063_1061, w_063_1064, w_063_1065, w_063_1066, w_063_1067, w_063_1069, w_063_1071, w_063_1072, w_063_1074, w_063_1077, w_063_1078, w_063_1079, w_063_1082, w_063_1083, w_063_1086, w_063_1088, w_063_1089, w_063_1090, w_063_1091, w_063_1097, w_063_1099, w_063_1100, w_063_1101, w_063_1102, w_063_1104, w_063_1105, w_063_1107, w_063_1109, w_063_1112, w_063_1113, w_063_1115, w_063_1116, w_063_1117, w_063_1118, w_063_1120, w_063_1121, w_063_1124, w_063_1128, w_063_1130, w_063_1131, w_063_1132, w_063_1133, w_063_1134, w_063_1137, w_063_1139, w_063_1142, w_063_1144, w_063_1145, w_063_1149, w_063_1150, w_063_1151, w_063_1152, w_063_1153, w_063_1154, w_063_1155, w_063_1156, w_063_1157, w_063_1159, w_063_1160, w_063_1162, w_063_1163, w_063_1164, w_063_1165, w_063_1168, w_063_1169, w_063_1170, w_063_1171, w_063_1172, w_063_1173, w_063_1174, w_063_1175, w_063_1176, w_063_1177, w_063_1178, w_063_1180, w_063_1181, w_063_1182, w_063_1184, w_063_1185, w_063_1186, w_063_1187, w_063_1189, w_063_1191, w_063_1193, w_063_1195, w_063_1196, w_063_1197, w_063_1198, w_063_1199, w_063_1200, w_063_1201, w_063_1202, w_063_1203, w_063_1204, w_063_1206, w_063_1207, w_063_1208, w_063_1209, w_063_1210, w_063_1211, w_063_1213, w_063_1214, w_063_1217, w_063_1218, w_063_1220, w_063_1221, w_063_1223, w_063_1226, w_063_1227, w_063_1228, w_063_1231, w_063_1232, w_063_1233, w_063_1234, w_063_1238, w_063_1239, w_063_1240, w_063_1241, w_063_1242, w_063_1244, w_063_1245, w_063_1246, w_063_1248, w_063_1250, w_063_1251, w_063_1252, w_063_1253, w_063_1254, w_063_1255, w_063_1257, w_063_1258, w_063_1261, w_063_1263, w_063_1264, w_063_1265, w_063_1266, w_063_1268, w_063_1269, w_063_1270, w_063_1272, w_063_1274, w_063_1275, w_063_1276, w_063_1277, w_063_1278, w_063_1279, w_063_1280, w_063_1281, w_063_1284, w_063_1286, w_063_1287, w_063_1288, w_063_1289, w_063_1290, w_063_1291, w_063_1294, w_063_1295, w_063_1296, w_063_1298, w_063_1299, w_063_1300, w_063_1301, w_063_1303, w_063_1304, w_063_1305, w_063_1306, w_063_1307, w_063_1308, w_063_1311, w_063_1312, w_063_1313, w_063_1314, w_063_1315, w_063_1317, w_063_1319, w_063_1320, w_063_1323, w_063_1326, w_063_1328, w_063_1335, w_063_1336, w_063_1337, w_063_1339, w_063_1340, w_063_1341, w_063_1342, w_063_1343, w_063_1345, w_063_1347, w_063_1349, w_063_1350, w_063_1351, w_063_1352, w_063_1353, w_063_1354, w_063_1356, w_063_1357, w_063_1359, w_063_1360, w_063_1361, w_063_1366, w_063_1367, w_063_1368, w_063_1369, w_063_1370, w_063_1371, w_063_1372, w_063_1373, w_063_1374, w_063_1375, w_063_1377, w_063_1379, w_063_1381, w_063_1382, w_063_1383, w_063_1384, w_063_1385, w_063_1387, w_063_1388, w_063_1389, w_063_1390, w_063_1392, w_063_1394, w_063_1395, w_063_1399, w_063_1400, w_063_1401, w_063_1402, w_063_1403, w_063_1404, w_063_1405, w_063_1406, w_063_1410, w_063_1412, w_063_1413, w_063_1414, w_063_1415, w_063_1417, w_063_1418, w_063_1419, w_063_1420, w_063_1421, w_063_1422, w_063_1427, w_063_1428, w_063_1429, w_063_1430, w_063_1431, w_063_1432, w_063_1433, w_063_1439, w_063_1440, w_063_1444, w_063_1445, w_063_1446, w_063_1447, w_063_1449, w_063_1450, w_063_1451, w_063_1453, w_063_1457, w_063_1458, w_063_1459, w_063_1462, w_063_1463, w_063_1464, w_063_1466, w_063_1468, w_063_1470, w_063_1471, w_063_1473, w_063_1474, w_063_1476, w_063_1480, w_063_1481, w_063_1482, w_063_1484, w_063_1485, w_063_1486, w_063_1487, w_063_1488, w_063_1489, w_063_1490, w_063_1491, w_063_1494, w_063_1495, w_063_1496, w_063_1497, w_063_1501, w_063_1502, w_063_1503, w_063_1505, w_063_1506, w_063_1507, w_063_1509, w_063_1510, w_063_1512, w_063_1522, w_063_1530, w_063_1532, w_063_1539, w_063_1541, w_063_1543, w_063_1546, w_063_1551, w_063_1553, w_063_1555, w_063_1557, w_063_1559, w_063_1560, w_063_1563, w_063_1565, w_063_1566, w_063_1575, w_063_1577, w_063_1579, w_063_1582, w_063_1583, w_063_1584, w_063_1586, w_063_1587, w_063_1589, w_063_1590, w_063_1594, w_063_1595, w_063_1601, w_063_1607, w_063_1608, w_063_1609, w_063_1610, w_063_1614, w_063_1620, w_063_1623, w_063_1624, w_063_1625, w_063_1627, w_063_1630, w_063_1632, w_063_1635, w_063_1636, w_063_1639, w_063_1640, w_063_1641, w_063_1642, w_063_1643, w_063_1648, w_063_1650, w_063_1653, w_063_1656, w_063_1657, w_063_1668, w_063_1676, w_063_1681, w_063_1685, w_063_1686, w_063_1691, w_063_1697, w_063_1703, w_063_1704, w_063_1705, w_063_1706, w_063_1707, w_063_1709, w_063_1710, w_063_1713, w_063_1714, w_063_1715, w_063_1716, w_063_1717, w_063_1722, w_063_1724, w_063_1725, w_063_1726, w_063_1733, w_063_1735, w_063_1736, w_063_1739, w_063_1743, w_063_1749, w_063_1756, w_063_1763, w_063_1764, w_063_1765, w_063_1770, w_063_1774, w_063_1775, w_063_1777, w_063_1781, w_063_1782, w_063_1787, w_063_1788, w_063_1789, w_063_1792, w_063_1793, w_063_1799, w_063_1800, w_063_1801, w_063_1806, w_063_1808, w_063_1817, w_063_1822, w_063_1823, w_063_1824, w_063_1826, w_063_1828, w_063_1832, w_063_1833, w_063_1835, w_063_1836, w_063_1839, w_063_1845, w_063_1847, w_063_1849, w_063_1852, w_063_1853, w_063_1856, w_063_1857, w_063_1860, w_063_1862, w_063_1866, w_063_1867, w_063_1876, w_063_1877, w_063_1883, w_063_1888, w_063_1894, w_063_1895, w_063_1896, w_063_1899, w_063_1900, w_063_1903, w_063_1905, w_063_1910, w_063_1912, w_063_1914, w_063_1923, w_063_1924, w_063_1927, w_063_1928, w_063_1930, w_063_1932, w_063_1934, w_063_1936, w_063_1937, w_063_1939, w_063_1940, w_063_1942, w_063_1944, w_063_1945, w_063_1948, w_063_1949, w_063_1951, w_063_1952, w_063_1953, w_063_1958, w_063_1959, w_063_1960, w_063_1964, w_063_1984, w_063_1986, w_063_1991, w_063_1992, w_063_1993, w_063_1995, w_063_1999, w_063_2000, w_063_2004, w_063_2009, w_063_2017, w_063_2018, w_063_2022, w_063_2026, w_063_2028, w_063_2033, w_063_2034, w_063_2035, w_063_2036, w_063_2037, w_063_2039, w_063_2043, w_063_2044, w_063_2048, w_063_2049, w_063_2051, w_063_2052, w_063_2055, w_063_2056, w_063_2058, w_063_2061, w_063_2065, w_063_2067, w_063_2070, w_063_2071, w_063_2072, w_063_2073, w_063_2075, w_063_2077, w_063_2080, w_063_2086, w_063_2087, w_063_2092, w_063_2093, w_063_2097, w_063_2099, w_063_2101, w_063_2102, w_063_2105, w_063_2112, w_063_2114, w_063_2116, w_063_2120, w_063_2126, w_063_2129, w_063_2131, w_063_2133, w_063_2134, w_063_2136, w_063_2137, w_063_2139, w_063_2140, w_063_2143, w_063_2148, w_063_2153, w_063_2159, w_063_2161, w_063_2164, w_063_2165, w_063_2166, w_063_2167, w_063_2169, w_063_2172, w_063_2174, w_063_2175, w_063_2176, w_063_2177, w_063_2178, w_063_2182, w_063_2183, w_063_2188, w_063_2189, w_063_2190, w_063_2193, w_063_2197, w_063_2202, w_063_2206, w_063_2207, w_063_2208, w_063_2210, w_063_2214, w_063_2215, w_063_2218, w_063_2220, w_063_2222, w_063_2225, w_063_2229, w_063_2237, w_063_2242, w_063_2244, w_063_2246, w_063_2248, w_063_2251, w_063_2252, w_063_2253, w_063_2254, w_063_2259, w_063_2260, w_063_2261, w_063_2262, w_063_2264, w_063_2268, w_063_2269, w_063_2273, w_063_2275, w_063_2279, w_063_2281, w_063_2286, w_063_2288, w_063_2289, w_063_2293, w_063_2297, w_063_2298, w_063_2299, w_063_2303, w_063_2306, w_063_2307, w_063_2313, w_063_2314, w_063_2316, w_063_2322, w_063_2323, w_063_2327, w_063_2328, w_063_2330, w_063_2333, w_063_2335, w_063_2337, w_063_2341, w_063_2348, w_063_2352, w_063_2355, w_063_2360, w_063_2361, w_063_2362, w_063_2367, w_063_2374, w_063_2377, w_063_2383, w_063_2388, w_063_2391, w_063_2392, w_063_2393, w_063_2394, w_063_2396, w_063_2397, w_063_2400, w_063_2401, w_063_2402, w_063_2404, w_063_2406, w_063_2408, w_063_2410, w_063_2415, w_063_2420, w_063_2422, w_063_2423, w_063_2424, w_063_2425, w_063_2430, w_063_2433, w_063_2435, w_063_2437, w_063_2442, w_063_2443, w_063_2447, w_063_2450, w_063_2451, w_063_2452, w_063_2455, w_063_2456, w_063_2459, w_063_2461, w_063_2468, w_063_2470, w_063_2472, w_063_2473, w_063_2475, w_063_2476, w_063_2477, w_063_2478, w_063_2479, w_063_2481, w_063_2485, w_063_2488, w_063_2490, w_063_2491, w_063_2493, w_063_2494, w_063_2495, w_063_2498, w_063_2499, w_063_2500, w_063_2506, w_063_2510, w_063_2511, w_063_2513, w_063_2519, w_063_2520, w_063_2521, w_063_2525, w_063_2527, w_063_2529, w_063_2530, w_063_2533, w_063_2536, w_063_2537, w_063_2538, w_063_2543, w_063_2546, w_063_2552, w_063_2553, w_063_2555, w_063_2559, w_063_2560, w_063_2561, w_063_2565, w_063_2567, w_063_2569, w_063_2570, w_063_2571, w_063_2572, w_063_2574, w_063_2576, w_063_2577, w_063_2578, w_063_2579, w_063_2580, w_063_2582, w_063_2585, w_063_2590, w_063_2591, w_063_2592, w_063_2595, w_063_2596, w_063_2598, w_063_2600, w_063_2603, w_063_2604, w_063_2605, w_063_2608, w_063_2613, w_063_2615, w_063_2616, w_063_2617, w_063_2621, w_063_2624, w_063_2625, w_063_2626, w_063_2628, w_063_2629, w_063_2630, w_063_2632, w_063_2633, w_063_2635, w_063_2636, w_063_2637, w_063_2638, w_063_2639, w_063_2642, w_063_2645, w_063_2647, w_063_2648, w_063_2650, w_063_2652, w_063_2653, w_063_2655, w_063_2659, w_063_2663, w_063_2667, w_063_2668, w_063_2669, w_063_2670, w_063_2671, w_063_2675, w_063_2677, w_063_2679, w_063_2683, w_063_2688, w_063_2690, w_063_2691, w_063_2692, w_063_2693, w_063_2694, w_063_2695, w_063_2696, w_063_2698, w_063_2700, w_063_2702, w_063_2704, w_063_2708, w_063_2710, w_063_2713, w_063_2719, w_063_2720, w_063_2722, w_063_2725, w_063_2727, w_063_2728, w_063_2729, w_063_2730, w_063_2732, w_063_2734, w_063_2735, w_063_2736, w_063_2738, w_063_2739, w_063_2742, w_063_2746, w_063_2750, w_063_2751, w_063_2752, w_063_2754, w_063_2757, w_063_2758, w_063_2759, w_063_2762, w_063_2764, w_063_2767, w_063_2769, w_063_2770, w_063_2773, w_063_2774, w_063_2778, w_063_2779, w_063_2782, w_063_2783, w_063_2784, w_063_2785, w_063_2787, w_063_2790, w_063_2792, w_063_2794, w_063_2796, w_063_2800, w_063_2801, w_063_2803, w_063_2805, w_063_2807, w_063_2810, w_063_2812, w_063_2813, w_063_2819, w_063_2824, w_063_2827, w_063_2831, w_063_2832, w_063_2845, w_063_2846, w_063_2849, w_063_2850, w_063_2851, w_063_2853, w_063_2855, w_063_2859, w_063_2860, w_063_2861, w_063_2863, w_063_2865, w_063_2866, w_063_2867, w_063_2869, w_063_2870, w_063_2872, w_063_2873, w_063_2874, w_063_2875, w_063_2877, w_063_2878, w_063_2880, w_063_2881, w_063_2882, w_063_2888, w_063_2889, w_063_2890, w_063_2892, w_063_2893, w_063_2895, w_063_2896, w_063_2897, w_063_2898, w_063_2899, w_063_2907, w_063_2910, w_063_2913, w_063_2917, w_063_2918, w_063_2920, w_063_2923, w_063_2932, w_063_2934, w_063_2937, w_063_2939, w_063_2940, w_063_2941, w_063_2944, w_063_2947, w_063_2948, w_063_2954, w_063_2956, w_063_2957, w_063_2960, w_063_2966, w_063_2969, w_063_2972, w_063_2973, w_063_2976, w_063_2979, w_063_2980, w_063_2983, w_063_2984, w_063_2989, w_063_2991, w_063_2994, w_063_2995, w_063_3001, w_063_3004, w_063_3009, w_063_3011, w_063_3016, w_063_3017, w_063_3018, w_063_3019, w_063_3020, w_063_3022, w_063_3027, w_063_3038, w_063_3039, w_063_3040, w_063_3043, w_063_3045, w_063_3047, w_063_3048, w_063_3049, w_063_3052, w_063_3053, w_063_3054, w_063_3055, w_063_3060, w_063_3064, w_063_3070, w_063_3071, w_063_3072, w_063_3075, w_063_3078, w_063_3087, w_063_3089, w_063_3090, w_063_3091, w_063_3093, w_063_3094, w_063_3100, w_063_3104, w_063_3107, w_063_3108, w_063_3111, w_063_3113, w_063_3115, w_063_3118, w_063_3123, w_063_3128, w_063_3129, w_063_3130, w_063_3133, w_063_3134, w_063_3136, w_063_3137, w_063_3138, w_063_3139, w_063_3140, w_063_3141, w_063_3144, w_063_3146, w_063_3149, w_063_3152, w_063_3153, w_063_3154, w_063_3157, w_063_3166, w_063_3167, w_063_3169, w_063_3170, w_063_3171, w_063_3176, w_063_3177, w_063_3180, w_063_3186, w_063_3189, w_063_3190, w_063_3191, w_063_3195, w_063_3199, w_063_3202, w_063_3203, w_063_3204, w_063_3206, w_063_3210, w_063_3212, w_063_3213, w_063_3227, w_063_3229, w_063_3231, w_063_3234, w_063_3236, w_063_3237, w_063_3245, w_063_3246, w_063_3248, w_063_3250, w_063_3255, w_063_3256, w_063_3258, w_063_3260, w_063_3267, w_063_3272, w_063_3274, w_063_3275, w_063_3279, w_063_3285, w_063_3292, w_063_3294, w_063_3299, w_063_3300, w_063_3304, w_063_3306, w_063_3307, w_063_3309, w_063_3310, w_063_3311, w_063_3313, w_063_3314, w_063_3315, w_063_3317, w_063_3318, w_063_3319, w_063_3320, w_063_3321, w_063_3322, w_063_3323, w_063_3329, w_063_3330, w_063_3331, w_063_3336, w_063_3337, w_063_3341, w_063_3343, w_063_3346, w_063_3352, w_063_3353, w_063_3354, w_063_3357, w_063_3358, w_063_3360, w_063_3366, w_063_3367, w_063_3373, w_063_3375, w_063_3382, w_063_3387, w_063_3393, w_063_3394, w_063_3397, w_063_3398, w_063_3399, w_063_3400, w_063_3401, w_063_3402, w_063_3406, w_063_3408, w_063_3414, w_063_3415, w_063_3417, w_063_3425, w_063_3430, w_063_3431, w_063_3432, w_063_3433, w_063_3436, w_063_3438, w_063_3440, w_063_3447, w_063_3449, w_063_3452, w_063_3454, w_063_3455, w_063_3460, w_063_3462, w_063_3464, w_063_3465, w_063_3466, w_063_3468, w_063_3470, w_063_3472, w_063_3474, w_063_3475, w_063_3476, w_063_3477, w_063_3478, w_063_3480, w_063_3483, w_063_3484, w_063_3485;
  wire w_064_001, w_064_002, w_064_003, w_064_004, w_064_005, w_064_006, w_064_007, w_064_008, w_064_009, w_064_013, w_064_014, w_064_016, w_064_017, w_064_018, w_064_019, w_064_020, w_064_022, w_064_024, w_064_025, w_064_026, w_064_030, w_064_031, w_064_032, w_064_033, w_064_034, w_064_035, w_064_036, w_064_038, w_064_039, w_064_040, w_064_042, w_064_045, w_064_047, w_064_049, w_064_050, w_064_051, w_064_052, w_064_053, w_064_055, w_064_056, w_064_057, w_064_058, w_064_059, w_064_060, w_064_061, w_064_062, w_064_063, w_064_064, w_064_067, w_064_068, w_064_069, w_064_071, w_064_074, w_064_075, w_064_080, w_064_082, w_064_083, w_064_085, w_064_088, w_064_089, w_064_093, w_064_094, w_064_097, w_064_098, w_064_099, w_064_100, w_064_102, w_064_105, w_064_106, w_064_108, w_064_112, w_064_114, w_064_115, w_064_116, w_064_117, w_064_118, w_064_119, w_064_121, w_064_122, w_064_124, w_064_125, w_064_126, w_064_127, w_064_129, w_064_130, w_064_131, w_064_132, w_064_133, w_064_134, w_064_135, w_064_136, w_064_137, w_064_139, w_064_140, w_064_141, w_064_142, w_064_143, w_064_144, w_064_145, w_064_146, w_064_147, w_064_149, w_064_150, w_064_152, w_064_153, w_064_154, w_064_155, w_064_156, w_064_157, w_064_158, w_064_161, w_064_162, w_064_163, w_064_164, w_064_165, w_064_166, w_064_167, w_064_168, w_064_169, w_064_172, w_064_173, w_064_176, w_064_177, w_064_178, w_064_180, w_064_182, w_064_183, w_064_184, w_064_186, w_064_188, w_064_189, w_064_191, w_064_193, w_064_194, w_064_196, w_064_198, w_064_199, w_064_200, w_064_201, w_064_202, w_064_203, w_064_204, w_064_205, w_064_207, w_064_208, w_064_209, w_064_213, w_064_214, w_064_215, w_064_216, w_064_218, w_064_219, w_064_220, w_064_221, w_064_222, w_064_225, w_064_226, w_064_228, w_064_229, w_064_230, w_064_232, w_064_233, w_064_234, w_064_236, w_064_237, w_064_238, w_064_240, w_064_243, w_064_244, w_064_245, w_064_249, w_064_252, w_064_253, w_064_254, w_064_256, w_064_257, w_064_258, w_064_259, w_064_261, w_064_262, w_064_263, w_064_264, w_064_265, w_064_267, w_064_268, w_064_271, w_064_273, w_064_277, w_064_278, w_064_279, w_064_280, w_064_281, w_064_282, w_064_284, w_064_285, w_064_287, w_064_290, w_064_292, w_064_293, w_064_294, w_064_295, w_064_296, w_064_297, w_064_298, w_064_299, w_064_300, w_064_301, w_064_304, w_064_306, w_064_307, w_064_308, w_064_309, w_064_310, w_064_311, w_064_312, w_064_314, w_064_315, w_064_318, w_064_319, w_064_322, w_064_323, w_064_324, w_064_325, w_064_326, w_064_327, w_064_328, w_064_329, w_064_330, w_064_331, w_064_332, w_064_333, w_064_335, w_064_337, w_064_339, w_064_340, w_064_342, w_064_343, w_064_346, w_064_348, w_064_349, w_064_351, w_064_352, w_064_353, w_064_356, w_064_357, w_064_363, w_064_365, w_064_366, w_064_367, w_064_368, w_064_369, w_064_371, w_064_372, w_064_377, w_064_379, w_064_382, w_064_383, w_064_384, w_064_386, w_064_389, w_064_390, w_064_391, w_064_392, w_064_393, w_064_394, w_064_395, w_064_396, w_064_399, w_064_402, w_064_403, w_064_404, w_064_405, w_064_407, w_064_408, w_064_409, w_064_413, w_064_414, w_064_416, w_064_417, w_064_420, w_064_422, w_064_423, w_064_426, w_064_427, w_064_428, w_064_429, w_064_430, w_064_432, w_064_433, w_064_434, w_064_436, w_064_437, w_064_439, w_064_440, w_064_441, w_064_443, w_064_444, w_064_445, w_064_448, w_064_451, w_064_453, w_064_454, w_064_459, w_064_461, w_064_462, w_064_464, w_064_466, w_064_467, w_064_469, w_064_471, w_064_475, w_064_476, w_064_477, w_064_478, w_064_480, w_064_481, w_064_482, w_064_483, w_064_484, w_064_485, w_064_486, w_064_487, w_064_488, w_064_492, w_064_493, w_064_495, w_064_497, w_064_498, w_064_500, w_064_501, w_064_503, w_064_504, w_064_505, w_064_506, w_064_507, w_064_508, w_064_509, w_064_510, w_064_511, w_064_513, w_064_516, w_064_518, w_064_520, w_064_522, w_064_524, w_064_526, w_064_527, w_064_530, w_064_531, w_064_533, w_064_534, w_064_536, w_064_538, w_064_539, w_064_540, w_064_542, w_064_543, w_064_544, w_064_545, w_064_546, w_064_548, w_064_551, w_064_554, w_064_557, w_064_558, w_064_559, w_064_562, w_064_563, w_064_564, w_064_565, w_064_566, w_064_570, w_064_571, w_064_574, w_064_575, w_064_578, w_064_579, w_064_581, w_064_582, w_064_583, w_064_584, w_064_585, w_064_586, w_064_589, w_064_593, w_064_597, w_064_598, w_064_599, w_064_600, w_064_601, w_064_602, w_064_603, w_064_604, w_064_606, w_064_607, w_064_608, w_064_610, w_064_613, w_064_614, w_064_620, w_064_623, w_064_624, w_064_626, w_064_627, w_064_628, w_064_630, w_064_631, w_064_632, w_064_633, w_064_634, w_064_635, w_064_636, w_064_637, w_064_638, w_064_639, w_064_640, w_064_642, w_064_643, w_064_645, w_064_646, w_064_647, w_064_649, w_064_652, w_064_653, w_064_654, w_064_656, w_064_657, w_064_659, w_064_661, w_064_662, w_064_664, w_064_668, w_064_669, w_064_670, w_064_672, w_064_675, w_064_676, w_064_677, w_064_680, w_064_682, w_064_684, w_064_685, w_064_686, w_064_687, w_064_690, w_064_691, w_064_692, w_064_693, w_064_695, w_064_698, w_064_699, w_064_700, w_064_703, w_064_705, w_064_706, w_064_707, w_064_708, w_064_711, w_064_712, w_064_714, w_064_715, w_064_716, w_064_717, w_064_718, w_064_720, w_064_721, w_064_723, w_064_725, w_064_726, w_064_727, w_064_728, w_064_730, w_064_732, w_064_733, w_064_736, w_064_737, w_064_738, w_064_740, w_064_741, w_064_742, w_064_743, w_064_744, w_064_745, w_064_747, w_064_748, w_064_750, w_064_752, w_064_754, w_064_755, w_064_757, w_064_758, w_064_759, w_064_760, w_064_761, w_064_762, w_064_763, w_064_765, w_064_768, w_064_771, w_064_773, w_064_774, w_064_775, w_064_778, w_064_779, w_064_781, w_064_783, w_064_784, w_064_788, w_064_789, w_064_791, w_064_792, w_064_795, w_064_796, w_064_800, w_064_801, w_064_804, w_064_805, w_064_806, w_064_807, w_064_808, w_064_809, w_064_811, w_064_814, w_064_817, w_064_819, w_064_820, w_064_823, w_064_825, w_064_830, w_064_831, w_064_833, w_064_834, w_064_836, w_064_837, w_064_838, w_064_840, w_064_842, w_064_843, w_064_844, w_064_847, w_064_848, w_064_849, w_064_853, w_064_854, w_064_855, w_064_856, w_064_857, w_064_858, w_064_859, w_064_860, w_064_861, w_064_863, w_064_864, w_064_867, w_064_868, w_064_870, w_064_871, w_064_872, w_064_874, w_064_875, w_064_876, w_064_877, w_064_881, w_064_882, w_064_883, w_064_887, w_064_888, w_064_891, w_064_892, w_064_893, w_064_899, w_064_900, w_064_901, w_064_903, w_064_904, w_064_906, w_064_907, w_064_910, w_064_911, w_064_913, w_064_914, w_064_915, w_064_916, w_064_918, w_064_920, w_064_921, w_064_923, w_064_924, w_064_925, w_064_927, w_064_928, w_064_929, w_064_930, w_064_931, w_064_932, w_064_934, w_064_935, w_064_936, w_064_937, w_064_940, w_064_941, w_064_942, w_064_946, w_064_947, w_064_949, w_064_950, w_064_951, w_064_952, w_064_953, w_064_954, w_064_955, w_064_956, w_064_957, w_064_959, w_064_960, w_064_961, w_064_962, w_064_963, w_064_964, w_064_965, w_064_966, w_064_969, w_064_970, w_064_972, w_064_974, w_064_975, w_064_976, w_064_979, w_064_980, w_064_983, w_064_985, w_064_986, w_064_988, w_064_989, w_064_990, w_064_991, w_064_993, w_064_994, w_064_995, w_064_997, w_064_998, w_064_1000, w_064_1002, w_064_1003, w_064_1004, w_064_1005, w_064_1006, w_064_1010, w_064_1013, w_064_1014, w_064_1015, w_064_1017, w_064_1018, w_064_1019, w_064_1020, w_064_1021, w_064_1023, w_064_1024, w_064_1025, w_064_1028, w_064_1030, w_064_1031, w_064_1034, w_064_1035, w_064_1036, w_064_1039, w_064_1040, w_064_1043, w_064_1044, w_064_1045, w_064_1046, w_064_1048, w_064_1049, w_064_1051, w_064_1053, w_064_1054, w_064_1055, w_064_1056, w_064_1057, w_064_1058, w_064_1060, w_064_1061, w_064_1062, w_064_1063, w_064_1064, w_064_1065, w_064_1066, w_064_1067, w_064_1069, w_064_1072, w_064_1073, w_064_1074, w_064_1075, w_064_1076, w_064_1077, w_064_1079, w_064_1080, w_064_1081, w_064_1082, w_064_1083, w_064_1084, w_064_1086, w_064_1087, w_064_1088, w_064_1090, w_064_1091, w_064_1092, w_064_1093, w_064_1094, w_064_1095, w_064_1097, w_064_1099, w_064_1100, w_064_1101, w_064_1104, w_064_1105, w_064_1107, w_064_1108, w_064_1109, w_064_1110, w_064_1113, w_064_1115, w_064_1116, w_064_1118, w_064_1119, w_064_1123, w_064_1125, w_064_1126, w_064_1127, w_064_1128, w_064_1130, w_064_1131, w_064_1132, w_064_1133, w_064_1134, w_064_1137, w_064_1138, w_064_1139, w_064_1143, w_064_1144, w_064_1146, w_064_1147, w_064_1149, w_064_1150, w_064_1151, w_064_1153, w_064_1155, w_064_1156, w_064_1157, w_064_1158, w_064_1160, w_064_1162, w_064_1163, w_064_1164, w_064_1165, w_064_1167, w_064_1168, w_064_1170, w_064_1171, w_064_1172, w_064_1174, w_064_1175, w_064_1179, w_064_1180, w_064_1181, w_064_1182, w_064_1183, w_064_1184, w_064_1185, w_064_1186, w_064_1187, w_064_1188, w_064_1190, w_064_1191, w_064_1193, w_064_1195, w_064_1196, w_064_1198, w_064_1199, w_064_1202, w_064_1205, w_064_1207, w_064_1208, w_064_1210, w_064_1211, w_064_1212, w_064_1213, w_064_1215, w_064_1216, w_064_1220, w_064_1221, w_064_1222, w_064_1223, w_064_1224, w_064_1225, w_064_1226, w_064_1227, w_064_1228, w_064_1229, w_064_1230, w_064_1231, w_064_1232, w_064_1234, w_064_1235, w_064_1236, w_064_1237, w_064_1239, w_064_1240, w_064_1244, w_064_1245, w_064_1249, w_064_1250, w_064_1251, w_064_1255, w_064_1256, w_064_1257, w_064_1259, w_064_1260, w_064_1262, w_064_1263, w_064_1264, w_064_1266, w_064_1267, w_064_1268, w_064_1269, w_064_1272, w_064_1273, w_064_1274, w_064_1275, w_064_1276, w_064_1277, w_064_1278, w_064_1279, w_064_1281, w_064_1283, w_064_1284, w_064_1287, w_064_1288, w_064_1289, w_064_1291, w_064_1293, w_064_1295, w_064_1298, w_064_1299, w_064_1300, w_064_1301, w_064_1302, w_064_1304, w_064_1306, w_064_1308, w_064_1311, w_064_1312, w_064_1314, w_064_1316, w_064_1317, w_064_1318, w_064_1319, w_064_1320, w_064_1322, w_064_1323, w_064_1324, w_064_1327, w_064_1328, w_064_1329, w_064_1330, w_064_1331, w_064_1332, w_064_1333, w_064_1334, w_064_1336, w_064_1338, w_064_1340, w_064_1341, w_064_1343, w_064_1344, w_064_1345, w_064_1346, w_064_1347, w_064_1349, w_064_1351, w_064_1354, w_064_1356, w_064_1357, w_064_1358, w_064_1359, w_064_1360, w_064_1361, w_064_1362, w_064_1363, w_064_1364, w_064_1367, w_064_1368, w_064_1369, w_064_1370, w_064_1371, w_064_1372, w_064_1373, w_064_1376, w_064_1378, w_064_1379, w_064_1383, w_064_1384, w_064_1385, w_064_1388, w_064_1389, w_064_1394, w_064_1395, w_064_1396, w_064_1399, w_064_1400, w_064_1401, w_064_1402, w_064_1403, w_064_1408, w_064_1409, w_064_1411, w_064_1412, w_064_1413, w_064_1414, w_064_1415, w_064_1416, w_064_1417, w_064_1418, w_064_1419, w_064_1420, w_064_1421, w_064_1422, w_064_1424, w_064_1425, w_064_1426, w_064_1428, w_064_1429, w_064_1430, w_064_1431, w_064_1434, w_064_1436, w_064_1437, w_064_1438, w_064_1439, w_064_1441, w_064_1442, w_064_1444, w_064_1446, w_064_1447, w_064_1448, w_064_1450, w_064_1451, w_064_1452, w_064_1456, w_064_1457, w_064_1459, w_064_1460, w_064_1462, w_064_1463, w_064_1467, w_064_1468, w_064_1470, w_064_1473, w_064_1474, w_064_1475, w_064_1476, w_064_1480, w_064_1482, w_064_1485, w_064_1486, w_064_1489, w_064_1490, w_064_1491, w_064_1493, w_064_1494, w_064_1496, w_064_1497, w_064_1498, w_064_1499, w_064_1500, w_064_1503, w_064_1504, w_064_1505, w_064_1506, w_064_1509, w_064_1511, w_064_1514, w_064_1515, w_064_1517, w_064_1518, w_064_1519, w_064_1520, w_064_1521, w_064_1522, w_064_1523, w_064_1525, w_064_1526, w_064_1527, w_064_1528, w_064_1529, w_064_1530, w_064_1531, w_064_1533, w_064_1534, w_064_1536, w_064_1542, w_064_1544, w_064_1547, w_064_1551, w_064_1556, w_064_1557, w_064_1558, w_064_1563, w_064_1565, w_064_1566, w_064_1568, w_064_1573, w_064_1577, w_064_1578, w_064_1579, w_064_1581, w_064_1584, w_064_1589, w_064_1593, w_064_1596, w_064_1599, w_064_1602, w_064_1603, w_064_1607, w_064_1615, w_064_1617, w_064_1621, w_064_1628, w_064_1631, w_064_1633, w_064_1639, w_064_1640, w_064_1643, w_064_1644, w_064_1645, w_064_1648, w_064_1649, w_064_1650, w_064_1651, w_064_1655, w_064_1661, w_064_1663, w_064_1664, w_064_1665, w_064_1669, w_064_1670, w_064_1671, w_064_1672, w_064_1680, w_064_1682, w_064_1683, w_064_1686, w_064_1692, w_064_1693, w_064_1701, w_064_1702, w_064_1706, w_064_1707, w_064_1708, w_064_1709, w_064_1710, w_064_1713, w_064_1715, w_064_1718, w_064_1719, w_064_1721, w_064_1724, w_064_1728, w_064_1729, w_064_1730, w_064_1734, w_064_1736, w_064_1737, w_064_1738, w_064_1739, w_064_1740, w_064_1743, w_064_1745, w_064_1748, w_064_1753, w_064_1754, w_064_1757, w_064_1762, w_064_1764, w_064_1765, w_064_1766, w_064_1769, w_064_1771, w_064_1773, w_064_1774, w_064_1779, w_064_1786, w_064_1789, w_064_1791, w_064_1792, w_064_1793, w_064_1795, w_064_1797, w_064_1801, w_064_1802, w_064_1803, w_064_1805, w_064_1806, w_064_1812, w_064_1814, w_064_1815, w_064_1817, w_064_1819, w_064_1820, w_064_1822, w_064_1823, w_064_1824, w_064_1825, w_064_1827, w_064_1828, w_064_1830, w_064_1834, w_064_1836, w_064_1838, w_064_1839, w_064_1841, w_064_1843, w_064_1844, w_064_1847, w_064_1848, w_064_1849, w_064_1850, w_064_1851, w_064_1853, w_064_1858, w_064_1862, w_064_1863, w_064_1864, w_064_1867, w_064_1869, w_064_1873, w_064_1877, w_064_1886, w_064_1891, w_064_1894, w_064_1904, w_064_1905, w_064_1906, w_064_1917, w_064_1918, w_064_1919, w_064_1922, w_064_1927, w_064_1930, w_064_1931, w_064_1935, w_064_1937, w_064_1938, w_064_1939, w_064_1940, w_064_1944, w_064_1945, w_064_1946, w_064_1949, w_064_1950, w_064_1956, w_064_1964, w_064_1965, w_064_1969, w_064_1971, w_064_1976, w_064_1977, w_064_1979, w_064_1983, w_064_1984, w_064_1985, w_064_1986, w_064_1987, w_064_1988, w_064_1991, w_064_1992, w_064_1994, w_064_1995, w_064_1996, w_064_1997, w_064_2001, w_064_2002, w_064_2015, w_064_2016, w_064_2019, w_064_2022, w_064_2023, w_064_2026, w_064_2027, w_064_2029, w_064_2030, w_064_2033, w_064_2036, w_064_2037, w_064_2040, w_064_2044, w_064_2047, w_064_2049, w_064_2053, w_064_2056, w_064_2057, w_064_2058, w_064_2060, w_064_2061, w_064_2065, w_064_2068, w_064_2069, w_064_2075, w_064_2078, w_064_2079, w_064_2081, w_064_2082, w_064_2084, w_064_2085, w_064_2092, w_064_2093, w_064_2098, w_064_2101, w_064_2102, w_064_2103, w_064_2104, w_064_2105, w_064_2107, w_064_2108, w_064_2111, w_064_2115, w_064_2116, w_064_2118, w_064_2119, w_064_2120, w_064_2121, w_064_2122, w_064_2123, w_064_2127, w_064_2129, w_064_2130, w_064_2131, w_064_2132, w_064_2133, w_064_2148, w_064_2149, w_064_2150, w_064_2151, w_064_2152, w_064_2157, w_064_2159, w_064_2162, w_064_2163, w_064_2166, w_064_2168, w_064_2170, w_064_2171, w_064_2174, w_064_2176, w_064_2177, w_064_2179, w_064_2181, w_064_2182, w_064_2185, w_064_2186, w_064_2187, w_064_2193, w_064_2194, w_064_2195, w_064_2198, w_064_2199, w_064_2203, w_064_2205, w_064_2207, w_064_2208, w_064_2210, w_064_2216, w_064_2217, w_064_2218, w_064_2220, w_064_2221, w_064_2223, w_064_2225, w_064_2226, w_064_2235, w_064_2237, w_064_2238, w_064_2241, w_064_2242, w_064_2243, w_064_2248, w_064_2250, w_064_2256, w_064_2260, w_064_2261, w_064_2262, w_064_2264, w_064_2265, w_064_2267, w_064_2268, w_064_2271, w_064_2272, w_064_2274, w_064_2277, w_064_2280, w_064_2281, w_064_2282, w_064_2283, w_064_2284, w_064_2285, w_064_2286, w_064_2287, w_064_2289, w_064_2290, w_064_2291, w_064_2294, w_064_2297, w_064_2298, w_064_2304, w_064_2305, w_064_2310, w_064_2313, w_064_2314, w_064_2316, w_064_2317, w_064_2320, w_064_2324, w_064_2326, w_064_2331, w_064_2332, w_064_2333, w_064_2334, w_064_2337, w_064_2340, w_064_2341, w_064_2342, w_064_2344, w_064_2345, w_064_2348, w_064_2349, w_064_2350, w_064_2353, w_064_2354, w_064_2361, w_064_2363, w_064_2366, w_064_2371, w_064_2373, w_064_2378, w_064_2384, w_064_2385, w_064_2388, w_064_2389, w_064_2391, w_064_2392, w_064_2395, w_064_2397, w_064_2400, w_064_2402, w_064_2406, w_064_2408, w_064_2409, w_064_2410, w_064_2412, w_064_2414, w_064_2415, w_064_2419, w_064_2420, w_064_2421, w_064_2429, w_064_2431, w_064_2432, w_064_2433, w_064_2438, w_064_2443, w_064_2445, w_064_2447, w_064_2448, w_064_2451, w_064_2452, w_064_2453, w_064_2462, w_064_2465, w_064_2467, w_064_2470, w_064_2472, w_064_2473, w_064_2474, w_064_2476, w_064_2481, w_064_2483, w_064_2484, w_064_2485, w_064_2487, w_064_2488, w_064_2490, w_064_2492, w_064_2493, w_064_2498, w_064_2500, w_064_2503, w_064_2504, w_064_2505, w_064_2506, w_064_2507, w_064_2509, w_064_2512, w_064_2517, w_064_2519, w_064_2520, w_064_2521, w_064_2524, w_064_2525, w_064_2530, w_064_2534, w_064_2536, w_064_2537, w_064_2538, w_064_2539, w_064_2540, w_064_2542, w_064_2546, w_064_2549, w_064_2551, w_064_2555, w_064_2557, w_064_2560, w_064_2561, w_064_2565, w_064_2566, w_064_2570, w_064_2575, w_064_2576, w_064_2577, w_064_2579, w_064_2580, w_064_2581, w_064_2583, w_064_2584, w_064_2585, w_064_2587, w_064_2588, w_064_2591, w_064_2592, w_064_2596, w_064_2597, w_064_2598, w_064_2600, w_064_2603, w_064_2607, w_064_2614, w_064_2616, w_064_2618, w_064_2620, w_064_2624, w_064_2627, w_064_2628, w_064_2631, w_064_2632, w_064_2634, w_064_2636, w_064_2638, w_064_2644, w_064_2646, w_064_2647, w_064_2648, w_064_2649, w_064_2651, w_064_2653, w_064_2655, w_064_2659, w_064_2666, w_064_2669, w_064_2679, w_064_2683, w_064_2686, w_064_2690, w_064_2691, w_064_2695, w_064_2696, w_064_2697, w_064_2701, w_064_2706, w_064_2712, w_064_2717, w_064_2720, w_064_2723, w_064_2724, w_064_2725, w_064_2728, w_064_2730, w_064_2738, w_064_2741, w_064_2743, w_064_2744, w_064_2750, w_064_2755, w_064_2756, w_064_2757, w_064_2762, w_064_2763, w_064_2765, w_064_2770, w_064_2775, w_064_2776, w_064_2779, w_064_2780, w_064_2781, w_064_2782, w_064_2783, w_064_2786, w_064_2787, w_064_2794, w_064_2795, w_064_2797, w_064_2798, w_064_2801, w_064_2804, w_064_2805, w_064_2811, w_064_2815, w_064_2816, w_064_2820, w_064_2821, w_064_2822, w_064_2823, w_064_2824, w_064_2827, w_064_2831, w_064_2832, w_064_2833, w_064_2834, w_064_2835, w_064_2836, w_064_2837, w_064_2838, w_064_2839, w_064_2840, w_064_2842, w_064_2843, w_064_2845, w_064_2847, w_064_2849, w_064_2855, w_064_2856, w_064_2858, w_064_2859, w_064_2862, w_064_2870, w_064_2875, w_064_2879, w_064_2883, w_064_2885, w_064_2887, w_064_2890, w_064_2891, w_064_2896, w_064_2898, w_064_2900, w_064_2901, w_064_2902, w_064_2904, w_064_2905, w_064_2907, w_064_2911, w_064_2914, w_064_2915, w_064_2918, w_064_2922, w_064_2923, w_064_2924, w_064_2926, w_064_2928, w_064_2932, w_064_2934, w_064_2935, w_064_2939, w_064_2942, w_064_2944, w_064_2946, w_064_2948, w_064_2950, w_064_2953, w_064_2955, w_064_2956, w_064_2957, w_064_2964, w_064_2965, w_064_2966, w_064_2970, w_064_2972, w_064_2974, w_064_2976, w_064_2977, w_064_2979, w_064_2981, w_064_2982, w_064_2983, w_064_2984, w_064_2990, w_064_2991, w_064_2993, w_064_2995, w_064_2999, w_064_3001, w_064_3007, w_064_3008, w_064_3010, w_064_3014, w_064_3019, w_064_3020, w_064_3024, w_064_3029, w_064_3030, w_064_3032, w_064_3034, w_064_3042, w_064_3044, w_064_3048, w_064_3049, w_064_3050, w_064_3053, w_064_3061, w_064_3076, w_064_3077, w_064_3080, w_064_3083, w_064_3089, w_064_3090, w_064_3091, w_064_3092, w_064_3097, w_064_3098, w_064_3101, w_064_3102, w_064_3116, w_064_3118, w_064_3121, w_064_3122, w_064_3123, w_064_3124, w_064_3125, w_064_3131, w_064_3133, w_064_3135, w_064_3136, w_064_3137, w_064_3138, w_064_3141, w_064_3143, w_064_3144, w_064_3150, w_064_3151, w_064_3153, w_064_3159, w_064_3161, w_064_3162, w_064_3166, w_064_3168, w_064_3169, w_064_3170, w_064_3174, w_064_3176, w_064_3178, w_064_3179, w_064_3180, w_064_3181, w_064_3183, w_064_3184, w_064_3186, w_064_3188, w_064_3193, w_064_3199, w_064_3202, w_064_3204, w_064_3207, w_064_3208, w_064_3210, w_064_3211, w_064_3213, w_064_3215, w_064_3218, w_064_3219, w_064_3221, w_064_3222, w_064_3226, w_064_3228, w_064_3229, w_064_3233, w_064_3234, w_064_3238, w_064_3240, w_064_3241, w_064_3242, w_064_3247, w_064_3248, w_064_3250, w_064_3252, w_064_3253, w_064_3254, w_064_3257, w_064_3261, w_064_3262, w_064_3264, w_064_3265, w_064_3266, w_064_3267, w_064_3270, w_064_3272, w_064_3274, w_064_3275, w_064_3277, w_064_3278, w_064_3279, w_064_3281, w_064_3282, w_064_3286, w_064_3287, w_064_3289, w_064_3291, w_064_3292, w_064_3295, w_064_3296, w_064_3299, w_064_3303, w_064_3305, w_064_3310, w_064_3320, w_064_3321, w_064_3323, w_064_3325, w_064_3326, w_064_3329, w_064_3330, w_064_3333, w_064_3336, w_064_3338, w_064_3339, w_064_3340, w_064_3345, w_064_3351, w_064_3354, w_064_3356, w_064_3357, w_064_3361, w_064_3365, w_064_3367, w_064_3368, w_064_3371, w_064_3372, w_064_3374, w_064_3377, w_064_3379, w_064_3380, w_064_3385, w_064_3386, w_064_3389, w_064_3390, w_064_3399, w_064_3400, w_064_3405, w_064_3406, w_064_3407, w_064_3410, w_064_3414, w_064_3422, w_064_3424, w_064_3428, w_064_3429, w_064_3432, w_064_3433, w_064_3434, w_064_3438, w_064_3440, w_064_3441, w_064_3442, w_064_3443, w_064_3448, w_064_3449, w_064_3450, w_064_3451, w_064_3457, w_064_3460, w_064_3461, w_064_3463, w_064_3464, w_064_3466, w_064_3468;
  wire w_065_000, w_065_001, w_065_002, w_065_003, w_065_004, w_065_005, w_065_006, w_065_007, w_065_008, w_065_009, w_065_010, w_065_011, w_065_012, w_065_013, w_065_014, w_065_015, w_065_016, w_065_017, w_065_018, w_065_019, w_065_020, w_065_021, w_065_022, w_065_023, w_065_024, w_065_025, w_065_026, w_065_027, w_065_028, w_065_029, w_065_030, w_065_031, w_065_032, w_065_033, w_065_034, w_065_035, w_065_036, w_065_037, w_065_038, w_065_039, w_065_040, w_065_041, w_065_042, w_065_043, w_065_044, w_065_045, w_065_046, w_065_047, w_065_048, w_065_049, w_065_050, w_065_051, w_065_052, w_065_053, w_065_054, w_065_055, w_065_056, w_065_057, w_065_058, w_065_059, w_065_060, w_065_061, w_065_062, w_065_063, w_065_064, w_065_065, w_065_066, w_065_067, w_065_068, w_065_069, w_065_070, w_065_071, w_065_072, w_065_073, w_065_074, w_065_075, w_065_076, w_065_077, w_065_078, w_065_079, w_065_080, w_065_081, w_065_082, w_065_083, w_065_084, w_065_085, w_065_086, w_065_087, w_065_088, w_065_089, w_065_090, w_065_091, w_065_092, w_065_093, w_065_094, w_065_095, w_065_096, w_065_097, w_065_098, w_065_099, w_065_100, w_065_101, w_065_102, w_065_103, w_065_104, w_065_105, w_065_106, w_065_107, w_065_108, w_065_109, w_065_110, w_065_111, w_065_112, w_065_113, w_065_114, w_065_115, w_065_116, w_065_117, w_065_118;
  wire w_066_000, w_066_002, w_066_004, w_066_005, w_066_006, w_066_007, w_066_008, w_066_009, w_066_010, w_066_012, w_066_013, w_066_014, w_066_015, w_066_016, w_066_021, w_066_022, w_066_024, w_066_027, w_066_029, w_066_030, w_066_031, w_066_032, w_066_033, w_066_034, w_066_035, w_066_036, w_066_039, w_066_041, w_066_043, w_066_044, w_066_047, w_066_048, w_066_049, w_066_050, w_066_051, w_066_052, w_066_053, w_066_054, w_066_056, w_066_057, w_066_065, w_066_066, w_066_067, w_066_069, w_066_073, w_066_074, w_066_077, w_066_079, w_066_082, w_066_084, w_066_085, w_066_087, w_066_088, w_066_089, w_066_093, w_066_094, w_066_097, w_066_098, w_066_100, w_066_101, w_066_102, w_066_103, w_066_105, w_066_106, w_066_108, w_066_111, w_066_113, w_066_115, w_066_116, w_066_118, w_066_120, w_066_121, w_066_123, w_066_124, w_066_125, w_066_126, w_066_127, w_066_128, w_066_129, w_066_130, w_066_133, w_066_134, w_066_135, w_066_136, w_066_138, w_066_139, w_066_140, w_066_141, w_066_142, w_066_143, w_066_144, w_066_145, w_066_146, w_066_148, w_066_150, w_066_151, w_066_152, w_066_153, w_066_154, w_066_157, w_066_159, w_066_160, w_066_163, w_066_164, w_066_167, w_066_168, w_066_169, w_066_170, w_066_171, w_066_172, w_066_174, w_066_176, w_066_177, w_066_179, w_066_180, w_066_182, w_066_183, w_066_184, w_066_185, w_066_187, w_066_188, w_066_189, w_066_191, w_066_192, w_066_194, w_066_197, w_066_198, w_066_200, w_066_201, w_066_202, w_066_203, w_066_204, w_066_206, w_066_209, w_066_210, w_066_213, w_066_214, w_066_215, w_066_217, w_066_218, w_066_219, w_066_221, w_066_224, w_066_226, w_066_228, w_066_230, w_066_231, w_066_232, w_066_233, w_066_234, w_066_239, w_066_241, w_066_242, w_066_243, w_066_244, w_066_248, w_066_249, w_066_250, w_066_251, w_066_252, w_066_254, w_066_255, w_066_256, w_066_257, w_066_259, w_066_260, w_066_261, w_066_262, w_066_263, w_066_264, w_066_266, w_066_267, w_066_268, w_066_269, w_066_271, w_066_272, w_066_274, w_066_275, w_066_277, w_066_281, w_066_282, w_066_286, w_066_287, w_066_288, w_066_289, w_066_290, w_066_291, w_066_292, w_066_293, w_066_295, w_066_296, w_066_298, w_066_299, w_066_300, w_066_301, w_066_304, w_066_305, w_066_306, w_066_307, w_066_308, w_066_309, w_066_310, w_066_312, w_066_313, w_066_314, w_066_315, w_066_316, w_066_317, w_066_318, w_066_319, w_066_320, w_066_321, w_066_323, w_066_325, w_066_326, w_066_327, w_066_330, w_066_331, w_066_333, w_066_336, w_066_337, w_066_339, w_066_340, w_066_341, w_066_342, w_066_344, w_066_346, w_066_347, w_066_348, w_066_351, w_066_352, w_066_353, w_066_354, w_066_359, w_066_364, w_066_365, w_066_366, w_066_367, w_066_368, w_066_369, w_066_372, w_066_373, w_066_374, w_066_377, w_066_380, w_066_381, w_066_382, w_066_384, w_066_385, w_066_386, w_066_387, w_066_389, w_066_391, w_066_393, w_066_394, w_066_397, w_066_398, w_066_399, w_066_401, w_066_404, w_066_407, w_066_409, w_066_411, w_066_412, w_066_415, w_066_416, w_066_417, w_066_419, w_066_422, w_066_424, w_066_426, w_066_427, w_066_428, w_066_429, w_066_430, w_066_431, w_066_433, w_066_434, w_066_442, w_066_444, w_066_445, w_066_446, w_066_447, w_066_448, w_066_449, w_066_451, w_066_453, w_066_454, w_066_455, w_066_457, w_066_458, w_066_459, w_066_460, w_066_462, w_066_463, w_066_465, w_066_466, w_066_467, w_066_469, w_066_471, w_066_472, w_066_473, w_066_475, w_066_479, w_066_481, w_066_482, w_066_483, w_066_484, w_066_486, w_066_487, w_066_491, w_066_492, w_066_493, w_066_494, w_066_497, w_066_498, w_066_499, w_066_500, w_066_502, w_066_506, w_066_507, w_066_510, w_066_512, w_066_513, w_066_514, w_066_515, w_066_516, w_066_518, w_066_522, w_066_523, w_066_524, w_066_525, w_066_526, w_066_527, w_066_529, w_066_531, w_066_534, w_066_535, w_066_537, w_066_538, w_066_540, w_066_541, w_066_542, w_066_546, w_066_547, w_066_548, w_066_549, w_066_550, w_066_552, w_066_553, w_066_556, w_066_560, w_066_562, w_066_565, w_066_566, w_066_568, w_066_569, w_066_571, w_066_572, w_066_574, w_066_575, w_066_576, w_066_580, w_066_581, w_066_582, w_066_583, w_066_585, w_066_586, w_066_591, w_066_592, w_066_593, w_066_594, w_066_595, w_066_597, w_066_600, w_066_601, w_066_602, w_066_603, w_066_606, w_066_609, w_066_611, w_066_613, w_066_614, w_066_615, w_066_619, w_066_620, w_066_621, w_066_622, w_066_624, w_066_627, w_066_629, w_066_630, w_066_631, w_066_632, w_066_633, w_066_634, w_066_635, w_066_637, w_066_638, w_066_639, w_066_640, w_066_641, w_066_643, w_066_646, w_066_647, w_066_648, w_066_649, w_066_651, w_066_652, w_066_653, w_066_655, w_066_657, w_066_658, w_066_661, w_066_663, w_066_666, w_066_668, w_066_669, w_066_670, w_066_671, w_066_675, w_066_676, w_066_678, w_066_679, w_066_680, w_066_682, w_066_684, w_066_686, w_066_689, w_066_694, w_066_697, w_066_698, w_066_703, w_066_704, w_066_705, w_066_706, w_066_708, w_066_709, w_066_710, w_066_711, w_066_712, w_066_713, w_066_714, w_066_716, w_066_717, w_066_718, w_066_720, w_066_721, w_066_723, w_066_724, w_066_727, w_066_728, w_066_729, w_066_730, w_066_731, w_066_732, w_066_734, w_066_737, w_066_738, w_066_740, w_066_741, w_066_742, w_066_744, w_066_745, w_066_746, w_066_747, w_066_750, w_066_752, w_066_754, w_066_755, w_066_756, w_066_757, w_066_758, w_066_759, w_066_760, w_066_761, w_066_764, w_066_765, w_066_767, w_066_768, w_066_769, w_066_770, w_066_771, w_066_773, w_066_774, w_066_776, w_066_780, w_066_781, w_066_782, w_066_784, w_066_785, w_066_786, w_066_788, w_066_789, w_066_790, w_066_791, w_066_792, w_066_793, w_066_794, w_066_796, w_066_797, w_066_798, w_066_799, w_066_800, w_066_802, w_066_803, w_066_804, w_066_805, w_066_806, w_066_807, w_066_808, w_066_809, w_066_810, w_066_811, w_066_812, w_066_813, w_066_814, w_066_815, w_066_816, w_066_818, w_066_819, w_066_822, w_066_823, w_066_826, w_066_827, w_066_828, w_066_831, w_066_832, w_066_833, w_066_834, w_066_835, w_066_836, w_066_837, w_066_838, w_066_841, w_066_842, w_066_843, w_066_844, w_066_845, w_066_846, w_066_848, w_066_849, w_066_850, w_066_851, w_066_852, w_066_853, w_066_854, w_066_855, w_066_856, w_066_857, w_066_859, w_066_864, w_066_865, w_066_866, w_066_868, w_066_871, w_066_872, w_066_874, w_066_875, w_066_877, w_066_880, w_066_881, w_066_882, w_066_883, w_066_884, w_066_885, w_066_886, w_066_888, w_066_890, w_066_892, w_066_895, w_066_897, w_066_900, w_066_902, w_066_903, w_066_907, w_066_909, w_066_910, w_066_911, w_066_912, w_066_913, w_066_914, w_066_916, w_066_919, w_066_921, w_066_922, w_066_925, w_066_926, w_066_927, w_066_928, w_066_929, w_066_931, w_066_932, w_066_933, w_066_935, w_066_936, w_066_937, w_066_939, w_066_940, w_066_941, w_066_942, w_066_943, w_066_945, w_066_946, w_066_948, w_066_951, w_066_952, w_066_953, w_066_954, w_066_955, w_066_957, w_066_959, w_066_962, w_066_965, w_066_967, w_066_968, w_066_969, w_066_972, w_066_973, w_066_974, w_066_975, w_066_976, w_066_980, w_066_981, w_066_982, w_066_983, w_066_991, w_066_992, w_066_993, w_066_994, w_066_995, w_066_996, w_066_997, w_066_1002, w_066_1003, w_066_1004, w_066_1005, w_066_1006, w_066_1009, w_066_1010, w_066_1011, w_066_1013, w_066_1014, w_066_1019, w_066_1021, w_066_1022, w_066_1025, w_066_1026, w_066_1028, w_066_1030, w_066_1031, w_066_1032, w_066_1035, w_066_1037, w_066_1038, w_066_1039, w_066_1040, w_066_1043, w_066_1046, w_066_1047, w_066_1050, w_066_1052, w_066_1058, w_066_1059, w_066_1062, w_066_1063, w_066_1064, w_066_1066, w_066_1067, w_066_1068, w_066_1069, w_066_1070, w_066_1071, w_066_1072, w_066_1073, w_066_1074, w_066_1075, w_066_1076, w_066_1077, w_066_1078, w_066_1079, w_066_1083, w_066_1086, w_066_1087, w_066_1088, w_066_1090, w_066_1091, w_066_1095, w_066_1097, w_066_1098, w_066_1099, w_066_1100, w_066_1102, w_066_1103, w_066_1104, w_066_1105, w_066_1108, w_066_1110, w_066_1111, w_066_1112, w_066_1114, w_066_1116, w_066_1120, w_066_1121, w_066_1123, w_066_1124, w_066_1127, w_066_1129, w_066_1130, w_066_1131, w_066_1134, w_066_1136, w_066_1138, w_066_1140, w_066_1144, w_066_1146, w_066_1147, w_066_1148, w_066_1150, w_066_1151, w_066_1154, w_066_1157, w_066_1158, w_066_1164, w_066_1170, w_066_1172, w_066_1174, w_066_1175, w_066_1176, w_066_1177, w_066_1178, w_066_1179, w_066_1180, w_066_1183, w_066_1184, w_066_1185, w_066_1186, w_066_1187, w_066_1188, w_066_1190, w_066_1194, w_066_1195, w_066_1197, w_066_1198, w_066_1199, w_066_1200, w_066_1201, w_066_1202, w_066_1205, w_066_1206, w_066_1208, w_066_1209, w_066_1210, w_066_1211, w_066_1212, w_066_1213, w_066_1214, w_066_1216, w_066_1219, w_066_1220, w_066_1221, w_066_1224, w_066_1225, w_066_1226, w_066_1228, w_066_1229, w_066_1230, w_066_1235, w_066_1237, w_066_1238, w_066_1239, w_066_1241, w_066_1243, w_066_1245, w_066_1247, w_066_1248, w_066_1249, w_066_1253, w_066_1254, w_066_1255, w_066_1256, w_066_1258, w_066_1260, w_066_1262, w_066_1264, w_066_1265, w_066_1268, w_066_1269, w_066_1270, w_066_1273, w_066_1274, w_066_1275, w_066_1276, w_066_1277, w_066_1278, w_066_1281, w_066_1282, w_066_1285, w_066_1288, w_066_1290, w_066_1291, w_066_1293, w_066_1295, w_066_1298, w_066_1299, w_066_1300, w_066_1302, w_066_1303, w_066_1304, w_066_1305, w_066_1306, w_066_1307, w_066_1308, w_066_1309, w_066_1314, w_066_1316, w_066_1317, w_066_1319, w_066_1320, w_066_1322, w_066_1325, w_066_1326, w_066_1327, w_066_1331, w_066_1335, w_066_1336, w_066_1337, w_066_1338, w_066_1339, w_066_1340, w_066_1342, w_066_1345, w_066_1347, w_066_1348, w_066_1350, w_066_1351, w_066_1354, w_066_1356, w_066_1357, w_066_1358, w_066_1359, w_066_1360, w_066_1361, w_066_1365, w_066_1366, w_066_1367, w_066_1368, w_066_1369, w_066_1370, w_066_1371, w_066_1372, w_066_1374, w_066_1377, w_066_1378, w_066_1381, w_066_1382, w_066_1384, w_066_1387, w_066_1389, w_066_1390, w_066_1391, w_066_1393, w_066_1394, w_066_1395, w_066_1396, w_066_1398, w_066_1399, w_066_1400, w_066_1404, w_066_1407, w_066_1408, w_066_1410, w_066_1411, w_066_1412, w_066_1413, w_066_1415, w_066_1416, w_066_1417, w_066_1419, w_066_1420, w_066_1421, w_066_1422, w_066_1423, w_066_1424, w_066_1425, w_066_1427, w_066_1428, w_066_1429, w_066_1430, w_066_1431, w_066_1433, w_066_1434, w_066_1436, w_066_1437, w_066_1440, w_066_1442, w_066_1443, w_066_1446, w_066_1449, w_066_1450, w_066_1452, w_066_1454, w_066_1457, w_066_1460, w_066_1461, w_066_1463, w_066_1464, w_066_1465, w_066_1466, w_066_1468, w_066_1469, w_066_1470, w_066_1471, w_066_1473, w_066_1477, w_066_1479, w_066_1480, w_066_1484, w_066_1485, w_066_1488, w_066_1490, w_066_1491, w_066_1493, w_066_1494, w_066_1496, w_066_1498, w_066_1499, w_066_1500, w_066_1501, w_066_1502, w_066_1503, w_066_1504, w_066_1505, w_066_1506, w_066_1510, w_066_1512, w_066_1513, w_066_1514, w_066_1515, w_066_1516, w_066_1517, w_066_1518, w_066_1521, w_066_1522, w_066_1525, w_066_1526, w_066_1528, w_066_1530, w_066_1532, w_066_1533, w_066_1534, w_066_1535, w_066_1536, w_066_1538, w_066_1540, w_066_1541, w_066_1542, w_066_1544, w_066_1545, w_066_1546, w_066_1547, w_066_1549, w_066_1550, w_066_1551, w_066_1554, w_066_1555, w_066_1557, w_066_1558, w_066_1559, w_066_1560, w_066_1561, w_066_1563, w_066_1564, w_066_1567, w_066_1569, w_066_1572, w_066_1573, w_066_1577, w_066_1579, w_066_1582, w_066_1583, w_066_1587, w_066_1589, w_066_1590, w_066_1591, w_066_1592, w_066_1596, w_066_1597, w_066_1599, w_066_1600, w_066_1602, w_066_1603, w_066_1605, w_066_1606, w_066_1607, w_066_1611, w_066_1612, w_066_1613, w_066_1615, w_066_1618, w_066_1619, w_066_1621, w_066_1624, w_066_1625, w_066_1628, w_066_1629, w_066_1631, w_066_1633, w_066_1634, w_066_1635, w_066_1636, w_066_1638, w_066_1639, w_066_1641, w_066_1646, w_066_1647, w_066_1650, w_066_1655, w_066_1656, w_066_1657, w_066_1659, w_066_1661, w_066_1663, w_066_1664, w_066_1667, w_066_1668, w_066_1671, w_066_1674, w_066_1677, w_066_1679, w_066_1680, w_066_1682, w_066_1683, w_066_1684, w_066_1686, w_066_1687, w_066_1688, w_066_1689, w_066_1691, w_066_1695, w_066_1696, w_066_1697, w_066_1700, w_066_1701, w_066_1704, w_066_1709, w_066_1710, w_066_1713, w_066_1714, w_066_1715, w_066_1716, w_066_1717, w_066_1718, w_066_1722, w_066_1725, w_066_1727, w_066_1731, w_066_1732, w_066_1735, w_066_1736, w_066_1739, w_066_1740, w_066_1741, w_066_1742, w_066_1744, w_066_1745, w_066_1746, w_066_1747, w_066_1748, w_066_1749, w_066_1750, w_066_1753, w_066_1755, w_066_1756, w_066_1757, w_066_1758, w_066_1759, w_066_1760, w_066_1762, w_066_1763, w_066_1764, w_066_1765, w_066_1767, w_066_1768, w_066_1769, w_066_1770, w_066_1771, w_066_1772, w_066_1773, w_066_1775, w_066_1776, w_066_1778, w_066_1779, w_066_1782, w_066_1784, w_066_1785, w_066_1786, w_066_1789, w_066_1790, w_066_1791, w_066_1792, w_066_1795, w_066_1796, w_066_1797, w_066_1801, w_066_1802, w_066_1803, w_066_1804, w_066_1806, w_066_1807, w_066_1808, w_066_1809, w_066_1810, w_066_1812, w_066_1813, w_066_1814, w_066_1817, w_066_1820, w_066_1821, w_066_1822, w_066_1828, w_066_1830, w_066_1832, w_066_1833, w_066_1834, w_066_1837, w_066_1838, w_066_1839, w_066_1840, w_066_1841, w_066_1842, w_066_1844, w_066_1845, w_066_1849, w_066_1850, w_066_1851, w_066_1852, w_066_1853, w_066_1856, w_066_1857, w_066_1858, w_066_1859, w_066_1860, w_066_1861, w_066_1862, w_066_1863, w_066_1866, w_066_1868, w_066_1869, w_066_1870, w_066_1872, w_066_1873, w_066_1875, w_066_1880, w_066_1881, w_066_1882, w_066_1885, w_066_1888, w_066_1889, w_066_1890, w_066_1892, w_066_1893, w_066_1895, w_066_1896, w_066_1897, w_066_1900, w_066_1901, w_066_1902, w_066_1904, w_066_1905, w_066_1906, w_066_1907, w_066_1908, w_066_1909, w_066_1910, w_066_1911, w_066_1912, w_066_1914, w_066_1915, w_066_1916, w_066_1918, w_066_1919, w_066_1922, w_066_1923, w_066_1925, w_066_1926, w_066_1928, w_066_1930, w_066_1932, w_066_1933, w_066_1935, w_066_1937, w_066_1938, w_066_1939, w_066_1940, w_066_1941, w_066_1943, w_066_1945, w_066_1947, w_066_1950, w_066_1951, w_066_1952, w_066_1953, w_066_1957, w_066_1958, w_066_1962, w_066_1963, w_066_1964, w_066_1965, w_066_1966, w_066_1969, w_066_1971, w_066_1972, w_066_1974, w_066_1977, w_066_1979, w_066_1980, w_066_1981, w_066_1982, w_066_1983, w_066_1984, w_066_1985, w_066_1986, w_066_1987, w_066_1992, w_066_1997, w_066_1998, w_066_2001, w_066_2002, w_066_2003, w_066_2004, w_066_2005, w_066_2007, w_066_2009, w_066_2013, w_066_2014, w_066_2015, w_066_2016, w_066_2017, w_066_2018, w_066_2019, w_066_2020, w_066_2021, w_066_2024, w_066_2025, w_066_2026, w_066_2027, w_066_2028, w_066_2032, w_066_2033, w_066_2034, w_066_2035, w_066_2036, w_066_2037, w_066_2038, w_066_2039, w_066_2040, w_066_2041, w_066_2042, w_066_2044, w_066_2046, w_066_2048, w_066_2049, w_066_2051, w_066_2054, w_066_2055, w_066_2057, w_066_2058, w_066_2059, w_066_2060, w_066_2062, w_066_2063, w_066_2065, w_066_2067, w_066_2068, w_066_2071, w_066_2074, w_066_2075, w_066_2076, w_066_2079, w_066_2082, w_066_2083, w_066_2084, w_066_2085, w_066_2086, w_066_2087, w_066_2088, w_066_2089, w_066_2091, w_066_2092, w_066_2093, w_066_2094, w_066_2095, w_066_2097, w_066_2098, w_066_2099, w_066_2101, w_066_2102, w_066_2105, w_066_2106, w_066_2107, w_066_2108, w_066_2109, w_066_2111, w_066_2113, w_066_2117, w_066_2120, w_066_2122, w_066_2126, w_066_2127, w_066_2132, w_066_2133, w_066_2134, w_066_2138, w_066_2139, w_066_2140, w_066_2141, w_066_2146, w_066_2147, w_066_2148, w_066_2150, w_066_2152, w_066_2154, w_066_2155, w_066_2157, w_066_2161, w_066_2162, w_066_2164, w_066_2165, w_066_2166, w_066_2167, w_066_2168, w_066_2170, w_066_2171, w_066_2173, w_066_2175, w_066_2176, w_066_2180, w_066_2183, w_066_2184, w_066_2189, w_066_2190, w_066_2192, w_066_2196, w_066_2198, w_066_2205, w_066_2209, w_066_2211, w_066_2212, w_066_2215, w_066_2216, w_066_2219, w_066_2228, w_066_2229, w_066_2231, w_066_2235, w_066_2238, w_066_2239, w_066_2243, w_066_2244, w_066_2247, w_066_2249, w_066_2251, w_066_2252, w_066_2253, w_066_2259, w_066_2263, w_066_2265, w_066_2268, w_066_2274, w_066_2275, w_066_2278, w_066_2284, w_066_2286, w_066_2295, w_066_2299, w_066_2300, w_066_2301, w_066_2302, w_066_2306, w_066_2307, w_066_2308, w_066_2312, w_066_2316, w_066_2317, w_066_2319, w_066_2321, w_066_2327, w_066_2330, w_066_2331, w_066_2332, w_066_2333, w_066_2335, w_066_2337, w_066_2339, w_066_2340, w_066_2347, w_066_2351, w_066_2355, w_066_2357, w_066_2358, w_066_2359, w_066_2360, w_066_2361, w_066_2362, w_066_2364, w_066_2366, w_066_2368, w_066_2369, w_066_2378, w_066_2379, w_066_2380, w_066_2381, w_066_2382, w_066_2386, w_066_2387, w_066_2397, w_066_2399, w_066_2405, w_066_2410, w_066_2412, w_066_2415, w_066_2420, w_066_2423, w_066_2425, w_066_2426, w_066_2433, w_066_2435, w_066_2438, w_066_2440, w_066_2442, w_066_2445, w_066_2454, w_066_2457, w_066_2459, w_066_2460, w_066_2463, w_066_2464, w_066_2465, w_066_2467, w_066_2468, w_066_2469, w_066_2471, w_066_2472, w_066_2473, w_066_2475, w_066_2476, w_066_2479, w_066_2485, w_066_2488, w_066_2492, w_066_2494, w_066_2503, w_066_2506, w_066_2510, w_066_2511, w_066_2517, w_066_2519, w_066_2523, w_066_2526, w_066_2531, w_066_2532, w_066_2533, w_066_2534, w_066_2537, w_066_2538, w_066_2539, w_066_2543, w_066_2552, w_066_2554, w_066_2556, w_066_2557, w_066_2558, w_066_2559, w_066_2561, w_066_2564, w_066_2570, w_066_2574, w_066_2576, w_066_2577, w_066_2578, w_066_2581, w_066_2582, w_066_2584, w_066_2588, w_066_2594, w_066_2597, w_066_2605, w_066_2609, w_066_2617, w_066_2618, w_066_2622, w_066_2623, w_066_2625, w_066_2627, w_066_2633, w_066_2636, w_066_2644, w_066_2645, w_066_2646, w_066_2651, w_066_2653, w_066_2656, w_066_2659, w_066_2665, w_066_2667, w_066_2669, w_066_2670, w_066_2671, w_066_2672, w_066_2676, w_066_2679, w_066_2680, w_066_2685, w_066_2686, w_066_2692, w_066_2695, w_066_2697, w_066_2700, w_066_2701, w_066_2702, w_066_2706, w_066_2708, w_066_2710, w_066_2713, w_066_2714, w_066_2717, w_066_2719, w_066_2720, w_066_2722, w_066_2725, w_066_2729, w_066_2734, w_066_2735, w_066_2740, w_066_2743, w_066_2746, w_066_2748, w_066_2749, w_066_2750, w_066_2753, w_066_2755, w_066_2758, w_066_2759, w_066_2761, w_066_2762, w_066_2763, w_066_2765, w_066_2766, w_066_2768, w_066_2777, w_066_2778, w_066_2779, w_066_2784, w_066_2791, w_066_2792, w_066_2794, w_066_2798, w_066_2802, w_066_2804, w_066_2806, w_066_2808, w_066_2809, w_066_2811, w_066_2814, w_066_2818, w_066_2824, w_066_2834, w_066_2838, w_066_2840, w_066_2843, w_066_2845, w_066_2846, w_066_2847, w_066_2849, w_066_2850, w_066_2854, w_066_2855, w_066_2856, w_066_2857, w_066_2858, w_066_2859, w_066_2860, w_066_2861, w_066_2865, w_066_2866, w_066_2867, w_066_2868, w_066_2869, w_066_2871;
  wire w_067_001, w_067_003, w_067_004, w_067_005, w_067_007, w_067_008, w_067_011, w_067_012, w_067_015, w_067_016, w_067_017, w_067_018, w_067_019, w_067_020, w_067_021, w_067_022, w_067_023, w_067_024, w_067_025, w_067_026, w_067_033, w_067_034, w_067_035, w_067_036, w_067_037, w_067_038, w_067_039, w_067_040, w_067_043, w_067_044, w_067_046, w_067_047, w_067_050, w_067_053, w_067_055, w_067_056, w_067_057, w_067_059, w_067_060, w_067_061, w_067_064, w_067_069, w_067_070, w_067_072, w_067_073, w_067_074, w_067_076, w_067_077, w_067_078, w_067_079, w_067_080, w_067_081, w_067_082, w_067_085, w_067_086, w_067_087, w_067_088, w_067_089, w_067_090, w_067_092, w_067_093, w_067_095, w_067_096, w_067_097, w_067_100, w_067_101, w_067_102, w_067_103, w_067_104, w_067_105, w_067_106, w_067_109, w_067_117, w_067_119, w_067_120, w_067_121, w_067_123, w_067_125, w_067_129, w_067_131, w_067_132, w_067_133, w_067_134, w_067_135, w_067_137, w_067_142, w_067_143, w_067_149, w_067_151, w_067_153, w_067_154, w_067_158, w_067_159, w_067_161, w_067_164, w_067_169, w_067_170, w_067_171, w_067_172, w_067_173, w_067_174, w_067_175, w_067_178, w_067_183, w_067_189, w_067_192, w_067_194, w_067_197, w_067_201, w_067_203, w_067_209, w_067_210, w_067_211, w_067_219, w_067_225, w_067_232, w_067_234, w_067_235, w_067_242, w_067_244, w_067_245, w_067_247, w_067_249, w_067_251, w_067_252, w_067_254, w_067_257, w_067_261, w_067_264, w_067_268, w_067_269, w_067_271, w_067_272, w_067_275, w_067_276, w_067_281, w_067_282, w_067_284, w_067_285, w_067_286, w_067_295, w_067_297, w_067_302, w_067_304, w_067_305, w_067_313, w_067_316, w_067_318, w_067_320, w_067_324, w_067_325, w_067_328, w_067_329, w_067_334, w_067_342, w_067_348, w_067_352, w_067_354, w_067_355, w_067_358, w_067_359, w_067_364, w_067_367, w_067_368, w_067_372, w_067_373, w_067_376, w_067_377, w_067_383, w_067_386, w_067_387, w_067_388, w_067_395, w_067_396, w_067_397, w_067_405, w_067_407, w_067_408, w_067_415, w_067_418, w_067_419, w_067_420, w_067_422, w_067_424, w_067_429, w_067_436, w_067_438, w_067_439, w_067_440, w_067_442, w_067_443, w_067_449, w_067_450, w_067_459, w_067_463, w_067_465, w_067_470, w_067_472, w_067_476, w_067_480, w_067_483, w_067_484, w_067_485, w_067_487, w_067_491, w_067_493, w_067_495, w_067_499, w_067_500, w_067_503, w_067_505, w_067_506, w_067_511, w_067_512, w_067_513, w_067_514, w_067_515, w_067_516, w_067_520, w_067_521, w_067_529, w_067_531, w_067_536, w_067_537, w_067_540, w_067_542, w_067_543, w_067_544, w_067_546, w_067_549, w_067_550, w_067_551, w_067_552, w_067_553, w_067_555, w_067_556, w_067_557, w_067_558, w_067_560, w_067_561, w_067_563, w_067_567, w_067_572, w_067_574, w_067_576, w_067_580, w_067_581, w_067_585, w_067_589, w_067_590, w_067_591, w_067_592, w_067_593, w_067_594, w_067_595, w_067_598, w_067_601, w_067_602, w_067_603, w_067_605, w_067_606, w_067_607, w_067_611, w_067_617, w_067_619, w_067_621, w_067_625, w_067_626, w_067_627, w_067_631, w_067_635, w_067_639, w_067_640, w_067_644, w_067_647, w_067_648, w_067_650, w_067_656, w_067_660, w_067_667, w_067_669, w_067_675, w_067_676, w_067_681, w_067_686, w_067_689, w_067_695, w_067_696, w_067_699, w_067_702, w_067_705, w_067_707, w_067_709, w_067_711, w_067_718, w_067_721, w_067_722, w_067_724, w_067_725, w_067_727, w_067_729, w_067_732, w_067_733, w_067_735, w_067_736, w_067_738, w_067_739, w_067_741, w_067_744, w_067_746, w_067_748, w_067_750, w_067_768, w_067_770, w_067_773, w_067_775, w_067_778, w_067_782, w_067_783, w_067_784, w_067_785, w_067_787, w_067_789, w_067_794, w_067_795, w_067_797, w_067_798, w_067_799, w_067_802, w_067_809, w_067_812, w_067_814, w_067_815, w_067_818, w_067_820, w_067_823, w_067_824, w_067_828, w_067_831, w_067_834, w_067_840, w_067_843, w_067_846, w_067_847, w_067_853, w_067_855, w_067_856, w_067_857, w_067_859, w_067_861, w_067_865, w_067_869, w_067_876, w_067_878, w_067_881, w_067_882, w_067_884, w_067_893, w_067_896, w_067_901, w_067_902, w_067_909, w_067_910, w_067_915, w_067_918, w_067_922, w_067_924, w_067_929, w_067_932, w_067_933, w_067_936, w_067_938, w_067_945, w_067_948, w_067_949, w_067_950, w_067_952, w_067_956, w_067_957, w_067_958, w_067_961, w_067_962, w_067_964, w_067_966, w_067_972, w_067_975, w_067_976, w_067_983, w_067_987, w_067_992, w_067_993, w_067_994, w_067_996, w_067_999, w_067_1000, w_067_1001, w_067_1003, w_067_1007, w_067_1009, w_067_1010, w_067_1013, w_067_1016, w_067_1018, w_067_1020, w_067_1021, w_067_1022, w_067_1024, w_067_1028, w_067_1029, w_067_1032, w_067_1037, w_067_1043, w_067_1045, w_067_1046, w_067_1047, w_067_1048, w_067_1049, w_067_1050, w_067_1053, w_067_1054, w_067_1056, w_067_1061, w_067_1063, w_067_1066, w_067_1067, w_067_1071, w_067_1072, w_067_1076, w_067_1077, w_067_1085, w_067_1089, w_067_1091, w_067_1092, w_067_1093, w_067_1094, w_067_1096, w_067_1099, w_067_1100, w_067_1101, w_067_1103, w_067_1104, w_067_1113, w_067_1118, w_067_1119, w_067_1120, w_067_1132, w_067_1135, w_067_1137, w_067_1141, w_067_1143, w_067_1144, w_067_1147, w_067_1152, w_067_1154, w_067_1156, w_067_1158, w_067_1160, w_067_1163, w_067_1169, w_067_1171, w_067_1172, w_067_1173, w_067_1177, w_067_1178, w_067_1181, w_067_1183, w_067_1186, w_067_1187, w_067_1190, w_067_1192, w_067_1196, w_067_1199, w_067_1200, w_067_1204, w_067_1205, w_067_1208, w_067_1209, w_067_1212, w_067_1213, w_067_1216, w_067_1217, w_067_1222, w_067_1231, w_067_1233, w_067_1235, w_067_1236, w_067_1239, w_067_1240, w_067_1250, w_067_1254, w_067_1256, w_067_1268, w_067_1274, w_067_1275, w_067_1276, w_067_1279, w_067_1280, w_067_1288, w_067_1289, w_067_1290, w_067_1291, w_067_1293, w_067_1298, w_067_1299, w_067_1303, w_067_1306, w_067_1307, w_067_1308, w_067_1309, w_067_1313, w_067_1316, w_067_1317, w_067_1318, w_067_1322, w_067_1324, w_067_1325, w_067_1328, w_067_1330, w_067_1331, w_067_1333, w_067_1334, w_067_1336, w_067_1338, w_067_1340, w_067_1341, w_067_1343, w_067_1344, w_067_1345, w_067_1346, w_067_1348, w_067_1351, w_067_1354, w_067_1355, w_067_1357, w_067_1360, w_067_1362, w_067_1365, w_067_1366, w_067_1370, w_067_1374, w_067_1378, w_067_1383, w_067_1384, w_067_1385, w_067_1388, w_067_1390, w_067_1391, w_067_1392, w_067_1396, w_067_1397, w_067_1400, w_067_1402, w_067_1403, w_067_1404, w_067_1408, w_067_1409, w_067_1410, w_067_1411, w_067_1412, w_067_1414, w_067_1421, w_067_1424, w_067_1425, w_067_1427, w_067_1428, w_067_1429, w_067_1432, w_067_1434, w_067_1435, w_067_1437, w_067_1439, w_067_1440, w_067_1441, w_067_1442, w_067_1444, w_067_1445, w_067_1448, w_067_1451, w_067_1457, w_067_1459, w_067_1460, w_067_1464, w_067_1466, w_067_1468, w_067_1471, w_067_1472, w_067_1473, w_067_1475, w_067_1477, w_067_1480, w_067_1481, w_067_1485, w_067_1487, w_067_1491, w_067_1492, w_067_1494, w_067_1495, w_067_1497, w_067_1499, w_067_1501, w_067_1506, w_067_1508, w_067_1510, w_067_1511, w_067_1512, w_067_1514, w_067_1515, w_067_1517, w_067_1520, w_067_1521, w_067_1523, w_067_1524, w_067_1525, w_067_1526, w_067_1528, w_067_1529, w_067_1531, w_067_1533, w_067_1535, w_067_1537, w_067_1544, w_067_1545, w_067_1546, w_067_1547, w_067_1549, w_067_1550, w_067_1552, w_067_1561, w_067_1564, w_067_1568, w_067_1571, w_067_1577, w_067_1578, w_067_1579, w_067_1580, w_067_1585, w_067_1591, w_067_1592, w_067_1593, w_067_1594, w_067_1597, w_067_1598, w_067_1599, w_067_1601, w_067_1608, w_067_1609, w_067_1610, w_067_1613, w_067_1615, w_067_1621, w_067_1622, w_067_1624, w_067_1627, w_067_1630, w_067_1636, w_067_1639, w_067_1642, w_067_1648, w_067_1649, w_067_1652, w_067_1656, w_067_1657, w_067_1658, w_067_1659, w_067_1661, w_067_1662, w_067_1663, w_067_1666, w_067_1667, w_067_1668, w_067_1676, w_067_1678, w_067_1679, w_067_1684, w_067_1692, w_067_1694, w_067_1699, w_067_1701, w_067_1705, w_067_1707, w_067_1708, w_067_1710, w_067_1711, w_067_1716, w_067_1717, w_067_1719, w_067_1721, w_067_1722, w_067_1723, w_067_1724, w_067_1729, w_067_1732, w_067_1735, w_067_1736, w_067_1743, w_067_1747, w_067_1751, w_067_1752, w_067_1757, w_067_1758, w_067_1759, w_067_1761, w_067_1765, w_067_1767, w_067_1768, w_067_1772, w_067_1773, w_067_1778, w_067_1786, w_067_1789, w_067_1793, w_067_1795, w_067_1796, w_067_1798, w_067_1805, w_067_1806, w_067_1807, w_067_1808, w_067_1809, w_067_1810, w_067_1817, w_067_1822, w_067_1823, w_067_1824, w_067_1826, w_067_1827, w_067_1830, w_067_1832, w_067_1834, w_067_1835, w_067_1836, w_067_1840, w_067_1844, w_067_1847, w_067_1849, w_067_1855, w_067_1859, w_067_1863, w_067_1866, w_067_1871, w_067_1872, w_067_1873, w_067_1888, w_067_1891, w_067_1892, w_067_1894, w_067_1896, w_067_1905, w_067_1906, w_067_1908, w_067_1909, w_067_1912, w_067_1914, w_067_1917, w_067_1919, w_067_1920, w_067_1921, w_067_1922, w_067_1923, w_067_1924, w_067_1926, w_067_1936, w_067_1940, w_067_1945, w_067_1948, w_067_1951, w_067_1953, w_067_1956, w_067_1959, w_067_1960, w_067_1961, w_067_1962, w_067_1965, w_067_1972, w_067_1973, w_067_1975, w_067_1976, w_067_1978, w_067_1979, w_067_1982, w_067_1984, w_067_1989, w_067_1990, w_067_1991, w_067_1999, w_067_2002, w_067_2011, w_067_2015, w_067_2017, w_067_2018, w_067_2019, w_067_2020, w_067_2023, w_067_2029, w_067_2030, w_067_2031, w_067_2033, w_067_2034, w_067_2036, w_067_2038, w_067_2042, w_067_2048, w_067_2049, w_067_2057, w_067_2066, w_067_2069, w_067_2071, w_067_2072, w_067_2073, w_067_2075, w_067_2076, w_067_2081, w_067_2082, w_067_2083, w_067_2084, w_067_2087, w_067_2089, w_067_2090, w_067_2091, w_067_2092, w_067_2093, w_067_2094, w_067_2099, w_067_2104, w_067_2108, w_067_2109, w_067_2111, w_067_2115, w_067_2116, w_067_2118, w_067_2119, w_067_2121, w_067_2122, w_067_2126, w_067_2127, w_067_2134, w_067_2138, w_067_2139, w_067_2142, w_067_2144, w_067_2145, w_067_2154, w_067_2155, w_067_2159, w_067_2162, w_067_2163, w_067_2165, w_067_2168, w_067_2176, w_067_2178, w_067_2181, w_067_2182, w_067_2183, w_067_2188, w_067_2189, w_067_2191, w_067_2194, w_067_2198, w_067_2199, w_067_2211, w_067_2214, w_067_2215, w_067_2216, w_067_2221, w_067_2222, w_067_2223, w_067_2227, w_067_2229, w_067_2230, w_067_2232, w_067_2235, w_067_2237, w_067_2248, w_067_2250, w_067_2251, w_067_2253, w_067_2254, w_067_2255, w_067_2256, w_067_2259, w_067_2261, w_067_2263, w_067_2265, w_067_2269, w_067_2277, w_067_2278, w_067_2279, w_067_2284, w_067_2287, w_067_2291, w_067_2292, w_067_2294, w_067_2296, w_067_2297, w_067_2299, w_067_2300, w_067_2302, w_067_2306, w_067_2307, w_067_2308, w_067_2309, w_067_2311, w_067_2312, w_067_2313, w_067_2314, w_067_2316, w_067_2318, w_067_2322, w_067_2324, w_067_2325, w_067_2328, w_067_2331, w_067_2333, w_067_2336, w_067_2337, w_067_2340, w_067_2341, w_067_2342, w_067_2343, w_067_2352, w_067_2354, w_067_2356, w_067_2358, w_067_2359, w_067_2360, w_067_2361, w_067_2362, w_067_2363, w_067_2364, w_067_2365, w_067_2367, w_067_2368, w_067_2369, w_067_2373, w_067_2376, w_067_2378, w_067_2381, w_067_2387, w_067_2389, w_067_2390, w_067_2391, w_067_2393, w_067_2394, w_067_2396, w_067_2400, w_067_2404, w_067_2408, w_067_2410, w_067_2412, w_067_2417, w_067_2418, w_067_2419, w_067_2420, w_067_2423, w_067_2427, w_067_2429, w_067_2431, w_067_2437, w_067_2440, w_067_2441, w_067_2444, w_067_2446, w_067_2456, w_067_2472, w_067_2473, w_067_2475, w_067_2480, w_067_2483, w_067_2485, w_067_2488, w_067_2489, w_067_2494, w_067_2495, w_067_2496, w_067_2497, w_067_2498, w_067_2503, w_067_2513, w_067_2515, w_067_2516, w_067_2518, w_067_2519, w_067_2521, w_067_2522, w_067_2525, w_067_2528, w_067_2529, w_067_2531, w_067_2535, w_067_2536, w_067_2537, w_067_2539, w_067_2540, w_067_2542, w_067_2543, w_067_2545, w_067_2547, w_067_2554, w_067_2555, w_067_2556, w_067_2558, w_067_2559, w_067_2562, w_067_2563, w_067_2564, w_067_2566, w_067_2567, w_067_2571, w_067_2572, w_067_2574, w_067_2575, w_067_2578, w_067_2579, w_067_2582, w_067_2583, w_067_2592, w_067_2598, w_067_2601, w_067_2604, w_067_2605, w_067_2608, w_067_2610, w_067_2611, w_067_2613, w_067_2615, w_067_2620, w_067_2630, w_067_2631, w_067_2633, w_067_2634, w_067_2637, w_067_2638, w_067_2643, w_067_2644, w_067_2648, w_067_2650, w_067_2651, w_067_2652, w_067_2654, w_067_2655, w_067_2656, w_067_2663, w_067_2665, w_067_2666, w_067_2671, w_067_2672, w_067_2673, w_067_2677, w_067_2678, w_067_2679, w_067_2680, w_067_2681, w_067_2683, w_067_2686, w_067_2688, w_067_2689, w_067_2690, w_067_2696, w_067_2699, w_067_2706, w_067_2710, w_067_2712, w_067_2713, w_067_2714, w_067_2715, w_067_2722, w_067_2723, w_067_2730, w_067_2735, w_067_2739, w_067_2742, w_067_2744, w_067_2747, w_067_2750, w_067_2752, w_067_2754, w_067_2757, w_067_2759, w_067_2761, w_067_2764, w_067_2765, w_067_2768, w_067_2770, w_067_2771, w_067_2775, w_067_2782, w_067_2785, w_067_2791, w_067_2794, w_067_2798, w_067_2799, w_067_2800, w_067_2802, w_067_2804, w_067_2807, w_067_2810, w_067_2814, w_067_2819, w_067_2825, w_067_2836, w_067_2837, w_067_2838, w_067_2844, w_067_2845, w_067_2846, w_067_2849, w_067_2850, w_067_2852, w_067_2855, w_067_2856, w_067_2859, w_067_2861, w_067_2862, w_067_2867, w_067_2869, w_067_2871, w_067_2872, w_067_2874, w_067_2878, w_067_2884, w_067_2885, w_067_2887, w_067_2891, w_067_2896, w_067_2897, w_067_2900, w_067_2901, w_067_2902, w_067_2903, w_067_2905, w_067_2909, w_067_2910, w_067_2911, w_067_2916, w_067_2922, w_067_2923, w_067_2925, w_067_2933, w_067_2935, w_067_2937, w_067_2938, w_067_2939, w_067_2940, w_067_2941, w_067_2943, w_067_2948, w_067_2949, w_067_2953, w_067_2954, w_067_2955, w_067_2956, w_067_2958, w_067_2960, w_067_2963, w_067_2965, w_067_2966, w_067_2971, w_067_2974, w_067_2977, w_067_2979, w_067_2980, w_067_2987, w_067_2991, w_067_2993, w_067_2994, w_067_2996, w_067_2999, w_067_3001, w_067_3006, w_067_3007, w_067_3008, w_067_3013, w_067_3014, w_067_3015, w_067_3016, w_067_3018, w_067_3019, w_067_3021, w_067_3027, w_067_3028, w_067_3029, w_067_3030, w_067_3031, w_067_3036, w_067_3037, w_067_3038, w_067_3041, w_067_3043, w_067_3046, w_067_3048, w_067_3054, w_067_3055, w_067_3057, w_067_3062, w_067_3065, w_067_3066, w_067_3072, w_067_3073, w_067_3074, w_067_3075, w_067_3084, w_067_3086, w_067_3092, w_067_3093, w_067_3094, w_067_3100, w_067_3102, w_067_3104, w_067_3105, w_067_3107, w_067_3110, w_067_3112, w_067_3114, w_067_3123, w_067_3126, w_067_3128, w_067_3129, w_067_3132, w_067_3134, w_067_3135, w_067_3137, w_067_3140, w_067_3142, w_067_3144, w_067_3159, w_067_3160, w_067_3162, w_067_3166, w_067_3170, w_067_3172, w_067_3173, w_067_3178, w_067_3179, w_067_3180, w_067_3185, w_067_3187, w_067_3189, w_067_3190, w_067_3191, w_067_3193, w_067_3194, w_067_3198, w_067_3203, w_067_3204, w_067_3206, w_067_3207, w_067_3210, w_067_3214, w_067_3215, w_067_3226, w_067_3227, w_067_3232, w_067_3233, w_067_3241, w_067_3242, w_067_3243, w_067_3253, w_067_3255, w_067_3256, w_067_3259, w_067_3260, w_067_3265, w_067_3266, w_067_3269, w_067_3273, w_067_3279, w_067_3280, w_067_3282, w_067_3283, w_067_3285, w_067_3288, w_067_3292, w_067_3293, w_067_3295, w_067_3296, w_067_3298, w_067_3299, w_067_3300, w_067_3302, w_067_3303, w_067_3304, w_067_3308, w_067_3311, w_067_3313, w_067_3316, w_067_3321, w_067_3323, w_067_3329, w_067_3330, w_067_3331, w_067_3332, w_067_3333, w_067_3334, w_067_3337, w_067_3340, w_067_3346, w_067_3349, w_067_3350, w_067_3351, w_067_3353, w_067_3355, w_067_3356, w_067_3357, w_067_3363, w_067_3366, w_067_3368, w_067_3369, w_067_3373, w_067_3378, w_067_3380, w_067_3381, w_067_3383, w_067_3386, w_067_3388, w_067_3391, w_067_3392, w_067_3394, w_067_3398, w_067_3399, w_067_3400, w_067_3401, w_067_3402, w_067_3404, w_067_3405, w_067_3410, w_067_3412, w_067_3413, w_067_3418, w_067_3423, w_067_3424, w_067_3425, w_067_3426, w_067_3427, w_067_3429, w_067_3433, w_067_3435, w_067_3440, w_067_3442, w_067_3443, w_067_3445, w_067_3446, w_067_3447, w_067_3448, w_067_3450, w_067_3454, w_067_3455, w_067_3458, w_067_3461, w_067_3465, w_067_3466, w_067_3473, w_067_3474, w_067_3476, w_067_3478, w_067_3479, w_067_3480, w_067_3481, w_067_3484, w_067_3487, w_067_3491, w_067_3495, w_067_3500, w_067_3501, w_067_3502, w_067_3504, w_067_3505, w_067_3509, w_067_3513, w_067_3516, w_067_3521, w_067_3526, w_067_3527, w_067_3528, w_067_3529, w_067_3530, w_067_3531, w_067_3532, w_067_3533, w_067_3534, w_067_3536, w_067_3544, w_067_3546, w_067_3547, w_067_3548, w_067_3549, w_067_3551, w_067_3556, w_067_3558, w_067_3559, w_067_3562, w_067_3568, w_067_3570, w_067_3573, w_067_3576, w_067_3578, w_067_3580, w_067_3581, w_067_3582, w_067_3583, w_067_3584, w_067_3585, w_067_3586, w_067_3587, w_067_3590, w_067_3592, w_067_3593, w_067_3594, w_067_3595, w_067_3599, w_067_3601, w_067_3602, w_067_3604, w_067_3605, w_067_3612, w_067_3616, w_067_3617, w_067_3619, w_067_3626, w_067_3627, w_067_3628, w_067_3629, w_067_3630, w_067_3632, w_067_3633, w_067_3635, w_067_3639, w_067_3640, w_067_3641, w_067_3642, w_067_3644, w_067_3650, w_067_3652, w_067_3654, w_067_3656, w_067_3657, w_067_3665, w_067_3666, w_067_3668, w_067_3674, w_067_3675, w_067_3677, w_067_3682, w_067_3683, w_067_3686, w_067_3690, w_067_3691, w_067_3694, w_067_3695, w_067_3696, w_067_3700, w_067_3703, w_067_3705, w_067_3710, w_067_3712, w_067_3713, w_067_3716, w_067_3721, w_067_3722, w_067_3724, w_067_3725, w_067_3726, w_067_3728, w_067_3735, w_067_3741, w_067_3743, w_067_3744, w_067_3745, w_067_3747, w_067_3749, w_067_3750, w_067_3756, w_067_3759, w_067_3760, w_067_3761, w_067_3763, w_067_3766, w_067_3768, w_067_3769, w_067_3771, w_067_3775, w_067_3776, w_067_3777, w_067_3779, w_067_3780, w_067_3783, w_067_3784, w_067_3785, w_067_3786, w_067_3787, w_067_3789, w_067_3793, w_067_3795, w_067_3797, w_067_3799, w_067_3803, w_067_3805, w_067_3806, w_067_3807, w_067_3811, w_067_3814, w_067_3816, w_067_3817, w_067_3826, w_067_3830, w_067_3832, w_067_3835, w_067_3839, w_067_3844, w_067_3845, w_067_3846, w_067_3848, w_067_3851, w_067_3852, w_067_3854, w_067_3855, w_067_3861, w_067_3863, w_067_3868, w_067_3869, w_067_3870, w_067_3873, w_067_3874, w_067_3875, w_067_3880, w_067_3881, w_067_3895, w_067_3896, w_067_3897, w_067_3898, w_067_3902, w_067_3905, w_067_3906, w_067_3908, w_067_3913, w_067_3914, w_067_3915, w_067_3917, w_067_3918, w_067_3922, w_067_3926, w_067_3927, w_067_3932, w_067_3933, w_067_3934, w_067_3935, w_067_3940, w_067_3942, w_067_3943, w_067_3947, w_067_3948, w_067_3949, w_067_3950, w_067_3953, w_067_3961, w_067_3966, w_067_3968, w_067_3969, w_067_3971, w_067_3975, w_067_3977, w_067_3980, w_067_3981, w_067_3983, w_067_3984, w_067_3985, w_067_3996, w_067_3997, w_067_4003, w_067_4004, w_067_4005, w_067_4006, w_067_4007, w_067_4009, w_067_4010, w_067_4014, w_067_4016, w_067_4018, w_067_4026, w_067_4028, w_067_4029, w_067_4034, w_067_4037, w_067_4039, w_067_4040, w_067_4043, w_067_4044, w_067_4045, w_067_4046, w_067_4049, w_067_4050, w_067_4051, w_067_4052, w_067_4055, w_067_4056, w_067_4061, w_067_4063, w_067_4064, w_067_4069, w_067_4070, w_067_4079, w_067_4080, w_067_4081, w_067_4083, w_067_4086, w_067_4089, w_067_4090, w_067_4092, w_067_4093, w_067_4095, w_067_4096, w_067_4098, w_067_4100, w_067_4103, w_067_4104, w_067_4105, w_067_4106, w_067_4107, w_067_4110, w_067_4113, w_067_4116, w_067_4117, w_067_4128, w_067_4132, w_067_4134, w_067_4142, w_067_4144, w_067_4150, w_067_4152, w_067_4159, w_067_4163, w_067_4165, w_067_4166, w_067_4170, w_067_4172, w_067_4173, w_067_4175, w_067_4177, w_067_4178, w_067_4185, w_067_4186, w_067_4189, w_067_4193, w_067_4196, w_067_4198, w_067_4203, w_067_4204, w_067_4206, w_067_4207, w_067_4209, w_067_4211, w_067_4214, w_067_4218, w_067_4219, w_067_4220, w_067_4223, w_067_4224, w_067_4241, w_067_4242, w_067_4245, w_067_4251, w_067_4256, w_067_4257, w_067_4259, w_067_4260, w_067_4264, w_067_4272, w_067_4273, w_067_4274, w_067_4281, w_067_4282, w_067_4287, w_067_4288, w_067_4295, w_067_4299, w_067_4300, w_067_4307, w_067_4308, w_067_4309, w_067_4310, w_067_4313, w_067_4319, w_067_4320, w_067_4322, w_067_4328, w_067_4331, w_067_4339, w_067_4340, w_067_4342, w_067_4343, w_067_4344, w_067_4346, w_067_4347, w_067_4350, w_067_4351, w_067_4352, w_067_4356, w_067_4357, w_067_4362, w_067_4364, w_067_4365, w_067_4369, w_067_4372, w_067_4375, w_067_4377, w_067_4382, w_067_4385, w_067_4389, w_067_4394, w_067_4398, w_067_4399, w_067_4405, w_067_4408, w_067_4409, w_067_4410, w_067_4413, w_067_4414, w_067_4415, w_067_4417, w_067_4418, w_067_4422, w_067_4423, w_067_4424, w_067_4426, w_067_4429, w_067_4430, w_067_4433, w_067_4436, w_067_4438, w_067_4439, w_067_4440, w_067_4442, w_067_4444, w_067_4447, w_067_4448, w_067_4449, w_067_4453, w_067_4455, w_067_4460, w_067_4463, w_067_4464, w_067_4467, w_067_4470, w_067_4473, w_067_4475, w_067_4477, w_067_4482, w_067_4487, w_067_4488, w_067_4489, w_067_4491, w_067_4498, w_067_4499, w_067_4505, w_067_4509, w_067_4511, w_067_4512, w_067_4516, w_067_4517, w_067_4518, w_067_4519, w_067_4520, w_067_4524, w_067_4528, w_067_4531, w_067_4533, w_067_4538, w_067_4539, w_067_4540, w_067_4541, w_067_4542, w_067_4544, w_067_4552, w_067_4556, w_067_4557, w_067_4559, w_067_4560, w_067_4562, w_067_4570, w_067_4573, w_067_4574, w_067_4575, w_067_4576, w_067_4577, w_067_4578, w_067_4583, w_067_4584, w_067_4590, w_067_4593, w_067_4596, w_067_4597, w_067_4598, w_067_4605, w_067_4609, w_067_4613, w_067_4614, w_067_4616, w_067_4618, w_067_4619, w_067_4621, w_067_4625, w_067_4626, w_067_4627, w_067_4629, w_067_4631, w_067_4632, w_067_4633, w_067_4634, w_067_4636, w_067_4637, w_067_4640, w_067_4645, w_067_4647, w_067_4649, w_067_4650, w_067_4651, w_067_4653, w_067_4655, w_067_4656, w_067_4657, w_067_4658, w_067_4659, w_067_4661, w_067_4662, w_067_4668, w_067_4670, w_067_4672, w_067_4674, w_067_4677, w_067_4684, w_067_4686, w_067_4687, w_067_4692, w_067_4696, w_067_4700, w_067_4704, w_067_4707, w_067_4710, w_067_4716, w_067_4718, w_067_4719, w_067_4720, w_067_4721, w_067_4725, w_067_4733, w_067_4736, w_067_4741, w_067_4742, w_067_4744, w_067_4746, w_067_4748, w_067_4750, w_067_4755, w_067_4756, w_067_4757, w_067_4758, w_067_4761, w_067_4762, w_067_4772, w_067_4773, w_067_4775, w_067_4778, w_067_4779, w_067_4783, w_067_4785, w_067_4787, w_067_4788, w_067_4792, w_067_4794, w_067_4795, w_067_4797, w_067_4799, w_067_4802, w_067_4804, w_067_4807, w_067_4809, w_067_4810, w_067_4812, w_067_4813, w_067_4814, w_067_4816, w_067_4817, w_067_4823, w_067_4825, w_067_4830, w_067_4833, w_067_4834, w_067_4836, w_067_4838, w_067_4839, w_067_4841, w_067_4842, w_067_4846, w_067_4849, w_067_4850, w_067_4853, w_067_4854, w_067_4856, w_067_4858, w_067_4861, w_067_4862, w_067_4866, w_067_4871, w_067_4875, w_067_4876, w_067_4879, w_067_4880, w_067_4881, w_067_4884, w_067_4885;
  wire w_068_001, w_068_004, w_068_005, w_068_006, w_068_009, w_068_011, w_068_012, w_068_013, w_068_016, w_068_017, w_068_020, w_068_021, w_068_022, w_068_023, w_068_027, w_068_030, w_068_031, w_068_032, w_068_033, w_068_034, w_068_035, w_068_036, w_068_037, w_068_038, w_068_040, w_068_041, w_068_042, w_068_043, w_068_044, w_068_045, w_068_047, w_068_048, w_068_049, w_068_051, w_068_053, w_068_054, w_068_056, w_068_057, w_068_059, w_068_060, w_068_061, w_068_062, w_068_064, w_068_066, w_068_067, w_068_068, w_068_071, w_068_073, w_068_075, w_068_076, w_068_080, w_068_082, w_068_084, w_068_085, w_068_087, w_068_091, w_068_094, w_068_095, w_068_096, w_068_097, w_068_098, w_068_101, w_068_102, w_068_106, w_068_107, w_068_108, w_068_109, w_068_110, w_068_114, w_068_116, w_068_117, w_068_118, w_068_119, w_068_120, w_068_121, w_068_122, w_068_123, w_068_124, w_068_125, w_068_128, w_068_129, w_068_130, w_068_132, w_068_133, w_068_134, w_068_135, w_068_136, w_068_138, w_068_142, w_068_143, w_068_145, w_068_146, w_068_148, w_068_149, w_068_153, w_068_154, w_068_156, w_068_158, w_068_163, w_068_164, w_068_165, w_068_166, w_068_167, w_068_168, w_068_169, w_068_171, w_068_172, w_068_173, w_068_175, w_068_176, w_068_178, w_068_179, w_068_183, w_068_184, w_068_185, w_068_186, w_068_187, w_068_188, w_068_189, w_068_190, w_068_192, w_068_193, w_068_195, w_068_196, w_068_198, w_068_199, w_068_201, w_068_202, w_068_204, w_068_205, w_068_206, w_068_208, w_068_212, w_068_213, w_068_214, w_068_216, w_068_218, w_068_219, w_068_220, w_068_223, w_068_230, w_068_231, w_068_234, w_068_237, w_068_238, w_068_242, w_068_243, w_068_244, w_068_246, w_068_247, w_068_248, w_068_251, w_068_253, w_068_254, w_068_257, w_068_260, w_068_262, w_068_263, w_068_264, w_068_266, w_068_267, w_068_268, w_068_269, w_068_270, w_068_272, w_068_273, w_068_275, w_068_277, w_068_278, w_068_279, w_068_280, w_068_282, w_068_283, w_068_284, w_068_285, w_068_287, w_068_288, w_068_289, w_068_290, w_068_291, w_068_292, w_068_294, w_068_296, w_068_298, w_068_299, w_068_300, w_068_301, w_068_302, w_068_303, w_068_304, w_068_305, w_068_307, w_068_308, w_068_309, w_068_310, w_068_313, w_068_314, w_068_315, w_068_316, w_068_317, w_068_318, w_068_319, w_068_321, w_068_323, w_068_324, w_068_325, w_068_327, w_068_328, w_068_330, w_068_332, w_068_333, w_068_334, w_068_339, w_068_340, w_068_341, w_068_347, w_068_348, w_068_349, w_068_350, w_068_354, w_068_356, w_068_357, w_068_358, w_068_359, w_068_362, w_068_364, w_068_365, w_068_367, w_068_368, w_068_370, w_068_372, w_068_373, w_068_375, w_068_376, w_068_378, w_068_379, w_068_380, w_068_381, w_068_382, w_068_383, w_068_385, w_068_386, w_068_388, w_068_389, w_068_390, w_068_391, w_068_393, w_068_396, w_068_398, w_068_400, w_068_402, w_068_403, w_068_404, w_068_409, w_068_410, w_068_411, w_068_412, w_068_413, w_068_421, w_068_422, w_068_423, w_068_425, w_068_428, w_068_430, w_068_431, w_068_433, w_068_436, w_068_437, w_068_438, w_068_439, w_068_444, w_068_448, w_068_450, w_068_454, w_068_455, w_068_459, w_068_460, w_068_464, w_068_467, w_068_470, w_068_473, w_068_474, w_068_475, w_068_476, w_068_477, w_068_482, w_068_487, w_068_489, w_068_491, w_068_494, w_068_495, w_068_496, w_068_497, w_068_498, w_068_499, w_068_501, w_068_505, w_068_507, w_068_510, w_068_514, w_068_516, w_068_522, w_068_524, w_068_529, w_068_532, w_068_538, w_068_539, w_068_542, w_068_543, w_068_544, w_068_547, w_068_550, w_068_554, w_068_556, w_068_557, w_068_558, w_068_561, w_068_562, w_068_565, w_068_568, w_068_569, w_068_570, w_068_571, w_068_575, w_068_579, w_068_583, w_068_584, w_068_586, w_068_590, w_068_594, w_068_595, w_068_596, w_068_597, w_068_599, w_068_601, w_068_603, w_068_609, w_068_610, w_068_611, w_068_612, w_068_617, w_068_622, w_068_624, w_068_625, w_068_627, w_068_628, w_068_629, w_068_630, w_068_631, w_068_634, w_068_636, w_068_639, w_068_640, w_068_642, w_068_647, w_068_650, w_068_653, w_068_654, w_068_655, w_068_657, w_068_659, w_068_660, w_068_663, w_068_664, w_068_665, w_068_668, w_068_670, w_068_671, w_068_678, w_068_682, w_068_684, w_068_685, w_068_686, w_068_689, w_068_693, w_068_702, w_068_705, w_068_708, w_068_713, w_068_715, w_068_716, w_068_719, w_068_720, w_068_727, w_068_728, w_068_732, w_068_734, w_068_738, w_068_739, w_068_740, w_068_741, w_068_742, w_068_743, w_068_749, w_068_750, w_068_752, w_068_757, w_068_759, w_068_760, w_068_762, w_068_770, w_068_776, w_068_777, w_068_779, w_068_781, w_068_784, w_068_785, w_068_789, w_068_793, w_068_795, w_068_804, w_068_805, w_068_807, w_068_808, w_068_809, w_068_812, w_068_816, w_068_818, w_068_820, w_068_822, w_068_827, w_068_832, w_068_838, w_068_839, w_068_841, w_068_844, w_068_857, w_068_859, w_068_861, w_068_864, w_068_865, w_068_867, w_068_868, w_068_870, w_068_872, w_068_876, w_068_880, w_068_882, w_068_887, w_068_890, w_068_891, w_068_896, w_068_898, w_068_899, w_068_900, w_068_902, w_068_905, w_068_907, w_068_910, w_068_913, w_068_914, w_068_918, w_068_921, w_068_923, w_068_924, w_068_926, w_068_928, w_068_931, w_068_933, w_068_934, w_068_935, w_068_936, w_068_939, w_068_940, w_068_941, w_068_943, w_068_947, w_068_948, w_068_951, w_068_957, w_068_958, w_068_964, w_068_967, w_068_968, w_068_971, w_068_972, w_068_973, w_068_976, w_068_977, w_068_986, w_068_990, w_068_991, w_068_996, w_068_999, w_068_1000, w_068_1002, w_068_1010, w_068_1011, w_068_1014, w_068_1015, w_068_1025, w_068_1028, w_068_1031, w_068_1033, w_068_1034, w_068_1041, w_068_1042, w_068_1043, w_068_1059, w_068_1060, w_068_1061, w_068_1062, w_068_1064, w_068_1065, w_068_1066, w_068_1068, w_068_1069, w_068_1072, w_068_1076, w_068_1077, w_068_1078, w_068_1083, w_068_1085, w_068_1089, w_068_1092, w_068_1094, w_068_1095, w_068_1104, w_068_1105, w_068_1106, w_068_1111, w_068_1114, w_068_1120, w_068_1128, w_068_1131, w_068_1133, w_068_1135, w_068_1136, w_068_1138, w_068_1140, w_068_1146, w_068_1148, w_068_1149, w_068_1151, w_068_1153, w_068_1154, w_068_1156, w_068_1157, w_068_1159, w_068_1173, w_068_1174, w_068_1178, w_068_1181, w_068_1182, w_068_1184, w_068_1186, w_068_1189, w_068_1191, w_068_1196, w_068_1198, w_068_1199, w_068_1201, w_068_1202, w_068_1203, w_068_1204, w_068_1210, w_068_1214, w_068_1218, w_068_1219, w_068_1226, w_068_1227, w_068_1228, w_068_1230, w_068_1234, w_068_1235, w_068_1239, w_068_1243, w_068_1245, w_068_1246, w_068_1247, w_068_1248, w_068_1250, w_068_1258, w_068_1263, w_068_1265, w_068_1266, w_068_1268, w_068_1271, w_068_1273, w_068_1274, w_068_1275, w_068_1276, w_068_1277, w_068_1281, w_068_1282, w_068_1283, w_068_1287, w_068_1289, w_068_1292, w_068_1298, w_068_1300, w_068_1301, w_068_1305, w_068_1309, w_068_1310, w_068_1311, w_068_1312, w_068_1315, w_068_1317, w_068_1318, w_068_1321, w_068_1323, w_068_1328, w_068_1329, w_068_1330, w_068_1333, w_068_1334, w_068_1337, w_068_1339, w_068_1340, w_068_1341, w_068_1343, w_068_1350, w_068_1351, w_068_1357, w_068_1358, w_068_1361, w_068_1365, w_068_1372, w_068_1377, w_068_1379, w_068_1380, w_068_1381, w_068_1394, w_068_1397, w_068_1398, w_068_1399, w_068_1400, w_068_1403, w_068_1411, w_068_1412, w_068_1413, w_068_1414, w_068_1418, w_068_1420, w_068_1424, w_068_1426, w_068_1427, w_068_1429, w_068_1434, w_068_1435, w_068_1439, w_068_1444, w_068_1445, w_068_1448, w_068_1450, w_068_1454, w_068_1455, w_068_1456, w_068_1459, w_068_1461, w_068_1467, w_068_1468, w_068_1469, w_068_1470, w_068_1473, w_068_1477, w_068_1479, w_068_1481, w_068_1483, w_068_1488, w_068_1489, w_068_1496, w_068_1504, w_068_1505, w_068_1507, w_068_1509, w_068_1510, w_068_1511, w_068_1512, w_068_1515, w_068_1517, w_068_1522, w_068_1523, w_068_1526, w_068_1529, w_068_1530, w_068_1534, w_068_1536, w_068_1541, w_068_1542, w_068_1543, w_068_1549, w_068_1554, w_068_1556, w_068_1560, w_068_1562, w_068_1566, w_068_1567, w_068_1568, w_068_1569, w_068_1570, w_068_1571, w_068_1573, w_068_1574, w_068_1576, w_068_1579, w_068_1580, w_068_1583, w_068_1584, w_068_1587, w_068_1588, w_068_1592, w_068_1601, w_068_1602, w_068_1603, w_068_1608, w_068_1613, w_068_1615, w_068_1617, w_068_1621, w_068_1622, w_068_1624, w_068_1625, w_068_1632, w_068_1634, w_068_1636, w_068_1637, w_068_1638, w_068_1642, w_068_1645, w_068_1648, w_068_1651, w_068_1652, w_068_1654, w_068_1656, w_068_1657, w_068_1659, w_068_1660, w_068_1661, w_068_1663, w_068_1668, w_068_1669, w_068_1672, w_068_1673, w_068_1675, w_068_1679, w_068_1680, w_068_1682, w_068_1683, w_068_1684, w_068_1693, w_068_1697, w_068_1700, w_068_1702, w_068_1704, w_068_1707, w_068_1709, w_068_1711, w_068_1716, w_068_1719, w_068_1725, w_068_1727, w_068_1728, w_068_1732, w_068_1735, w_068_1736, w_068_1739, w_068_1740, w_068_1744, w_068_1750, w_068_1754, w_068_1757, w_068_1760, w_068_1762, w_068_1769, w_068_1771, w_068_1773, w_068_1776, w_068_1777, w_068_1778, w_068_1780, w_068_1781, w_068_1782, w_068_1784, w_068_1785, w_068_1787, w_068_1791, w_068_1793, w_068_1795, w_068_1798, w_068_1799, w_068_1800, w_068_1803, w_068_1804, w_068_1806, w_068_1808, w_068_1809, w_068_1817, w_068_1818, w_068_1820, w_068_1822, w_068_1829, w_068_1831, w_068_1832, w_068_1834, w_068_1836, w_068_1839, w_068_1840, w_068_1841, w_068_1843, w_068_1846, w_068_1848, w_068_1849, w_068_1851, w_068_1853, w_068_1854, w_068_1857, w_068_1858, w_068_1859, w_068_1861, w_068_1865, w_068_1870, w_068_1872, w_068_1875, w_068_1879, w_068_1881, w_068_1884, w_068_1887, w_068_1888, w_068_1891, w_068_1897, w_068_1899, w_068_1901, w_068_1905, w_068_1909, w_068_1911, w_068_1917, w_068_1918, w_068_1921, w_068_1922, w_068_1923, w_068_1924, w_068_1925, w_068_1927, w_068_1929, w_068_1932, w_068_1934, w_068_1937, w_068_1938, w_068_1942, w_068_1946, w_068_1947, w_068_1948, w_068_1952, w_068_1957, w_068_1958, w_068_1964, w_068_1966, w_068_1972, w_068_1974, w_068_1975, w_068_1976, w_068_1977, w_068_1979, w_068_1980, w_068_1982, w_068_1988, w_068_1989, w_068_1990, w_068_1991, w_068_1993, w_068_1994, w_068_1998, w_068_2007, w_068_2008, w_068_2009, w_068_2013, w_068_2016, w_068_2017, w_068_2020, w_068_2025, w_068_2026, w_068_2029, w_068_2037, w_068_2040, w_068_2041, w_068_2042, w_068_2048, w_068_2049, w_068_2050, w_068_2051, w_068_2052, w_068_2054, w_068_2056, w_068_2057, w_068_2064, w_068_2067, w_068_2072, w_068_2073, w_068_2074, w_068_2075, w_068_2078, w_068_2083, w_068_2084, w_068_2085, w_068_2087, w_068_2089, w_068_2090, w_068_2096, w_068_2098, w_068_2099, w_068_2102, w_068_2103, w_068_2105, w_068_2111, w_068_2115, w_068_2116, w_068_2120, w_068_2121, w_068_2127, w_068_2128, w_068_2129, w_068_2130, w_068_2131, w_068_2134, w_068_2136, w_068_2137, w_068_2138, w_068_2144, w_068_2146, w_068_2149, w_068_2151, w_068_2152, w_068_2159, w_068_2162, w_068_2163, w_068_2166, w_068_2168, w_068_2172, w_068_2173, w_068_2176, w_068_2177, w_068_2178, w_068_2180, w_068_2181, w_068_2185, w_068_2188, w_068_2189, w_068_2190, w_068_2196, w_068_2197, w_068_2199, w_068_2203, w_068_2205, w_068_2209, w_068_2214, w_068_2219, w_068_2227, w_068_2229, w_068_2233, w_068_2234, w_068_2235, w_068_2238, w_068_2239, w_068_2240, w_068_2242, w_068_2244, w_068_2245, w_068_2248, w_068_2249, w_068_2253, w_068_2254, w_068_2255, w_068_2257, w_068_2259, w_068_2260, w_068_2261, w_068_2266, w_068_2269, w_068_2270, w_068_2271, w_068_2272, w_068_2275, w_068_2277, w_068_2279, w_068_2281, w_068_2283, w_068_2285, w_068_2286, w_068_2288, w_068_2290, w_068_2292, w_068_2293, w_068_2295, w_068_2297, w_068_2299, w_068_2302, w_068_2304, w_068_2308, w_068_2309, w_068_2313, w_068_2316, w_068_2317, w_068_2318, w_068_2320, w_068_2325, w_068_2329, w_068_2330, w_068_2335, w_068_2336, w_068_2341, w_068_2343, w_068_2344, w_068_2345, w_068_2347, w_068_2349, w_068_2355, w_068_2357, w_068_2358, w_068_2360, w_068_2361, w_068_2364, w_068_2367, w_068_2370, w_068_2373, w_068_2374, w_068_2375, w_068_2376, w_068_2379, w_068_2380, w_068_2384, w_068_2385, w_068_2390, w_068_2391, w_068_2392, w_068_2393, w_068_2394, w_068_2397, w_068_2401, w_068_2402, w_068_2403, w_068_2405, w_068_2408, w_068_2411, w_068_2412, w_068_2415, w_068_2418, w_068_2421, w_068_2422, w_068_2424, w_068_2425, w_068_2426, w_068_2428, w_068_2430, w_068_2434, w_068_2435, w_068_2437, w_068_2438, w_068_2440, w_068_2441, w_068_2444, w_068_2445, w_068_2449, w_068_2451, w_068_2457, w_068_2458, w_068_2460, w_068_2461, w_068_2462, w_068_2463, w_068_2470, w_068_2475, w_068_2480, w_068_2487, w_068_2490, w_068_2491, w_068_2493, w_068_2494, w_068_2495, w_068_2497, w_068_2500, w_068_2502, w_068_2511, w_068_2513, w_068_2514, w_068_2515, w_068_2519, w_068_2520, w_068_2522, w_068_2528, w_068_2531, w_068_2533, w_068_2535, w_068_2536, w_068_2538, w_068_2541, w_068_2542, w_068_2544, w_068_2547, w_068_2549, w_068_2558, w_068_2560, w_068_2561, w_068_2563, w_068_2564, w_068_2567, w_068_2568, w_068_2572, w_068_2573, w_068_2574, w_068_2576, w_068_2577, w_068_2578, w_068_2590, w_068_2592, w_068_2593, w_068_2596, w_068_2597, w_068_2603, w_068_2605, w_068_2607, w_068_2610, w_068_2612, w_068_2613, w_068_2617, w_068_2618, w_068_2623, w_068_2624, w_068_2629, w_068_2632, w_068_2638, w_068_2639, w_068_2642, w_068_2643, w_068_2646, w_068_2649, w_068_2650, w_068_2652, w_068_2656, w_068_2658, w_068_2659, w_068_2661, w_068_2662, w_068_2663, w_068_2664, w_068_2665, w_068_2666, w_068_2669, w_068_2673, w_068_2681, w_068_2684, w_068_2688, w_068_2689, w_068_2690, w_068_2698, w_068_2701, w_068_2702, w_068_2704, w_068_2708, w_068_2711, w_068_2716, w_068_2720, w_068_2721, w_068_2730, w_068_2731, w_068_2734, w_068_2737, w_068_2739, w_068_2744, w_068_2747, w_068_2751, w_068_2752, w_068_2753, w_068_2755, w_068_2758, w_068_2759, w_068_2760, w_068_2763, w_068_2767, w_068_2769, w_068_2770, w_068_2771, w_068_2772, w_068_2777, w_068_2783, w_068_2786, w_068_2787, w_068_2791, w_068_2794, w_068_2800, w_068_2801, w_068_2804, w_068_2805, w_068_2807, w_068_2811, w_068_2813, w_068_2817, w_068_2820, w_068_2824, w_068_2825, w_068_2827, w_068_2828, w_068_2830, w_068_2831, w_068_2834, w_068_2840, w_068_2842, w_068_2847, w_068_2850, w_068_2852, w_068_2857, w_068_2858, w_068_2860, w_068_2861, w_068_2865, w_068_2868, w_068_2870, w_068_2871, w_068_2874, w_068_2875, w_068_2876, w_068_2877, w_068_2881, w_068_2885, w_068_2886, w_068_2888, w_068_2889, w_068_2892, w_068_2893, w_068_2897, w_068_2898, w_068_2901, w_068_2902, w_068_2903, w_068_2906, w_068_2907, w_068_2908, w_068_2909, w_068_2910, w_068_2911, w_068_2912, w_068_2913, w_068_2915, w_068_2917, w_068_2920, w_068_2921, w_068_2925, w_068_2926, w_068_2929, w_068_2930, w_068_2931, w_068_2932, w_068_2934, w_068_2937, w_068_2941, w_068_2948, w_068_2953, w_068_2955, w_068_2957, w_068_2958, w_068_2959, w_068_2961, w_068_2962, w_068_2966, w_068_2969, w_068_2975, w_068_2976, w_068_2979, w_068_2982, w_068_2988, w_068_2991, w_068_2992, w_068_3000, w_068_3002, w_068_3004, w_068_3006, w_068_3007, w_068_3008, w_068_3009, w_068_3010, w_068_3011, w_068_3016, w_068_3019, w_068_3023, w_068_3027, w_068_3028, w_068_3029, w_068_3030, w_068_3031, w_068_3032, w_068_3034, w_068_3036, w_068_3037, w_068_3039, w_068_3045, w_068_3048, w_068_3051, w_068_3055, w_068_3056, w_068_3058, w_068_3059, w_068_3060, w_068_3061, w_068_3063, w_068_3065, w_068_3066, w_068_3067, w_068_3068, w_068_3069, w_068_3071, w_068_3072, w_068_3075, w_068_3081, w_068_3082, w_068_3083, w_068_3088, w_068_3090, w_068_3091, w_068_3097, w_068_3098, w_068_3100, w_068_3101, w_068_3102, w_068_3103, w_068_3104, w_068_3106, w_068_3109, w_068_3110, w_068_3112, w_068_3117, w_068_3120, w_068_3121, w_068_3123, w_068_3124, w_068_3125, w_068_3126, w_068_3127, w_068_3130, w_068_3133, w_068_3135, w_068_3136, w_068_3138, w_068_3139, w_068_3140, w_068_3147, w_068_3151, w_068_3152, w_068_3154, w_068_3156, w_068_3159, w_068_3160, w_068_3164, w_068_3166, w_068_3169, w_068_3173, w_068_3175, w_068_3177, w_068_3180, w_068_3181, w_068_3182, w_068_3184, w_068_3187, w_068_3190, w_068_3191, w_068_3192, w_068_3195, w_068_3196, w_068_3200, w_068_3201, w_068_3203, w_068_3208, w_068_3213, w_068_3215, w_068_3216, w_068_3218, w_068_3219, w_068_3220, w_068_3228, w_068_3230, w_068_3231, w_068_3232, w_068_3235, w_068_3236, w_068_3237, w_068_3244, w_068_3250, w_068_3251, w_068_3255, w_068_3261, w_068_3265, w_068_3266, w_068_3280, w_068_3285, w_068_3288, w_068_3289, w_068_3296, w_068_3299, w_068_3302, w_068_3303, w_068_3308, w_068_3309, w_068_3316, w_068_3321, w_068_3325, w_068_3329, w_068_3333, w_068_3335, w_068_3337, w_068_3340, w_068_3342, w_068_3344, w_068_3345, w_068_3346, w_068_3347, w_068_3352, w_068_3354, w_068_3355, w_068_3361, w_068_3362, w_068_3363, w_068_3368, w_068_3370, w_068_3374, w_068_3377, w_068_3378, w_068_3379, w_068_3387, w_068_3389, w_068_3390, w_068_3392, w_068_3394, w_068_3397, w_068_3398, w_068_3399, w_068_3400, w_068_3402, w_068_3409, w_068_3412, w_068_3416, w_068_3417, w_068_3422, w_068_3425, w_068_3426, w_068_3427, w_068_3430, w_068_3432, w_068_3437, w_068_3442, w_068_3444, w_068_3446, w_068_3447, w_068_3449, w_068_3451, w_068_3458, w_068_3461, w_068_3470, w_068_3471, w_068_3478, w_068_3479, w_068_3482, w_068_3483, w_068_3484, w_068_3490, w_068_3491, w_068_3492, w_068_3495, w_068_3498, w_068_3500, w_068_3504, w_068_3505, w_068_3507, w_068_3511, w_068_3514, w_068_3515, w_068_3516, w_068_3531, w_068_3533, w_068_3535, w_068_3536, w_068_3538, w_068_3540, w_068_3541, w_068_3542, w_068_3546, w_068_3547, w_068_3551, w_068_3556, w_068_3559, w_068_3564, w_068_3565, w_068_3566, w_068_3572, w_068_3573, w_068_3578, w_068_3584, w_068_3586, w_068_3591, w_068_3592, w_068_3596, w_068_3597, w_068_3606, w_068_3608, w_068_3609, w_068_3611, w_068_3613, w_068_3614, w_068_3615, w_068_3616, w_068_3619, w_068_3620, w_068_3621, w_068_3622, w_068_3625, w_068_3626, w_068_3637, w_068_3638, w_068_3645, w_068_3646, w_068_3650, w_068_3654, w_068_3655, w_068_3658, w_068_3662, w_068_3663, w_068_3664, w_068_3667, w_068_3668, w_068_3671, w_068_3674, w_068_3681, w_068_3682, w_068_3683, w_068_3686, w_068_3687, w_068_3689, w_068_3692, w_068_3693, w_068_3698, w_068_3705, w_068_3707, w_068_3709, w_068_3718, w_068_3719, w_068_3720, w_068_3721, w_068_3722, w_068_3725, w_068_3727, w_068_3728, w_068_3729, w_068_3732, w_068_3733, w_068_3738, w_068_3739, w_068_3744, w_068_3746, w_068_3755, w_068_3756, w_068_3759, w_068_3760, w_068_3762, w_068_3769, w_068_3771, w_068_3773, w_068_3775, w_068_3776, w_068_3777, w_068_3778, w_068_3779, w_068_3780, w_068_3781, w_068_3782, w_068_3783, w_068_3788, w_068_3790, w_068_3791, w_068_3793, w_068_3794, w_068_3795, w_068_3796, w_068_3799, w_068_3800, w_068_3802, w_068_3803, w_068_3808, w_068_3809, w_068_3810, w_068_3813, w_068_3814, w_068_3817, w_068_3822, w_068_3825, w_068_3826, w_068_3836, w_068_3840, w_068_3842, w_068_3843, w_068_3844, w_068_3845, w_068_3846, w_068_3851, w_068_3852, w_068_3853, w_068_3864, w_068_3865, w_068_3868, w_068_3870, w_068_3872, w_068_3873, w_068_3874, w_068_3880, w_068_3882, w_068_3889, w_068_3892, w_068_3893, w_068_3895, w_068_3900, w_068_3902, w_068_3904, w_068_3905, w_068_3907, w_068_3909, w_068_3911, w_068_3913, w_068_3914, w_068_3921, w_068_3922, w_068_3935, w_068_3936, w_068_3937, w_068_3938, w_068_3940, w_068_3941, w_068_3943, w_068_3944, w_068_3945, w_068_3947, w_068_3951, w_068_3957, w_068_3960, w_068_3962, w_068_3966, w_068_3969, w_068_3970, w_068_3976, w_068_3977, w_068_3978, w_068_3979, w_068_3980, w_068_3981, w_068_3983, w_068_3984, w_068_3985, w_068_3986, w_068_3990, w_068_3991, w_068_3995, w_068_3996, w_068_3998, w_068_4001, w_068_4014, w_068_4016, w_068_4017, w_068_4018, w_068_4021, w_068_4022, w_068_4025, w_068_4030, w_068_4031, w_068_4033, w_068_4036, w_068_4037, w_068_4038, w_068_4040, w_068_4042, w_068_4045, w_068_4046, w_068_4048, w_068_4051, w_068_4052, w_068_4053, w_068_4056, w_068_4057, w_068_4059, w_068_4061, w_068_4063, w_068_4065, w_068_4066, w_068_4068, w_068_4070, w_068_4071, w_068_4083, w_068_4088, w_068_4092, w_068_4093, w_068_4094, w_068_4095, w_068_4097, w_068_4104, w_068_4108, w_068_4114, w_068_4115, w_068_4122, w_068_4124, w_068_4132, w_068_4134, w_068_4138, w_068_4140, w_068_4141, w_068_4142, w_068_4144, w_068_4145, w_068_4147, w_068_4150, w_068_4152, w_068_4153, w_068_4155, w_068_4158, w_068_4159, w_068_4160, w_068_4161, w_068_4162, w_068_4165, w_068_4169, w_068_4175, w_068_4178, w_068_4180, w_068_4191, w_068_4195, w_068_4197, w_068_4205, w_068_4206, w_068_4211, w_068_4212, w_068_4219, w_068_4220, w_068_4222, w_068_4226, w_068_4227, w_068_4229, w_068_4231, w_068_4233, w_068_4236, w_068_4237, w_068_4239, w_068_4240, w_068_4243, w_068_4251, w_068_4253, w_068_4256, w_068_4267, w_068_4271, w_068_4272, w_068_4274, w_068_4275, w_068_4277, w_068_4281, w_068_4282, w_068_4283, w_068_4284, w_068_4290, w_068_4292, w_068_4293, w_068_4294, w_068_4297, w_068_4301, w_068_4303, w_068_4304, w_068_4307, w_068_4311, w_068_4312, w_068_4315, w_068_4316, w_068_4317, w_068_4318, w_068_4319, w_068_4320, w_068_4321, w_068_4322, w_068_4325, w_068_4327, w_068_4328, w_068_4329, w_068_4331, w_068_4332, w_068_4333, w_068_4335, w_068_4337, w_068_4338, w_068_4339, w_068_4341, w_068_4343, w_068_4345, w_068_4346, w_068_4348, w_068_4350, w_068_4353, w_068_4358, w_068_4360, w_068_4361, w_068_4365, w_068_4367, w_068_4369, w_068_4372, w_068_4373, w_068_4374, w_068_4375, w_068_4380, w_068_4382, w_068_4385, w_068_4389, w_068_4390, w_068_4391, w_068_4394, w_068_4396, w_068_4404, w_068_4411, w_068_4414, w_068_4418, w_068_4432, w_068_4435, w_068_4439, w_068_4440, w_068_4441, w_068_4444, w_068_4448, w_068_4454, w_068_4455, w_068_4457, w_068_4459, w_068_4460, w_068_4461, w_068_4462, w_068_4466, w_068_4468, w_068_4469, w_068_4472, w_068_4474, w_068_4476, w_068_4478, w_068_4480, w_068_4481, w_068_4483, w_068_4484, w_068_4485, w_068_4486, w_068_4487, w_068_4488, w_068_4489, w_068_4492, w_068_4493, w_068_4496, w_068_4499, w_068_4501, w_068_4505, w_068_4507, w_068_4510, w_068_4511, w_068_4512, w_068_4515, w_068_4516, w_068_4519, w_068_4520, w_068_4526, w_068_4531, w_068_4532, w_068_4536, w_068_4537, w_068_4542, w_068_4544, w_068_4550, w_068_4554, w_068_4555, w_068_4557, w_068_4560, w_068_4564, w_068_4568, w_068_4569, w_068_4573, w_068_4575, w_068_4576, w_068_4582, w_068_4583, w_068_4584;
  wire w_069_000, w_069_001, w_069_002, w_069_003, w_069_005, w_069_006, w_069_008, w_069_009, w_069_010, w_069_011, w_069_012, w_069_013, w_069_014, w_069_016, w_069_017, w_069_018, w_069_019, w_069_020, w_069_021, w_069_022, w_069_023, w_069_024, w_069_025, w_069_026, w_069_027, w_069_028, w_069_029, w_069_030, w_069_031, w_069_032, w_069_033, w_069_034, w_069_035, w_069_036, w_069_037, w_069_039, w_069_040, w_069_041, w_069_042, w_069_043, w_069_044, w_069_045, w_069_046, w_069_047, w_069_048, w_069_049, w_069_050, w_069_051, w_069_052, w_069_053, w_069_054, w_069_055, w_069_056, w_069_057, w_069_058, w_069_060, w_069_061, w_069_062, w_069_063, w_069_064, w_069_065, w_069_066, w_069_067, w_069_068, w_069_069, w_069_070, w_069_071, w_069_072, w_069_073, w_069_074, w_069_075, w_069_076, w_069_077, w_069_078, w_069_080, w_069_081, w_069_082, w_069_083, w_069_084, w_069_085, w_069_086, w_069_087, w_069_089, w_069_090, w_069_091, w_069_092, w_069_093, w_069_094, w_069_095, w_069_096, w_069_097, w_069_098, w_069_099, w_069_100, w_069_101, w_069_102, w_069_103, w_069_104, w_069_105, w_069_106, w_069_107, w_069_108, w_069_109, w_069_110, w_069_112, w_069_113, w_069_115, w_069_116, w_069_117, w_069_118, w_069_119, w_069_120, w_069_121, w_069_122, w_069_123, w_069_124, w_069_125, w_069_126, w_069_128, w_069_129, w_069_130, w_069_131, w_069_132, w_069_133, w_069_134, w_069_135, w_069_136, w_069_137, w_069_138, w_069_139, w_069_140, w_069_141, w_069_142, w_069_143, w_069_144, w_069_145, w_069_146, w_069_148, w_069_149, w_069_150, w_069_151, w_069_152, w_069_153, w_069_154, w_069_155, w_069_156, w_069_157, w_069_158, w_069_159, w_069_160, w_069_161, w_069_162, w_069_163, w_069_164, w_069_165, w_069_166, w_069_167, w_069_168, w_069_169, w_069_170, w_069_171, w_069_172, w_069_173, w_069_174, w_069_175, w_069_176, w_069_177, w_069_178, w_069_179, w_069_181, w_069_182, w_069_183, w_069_184, w_069_185, w_069_186, w_069_187, w_069_188, w_069_189, w_069_190, w_069_191, w_069_192, w_069_193, w_069_194, w_069_195, w_069_196, w_069_197, w_069_198, w_069_199, w_069_200, w_069_201, w_069_202, w_069_203, w_069_204, w_069_206, w_069_207, w_069_208, w_069_209, w_069_210, w_069_211, w_069_212, w_069_213, w_069_214, w_069_215, w_069_216, w_069_217, w_069_218, w_069_219, w_069_220, w_069_221, w_069_222, w_069_223, w_069_225, w_069_226, w_069_227, w_069_228, w_069_229, w_069_230, w_069_231, w_069_232, w_069_233, w_069_234, w_069_235, w_069_236, w_069_237, w_069_238, w_069_239, w_069_240, w_069_241, w_069_242, w_069_243, w_069_244, w_069_245, w_069_246, w_069_248, w_069_249, w_069_251, w_069_252, w_069_253, w_069_254, w_069_255, w_069_256, w_069_257, w_069_258, w_069_259, w_069_260, w_069_261, w_069_262, w_069_263, w_069_264, w_069_265, w_069_266, w_069_267, w_069_268, w_069_269, w_069_270, w_069_271, w_069_272, w_069_274, w_069_275, w_069_276, w_069_277, w_069_278, w_069_279, w_069_280, w_069_281, w_069_282, w_069_283, w_069_284, w_069_285, w_069_286, w_069_287, w_069_288, w_069_289, w_069_290, w_069_291, w_069_292, w_069_293, w_069_294, w_069_295, w_069_296, w_069_297, w_069_298, w_069_299, w_069_300, w_069_301, w_069_302, w_069_303, w_069_304, w_069_305, w_069_306, w_069_307, w_069_308, w_069_309, w_069_310, w_069_311, w_069_312, w_069_313, w_069_314, w_069_315, w_069_316, w_069_317, w_069_318, w_069_319, w_069_320, w_069_321, w_069_322, w_069_324, w_069_325, w_069_326, w_069_327, w_069_328, w_069_329, w_069_330, w_069_331, w_069_332, w_069_333, w_069_334, w_069_335, w_069_336, w_069_337, w_069_338, w_069_339, w_069_340, w_069_341, w_069_342, w_069_343, w_069_344, w_069_345, w_069_346, w_069_347, w_069_348, w_069_349, w_069_350, w_069_351, w_069_352, w_069_353, w_069_354, w_069_355, w_069_356, w_069_357, w_069_358, w_069_359, w_069_360, w_069_361, w_069_362, w_069_363, w_069_364, w_069_365, w_069_366, w_069_367, w_069_368, w_069_369, w_069_370, w_069_371, w_069_372, w_069_373, w_069_374, w_069_375, w_069_376, w_069_377, w_069_378, w_069_379, w_069_380, w_069_381, w_069_382, w_069_383, w_069_384, w_069_385, w_069_386, w_069_387, w_069_388, w_069_389, w_069_390, w_069_391, w_069_392, w_069_393, w_069_394, w_069_395, w_069_396, w_069_397, w_069_399, w_069_400, w_069_401, w_069_402, w_069_403, w_069_404, w_069_405, w_069_406, w_069_407, w_069_408, w_069_409, w_069_410, w_069_411, w_069_412, w_069_413, w_069_414, w_069_415, w_069_416, w_069_417, w_069_418, w_069_419, w_069_420, w_069_421, w_069_422, w_069_423, w_069_424, w_069_425, w_069_427, w_069_428, w_069_429, w_069_430, w_069_431, w_069_432, w_069_433, w_069_434, w_069_435, w_069_436, w_069_438, w_069_439, w_069_440, w_069_441, w_069_442, w_069_443, w_069_444, w_069_445, w_069_446, w_069_447, w_069_448, w_069_449, w_069_450, w_069_451, w_069_452, w_069_453, w_069_454, w_069_455, w_069_456, w_069_457, w_069_458, w_069_459, w_069_460, w_069_461, w_069_462, w_069_463, w_069_464, w_069_465, w_069_466, w_069_467, w_069_468, w_069_469, w_069_470, w_069_471, w_069_472, w_069_473, w_069_474, w_069_475, w_069_476, w_069_477, w_069_478, w_069_479, w_069_481, w_069_482, w_069_483, w_069_484, w_069_485, w_069_486, w_069_487, w_069_488, w_069_489, w_069_490, w_069_491, w_069_492, w_069_493, w_069_494, w_069_495, w_069_496, w_069_497, w_069_498, w_069_499, w_069_500, w_069_501, w_069_502, w_069_503, w_069_504, w_069_505, w_069_506, w_069_507, w_069_508, w_069_509, w_069_510, w_069_511, w_069_512, w_069_513, w_069_514, w_069_515, w_069_516, w_069_517, w_069_518, w_069_519, w_069_520, w_069_521, w_069_522, w_069_523, w_069_524, w_069_525, w_069_526, w_069_527, w_069_528, w_069_529, w_069_530, w_069_531, w_069_532, w_069_533, w_069_534, w_069_535, w_069_536, w_069_537, w_069_538, w_069_539, w_069_540, w_069_541, w_069_542, w_069_543, w_069_544, w_069_545, w_069_546, w_069_547, w_069_548, w_069_550, w_069_551, w_069_552, w_069_553, w_069_554, w_069_555, w_069_556, w_069_557, w_069_558, w_069_559, w_069_560, w_069_561, w_069_562, w_069_563, w_069_564, w_069_565, w_069_566, w_069_567, w_069_568, w_069_569, w_069_570, w_069_571, w_069_572, w_069_573, w_069_574, w_069_575, w_069_576, w_069_577, w_069_578, w_069_579, w_069_580, w_069_581, w_069_582, w_069_583, w_069_584, w_069_585, w_069_586, w_069_587, w_069_588, w_069_589, w_069_590, w_069_591, w_069_592, w_069_594, w_069_595, w_069_596, w_069_597, w_069_598, w_069_599, w_069_600, w_069_601, w_069_602, w_069_603, w_069_604, w_069_606, w_069_607, w_069_608, w_069_610, w_069_611, w_069_612, w_069_613, w_069_614, w_069_615, w_069_616, w_069_617, w_069_618, w_069_619, w_069_620, w_069_621, w_069_622, w_069_623, w_069_624, w_069_625, w_069_626, w_069_627, w_069_628, w_069_629, w_069_630, w_069_631, w_069_632, w_069_633, w_069_634, w_069_635, w_069_636, w_069_637, w_069_638, w_069_639, w_069_640, w_069_641, w_069_642, w_069_643, w_069_645, w_069_646, w_069_647, w_069_648, w_069_649, w_069_650, w_069_651, w_069_652, w_069_653, w_069_654, w_069_655, w_069_656, w_069_657, w_069_658, w_069_659, w_069_660, w_069_661, w_069_662, w_069_663, w_069_664, w_069_665, w_069_666, w_069_667, w_069_668, w_069_669, w_069_670, w_069_671, w_069_672, w_069_673, w_069_674, w_069_675, w_069_676, w_069_677, w_069_678, w_069_679, w_069_680, w_069_681, w_069_682, w_069_683, w_069_685, w_069_686, w_069_687, w_069_688, w_069_689, w_069_690, w_069_691, w_069_692, w_069_693, w_069_694, w_069_695, w_069_696, w_069_697, w_069_698, w_069_699, w_069_700, w_069_701, w_069_702, w_069_703, w_069_704, w_069_705, w_069_706, w_069_707, w_069_708, w_069_709, w_069_710, w_069_711, w_069_712, w_069_714, w_069_715, w_069_716, w_069_717;
  wire w_070_000, w_070_001, w_070_002, w_070_003, w_070_004, w_070_005, w_070_007, w_070_008, w_070_009, w_070_010, w_070_012, w_070_013, w_070_014, w_070_015, w_070_016, w_070_017, w_070_018, w_070_021, w_070_022, w_070_024, w_070_025, w_070_026, w_070_027, w_070_028, w_070_029, w_070_031, w_070_032, w_070_034, w_070_036, w_070_037, w_070_038, w_070_039, w_070_040, w_070_041, w_070_042, w_070_043, w_070_044, w_070_046, w_070_049, w_070_050, w_070_051, w_070_052, w_070_054, w_070_056, w_070_057, w_070_059, w_070_060, w_070_061, w_070_064, w_070_065, w_070_066, w_070_067, w_070_068, w_070_069, w_070_070, w_070_071, w_070_072, w_070_073, w_070_074, w_070_075, w_070_076, w_070_078, w_070_079, w_070_080, w_070_081, w_070_082, w_070_083, w_070_084, w_070_085, w_070_087, w_070_089, w_070_091, w_070_092, w_070_093, w_070_094, w_070_095, w_070_096, w_070_097, w_070_099, w_070_100, w_070_101, w_070_102, w_070_103, w_070_104, w_070_105, w_070_107, w_070_109, w_070_110, w_070_111, w_070_112, w_070_113, w_070_114, w_070_115, w_070_116, w_070_117, w_070_118, w_070_120, w_070_121, w_070_122, w_070_123, w_070_124, w_070_125, w_070_126, w_070_131, w_070_132, w_070_134, w_070_136, w_070_137, w_070_139, w_070_140, w_070_143, w_070_145, w_070_146, w_070_147, w_070_148, w_070_149, w_070_150, w_070_151, w_070_152, w_070_154, w_070_155, w_070_157, w_070_158, w_070_159, w_070_160, w_070_161, w_070_162, w_070_163, w_070_165, w_070_167, w_070_168, w_070_169, w_070_170, w_070_172, w_070_173, w_070_174, w_070_175, w_070_176, w_070_177, w_070_179, w_070_181, w_070_183, w_070_184, w_070_185, w_070_186, w_070_187, w_070_188, w_070_189, w_070_191, w_070_192, w_070_196, w_070_197, w_070_198, w_070_199, w_070_201, w_070_204, w_070_205, w_070_206, w_070_207, w_070_209, w_070_211, w_070_212, w_070_214, w_070_216, w_070_217, w_070_219, w_070_220, w_070_223, w_070_224, w_070_225, w_070_227, w_070_228, w_070_229, w_070_230, w_070_231, w_070_232, w_070_233, w_070_234, w_070_235, w_070_236, w_070_237, w_070_238, w_070_239, w_070_240, w_070_241, w_070_242, w_070_244, w_070_247, w_070_248, w_070_249, w_070_250, w_070_251, w_070_252, w_070_255, w_070_256, w_070_258, w_070_259, w_070_260, w_070_261, w_070_262, w_070_263, w_070_264, w_070_265, w_070_266, w_070_267, w_070_273, w_070_274, w_070_275, w_070_276, w_070_277, w_070_278, w_070_280, w_070_281, w_070_282, w_070_283, w_070_285, w_070_286, w_070_289, w_070_290, w_070_291, w_070_292, w_070_293, w_070_294, w_070_295, w_070_297, w_070_298, w_070_299, w_070_300, w_070_301, w_070_303, w_070_305, w_070_306, w_070_307, w_070_308, w_070_309, w_070_312, w_070_314, w_070_315, w_070_316, w_070_318, w_070_320, w_070_321, w_070_322, w_070_323, w_070_324, w_070_325, w_070_326, w_070_327, w_070_328, w_070_329, w_070_330, w_070_331, w_070_334, w_070_335, w_070_336, w_070_337, w_070_339, w_070_340, w_070_341, w_070_342, w_070_343, w_070_344, w_070_346, w_070_347, w_070_348, w_070_350, w_070_351, w_070_352, w_070_353, w_070_354, w_070_355, w_070_356, w_070_357, w_070_358, w_070_359, w_070_360, w_070_364, w_070_365, w_070_368, w_070_369, w_070_370, w_070_371, w_070_373, w_070_374, w_070_375, w_070_376, w_070_377, w_070_378, w_070_379, w_070_380, w_070_381, w_070_383, w_070_384, w_070_385, w_070_386, w_070_388, w_070_390, w_070_394, w_070_395, w_070_397, w_070_398, w_070_399, w_070_400, w_070_401, w_070_402, w_070_403, w_070_404, w_070_405, w_070_406, w_070_408, w_070_410, w_070_415, w_070_416, w_070_417, w_070_418, w_070_419, w_070_420, w_070_421, w_070_423, w_070_424, w_070_426, w_070_429, w_070_430, w_070_431, w_070_432, w_070_433, w_070_434, w_070_436, w_070_438, w_070_439, w_070_440, w_070_441, w_070_443, w_070_444, w_070_445, w_070_446, w_070_448, w_070_449, w_070_450, w_070_456, w_070_458, w_070_459, w_070_460, w_070_461, w_070_462, w_070_463, w_070_464, w_070_466, w_070_469, w_070_470, w_070_471, w_070_472, w_070_473, w_070_475, w_070_477, w_070_478, w_070_480, w_070_481, w_070_483, w_070_484, w_070_485, w_070_486, w_070_488, w_070_489, w_070_491, w_070_493, w_070_494, w_070_495, w_070_497, w_070_498, w_070_499, w_070_500, w_070_501, w_070_505, w_070_506, w_070_507, w_070_508, w_070_509, w_070_510, w_070_511, w_070_512, w_070_513, w_070_514, w_070_515, w_070_516, w_070_517, w_070_518, w_070_519, w_070_520, w_070_522, w_070_523, w_070_524, w_070_526, w_070_527, w_070_528, w_070_530, w_070_531, w_070_532, w_070_533, w_070_535, w_070_536, w_070_539, w_070_540, w_070_542, w_070_543, w_070_544, w_070_545, w_070_547, w_070_548, w_070_550, w_070_551, w_070_552, w_070_554, w_070_555, w_070_556, w_070_559, w_070_560, w_070_561, w_070_562, w_070_563, w_070_564, w_070_565, w_070_567, w_070_569, w_070_572, w_070_573, w_070_575, w_070_576, w_070_577, w_070_579, w_070_580, w_070_581, w_070_583, w_070_585, w_070_587, w_070_588, w_070_591, w_070_592, w_070_593, w_070_594, w_070_595, w_070_597, w_070_598, w_070_600, w_070_601, w_070_602, w_070_603, w_070_604, w_070_605, w_070_607, w_070_608, w_070_609, w_070_612, w_070_613, w_070_615, w_070_616, w_070_618, w_070_619, w_070_620, w_070_621, w_070_622, w_070_623, w_070_624, w_070_625, w_070_626, w_070_627, w_070_629, w_070_630, w_070_631, w_070_632, w_070_633, w_070_634, w_070_635, w_070_636, w_070_637, w_070_638, w_070_639, w_070_640, w_070_641, w_070_642, w_070_644, w_070_645, w_070_647, w_070_648, w_070_649, w_070_650, w_070_651, w_070_652, w_070_653, w_070_655, w_070_656, w_070_658, w_070_659, w_070_660, w_070_662, w_070_663, w_070_664, w_070_665, w_070_666, w_070_668, w_070_669, w_070_670, w_070_672, w_070_673, w_070_674, w_070_675, w_070_676, w_070_677, w_070_678, w_070_679, w_070_680, w_070_684, w_070_686, w_070_687, w_070_689, w_070_691, w_070_694, w_070_695, w_070_696, w_070_698, w_070_699, w_070_700, w_070_701, w_070_702, w_070_703, w_070_704, w_070_705, w_070_706, w_070_707, w_070_708, w_070_709, w_070_710, w_070_712, w_070_714, w_070_715, w_070_716, w_070_717, w_070_718, w_070_719, w_070_720, w_070_721, w_070_722, w_070_723, w_070_724, w_070_726, w_070_727, w_070_728, w_070_730, w_070_731, w_070_732, w_070_733, w_070_734, w_070_735, w_070_736, w_070_737, w_070_738, w_070_739, w_070_740, w_070_741, w_070_742, w_070_743, w_070_744, w_070_745, w_070_746, w_070_747, w_070_748, w_070_749, w_070_752, w_070_753, w_070_754, w_070_755, w_070_756, w_070_757, w_070_758, w_070_760, w_070_763, w_070_764, w_070_766, w_070_770, w_070_771, w_070_772, w_070_774, w_070_776, w_070_780, w_070_781, w_070_782, w_070_784, w_070_785, w_070_786, w_070_788, w_070_789, w_070_790, w_070_791, w_070_792, w_070_793, w_070_795, w_070_796, w_070_797, w_070_798, w_070_799, w_070_800, w_070_801, w_070_802, w_070_803, w_070_804, w_070_806, w_070_807, w_070_808, w_070_809, w_070_810, w_070_811, w_070_812, w_070_813, w_070_814, w_070_815, w_070_816, w_070_818, w_070_821, w_070_824, w_070_826, w_070_827, w_070_828, w_070_829, w_070_830, w_070_831, w_070_834, w_070_835, w_070_836, w_070_837, w_070_838, w_070_839, w_070_840, w_070_842, w_070_843, w_070_844, w_070_847, w_070_848, w_070_849, w_070_850, w_070_851, w_070_854, w_070_855, w_070_856, w_070_857, w_070_858, w_070_859, w_070_860, w_070_862, w_070_863, w_070_865, w_070_866, w_070_867, w_070_868, w_070_869, w_070_870, w_070_872, w_070_873, w_070_874, w_070_875, w_070_877, w_070_878, w_070_879, w_070_881, w_070_882, w_070_883, w_070_884, w_070_885, w_070_886, w_070_887, w_070_890, w_070_891, w_070_892, w_070_894, w_070_895, w_070_896, w_070_897, w_070_898, w_070_899, w_070_900, w_070_901, w_070_902, w_070_903, w_070_904, w_070_905, w_070_906, w_070_907, w_070_908, w_070_910, w_070_911, w_070_912, w_070_913, w_070_914, w_070_915, w_070_916, w_070_918, w_070_919, w_070_920, w_070_921, w_070_922, w_070_923, w_070_924, w_070_925, w_070_926, w_070_927, w_070_928, w_070_930, w_070_931, w_070_932, w_070_933, w_070_934, w_070_935, w_070_936, w_070_937, w_070_938, w_070_939, w_070_943, w_070_945, w_070_946, w_070_948, w_070_950, w_070_951, w_070_953, w_070_954, w_070_955, w_070_956, w_070_957, w_070_959, w_070_960, w_070_961, w_070_962, w_070_963, w_070_964, w_070_965, w_070_966, w_070_969, w_070_970, w_070_973, w_070_975, w_070_976, w_070_977, w_070_979, w_070_980, w_070_981, w_070_982, w_070_983, w_070_984, w_070_986, w_070_987, w_070_989, w_070_990, w_070_992, w_070_994, w_070_995, w_070_996, w_070_997, w_070_998, w_070_999, w_070_1000, w_070_1001, w_070_1002, w_070_1003, w_070_1004, w_070_1005, w_070_1006, w_070_1007, w_070_1010, w_070_1012, w_070_1013, w_070_1014, w_070_1017, w_070_1018, w_070_1019, w_070_1022, w_070_1025, w_070_1027, w_070_1028, w_070_1030, w_070_1031, w_070_1032, w_070_1033, w_070_1034, w_070_1036, w_070_1037, w_070_1041, w_070_1042, w_070_1047, w_070_1049, w_070_1050, w_070_1053, w_070_1054, w_070_1057, w_070_1058, w_070_1059, w_070_1061, w_070_1065, w_070_1066, w_070_1067, w_070_1068, w_070_1069, w_070_1070, w_070_1071, w_070_1072, w_070_1073, w_070_1074, w_070_1075, w_070_1077, w_070_1082, w_070_1088, w_070_1089, w_070_1092, w_070_1093, w_070_1094, w_070_1096, w_070_1097, w_070_1101, w_070_1103, w_070_1105, w_070_1106, w_070_1107, w_070_1110, w_070_1112, w_070_1115, w_070_1116, w_070_1117, w_070_1119, w_070_1123, w_070_1125, w_070_1127, w_070_1129, w_070_1130, w_070_1131, w_070_1134, w_070_1135, w_070_1136, w_070_1138, w_070_1139, w_070_1141, w_070_1142, w_070_1149, w_070_1153, w_070_1154, w_070_1155, w_070_1158, w_070_1160, w_070_1161, w_070_1163, w_070_1164, w_070_1165, w_070_1166, w_070_1167, w_070_1168, w_070_1169, w_070_1170, w_070_1171, w_070_1172, w_070_1173, w_070_1175, w_070_1177, w_070_1178, w_070_1179, w_070_1180, w_070_1181, w_070_1184, w_070_1185, w_070_1187, w_070_1188, w_070_1189, w_070_1191, w_070_1192, w_070_1193, w_070_1194, w_070_1195, w_070_1196, w_070_1197, w_070_1201, w_070_1204, w_070_1206, w_070_1207, w_070_1211, w_070_1214, w_070_1215, w_070_1216, w_070_1217, w_070_1218, w_070_1219, w_070_1221, w_070_1222, w_070_1224, w_070_1225, w_070_1226, w_070_1227, w_070_1230, w_070_1233, w_070_1234, w_070_1235, w_070_1237, w_070_1239, w_070_1240, w_070_1241, w_070_1242, w_070_1245, w_070_1246, w_070_1247, w_070_1248, w_070_1249, w_070_1250, w_070_1251, w_070_1252, w_070_1253, w_070_1254, w_070_1257, w_070_1260, w_070_1261, w_070_1262, w_070_1265, w_070_1266, w_070_1267, w_070_1270, w_070_1272, w_070_1277, w_070_1279, w_070_1280, w_070_1282, w_070_1283, w_070_1285, w_070_1288, w_070_1289, w_070_1290, w_070_1291, w_070_1292, w_070_1297, w_070_1301, w_070_1302, w_070_1303, w_070_1305, w_070_1307, w_070_1311, w_070_1312, w_070_1314, w_070_1315, w_070_1317, w_070_1320, w_070_1321, w_070_1322, w_070_1323, w_070_1326, w_070_1328, w_070_1332, w_070_1336, w_070_1339, w_070_1340, w_070_1341, w_070_1344, w_070_1348, w_070_1350, w_070_1351, w_070_1352, w_070_1353, w_070_1355, w_070_1356, w_070_1357, w_070_1360, w_070_1363, w_070_1365, w_070_1366, w_070_1367, w_070_1369, w_070_1371, w_070_1375, w_070_1376, w_070_1377, w_070_1378, w_070_1379, w_070_1380, w_070_1381, w_070_1382, w_070_1384, w_070_1385, w_070_1386, w_070_1388, w_070_1391, w_070_1393, w_070_1395, w_070_1397, w_070_1398, w_070_1399, w_070_1400, w_070_1402, w_070_1403, w_070_1404, w_070_1405, w_070_1406, w_070_1407, w_070_1409, w_070_1410, w_070_1411, w_070_1413, w_070_1415, w_070_1417, w_070_1418, w_070_1421, w_070_1423, w_070_1424, w_070_1425, w_070_1426, w_070_1435, w_070_1437, w_070_1439, w_070_1441, w_070_1442, w_070_1444, w_070_1447, w_070_1449, w_070_1450, w_070_1452, w_070_1454, w_070_1456, w_070_1459, w_070_1460, w_070_1462, w_070_1463, w_070_1465, w_070_1466, w_070_1468, w_070_1469, w_070_1470, w_070_1471, w_070_1472, w_070_1473, w_070_1474, w_070_1475, w_070_1476, w_070_1477, w_070_1478, w_070_1479, w_070_1480, w_070_1481, w_070_1482, w_070_1483, w_070_1484, w_070_1485, w_070_1486, w_070_1489, w_070_1490, w_070_1491, w_070_1492, w_070_1494, w_070_1495, w_070_1496, w_070_1498, w_070_1499, w_070_1500, w_070_1503, w_070_1505, w_070_1507, w_070_1508, w_070_1509, w_070_1510, w_070_1512, w_070_1513, w_070_1514, w_070_1515, w_070_1516, w_070_1517, w_070_1518, w_070_1520, w_070_1521, w_070_1522, w_070_1523, w_070_1527, w_070_1528, w_070_1529, w_070_1532, w_070_1535, w_070_1537, w_070_1544, w_070_1547, w_070_1549, w_070_1554, w_070_1555, w_070_1556, w_070_1559, w_070_1560, w_070_1561, w_070_1562, w_070_1567, w_070_1572, w_070_1573, w_070_1574, w_070_1575, w_070_1576, w_070_1577, w_070_1578, w_070_1580, w_070_1581, w_070_1583, w_070_1584, w_070_1588, w_070_1589, w_070_1590, w_070_1591, w_070_1592, w_070_1594, w_070_1600, w_070_1601, w_070_1604, w_070_1605, w_070_1606, w_070_1607, w_070_1609, w_070_1610, w_070_1611, w_070_1614, w_070_1615, w_070_1617, w_070_1618, w_070_1619, w_070_1620, w_070_1622, w_070_1624, w_070_1627, w_070_1628, w_070_1629, w_070_1630, w_070_1631, w_070_1632, w_070_1633, w_070_1634, w_070_1635, w_070_1636, w_070_1637, w_070_1639, w_070_1644, w_070_1645, w_070_1646, w_070_1647, w_070_1648, w_070_1649, w_070_1650, w_070_1651, w_070_1653, w_070_1654, w_070_1655, w_070_1656, w_070_1661, w_070_1664, w_070_1669, w_070_1670, w_070_1671, w_070_1672, w_070_1674, w_070_1675, w_070_1677, w_070_1678, w_070_1679, w_070_1680, w_070_1681, w_070_1684, w_070_1686, w_070_1688, w_070_1691, w_070_1692, w_070_1693, w_070_1695, w_070_1699, w_070_1701, w_070_1702, w_070_1703, w_070_1705, w_070_1707, w_070_1708, w_070_1710, w_070_1711, w_070_1712, w_070_1715, w_070_1716, w_070_1719, w_070_1721, w_070_1722, w_070_1723, w_070_1726, w_070_1727, w_070_1728, w_070_1730, w_070_1731, w_070_1733, w_070_1734, w_070_1736, w_070_1737, w_070_1739, w_070_1740, w_070_1742, w_070_1743, w_070_1745, w_070_1746, w_070_1747, w_070_1750, w_070_1754, w_070_1755, w_070_1758, w_070_1759, w_070_1760, w_070_1762, w_070_1763, w_070_1766, w_070_1768, w_070_1772, w_070_1774, w_070_1775, w_070_1776, w_070_1778, w_070_1779, w_070_1780, w_070_1782, w_070_1783, w_070_1785, w_070_1786, w_070_1787, w_070_1788, w_070_1789, w_070_1790, w_070_1791, w_070_1792, w_070_1793, w_070_1796, w_070_1797, w_070_1798, w_070_1800, w_070_1804, w_070_1805, w_070_1806, w_070_1809, w_070_1811, w_070_1812, w_070_1813, w_070_1815, w_070_1816, w_070_1819, w_070_1820, w_070_1822, w_070_1823, w_070_1824, w_070_1825, w_070_1826, w_070_1827, w_070_1828, w_070_1829, w_070_1831, w_070_1832, w_070_1833, w_070_1835, w_070_1836, w_070_1838, w_070_1839, w_070_1840, w_070_1844, w_070_1845, w_070_1846, w_070_1847, w_070_1849, w_070_1850, w_070_1851, w_070_1853, w_070_1855, w_070_1856, w_070_1857, w_070_1858, w_070_1860, w_070_1862, w_070_1863, w_070_1865, w_070_1867, w_070_1868, w_070_1870, w_070_1872, w_070_1875, w_070_1876, w_070_1880, w_070_1881, w_070_1885, w_070_1886, w_070_1889, w_070_1890, w_070_1891, w_070_1893, w_070_1894, w_070_1895, w_070_1897, w_070_1898, w_070_1899, w_070_1900, w_070_1901, w_070_1902, w_070_1906, w_070_1907, w_070_1908, w_070_1910, w_070_1911, w_070_1916, w_070_1917, w_070_1918, w_070_1919, w_070_1920, w_070_1922, w_070_1924, w_070_1926, w_070_1927, w_070_1932, w_070_1933, w_070_1934, w_070_1936, w_070_1938, w_070_1941, w_070_1942, w_070_1945, w_070_1946, w_070_1947, w_070_1948, w_070_1950, w_070_1952, w_070_1953, w_070_1956, w_070_1957, w_070_1958, w_070_1960, w_070_1962, w_070_1963, w_070_1964, w_070_1965, w_070_1966, w_070_1968, w_070_1970, w_070_1971, w_070_1974, w_070_1977, w_070_1979;
  wire w_071_000, w_071_003, w_071_004, w_071_005, w_071_007, w_071_008, w_071_009, w_071_010, w_071_011, w_071_012, w_071_013, w_071_014, w_071_016, w_071_017, w_071_019, w_071_020, w_071_021, w_071_024, w_071_025, w_071_026, w_071_027, w_071_030, w_071_032, w_071_033, w_071_035, w_071_036, w_071_037, w_071_038, w_071_039, w_071_040, w_071_041, w_071_042, w_071_043, w_071_044, w_071_045, w_071_047, w_071_048, w_071_049, w_071_050, w_071_053, w_071_054, w_071_055, w_071_056, w_071_057, w_071_058, w_071_059, w_071_060, w_071_061, w_071_062, w_071_063, w_071_064, w_071_066, w_071_067, w_071_069, w_071_070, w_071_071, w_071_073, w_071_074, w_071_075, w_071_076, w_071_077, w_071_078, w_071_079, w_071_080, w_071_081, w_071_082, w_071_084, w_071_086, w_071_087, w_071_089, w_071_090, w_071_091, w_071_092, w_071_095, w_071_097, w_071_098, w_071_099, w_071_100, w_071_101, w_071_103, w_071_105, w_071_106, w_071_108, w_071_110, w_071_111, w_071_112, w_071_114, w_071_115, w_071_116, w_071_117, w_071_118, w_071_119, w_071_120, w_071_123, w_071_124, w_071_126, w_071_128, w_071_129, w_071_131, w_071_132, w_071_134, w_071_136, w_071_137, w_071_138, w_071_140, w_071_143, w_071_144, w_071_145, w_071_146, w_071_147, w_071_148, w_071_151, w_071_152, w_071_155, w_071_158, w_071_159, w_071_163, w_071_165, w_071_168, w_071_172, w_071_175, w_071_176, w_071_178, w_071_179, w_071_180, w_071_181, w_071_182, w_071_184, w_071_185, w_071_186, w_071_187, w_071_189, w_071_192, w_071_193, w_071_194, w_071_195, w_071_196, w_071_197, w_071_198, w_071_199, w_071_201, w_071_202, w_071_203, w_071_208, w_071_209, w_071_211, w_071_213, w_071_215, w_071_217, w_071_219, w_071_222, w_071_223, w_071_225, w_071_227, w_071_228, w_071_229, w_071_231, w_071_232, w_071_234, w_071_236, w_071_237, w_071_238, w_071_239, w_071_240, w_071_243, w_071_245, w_071_246, w_071_247, w_071_248, w_071_249, w_071_250, w_071_252, w_071_254, w_071_257, w_071_258, w_071_259, w_071_260, w_071_262, w_071_264, w_071_267, w_071_268, w_071_274, w_071_276, w_071_277, w_071_278, w_071_280, w_071_282, w_071_287, w_071_288, w_071_289, w_071_290, w_071_291, w_071_292, w_071_297, w_071_298, w_071_299, w_071_301, w_071_303, w_071_306, w_071_308, w_071_309, w_071_312, w_071_313, w_071_315, w_071_317, w_071_321, w_071_322, w_071_323, w_071_327, w_071_329, w_071_331, w_071_333, w_071_334, w_071_336, w_071_337, w_071_338, w_071_341, w_071_342, w_071_343, w_071_344, w_071_346, w_071_347, w_071_348, w_071_349, w_071_351, w_071_352, w_071_354, w_071_355, w_071_356, w_071_357, w_071_360, w_071_361, w_071_364, w_071_365, w_071_366, w_071_368, w_071_370, w_071_371, w_071_373, w_071_376, w_071_378, w_071_379, w_071_380, w_071_384, w_071_385, w_071_386, w_071_387, w_071_391, w_071_393, w_071_394, w_071_398, w_071_399, w_071_401, w_071_402, w_071_403, w_071_404, w_071_405, w_071_406, w_071_408, w_071_409, w_071_410, w_071_411, w_071_417, w_071_418, w_071_419, w_071_424, w_071_426, w_071_428, w_071_431, w_071_432, w_071_434, w_071_435, w_071_437, w_071_439, w_071_440, w_071_441, w_071_443, w_071_444, w_071_446, w_071_448, w_071_449, w_071_450, w_071_454, w_071_455, w_071_456, w_071_457, w_071_458, w_071_459, w_071_460, w_071_461, w_071_463, w_071_464, w_071_465, w_071_466, w_071_467, w_071_468, w_071_471, w_071_472, w_071_474, w_071_476, w_071_478, w_071_479, w_071_480, w_071_482, w_071_485, w_071_486, w_071_487, w_071_488, w_071_489, w_071_491, w_071_492, w_071_494, w_071_499, w_071_501, w_071_503, w_071_505, w_071_506, w_071_507, w_071_508, w_071_509, w_071_514, w_071_515, w_071_517, w_071_518, w_071_519, w_071_520, w_071_523, w_071_524, w_071_525, w_071_526, w_071_529, w_071_530, w_071_532, w_071_533, w_071_534, w_071_535, w_071_536, w_071_537, w_071_539, w_071_541, w_071_542, w_071_547, w_071_548, w_071_552, w_071_554, w_071_559, w_071_564, w_071_565, w_071_566, w_071_568, w_071_569, w_071_571, w_071_573, w_071_574, w_071_576, w_071_577, w_071_578, w_071_580, w_071_583, w_071_584, w_071_586, w_071_587, w_071_588, w_071_589, w_071_592, w_071_593, w_071_595, w_071_597, w_071_598, w_071_601, w_071_609, w_071_610, w_071_611, w_071_612, w_071_615, w_071_617, w_071_619, w_071_620, w_071_621, w_071_622, w_071_623, w_071_626, w_071_627, w_071_628, w_071_629, w_071_630, w_071_632, w_071_633, w_071_634, w_071_635, w_071_637, w_071_641, w_071_642, w_071_643, w_071_646, w_071_647, w_071_650, w_071_651, w_071_654, w_071_656, w_071_658, w_071_659, w_071_660, w_071_661, w_071_662, w_071_663, w_071_664, w_071_665, w_071_666, w_071_667, w_071_669, w_071_670, w_071_671, w_071_673, w_071_674, w_071_678, w_071_679, w_071_681, w_071_682, w_071_683, w_071_684, w_071_685, w_071_686, w_071_687, w_071_689, w_071_690, w_071_691, w_071_694, w_071_695, w_071_696, w_071_697, w_071_698, w_071_702, w_071_703, w_071_704, w_071_706, w_071_707, w_071_708, w_071_709, w_071_711, w_071_713, w_071_714, w_071_715, w_071_716, w_071_717, w_071_718, w_071_720, w_071_721, w_071_723, w_071_726, w_071_732, w_071_734, w_071_735, w_071_736, w_071_737, w_071_738, w_071_739, w_071_740, w_071_742, w_071_743, w_071_744, w_071_745, w_071_747, w_071_748, w_071_749, w_071_750, w_071_751, w_071_753, w_071_754, w_071_756, w_071_757, w_071_758, w_071_759, w_071_760, w_071_762, w_071_763, w_071_764, w_071_765, w_071_769, w_071_770, w_071_771, w_071_772, w_071_773, w_071_775, w_071_777, w_071_780, w_071_781, w_071_785, w_071_786, w_071_789, w_071_795, w_071_797, w_071_800, w_071_801, w_071_802, w_071_803, w_071_804, w_071_806, w_071_807, w_071_808, w_071_812, w_071_813, w_071_814, w_071_815, w_071_816, w_071_817, w_071_821, w_071_822, w_071_825, w_071_828, w_071_830, w_071_834, w_071_837, w_071_840, w_071_842, w_071_843, w_071_844, w_071_849, w_071_850, w_071_853, w_071_855, w_071_857, w_071_858, w_071_859, w_071_860, w_071_863, w_071_864, w_071_867, w_071_868, w_071_870, w_071_871, w_071_874, w_071_875, w_071_876, w_071_877, w_071_878, w_071_880, w_071_882, w_071_883, w_071_884, w_071_888, w_071_889, w_071_891, w_071_893, w_071_894, w_071_895, w_071_897, w_071_898, w_071_899, w_071_903, w_071_905, w_071_908, w_071_910, w_071_915, w_071_917, w_071_918, w_071_920, w_071_922, w_071_925, w_071_926, w_071_928, w_071_929, w_071_930, w_071_932, w_071_933, w_071_934, w_071_935, w_071_938, w_071_939, w_071_940, w_071_942, w_071_943, w_071_944, w_071_945, w_071_947, w_071_948, w_071_950, w_071_952, w_071_955, w_071_958, w_071_959, w_071_960, w_071_961, w_071_962, w_071_965, w_071_966, w_071_969, w_071_970, w_071_973, w_071_974, w_071_975, w_071_976, w_071_979, w_071_980, w_071_981, w_071_985, w_071_986, w_071_987, w_071_988, w_071_989, w_071_992, w_071_994, w_071_997, w_071_998, w_071_1000, w_071_1001, w_071_1003, w_071_1004, w_071_1005, w_071_1006, w_071_1008, w_071_1009, w_071_1011, w_071_1014, w_071_1016, w_071_1018, w_071_1020, w_071_1021, w_071_1022, w_071_1023, w_071_1025, w_071_1026, w_071_1028, w_071_1029, w_071_1030, w_071_1033, w_071_1034, w_071_1036, w_071_1037, w_071_1038, w_071_1039, w_071_1040, w_071_1041, w_071_1042, w_071_1044, w_071_1045, w_071_1046, w_071_1047, w_071_1048, w_071_1050, w_071_1055, w_071_1056, w_071_1057, w_071_1058, w_071_1059, w_071_1060, w_071_1061, w_071_1062, w_071_1063, w_071_1065, w_071_1066, w_071_1067, w_071_1068, w_071_1070, w_071_1071, w_071_1072, w_071_1073, w_071_1076, w_071_1077, w_071_1079, w_071_1082, w_071_1083, w_071_1084, w_071_1085, w_071_1086, w_071_1087, w_071_1088, w_071_1090, w_071_1091, w_071_1094, w_071_1098, w_071_1100, w_071_1101, w_071_1102, w_071_1103, w_071_1105, w_071_1108, w_071_1109, w_071_1110, w_071_1113, w_071_1114, w_071_1115, w_071_1117, w_071_1118, w_071_1119, w_071_1120, w_071_1121, w_071_1122, w_071_1123, w_071_1124, w_071_1125, w_071_1126, w_071_1127, w_071_1128, w_071_1129, w_071_1131, w_071_1133, w_071_1134, w_071_1135, w_071_1137, w_071_1138, w_071_1140, w_071_1142, w_071_1144, w_071_1148, w_071_1149, w_071_1150, w_071_1152, w_071_1153, w_071_1155, w_071_1156, w_071_1157, w_071_1158, w_071_1161, w_071_1162, w_071_1164, w_071_1165, w_071_1166, w_071_1169, w_071_1170, w_071_1173, w_071_1175, w_071_1178, w_071_1180, w_071_1181, w_071_1182, w_071_1183, w_071_1184, w_071_1186, w_071_1187, w_071_1188, w_071_1193, w_071_1195, w_071_1196, w_071_1199, w_071_1200, w_071_1204, w_071_1205, w_071_1206, w_071_1207, w_071_1208, w_071_1210, w_071_1211, w_071_1212, w_071_1214, w_071_1215, w_071_1216, w_071_1218, w_071_1221, w_071_1222, w_071_1224, w_071_1225, w_071_1226, w_071_1227, w_071_1228, w_071_1230, w_071_1232, w_071_1233, w_071_1235, w_071_1239, w_071_1240, w_071_1241, w_071_1242, w_071_1243, w_071_1244, w_071_1246, w_071_1248, w_071_1250, w_071_1251, w_071_1253, w_071_1254, w_071_1255, w_071_1256, w_071_1258, w_071_1260, w_071_1262, w_071_1263, w_071_1264, w_071_1267, w_071_1268, w_071_1269, w_071_1270, w_071_1271, w_071_1272, w_071_1274, w_071_1275, w_071_1277, w_071_1279, w_071_1280, w_071_1281, w_071_1285, w_071_1286, w_071_1288, w_071_1289, w_071_1291, w_071_1292, w_071_1294, w_071_1295, w_071_1296, w_071_1297, w_071_1298, w_071_1300, w_071_1301, w_071_1302, w_071_1306, w_071_1307, w_071_1308, w_071_1310, w_071_1314, w_071_1315, w_071_1316, w_071_1318, w_071_1319, w_071_1321, w_071_1322, w_071_1323, w_071_1324, w_071_1326, w_071_1327, w_071_1329, w_071_1330, w_071_1331, w_071_1335, w_071_1336, w_071_1338, w_071_1339, w_071_1340, w_071_1342, w_071_1344, w_071_1346, w_071_1350, w_071_1351, w_071_1352, w_071_1354, w_071_1355, w_071_1357, w_071_1360, w_071_1361, w_071_1364, w_071_1366, w_071_1370, w_071_1373, w_071_1374, w_071_1375, w_071_1376, w_071_1377, w_071_1380, w_071_1382, w_071_1385, w_071_1386, w_071_1388, w_071_1389, w_071_1390, w_071_1391, w_071_1393, w_071_1394, w_071_1397, w_071_1398, w_071_1399, w_071_1401, w_071_1402, w_071_1403, w_071_1404, w_071_1405, w_071_1408, w_071_1409, w_071_1410, w_071_1411, w_071_1413, w_071_1414, w_071_1415, w_071_1416, w_071_1417, w_071_1418, w_071_1420, w_071_1425, w_071_1429, w_071_1430, w_071_1434, w_071_1435, w_071_1438, w_071_1441, w_071_1444, w_071_1447, w_071_1448, w_071_1450, w_071_1451, w_071_1454, w_071_1455, w_071_1456, w_071_1457, w_071_1459, w_071_1461, w_071_1467, w_071_1468, w_071_1470, w_071_1472, w_071_1473, w_071_1478, w_071_1479, w_071_1481, w_071_1482, w_071_1484, w_071_1486, w_071_1488, w_071_1489, w_071_1491, w_071_1493, w_071_1494, w_071_1500, w_071_1501, w_071_1504, w_071_1505, w_071_1507, w_071_1508, w_071_1510, w_071_1511, w_071_1512, w_071_1514, w_071_1515, w_071_1516, w_071_1520, w_071_1521, w_071_1522, w_071_1524, w_071_1525, w_071_1526, w_071_1531, w_071_1532, w_071_1533, w_071_1534, w_071_1536, w_071_1537, w_071_1538, w_071_1539, w_071_1541, w_071_1543, w_071_1547, w_071_1548, w_071_1551, w_071_1552, w_071_1554, w_071_1555, w_071_1556, w_071_1557, w_071_1558, w_071_1559, w_071_1560, w_071_1562, w_071_1564, w_071_1565, w_071_1566, w_071_1567, w_071_1568, w_071_1569, w_071_1572, w_071_1573, w_071_1575, w_071_1580, w_071_1581, w_071_1583, w_071_1584, w_071_1585, w_071_1587, w_071_1588, w_071_1590, w_071_1593, w_071_1596, w_071_1597, w_071_1599, w_071_1600, w_071_1602, w_071_1604, w_071_1606, w_071_1607, w_071_1609, w_071_1611, w_071_1613, w_071_1614, w_071_1617, w_071_1618, w_071_1619, w_071_1620, w_071_1623, w_071_1626, w_071_1627, w_071_1628, w_071_1629, w_071_1630, w_071_1631, w_071_1633, w_071_1634, w_071_1635, w_071_1636, w_071_1638, w_071_1639, w_071_1640, w_071_1642, w_071_1643, w_071_1647, w_071_1648, w_071_1649, w_071_1650, w_071_1651, w_071_1652, w_071_1656, w_071_1657, w_071_1659, w_071_1660, w_071_1661, w_071_1663, w_071_1667, w_071_1668, w_071_1669, w_071_1670, w_071_1671, w_071_1672, w_071_1673, w_071_1676, w_071_1678, w_071_1680, w_071_1681, w_071_1684, w_071_1685, w_071_1686, w_071_1687, w_071_1688, w_071_1689, w_071_1690, w_071_1691, w_071_1692, w_071_1693, w_071_1694, w_071_1696, w_071_1698, w_071_1699, w_071_1700, w_071_1701, w_071_1703, w_071_1704, w_071_1707, w_071_1709, w_071_1711, w_071_1712, w_071_1714, w_071_1716, w_071_1717, w_071_1718, w_071_1721, w_071_1722, w_071_1723, w_071_1724, w_071_1725, w_071_1726, w_071_1727, w_071_1729, w_071_1732, w_071_1733, w_071_1736, w_071_1741, w_071_1742, w_071_1744, w_071_1745, w_071_1746, w_071_1748, w_071_1749, w_071_1750, w_071_1753, w_071_1755, w_071_1757, w_071_1758, w_071_1759, w_071_1760, w_071_1762, w_071_1765, w_071_1766, w_071_1767, w_071_1769, w_071_1770, w_071_1771, w_071_1772, w_071_1773, w_071_1774, w_071_1775, w_071_1776, w_071_1777, w_071_1778, w_071_1779, w_071_1782, w_071_1783, w_071_1785, w_071_1787, w_071_1788, w_071_1789, w_071_1790, w_071_1792, w_071_1793, w_071_1794, w_071_1797, w_071_1798, w_071_1799, w_071_1801, w_071_1803, w_071_1804, w_071_1806, w_071_1807, w_071_1809, w_071_1813, w_071_1815, w_071_1816, w_071_1817, w_071_1818, w_071_1820, w_071_1821, w_071_1822, w_071_1823, w_071_1824, w_071_1825, w_071_1826, w_071_1827, w_071_1831, w_071_1832, w_071_1833, w_071_1834, w_071_1837, w_071_1844, w_071_1845, w_071_1847, w_071_1848, w_071_1850, w_071_1852, w_071_1854, w_071_1856, w_071_1857, w_071_1858, w_071_1859, w_071_1862, w_071_1863, w_071_1864, w_071_1866, w_071_1867, w_071_1868, w_071_1869, w_071_1871, w_071_1873, w_071_1874, w_071_1876, w_071_1877, w_071_1882, w_071_1883, w_071_1884, w_071_1885, w_071_1886, w_071_1887, w_071_1890, w_071_1891, w_071_1895, w_071_1898, w_071_1899, w_071_1900, w_071_1901, w_071_1902, w_071_1903, w_071_1906, w_071_1907, w_071_1910, w_071_1911, w_071_1912, w_071_1913, w_071_1915, w_071_1918, w_071_1919, w_071_1920, w_071_1922, w_071_1923, w_071_1924, w_071_1925, w_071_1926, w_071_1930, w_071_1931, w_071_1934, w_071_1938, w_071_1940, w_071_1942, w_071_1946, w_071_1947, w_071_1950, w_071_1951, w_071_1952, w_071_1953, w_071_1956, w_071_1957, w_071_1958, w_071_1959, w_071_1961, w_071_1964, w_071_1966, w_071_1968, w_071_1969, w_071_1970, w_071_1971, w_071_1974, w_071_1976, w_071_1978, w_071_1979, w_071_1981, w_071_1982, w_071_1984, w_071_1985, w_071_1986, w_071_1987, w_071_1988, w_071_1989, w_071_1990, w_071_1993, w_071_1994, w_071_1995, w_071_1996, w_071_1997, w_071_2000, w_071_2004, w_071_2006, w_071_2007, w_071_2008, w_071_2009, w_071_2010, w_071_2013, w_071_2014, w_071_2015, w_071_2016, w_071_2017, w_071_2020, w_071_2021, w_071_2023, w_071_2024, w_071_2025, w_071_2027, w_071_2028, w_071_2029, w_071_2030, w_071_2031, w_071_2032, w_071_2034, w_071_2035, w_071_2037, w_071_2041, w_071_2043, w_071_2046, w_071_2049, w_071_2050, w_071_2052, w_071_2053, w_071_2054, w_071_2055, w_071_2057, w_071_2058, w_071_2064, w_071_2065, w_071_2066, w_071_2068, w_071_2069, w_071_2070, w_071_2072, w_071_2074, w_071_2076, w_071_2079, w_071_2081, w_071_2082, w_071_2083, w_071_2086, w_071_2087, w_071_2088, w_071_2089, w_071_2090, w_071_2092, w_071_2094, w_071_2096, w_071_2097, w_071_2101, w_071_2102, w_071_2103, w_071_2104, w_071_2105, w_071_2107, w_071_2108, w_071_2109, w_071_2112, w_071_2115, w_071_2116, w_071_2117, w_071_2118, w_071_2120, w_071_2122, w_071_2126, w_071_2127, w_071_2128, w_071_2129, w_071_2130, w_071_2132, w_071_2134, w_071_2135, w_071_2136, w_071_2137, w_071_2138, w_071_2139, w_071_2141, w_071_2143, w_071_2145, w_071_2147, w_071_2148, w_071_2150, w_071_2151, w_071_2154, w_071_2155, w_071_2156, w_071_2157, w_071_2158, w_071_2165, w_071_2166, w_071_2167, w_071_2169, w_071_2170, w_071_2171, w_071_2174, w_071_2176, w_071_2177, w_071_2178, w_071_2179, w_071_2182, w_071_2183, w_071_2184, w_071_2185, w_071_2186, w_071_2188, w_071_2190, w_071_2191, w_071_2192, w_071_2194, w_071_2195, w_071_2197, w_071_2198, w_071_2199, w_071_2201, w_071_2202, w_071_2204, w_071_2208, w_071_2212, w_071_2213, w_071_2214, w_071_2215, w_071_2216, w_071_2217, w_071_2222, w_071_2223, w_071_2226, w_071_2227, w_071_2228, w_071_2229, w_071_2230, w_071_2232, w_071_2236, w_071_2239, w_071_2242, w_071_2243, w_071_2245, w_071_2246, w_071_2248, w_071_2249, w_071_2250, w_071_2252, w_071_2253, w_071_2254, w_071_2255, w_071_2260, w_071_2262, w_071_2263, w_071_2265, w_071_2266, w_071_2267, w_071_2271, w_071_2272, w_071_2273, w_071_2274, w_071_2276, w_071_2277, w_071_2282, w_071_2283, w_071_2285, w_071_2286, w_071_2287, w_071_2294, w_071_2295, w_071_2297, w_071_2298, w_071_2300, w_071_2301, w_071_2302, w_071_2304, w_071_2307, w_071_2308, w_071_2309, w_071_2311, w_071_2312, w_071_2313, w_071_2314, w_071_2319, w_071_2320, w_071_2321, w_071_2324, w_071_2328, w_071_2331, w_071_2332, w_071_2333, w_071_2334, w_071_2337, w_071_2339, w_071_2340, w_071_2343, w_071_2344, w_071_2346, w_071_2347, w_071_2349, w_071_2350, w_071_2354, w_071_2356, w_071_2357, w_071_2358, w_071_2359, w_071_2361, w_071_2374, w_071_2375, w_071_2377, w_071_2378, w_071_2379, w_071_2385, w_071_2386, w_071_2387, w_071_2388, w_071_2394, w_071_2397, w_071_2398, w_071_2399, w_071_2400, w_071_2404, w_071_2406, w_071_2407, w_071_2408, w_071_2409, w_071_2411, w_071_2412, w_071_2415, w_071_2416, w_071_2417, w_071_2420, w_071_2421, w_071_2423, w_071_2424, w_071_2426, w_071_2428, w_071_2430, w_071_2431, w_071_2433, w_071_2434, w_071_2435, w_071_2436, w_071_2437, w_071_2438, w_071_2439, w_071_2442, w_071_2443, w_071_2446, w_071_2448, w_071_2450, w_071_2452, w_071_2453, w_071_2454, w_071_2455, w_071_2456, w_071_2457, w_071_2458, w_071_2459, w_071_2460, w_071_2462, w_071_2464, w_071_2465, w_071_2466, w_071_2467, w_071_2468, w_071_2469, w_071_2470, w_071_2471, w_071_2473;
  wire w_072_000, w_072_001, w_072_002, w_072_003, w_072_004, w_072_005, w_072_006, w_072_007, w_072_008, w_072_009, w_072_010, w_072_011, w_072_013, w_072_014, w_072_015, w_072_016, w_072_017, w_072_018, w_072_019, w_072_020, w_072_021, w_072_022, w_072_023, w_072_024, w_072_025, w_072_026, w_072_027, w_072_028, w_072_029, w_072_030, w_072_031, w_072_032, w_072_035, w_072_036, w_072_037, w_072_038, w_072_039, w_072_040, w_072_042, w_072_043, w_072_044, w_072_045, w_072_046, w_072_047, w_072_048, w_072_049, w_072_050, w_072_051, w_072_052, w_072_053, w_072_054, w_072_055, w_072_056, w_072_057, w_072_058, w_072_059, w_072_060, w_072_061, w_072_062, w_072_063, w_072_064, w_072_065, w_072_066, w_072_067, w_072_068, w_072_069, w_072_070, w_072_071, w_072_072, w_072_073, w_072_074, w_072_075, w_072_076, w_072_077, w_072_078, w_072_079, w_072_080, w_072_081, w_072_082, w_072_083, w_072_084, w_072_085, w_072_086, w_072_087, w_072_088, w_072_089, w_072_090, w_072_091, w_072_092, w_072_093, w_072_094, w_072_095, w_072_096, w_072_097, w_072_098, w_072_099, w_072_100, w_072_101, w_072_102, w_072_103, w_072_104, w_072_105, w_072_106, w_072_107, w_072_108, w_072_109, w_072_110, w_072_111, w_072_112, w_072_113, w_072_114, w_072_115, w_072_116, w_072_117, w_072_118, w_072_119, w_072_120, w_072_121, w_072_122, w_072_123, w_072_124, w_072_125, w_072_126, w_072_127, w_072_128, w_072_129, w_072_130, w_072_131, w_072_132, w_072_133, w_072_134, w_072_135, w_072_136, w_072_137, w_072_138, w_072_139, w_072_140, w_072_141, w_072_142, w_072_143, w_072_144, w_072_145, w_072_146, w_072_147, w_072_148, w_072_149, w_072_150, w_072_151, w_072_152, w_072_153, w_072_154, w_072_155, w_072_156, w_072_157, w_072_158, w_072_159, w_072_160, w_072_161, w_072_162, w_072_163, w_072_164, w_072_165, w_072_166, w_072_167, w_072_168, w_072_169, w_072_170, w_072_171, w_072_172, w_072_173, w_072_174, w_072_175, w_072_176, w_072_177, w_072_178, w_072_179, w_072_180, w_072_181, w_072_182, w_072_183, w_072_184, w_072_185, w_072_186, w_072_188, w_072_189, w_072_190, w_072_191, w_072_192, w_072_193, w_072_194, w_072_195, w_072_196, w_072_197, w_072_198, w_072_199, w_072_200, w_072_201, w_072_202, w_072_203, w_072_204, w_072_205, w_072_206, w_072_207, w_072_208, w_072_209, w_072_210, w_072_211, w_072_212, w_072_213, w_072_214, w_072_215, w_072_216, w_072_217, w_072_218, w_072_219, w_072_220, w_072_221, w_072_222, w_072_223, w_072_224, w_072_225, w_072_226, w_072_227, w_072_228, w_072_229, w_072_230, w_072_231, w_072_232, w_072_233, w_072_234, w_072_235, w_072_236, w_072_237, w_072_238, w_072_239, w_072_240, w_072_241, w_072_242, w_072_243, w_072_244, w_072_245, w_072_246, w_072_247, w_072_248, w_072_249, w_072_250, w_072_251, w_072_252, w_072_253, w_072_254, w_072_255, w_072_256, w_072_258, w_072_259, w_072_260, w_072_261, w_072_262, w_072_263, w_072_264, w_072_265, w_072_266, w_072_268, w_072_269, w_072_270, w_072_271, w_072_272, w_072_273, w_072_274, w_072_275, w_072_276, w_072_277, w_072_278, w_072_280, w_072_281, w_072_282, w_072_283, w_072_284, w_072_285, w_072_286, w_072_287, w_072_288, w_072_289, w_072_290, w_072_291, w_072_292, w_072_293, w_072_294, w_072_295, w_072_296, w_072_297, w_072_298, w_072_299, w_072_300, w_072_301, w_072_302, w_072_303, w_072_304, w_072_305, w_072_306, w_072_307, w_072_308, w_072_309, w_072_310, w_072_311, w_072_312, w_072_313, w_072_314, w_072_315, w_072_316, w_072_318, w_072_319, w_072_320, w_072_321, w_072_322, w_072_323, w_072_324, w_072_325, w_072_326, w_072_327, w_072_329, w_072_330, w_072_331, w_072_332, w_072_333, w_072_334, w_072_335, w_072_336, w_072_337, w_072_338, w_072_339, w_072_340, w_072_341, w_072_342, w_072_343, w_072_344, w_072_345, w_072_346, w_072_347, w_072_348, w_072_349, w_072_350, w_072_351, w_072_352, w_072_353, w_072_354, w_072_355, w_072_356, w_072_357, w_072_358, w_072_359, w_072_360, w_072_361, w_072_362, w_072_363, w_072_364, w_072_365, w_072_366, w_072_367, w_072_368, w_072_369, w_072_370, w_072_371, w_072_372, w_072_373, w_072_374, w_072_375, w_072_376, w_072_377, w_072_379, w_072_380, w_072_381, w_072_382, w_072_383, w_072_384, w_072_385, w_072_386, w_072_387, w_072_388, w_072_389, w_072_390, w_072_391, w_072_392, w_072_393, w_072_394, w_072_395, w_072_396, w_072_397, w_072_398, w_072_399, w_072_401, w_072_402, w_072_403, w_072_404, w_072_405, w_072_407, w_072_409, w_072_410, w_072_411, w_072_412, w_072_413, w_072_414, w_072_415, w_072_416, w_072_417, w_072_418, w_072_419, w_072_420, w_072_421, w_072_422, w_072_423, w_072_424, w_072_426, w_072_427, w_072_428, w_072_429, w_072_430, w_072_431, w_072_432, w_072_433, w_072_434, w_072_435, w_072_436, w_072_437, w_072_438, w_072_439, w_072_440, w_072_441, w_072_442, w_072_443, w_072_444, w_072_445, w_072_446, w_072_447, w_072_448, w_072_449, w_072_450, w_072_451, w_072_452, w_072_453, w_072_454, w_072_455, w_072_456, w_072_457, w_072_458, w_072_459, w_072_461, w_072_462, w_072_464, w_072_465, w_072_466, w_072_467, w_072_468, w_072_469, w_072_470, w_072_471, w_072_472, w_072_473, w_072_474, w_072_475, w_072_476, w_072_477, w_072_478, w_072_479, w_072_480, w_072_481, w_072_482, w_072_483, w_072_484, w_072_486, w_072_487, w_072_488, w_072_489, w_072_490, w_072_491, w_072_492, w_072_493, w_072_494, w_072_495, w_072_496, w_072_497, w_072_498, w_072_499, w_072_500, w_072_501, w_072_502, w_072_503, w_072_504, w_072_505, w_072_506, w_072_507, w_072_508, w_072_509, w_072_510, w_072_512, w_072_513, w_072_514, w_072_515, w_072_516, w_072_517, w_072_518, w_072_519, w_072_520, w_072_521, w_072_522, w_072_523, w_072_524, w_072_525, w_072_526, w_072_527, w_072_528, w_072_529, w_072_530, w_072_531, w_072_532, w_072_533, w_072_534, w_072_535, w_072_536, w_072_537, w_072_538, w_072_539, w_072_540, w_072_541, w_072_542, w_072_543, w_072_544, w_072_545, w_072_546, w_072_547, w_072_548, w_072_549, w_072_550, w_072_551, w_072_552, w_072_553, w_072_555, w_072_556, w_072_557, w_072_558, w_072_559, w_072_561, w_072_562, w_072_563, w_072_564, w_072_565, w_072_566, w_072_567, w_072_568, w_072_569, w_072_570, w_072_571, w_072_572, w_072_573, w_072_574, w_072_575, w_072_576, w_072_577, w_072_578, w_072_579, w_072_580, w_072_581, w_072_582, w_072_583, w_072_584, w_072_585, w_072_586, w_072_587, w_072_588, w_072_589, w_072_590, w_072_591, w_072_592, w_072_593, w_072_594, w_072_595, w_072_596, w_072_597, w_072_598, w_072_599, w_072_600, w_072_601, w_072_602, w_072_603, w_072_604, w_072_605, w_072_606, w_072_607, w_072_608, w_072_609, w_072_610, w_072_611, w_072_612, w_072_613, w_072_614, w_072_615, w_072_616, w_072_617, w_072_618, w_072_619, w_072_620, w_072_621, w_072_622, w_072_623, w_072_624, w_072_625, w_072_626, w_072_627, w_072_629, w_072_630, w_072_631, w_072_632, w_072_633, w_072_634, w_072_635, w_072_636, w_072_637, w_072_639, w_072_640, w_072_641, w_072_642, w_072_643, w_072_644;
  wire w_073_000, w_073_001, w_073_004, w_073_005, w_073_007, w_073_008, w_073_009, w_073_011, w_073_013, w_073_019, w_073_022, w_073_023, w_073_024, w_073_025, w_073_026, w_073_029, w_073_030, w_073_033, w_073_034, w_073_035, w_073_036, w_073_037, w_073_040, w_073_044, w_073_047, w_073_048, w_073_050, w_073_051, w_073_052, w_073_055, w_073_056, w_073_057, w_073_058, w_073_060, w_073_061, w_073_062, w_073_064, w_073_065, w_073_070, w_073_074, w_073_076, w_073_079, w_073_080, w_073_081, w_073_082, w_073_083, w_073_084, w_073_086, w_073_087, w_073_089, w_073_091, w_073_093, w_073_094, w_073_095, w_073_097, w_073_098, w_073_100, w_073_101, w_073_102, w_073_104, w_073_105, w_073_108, w_073_109, w_073_112, w_073_113, w_073_115, w_073_119, w_073_120, w_073_124, w_073_125, w_073_127, w_073_129, w_073_130, w_073_132, w_073_133, w_073_136, w_073_137, w_073_138, w_073_140, w_073_142, w_073_144, w_073_145, w_073_148, w_073_150, w_073_151, w_073_152, w_073_154, w_073_155, w_073_156, w_073_157, w_073_158, w_073_159, w_073_160, w_073_161, w_073_162, w_073_163, w_073_164, w_073_168, w_073_169, w_073_172, w_073_173, w_073_179, w_073_181, w_073_182, w_073_183, w_073_184, w_073_186, w_073_187, w_073_189, w_073_190, w_073_191, w_073_192, w_073_194, w_073_195, w_073_196, w_073_197, w_073_200, w_073_202, w_073_203, w_073_204, w_073_206, w_073_209, w_073_210, w_073_213, w_073_214, w_073_215, w_073_218, w_073_219, w_073_221, w_073_224, w_073_226, w_073_227, w_073_228, w_073_229, w_073_230, w_073_233, w_073_234, w_073_238, w_073_239, w_073_240, w_073_241, w_073_242, w_073_244, w_073_245, w_073_247, w_073_248, w_073_249, w_073_250, w_073_252, w_073_254, w_073_256, w_073_258, w_073_259, w_073_260, w_073_261, w_073_263, w_073_264, w_073_265, w_073_267, w_073_268, w_073_271, w_073_272, w_073_276, w_073_278, w_073_279, w_073_281, w_073_282, w_073_284, w_073_285, w_073_286, w_073_287, w_073_290, w_073_291, w_073_292, w_073_293, w_073_294, w_073_295, w_073_299, w_073_300, w_073_301, w_073_303, w_073_305, w_073_306, w_073_308, w_073_309, w_073_314, w_073_315, w_073_316, w_073_319, w_073_321, w_073_323, w_073_324, w_073_325, w_073_327, w_073_328, w_073_329, w_073_330, w_073_331, w_073_332, w_073_333, w_073_338, w_073_339, w_073_340, w_073_343, w_073_345, w_073_346, w_073_347, w_073_348, w_073_351, w_073_352, w_073_353, w_073_356, w_073_358, w_073_361, w_073_364, w_073_365, w_073_368, w_073_370, w_073_371, w_073_373, w_073_376, w_073_377, w_073_380, w_073_381, w_073_383, w_073_385, w_073_386, w_073_387, w_073_390, w_073_395, w_073_396, w_073_398, w_073_400, w_073_402, w_073_403, w_073_404, w_073_406, w_073_408, w_073_409, w_073_410, w_073_412, w_073_414, w_073_416, w_073_419, w_073_421, w_073_423, w_073_424, w_073_425, w_073_426, w_073_429, w_073_430, w_073_432, w_073_433, w_073_434, w_073_435, w_073_438, w_073_439, w_073_442, w_073_444, w_073_446, w_073_447, w_073_449, w_073_450, w_073_451, w_073_452, w_073_454, w_073_455, w_073_456, w_073_457, w_073_458, w_073_461, w_073_463, w_073_466, w_073_467, w_073_468, w_073_469, w_073_470, w_073_473, w_073_475, w_073_476, w_073_478, w_073_479, w_073_480, w_073_481, w_073_482, w_073_484, w_073_487, w_073_491, w_073_492, w_073_493, w_073_494, w_073_495, w_073_496, w_073_498, w_073_500, w_073_501, w_073_506, w_073_507, w_073_509, w_073_512, w_073_515, w_073_516, w_073_518, w_073_520, w_073_522, w_073_524, w_073_525, w_073_527, w_073_529, w_073_532, w_073_535, w_073_536, w_073_537, w_073_540, w_073_542, w_073_543, w_073_544, w_073_546, w_073_547, w_073_548, w_073_550, w_073_551, w_073_552, w_073_553, w_073_554, w_073_556, w_073_557, w_073_559, w_073_564, w_073_565, w_073_566, w_073_571, w_073_572, w_073_573, w_073_574, w_073_576, w_073_579, w_073_580, w_073_583, w_073_585, w_073_586, w_073_587, w_073_589, w_073_591, w_073_594, w_073_596, w_073_598, w_073_599, w_073_600, w_073_601, w_073_602, w_073_604, w_073_607, w_073_608, w_073_611, w_073_612, w_073_617, w_073_618, w_073_619, w_073_620, w_073_621, w_073_622, w_073_623, w_073_624, w_073_625, w_073_627, w_073_631, w_073_632, w_073_633, w_073_634, w_073_636, w_073_638, w_073_640, w_073_641, w_073_644, w_073_645, w_073_646, w_073_649, w_073_653, w_073_655, w_073_656, w_073_657, w_073_658, w_073_659, w_073_660, w_073_664, w_073_665, w_073_666, w_073_667, w_073_668, w_073_670, w_073_672, w_073_674, w_073_676, w_073_677, w_073_681, w_073_688, w_073_689, w_073_690, w_073_692, w_073_693, w_073_695, w_073_696, w_073_697, w_073_702, w_073_703, w_073_704, w_073_706, w_073_708, w_073_709, w_073_711, w_073_713, w_073_715, w_073_716, w_073_717, w_073_719, w_073_720, w_073_723, w_073_725, w_073_726, w_073_727, w_073_728, w_073_729, w_073_731, w_073_733, w_073_734, w_073_736, w_073_737, w_073_738, w_073_739, w_073_740, w_073_741, w_073_742, w_073_745, w_073_746, w_073_747, w_073_748, w_073_749, w_073_751, w_073_755, w_073_756, w_073_759, w_073_760, w_073_761, w_073_763, w_073_764, w_073_765, w_073_769, w_073_770, w_073_772, w_073_773, w_073_774, w_073_775, w_073_776, w_073_777, w_073_780, w_073_782, w_073_783, w_073_788, w_073_789, w_073_792, w_073_794, w_073_795, w_073_796, w_073_797, w_073_798, w_073_799, w_073_800, w_073_802, w_073_804, w_073_809, w_073_812, w_073_813, w_073_814, w_073_815, w_073_816, w_073_817, w_073_818, w_073_820, w_073_821, w_073_823, w_073_825, w_073_828, w_073_830, w_073_831, w_073_833, w_073_834, w_073_835, w_073_836, w_073_838, w_073_840, w_073_842, w_073_843, w_073_845, w_073_849, w_073_851, w_073_852, w_073_853, w_073_854, w_073_855, w_073_856, w_073_857, w_073_858, w_073_860, w_073_862, w_073_863, w_073_864, w_073_865, w_073_867, w_073_869, w_073_870, w_073_871, w_073_872, w_073_875, w_073_876, w_073_877, w_073_878, w_073_880, w_073_881, w_073_883, w_073_885, w_073_886, w_073_888, w_073_889, w_073_892, w_073_893, w_073_897, w_073_900, w_073_901, w_073_902, w_073_903, w_073_904, w_073_905, w_073_907, w_073_908, w_073_910, w_073_911, w_073_912, w_073_913, w_073_914, w_073_916, w_073_917, w_073_918, w_073_920, w_073_921, w_073_922, w_073_926, w_073_927, w_073_930, w_073_931, w_073_933, w_073_934, w_073_935, w_073_936, w_073_938, w_073_939, w_073_940, w_073_941, w_073_943, w_073_946, w_073_947, w_073_948, w_073_951, w_073_952, w_073_955, w_073_956, w_073_957, w_073_960, w_073_961, w_073_963, w_073_964, w_073_965, w_073_967, w_073_968, w_073_969, w_073_970, w_073_971, w_073_974, w_073_976, w_073_977, w_073_979, w_073_980, w_073_982, w_073_983, w_073_984, w_073_987, w_073_988, w_073_991, w_073_992, w_073_994, w_073_995, w_073_997, w_073_1001, w_073_1003, w_073_1005, w_073_1006, w_073_1007, w_073_1010, w_073_1011, w_073_1012, w_073_1015, w_073_1016, w_073_1018, w_073_1019, w_073_1021, w_073_1023, w_073_1025, w_073_1029, w_073_1031, w_073_1040, w_073_1041, w_073_1043, w_073_1044, w_073_1045, w_073_1046, w_073_1047, w_073_1048, w_073_1049, w_073_1051, w_073_1052, w_073_1053, w_073_1054, w_073_1055, w_073_1058, w_073_1059, w_073_1060, w_073_1061, w_073_1064, w_073_1065, w_073_1066, w_073_1068, w_073_1069, w_073_1072, w_073_1073, w_073_1074, w_073_1077, w_073_1079, w_073_1081, w_073_1082, w_073_1083, w_073_1084, w_073_1085, w_073_1086, w_073_1090, w_073_1092, w_073_1093, w_073_1094, w_073_1099, w_073_1100, w_073_1101, w_073_1103, w_073_1108, w_073_1111, w_073_1112, w_073_1113, w_073_1114, w_073_1115, w_073_1117, w_073_1119, w_073_1120, w_073_1121, w_073_1122, w_073_1123, w_073_1124, w_073_1125, w_073_1126, w_073_1133, w_073_1134, w_073_1137, w_073_1138, w_073_1139, w_073_1142, w_073_1147, w_073_1148, w_073_1149, w_073_1150, w_073_1153, w_073_1155, w_073_1156, w_073_1161, w_073_1162, w_073_1164, w_073_1165, w_073_1166, w_073_1167, w_073_1168, w_073_1169, w_073_1170, w_073_1171, w_073_1172, w_073_1173, w_073_1174, w_073_1175, w_073_1178, w_073_1180, w_073_1182, w_073_1184, w_073_1186, w_073_1190, w_073_1193, w_073_1195, w_073_1197, w_073_1198, w_073_1199, w_073_1200, w_073_1201, w_073_1202, w_073_1203, w_073_1207, w_073_1208, w_073_1209, w_073_1210, w_073_1212, w_073_1214, w_073_1215, w_073_1216, w_073_1217, w_073_1219, w_073_1220, w_073_1222, w_073_1223, w_073_1224, w_073_1227, w_073_1228, w_073_1229, w_073_1230, w_073_1231, w_073_1232, w_073_1234, w_073_1235, w_073_1236, w_073_1239, w_073_1241, w_073_1242, w_073_1243, w_073_1245, w_073_1246, w_073_1247, w_073_1250, w_073_1251, w_073_1252, w_073_1255, w_073_1257, w_073_1258, w_073_1259, w_073_1260, w_073_1261, w_073_1262, w_073_1263, w_073_1264, w_073_1265, w_073_1266, w_073_1269, w_073_1271, w_073_1273, w_073_1274, w_073_1276, w_073_1278, w_073_1281, w_073_1283, w_073_1284, w_073_1285, w_073_1287, w_073_1290, w_073_1291, w_073_1292, w_073_1296, w_073_1297, w_073_1298, w_073_1303, w_073_1311, w_073_1313, w_073_1315, w_073_1317, w_073_1318, w_073_1321, w_073_1324, w_073_1325, w_073_1327, w_073_1328, w_073_1329, w_073_1331, w_073_1332, w_073_1333, w_073_1334, w_073_1338, w_073_1340, w_073_1341, w_073_1342, w_073_1343, w_073_1344, w_073_1346, w_073_1348, w_073_1351, w_073_1352, w_073_1353, w_073_1354, w_073_1355, w_073_1356, w_073_1357, w_073_1359, w_073_1360, w_073_1363, w_073_1364, w_073_1365, w_073_1367, w_073_1368, w_073_1369, w_073_1373, w_073_1375, w_073_1376, w_073_1379, w_073_1381, w_073_1383, w_073_1386, w_073_1387, w_073_1388, w_073_1389, w_073_1390, w_073_1391, w_073_1397, w_073_1407, w_073_1410, w_073_1412, w_073_1415, w_073_1417, w_073_1418, w_073_1419, w_073_1420, w_073_1421, w_073_1422, w_073_1423, w_073_1424, w_073_1429, w_073_1430, w_073_1431, w_073_1432, w_073_1433, w_073_1436, w_073_1437, w_073_1438, w_073_1439, w_073_1440, w_073_1441, w_073_1442, w_073_1444, w_073_1447, w_073_1448, w_073_1449, w_073_1450, w_073_1451, w_073_1452, w_073_1456, w_073_1457, w_073_1459, w_073_1460, w_073_1461, w_073_1462, w_073_1464, w_073_1465, w_073_1467, w_073_1470, w_073_1471, w_073_1472, w_073_1476, w_073_1477, w_073_1478, w_073_1480, w_073_1485, w_073_1487, w_073_1489, w_073_1492, w_073_1493, w_073_1494, w_073_1495, w_073_1498, w_073_1499, w_073_1500, w_073_1503, w_073_1509, w_073_1510, w_073_1512, w_073_1513, w_073_1514, w_073_1517, w_073_1519, w_073_1520, w_073_1522, w_073_1526, w_073_1528, w_073_1529, w_073_1530, w_073_1532, w_073_1534, w_073_1535, w_073_1536, w_073_1539, w_073_1540, w_073_1542, w_073_1543, w_073_1544, w_073_1545, w_073_1549, w_073_1551, w_073_1552, w_073_1555, w_073_1556, w_073_1557, w_073_1558, w_073_1560, w_073_1562, w_073_1563, w_073_1567, w_073_1568, w_073_1569, w_073_1570, w_073_1572, w_073_1573, w_073_1576, w_073_1578, w_073_1579, w_073_1581, w_073_1582, w_073_1583, w_073_1584, w_073_1585, w_073_1587, w_073_1588, w_073_1590, w_073_1592, w_073_1600, w_073_1602, w_073_1603, w_073_1604, w_073_1605, w_073_1607, w_073_1610, w_073_1615, w_073_1616, w_073_1617, w_073_1621, w_073_1623, w_073_1625, w_073_1626, w_073_1627, w_073_1631, w_073_1633, w_073_1634, w_073_1635, w_073_1639, w_073_1641, w_073_1642, w_073_1643, w_073_1646, w_073_1647, w_073_1648, w_073_1650, w_073_1652, w_073_1653, w_073_1655, w_073_1657, w_073_1663, w_073_1666, w_073_1669, w_073_1671, w_073_1677, w_073_1678, w_073_1682, w_073_1684, w_073_1690, w_073_1693, w_073_1694, w_073_1695, w_073_1698, w_073_1700, w_073_1701, w_073_1702, w_073_1705, w_073_1706, w_073_1708, w_073_1711, w_073_1712, w_073_1714, w_073_1722, w_073_1726, w_073_1728, w_073_1729, w_073_1730, w_073_1733, w_073_1734, w_073_1736, w_073_1738, w_073_1740, w_073_1750, w_073_1755, w_073_1758, w_073_1759, w_073_1761, w_073_1770, w_073_1777, w_073_1782, w_073_1783, w_073_1784, w_073_1786, w_073_1787, w_073_1790, w_073_1791, w_073_1794, w_073_1795, w_073_1806, w_073_1808, w_073_1811, w_073_1812, w_073_1813, w_073_1816, w_073_1817, w_073_1819, w_073_1822, w_073_1824, w_073_1825, w_073_1827, w_073_1829, w_073_1831, w_073_1833, w_073_1835, w_073_1841, w_073_1843, w_073_1849, w_073_1852, w_073_1855, w_073_1856, w_073_1859, w_073_1862, w_073_1864, w_073_1865, w_073_1866, w_073_1867, w_073_1868, w_073_1869, w_073_1870, w_073_1873, w_073_1874, w_073_1877, w_073_1881, w_073_1884, w_073_1886, w_073_1890, w_073_1892, w_073_1895, w_073_1899, w_073_1900, w_073_1901, w_073_1903, w_073_1905, w_073_1907, w_073_1908, w_073_1909, w_073_1912, w_073_1914, w_073_1915, w_073_1916, w_073_1917, w_073_1920, w_073_1921, w_073_1925, w_073_1929, w_073_1930, w_073_1933, w_073_1939, w_073_1940, w_073_1942, w_073_1947, w_073_1949, w_073_1950, w_073_1951, w_073_1954, w_073_1955, w_073_1957, w_073_1958, w_073_1959, w_073_1961, w_073_1964, w_073_1965, w_073_1967, w_073_1968, w_073_1971, w_073_1972, w_073_1974, w_073_1975, w_073_1982, w_073_1986, w_073_1989, w_073_1994, w_073_1999, w_073_2000, w_073_2001, w_073_2013, w_073_2015, w_073_2017, w_073_2025, w_073_2028, w_073_2031, w_073_2036, w_073_2037, w_073_2040, w_073_2051, w_073_2057, w_073_2058, w_073_2060, w_073_2062, w_073_2063, w_073_2065, w_073_2071, w_073_2072, w_073_2076, w_073_2077, w_073_2078, w_073_2079, w_073_2082, w_073_2083, w_073_2094, w_073_2098, w_073_2100, w_073_2110, w_073_2113, w_073_2121, w_073_2130, w_073_2131, w_073_2132, w_073_2133, w_073_2137, w_073_2142, w_073_2143, w_073_2158, w_073_2160, w_073_2162, w_073_2163, w_073_2166, w_073_2168, w_073_2171, w_073_2173, w_073_2175, w_073_2176, w_073_2178, w_073_2186, w_073_2196, w_073_2198, w_073_2200, w_073_2201, w_073_2204, w_073_2205, w_073_2210, w_073_2211, w_073_2222, w_073_2223, w_073_2231, w_073_2234, w_073_2236, w_073_2239, w_073_2240, w_073_2243, w_073_2244, w_073_2246, w_073_2251, w_073_2253, w_073_2254, w_073_2259, w_073_2260, w_073_2261, w_073_2265, w_073_2268, w_073_2269, w_073_2270, w_073_2271, w_073_2272, w_073_2273, w_073_2274, w_073_2275, w_073_2277, w_073_2284, w_073_2287, w_073_2290, w_073_2292, w_073_2297, w_073_2298, w_073_2299, w_073_2300, w_073_2302, w_073_2306, w_073_2307, w_073_2309, w_073_2319, w_073_2322, w_073_2323, w_073_2335, w_073_2337, w_073_2340, w_073_2341, w_073_2348, w_073_2349, w_073_2353, w_073_2364, w_073_2369, w_073_2370, w_073_2373, w_073_2374, w_073_2378, w_073_2383, w_073_2384, w_073_2389, w_073_2393, w_073_2395, w_073_2396, w_073_2397, w_073_2404, w_073_2410, w_073_2411, w_073_2412, w_073_2414, w_073_2416, w_073_2417, w_073_2418, w_073_2419, w_073_2420, w_073_2421, w_073_2424, w_073_2425, w_073_2428, w_073_2443, w_073_2444, w_073_2445, w_073_2449, w_073_2451, w_073_2453, w_073_2455, w_073_2458, w_073_2459, w_073_2462, w_073_2463, w_073_2466, w_073_2467, w_073_2468, w_073_2477, w_073_2478, w_073_2479, w_073_2481, w_073_2482, w_073_2493, w_073_2503, w_073_2504, w_073_2509, w_073_2510, w_073_2517, w_073_2520, w_073_2526, w_073_2527, w_073_2529, w_073_2531, w_073_2533, w_073_2539, w_073_2541, w_073_2542, w_073_2543, w_073_2544, w_073_2545, w_073_2549, w_073_2551, w_073_2557, w_073_2558, w_073_2560, w_073_2564, w_073_2565, w_073_2566, w_073_2567, w_073_2570, w_073_2571, w_073_2574, w_073_2575, w_073_2577, w_073_2582, w_073_2584, w_073_2585, w_073_2588, w_073_2589, w_073_2591, w_073_2594, w_073_2605, w_073_2610, w_073_2612, w_073_2613, w_073_2621, w_073_2623, w_073_2624, w_073_2626, w_073_2630, w_073_2635, w_073_2637, w_073_2644, w_073_2647, w_073_2649, w_073_2651, w_073_2654, w_073_2658, w_073_2663, w_073_2667, w_073_2668, w_073_2670, w_073_2672, w_073_2674, w_073_2679, w_073_2683, w_073_2685, w_073_2687, w_073_2690, w_073_2692, w_073_2695, w_073_2700, w_073_2702, w_073_2703, w_073_2704, w_073_2706, w_073_2707, w_073_2710, w_073_2712, w_073_2718, w_073_2720, w_073_2723, w_073_2725, w_073_2726, w_073_2727, w_073_2728, w_073_2729, w_073_2730, w_073_2733, w_073_2737, w_073_2738, w_073_2739, w_073_2740, w_073_2744, w_073_2746, w_073_2748, w_073_2752, w_073_2756, w_073_2759, w_073_2768, w_073_2774, w_073_2779, w_073_2780, w_073_2783, w_073_2784, w_073_2785, w_073_2792, w_073_2795, w_073_2799, w_073_2800, w_073_2801, w_073_2802, w_073_2804, w_073_2807, w_073_2811, w_073_2815, w_073_2819, w_073_2820, w_073_2822, w_073_2825, w_073_2836, w_073_2839, w_073_2845, w_073_2846, w_073_2847, w_073_2849, w_073_2850, w_073_2852, w_073_2853, w_073_2854, w_073_2855, w_073_2858, w_073_2859, w_073_2863, w_073_2870, w_073_2871, w_073_2877, w_073_2880, w_073_2882, w_073_2883, w_073_2885, w_073_2887, w_073_2891, w_073_2895, w_073_2897, w_073_2898, w_073_2900, w_073_2901, w_073_2902, w_073_2905, w_073_2907, w_073_2910, w_073_2911, w_073_2917, w_073_2919, w_073_2920, w_073_2922, w_073_2928, w_073_2939, w_073_2943, w_073_2948, w_073_2950, w_073_2951, w_073_2953, w_073_2954, w_073_2956, w_073_2957, w_073_2959, w_073_2962, w_073_2963, w_073_2964, w_073_2975, w_073_2982, w_073_2985, w_073_2986, w_073_2987, w_073_2989, w_073_2990, w_073_2991, w_073_2997, w_073_2999, w_073_3001, w_073_3002, w_073_3004, w_073_3006, w_073_3009, w_073_3017, w_073_3019, w_073_3021, w_073_3024, w_073_3028, w_073_3029, w_073_3031, w_073_3032, w_073_3034, w_073_3038, w_073_3039, w_073_3042, w_073_3045, w_073_3047, w_073_3050, w_073_3051, w_073_3053, w_073_3054, w_073_3056, w_073_3057, w_073_3061, w_073_3064, w_073_3067, w_073_3069, w_073_3071, w_073_3073, w_073_3074, w_073_3075, w_073_3083, w_073_3088, w_073_3092, w_073_3093, w_073_3095, w_073_3096, w_073_3100, w_073_3103, w_073_3104, w_073_3105, w_073_3110, w_073_3111, w_073_3112, w_073_3115, w_073_3117, w_073_3118, w_073_3123, w_073_3124, w_073_3127, w_073_3131, w_073_3132, w_073_3136, w_073_3140, w_073_3142, w_073_3147, w_073_3149, w_073_3151, w_073_3155, w_073_3164, w_073_3166, w_073_3168, w_073_3169, w_073_3170, w_073_3171, w_073_3173, w_073_3181, w_073_3182, w_073_3183, w_073_3185, w_073_3190, w_073_3191, w_073_3194, w_073_3197, w_073_3199, w_073_3201, w_073_3207, w_073_3208, w_073_3209, w_073_3212, w_073_3214, w_073_3215, w_073_3221, w_073_3223, w_073_3225, w_073_3230, w_073_3234, w_073_3239, w_073_3246, w_073_3248, w_073_3250, w_073_3252, w_073_3255, w_073_3259, w_073_3262, w_073_3268, w_073_3269, w_073_3270, w_073_3271, w_073_3272, w_073_3274, w_073_3275, w_073_3277, w_073_3281, w_073_3288, w_073_3293, w_073_3295, w_073_3299, w_073_3301, w_073_3302, w_073_3303, w_073_3304, w_073_3305, w_073_3310, w_073_3311, w_073_3318, w_073_3324, w_073_3333, w_073_3336, w_073_3342, w_073_3344, w_073_3347, w_073_3348, w_073_3352;
  wire w_074_001, w_074_002, w_074_004, w_074_005, w_074_008, w_074_009, w_074_010, w_074_011, w_074_012, w_074_014, w_074_015, w_074_016, w_074_017, w_074_018, w_074_019, w_074_020, w_074_021, w_074_022, w_074_023, w_074_024, w_074_025, w_074_026, w_074_028, w_074_030, w_074_031, w_074_032, w_074_033, w_074_034, w_074_035, w_074_036, w_074_037, w_074_038, w_074_039, w_074_042, w_074_045, w_074_046, w_074_048, w_074_049, w_074_051, w_074_056, w_074_057, w_074_058, w_074_059, w_074_060, w_074_062, w_074_063, w_074_064, w_074_066, w_074_067, w_074_070, w_074_071, w_074_072, w_074_073, w_074_074, w_074_075, w_074_078, w_074_079, w_074_081, w_074_082, w_074_083, w_074_085, w_074_087, w_074_088, w_074_089, w_074_090, w_074_091, w_074_092, w_074_093, w_074_094, w_074_095, w_074_096, w_074_098, w_074_099, w_074_100, w_074_102, w_074_106, w_074_108, w_074_111, w_074_114, w_074_115, w_074_117, w_074_118, w_074_119, w_074_120, w_074_121, w_074_123, w_074_124, w_074_125, w_074_126, w_074_127, w_074_128, w_074_130, w_074_131, w_074_132, w_074_133, w_074_135, w_074_136, w_074_137, w_074_138, w_074_139, w_074_140, w_074_141, w_074_142, w_074_143, w_074_144, w_074_146, w_074_147, w_074_149, w_074_150, w_074_152, w_074_153, w_074_154, w_074_155, w_074_156, w_074_157, w_074_158, w_074_159, w_074_160, w_074_161, w_074_162, w_074_163, w_074_164, w_074_166, w_074_168, w_074_169, w_074_170, w_074_172, w_074_173, w_074_176, w_074_177, w_074_179, w_074_180, w_074_181, w_074_182, w_074_183, w_074_185, w_074_186, w_074_187, w_074_188, w_074_190, w_074_191, w_074_192, w_074_193, w_074_194, w_074_195, w_074_197, w_074_199, w_074_201, w_074_202, w_074_203, w_074_204, w_074_205, w_074_206, w_074_207, w_074_208, w_074_210, w_074_211, w_074_213, w_074_214, w_074_215, w_074_217, w_074_218, w_074_219, w_074_220, w_074_221, w_074_222, w_074_223, w_074_224, w_074_225, w_074_226, w_074_227, w_074_229, w_074_230, w_074_232, w_074_233, w_074_235, w_074_236, w_074_237, w_074_238, w_074_239, w_074_240, w_074_242, w_074_243, w_074_244, w_074_246, w_074_248, w_074_249, w_074_251, w_074_253, w_074_254, w_074_255, w_074_256, w_074_257, w_074_258, w_074_259, w_074_260, w_074_262, w_074_264, w_074_267, w_074_268, w_074_270, w_074_271, w_074_272, w_074_273, w_074_274, w_074_275, w_074_276, w_074_277, w_074_278, w_074_279, w_074_280, w_074_281, w_074_282, w_074_283, w_074_284, w_074_285, w_074_286, w_074_287, w_074_288, w_074_289, w_074_290, w_074_291, w_074_292, w_074_293, w_074_294, w_074_295, w_074_296, w_074_298, w_074_299, w_074_300, w_074_303, w_074_304, w_074_305, w_074_306, w_074_307, w_074_308, w_074_311, w_074_312, w_074_313, w_074_314, w_074_315, w_074_317, w_074_318, w_074_319, w_074_321, w_074_322, w_074_325, w_074_326, w_074_327, w_074_328, w_074_329, w_074_330, w_074_331, w_074_332, w_074_333, w_074_334, w_074_335, w_074_336, w_074_337, w_074_338, w_074_339, w_074_342, w_074_343, w_074_344, w_074_345, w_074_347, w_074_348, w_074_349, w_074_350, w_074_351, w_074_352, w_074_353, w_074_354, w_074_355, w_074_356, w_074_358, w_074_359, w_074_360, w_074_362, w_074_365, w_074_366, w_074_369, w_074_370, w_074_371, w_074_372, w_074_373, w_074_374, w_074_375, w_074_376, w_074_381, w_074_382, w_074_383, w_074_384, w_074_385, w_074_386, w_074_387, w_074_388, w_074_389, w_074_390, w_074_391, w_074_393, w_074_394, w_074_395, w_074_396, w_074_397, w_074_400, w_074_401, w_074_402, w_074_403, w_074_404, w_074_406, w_074_407, w_074_408, w_074_409, w_074_411, w_074_412, w_074_414, w_074_415, w_074_416, w_074_418, w_074_419, w_074_421, w_074_423, w_074_424, w_074_425, w_074_427, w_074_428, w_074_429, w_074_430, w_074_431, w_074_432, w_074_434, w_074_435, w_074_436, w_074_438, w_074_439, w_074_440, w_074_441, w_074_442, w_074_443, w_074_445, w_074_446, w_074_447, w_074_448, w_074_450, w_074_451, w_074_453, w_074_454, w_074_455, w_074_456, w_074_459, w_074_460, w_074_461, w_074_462, w_074_463, w_074_465, w_074_466, w_074_467, w_074_468, w_074_469, w_074_470, w_074_473, w_074_475, w_074_476, w_074_477, w_074_481, w_074_482, w_074_483, w_074_484, w_074_485, w_074_486, w_074_487, w_074_489, w_074_490, w_074_491, w_074_492, w_074_494, w_074_495, w_074_496, w_074_497, w_074_498, w_074_499, w_074_500, w_074_502, w_074_503, w_074_504, w_074_506, w_074_507, w_074_511, w_074_512, w_074_513, w_074_514, w_074_515, w_074_516, w_074_517, w_074_518, w_074_519, w_074_520, w_074_522, w_074_525, w_074_526, w_074_527, w_074_528, w_074_529, w_074_530, w_074_532, w_074_534, w_074_535, w_074_536, w_074_537, w_074_538, w_074_539, w_074_540, w_074_541, w_074_542, w_074_543, w_074_544, w_074_545, w_074_546, w_074_547, w_074_548, w_074_549, w_074_550, w_074_551, w_074_552, w_074_553, w_074_554, w_074_556, w_074_557, w_074_558, w_074_559, w_074_560, w_074_563, w_074_564, w_074_565, w_074_566, w_074_569, w_074_570, w_074_572, w_074_573, w_074_574, w_074_575, w_074_576, w_074_577, w_074_578, w_074_580, w_074_581, w_074_582, w_074_584, w_074_585, w_074_586, w_074_587, w_074_589, w_074_591, w_074_593, w_074_594, w_074_595, w_074_596, w_074_598, w_074_599, w_074_600, w_074_602, w_074_603, w_074_605, w_074_606, w_074_607, w_074_608, w_074_609, w_074_610, w_074_612, w_074_613, w_074_614, w_074_615, w_074_616, w_074_618, w_074_620, w_074_621, w_074_622, w_074_623, w_074_625, w_074_628, w_074_629, w_074_631, w_074_632, w_074_633, w_074_635, w_074_636, w_074_637, w_074_638, w_074_639, w_074_640, w_074_641, w_074_643, w_074_645, w_074_646, w_074_647, w_074_648, w_074_651, w_074_654, w_074_655, w_074_656, w_074_657, w_074_658, w_074_659, w_074_660, w_074_662, w_074_664, w_074_666, w_074_667, w_074_668, w_074_671, w_074_672, w_074_673, w_074_674, w_074_676, w_074_678, w_074_679, w_074_681, w_074_682, w_074_683, w_074_684, w_074_685, w_074_688, w_074_689, w_074_691, w_074_694, w_074_697, w_074_698, w_074_700, w_074_702, w_074_703, w_074_704, w_074_705, w_074_707, w_074_709, w_074_710, w_074_712, w_074_713, w_074_715, w_074_716, w_074_718, w_074_720, w_074_721, w_074_722, w_074_723, w_074_724, w_074_725, w_074_726, w_074_728, w_074_730, w_074_731, w_074_734, w_074_735, w_074_736, w_074_738, w_074_739, w_074_740, w_074_743, w_074_744, w_074_745, w_074_746, w_074_749, w_074_750, w_074_751, w_074_752, w_074_753, w_074_754, w_074_755, w_074_757, w_074_758, w_074_759, w_074_764, w_074_765, w_074_766, w_074_767, w_074_769, w_074_770, w_074_771, w_074_772, w_074_773, w_074_774, w_074_775, w_074_776, w_074_777, w_074_779, w_074_781, w_074_782, w_074_783, w_074_784, w_074_785, w_074_786, w_074_787, w_074_788, w_074_789, w_074_790, w_074_791, w_074_792, w_074_793, w_074_794, w_074_796, w_074_797, w_074_799, w_074_801, w_074_802, w_074_803, w_074_804, w_074_805, w_074_808, w_074_809, w_074_812, w_074_813, w_074_816, w_074_818, w_074_819, w_074_820, w_074_822, w_074_824, w_074_825, w_074_827, w_074_828, w_074_829, w_074_832, w_074_833, w_074_835, w_074_837, w_074_839, w_074_840, w_074_841, w_074_842, w_074_843, w_074_845, w_074_846, w_074_847, w_074_848, w_074_850, w_074_851, w_074_852, w_074_853, w_074_854, w_074_858, w_074_859, w_074_860, w_074_862, w_074_863, w_074_864, w_074_865, w_074_867, w_074_868, w_074_872, w_074_873, w_074_874, w_074_875, w_074_876, w_074_878, w_074_879, w_074_880, w_074_881, w_074_882, w_074_883, w_074_884, w_074_885, w_074_886, w_074_887, w_074_889, w_074_891, w_074_893, w_074_894, w_074_895, w_074_897, w_074_898, w_074_900, w_074_901, w_074_902, w_074_903, w_074_904, w_074_905, w_074_907, w_074_908, w_074_909, w_074_910, w_074_911, w_074_912, w_074_913, w_074_914, w_074_915, w_074_916, w_074_917, w_074_918, w_074_920, w_074_921, w_074_922, w_074_923, w_074_924, w_074_925, w_074_926, w_074_927, w_074_928, w_074_929, w_074_932, w_074_933, w_074_934, w_074_936, w_074_937, w_074_938, w_074_940, w_074_942, w_074_943, w_074_944, w_074_946, w_074_947, w_074_948, w_074_949, w_074_950, w_074_951, w_074_952, w_074_954, w_074_955, w_074_957, w_074_959, w_074_960, w_074_961, w_074_962, w_074_963, w_074_964, w_074_966, w_074_968, w_074_969, w_074_970, w_074_971, w_074_972, w_074_973, w_074_974, w_074_975, w_074_977, w_074_978, w_074_979, w_074_981, w_074_982, w_074_984, w_074_985, w_074_986, w_074_987, w_074_988, w_074_989, w_074_990, w_074_992, w_074_994, w_074_998, w_074_999, w_074_1000, w_074_1001, w_074_1002, w_074_1004, w_074_1005, w_074_1006, w_074_1007, w_074_1009, w_074_1010, w_074_1011, w_074_1012, w_074_1013, w_074_1015, w_074_1017, w_074_1018, w_074_1019, w_074_1020, w_074_1021, w_074_1022, w_074_1023, w_074_1024, w_074_1025, w_074_1028, w_074_1030, w_074_1034, w_074_1035, w_074_1036, w_074_1037, w_074_1038, w_074_1039, w_074_1040, w_074_1041, w_074_1043, w_074_1044, w_074_1045, w_074_1046, w_074_1047, w_074_1048, w_074_1049, w_074_1052, w_074_1053, w_074_1054, w_074_1056, w_074_1057, w_074_1058, w_074_1059, w_074_1061, w_074_1062, w_074_1063, w_074_1064, w_074_1065, w_074_1068, w_074_1070, w_074_1071, w_074_1072, w_074_1073, w_074_1074, w_074_1075, w_074_1076, w_074_1077, w_074_1081, w_074_1082, w_074_1083, w_074_1084, w_074_1086, w_074_1087, w_074_1088, w_074_1090, w_074_1091, w_074_1092, w_074_1093, w_074_1094, w_074_1095, w_074_1096, w_074_1097, w_074_1099, w_074_1100, w_074_1101, w_074_1102, w_074_1103, w_074_1106, w_074_1107, w_074_1111, w_074_1112, w_074_1113, w_074_1115, w_074_1117, w_074_1118, w_074_1122, w_074_1124, w_074_1125, w_074_1126, w_074_1127, w_074_1128, w_074_1130, w_074_1131, w_074_1132, w_074_1133, w_074_1134, w_074_1135, w_074_1136, w_074_1139, w_074_1141, w_074_1142, w_074_1143, w_074_1145, w_074_1147, w_074_1148, w_074_1150, w_074_1151, w_074_1152, w_074_1153, w_074_1154, w_074_1155, w_074_1156, w_074_1157, w_074_1159, w_074_1160, w_074_1162, w_074_1164, w_074_1165, w_074_1166, w_074_1168, w_074_1170, w_074_1171, w_074_1174, w_074_1176, w_074_1179, w_074_1180, w_074_1183, w_074_1184, w_074_1185, w_074_1187, w_074_1189, w_074_1190, w_074_1191, w_074_1194, w_074_1196, w_074_1198, w_074_1199, w_074_1203, w_074_1204, w_074_1205, w_074_1207, w_074_1210, w_074_1211, w_074_1213, w_074_1215, w_074_1216, w_074_1219, w_074_1221, w_074_1223, w_074_1224, w_074_1225, w_074_1228, w_074_1230, w_074_1231, w_074_1232, w_074_1237, w_074_1238, w_074_1240, w_074_1243, w_074_1245, w_074_1248, w_074_1249, w_074_1251, w_074_1252, w_074_1257, w_074_1258, w_074_1259, w_074_1263, w_074_1266, w_074_1270, w_074_1272, w_074_1274, w_074_1275, w_074_1278, w_074_1280, w_074_1284, w_074_1287, w_074_1288, w_074_1289, w_074_1293, w_074_1294, w_074_1297, w_074_1298, w_074_1299, w_074_1300, w_074_1305, w_074_1307, w_074_1308, w_074_1309, w_074_1311, w_074_1312, w_074_1315, w_074_1316, w_074_1317, w_074_1318, w_074_1319, w_074_1320, w_074_1322, w_074_1323, w_074_1324, w_074_1325, w_074_1326, w_074_1327, w_074_1330, w_074_1331, w_074_1332, w_074_1333, w_074_1334, w_074_1335, w_074_1336, w_074_1337, w_074_1338, w_074_1341, w_074_1343, w_074_1346, w_074_1347, w_074_1348, w_074_1350, w_074_1351, w_074_1352, w_074_1353, w_074_1355, w_074_1357, w_074_1359, w_074_1360, w_074_1361, w_074_1362, w_074_1363, w_074_1364, w_074_1365, w_074_1366, w_074_1369, w_074_1370, w_074_1372, w_074_1373, w_074_1378, w_074_1380, w_074_1382, w_074_1384, w_074_1387, w_074_1388, w_074_1390, w_074_1391, w_074_1393, w_074_1395, w_074_1396, w_074_1397, w_074_1398, w_074_1399, w_074_1400, w_074_1401, w_074_1402, w_074_1403, w_074_1404, w_074_1405, w_074_1406, w_074_1408, w_074_1410, w_074_1413, w_074_1415, w_074_1416, w_074_1417, w_074_1419, w_074_1420, w_074_1425, w_074_1426, w_074_1428, w_074_1429, w_074_1432, w_074_1433, w_074_1436, w_074_1437, w_074_1438, w_074_1439, w_074_1440, w_074_1442, w_074_1444, w_074_1447, w_074_1449, w_074_1450, w_074_1451, w_074_1452, w_074_1453, w_074_1454, w_074_1457, w_074_1458, w_074_1460, w_074_1461, w_074_1462, w_074_1463, w_074_1464, w_074_1465, w_074_1467, w_074_1471, w_074_1472, w_074_1473, w_074_1474, w_074_1476, w_074_1477, w_074_1479, w_074_1480, w_074_1481, w_074_1482, w_074_1483, w_074_1484, w_074_1485, w_074_1486, w_074_1487, w_074_1488, w_074_1489, w_074_1491, w_074_1493, w_074_1496, w_074_1497, w_074_1498, w_074_1499, w_074_1500, w_074_1502, w_074_1503, w_074_1504, w_074_1508, w_074_1509, w_074_1510, w_074_1511, w_074_1512, w_074_1516, w_074_1517, w_074_1518, w_074_1519, w_074_1520, w_074_1521, w_074_1522, w_074_1523, w_074_1524, w_074_1525, w_074_1526, w_074_1527, w_074_1531, w_074_1534, w_074_1535, w_074_1537, w_074_1538, w_074_1540, w_074_1542, w_074_1544, w_074_1545, w_074_1547, w_074_1549, w_074_1551, w_074_1555, w_074_1556, w_074_1557, w_074_1558, w_074_1560, w_074_1561, w_074_1562, w_074_1563, w_074_1567, w_074_1569, w_074_1572, w_074_1573, w_074_1574, w_074_1575, w_074_1577, w_074_1580, w_074_1581, w_074_1583, w_074_1584, w_074_1585, w_074_1586, w_074_1587, w_074_1589, w_074_1592, w_074_1593, w_074_1594, w_074_1596, w_074_1598, w_074_1601, w_074_1603, w_074_1604, w_074_1605, w_074_1606, w_074_1607, w_074_1608, w_074_1609, w_074_1610, w_074_1611, w_074_1612, w_074_1614, w_074_1616, w_074_1617, w_074_1618, w_074_1619, w_074_1621, w_074_1622, w_074_1625, w_074_1626, w_074_1627, w_074_1632, w_074_1633, w_074_1634, w_074_1636, w_074_1637, w_074_1638, w_074_1639, w_074_1640, w_074_1644, w_074_1647, w_074_1649, w_074_1650, w_074_1651, w_074_1653, w_074_1654, w_074_1656, w_074_1657, w_074_1659, w_074_1660, w_074_1663, w_074_1664, w_074_1665, w_074_1666, w_074_1667, w_074_1668, w_074_1669, w_074_1671, w_074_1672, w_074_1673, w_074_1677, w_074_1679, w_074_1680, w_074_1681, w_074_1682, w_074_1685, w_074_1687, w_074_1688, w_074_1694, w_074_1696, w_074_1697, w_074_1699, w_074_1701, w_074_1702, w_074_1703, w_074_1705, w_074_1708, w_074_1709, w_074_1710, w_074_1711, w_074_1712, w_074_1713, w_074_1714, w_074_1717, w_074_1718, w_074_1721, w_074_1722, w_074_1723, w_074_1724, w_074_1725, w_074_1728, w_074_1729, w_074_1731, w_074_1732, w_074_1733, w_074_1737, w_074_1739, w_074_1740, w_074_1741, w_074_1742, w_074_1743, w_074_1745, w_074_1746, w_074_1747, w_074_1748, w_074_1749, w_074_1751, w_074_1752, w_074_1754, w_074_1757, w_074_1761, w_074_1762, w_074_1763, w_074_1766, w_074_1768, w_074_1769, w_074_1770, w_074_1771, w_074_1772, w_074_1774, w_074_1777, w_074_1778, w_074_1780, w_074_1781, w_074_1785, w_074_1787, w_074_1788, w_074_1790, w_074_1791, w_074_1792, w_074_1793, w_074_1795, w_074_1797, w_074_1799, w_074_1800, w_074_1801, w_074_1802, w_074_1806, w_074_1807, w_074_1808, w_074_1810, w_074_1811, w_074_1812, w_074_1813, w_074_1815, w_074_1816, w_074_1817, w_074_1819, w_074_1820, w_074_1824, w_074_1826, w_074_1830, w_074_1831, w_074_1833, w_074_1834, w_074_1837, w_074_1838, w_074_1839, w_074_1840, w_074_1843, w_074_1845, w_074_1846, w_074_1847, w_074_1848, w_074_1850, w_074_1851, w_074_1852, w_074_1853, w_074_1855, w_074_1856, w_074_1857, w_074_1863, w_074_1864, w_074_1865, w_074_1866, w_074_1867, w_074_1868, w_074_1869, w_074_1870, w_074_1871, w_074_1872, w_074_1875, w_074_1878, w_074_1879, w_074_1880, w_074_1881, w_074_1882, w_074_1883, w_074_1884, w_074_1885, w_074_1886, w_074_1887, w_074_1892, w_074_1893, w_074_1895, w_074_1897, w_074_1901, w_074_1902, w_074_1904, w_074_1905, w_074_1910, w_074_1915, w_074_1916, w_074_1917, w_074_1918, w_074_1920, w_074_1921, w_074_1923, w_074_1926, w_074_1927, w_074_1928, w_074_1930, w_074_1931, w_074_1932, w_074_1938, w_074_1943, w_074_1944, w_074_1945, w_074_1947, w_074_1950;
  wire w_075_000, w_075_001, w_075_002, w_075_003, w_075_004, w_075_005, w_075_006, w_075_007, w_075_008, w_075_009, w_075_010, w_075_011, w_075_012, w_075_013, w_075_014, w_075_015, w_075_016, w_075_017, w_075_018, w_075_019, w_075_020, w_075_021, w_075_022, w_075_023, w_075_024, w_075_025, w_075_026, w_075_027, w_075_028, w_075_029, w_075_030, w_075_031, w_075_032, w_075_033, w_075_034, w_075_035, w_075_036, w_075_037, w_075_038, w_075_039, w_075_040, w_075_041, w_075_042, w_075_043, w_075_044, w_075_045, w_075_046, w_075_047, w_075_048, w_075_049, w_075_050, w_075_051, w_075_052, w_075_053, w_075_054, w_075_055, w_075_056, w_075_057, w_075_058, w_075_059, w_075_060, w_075_061, w_075_062, w_075_063, w_075_064, w_075_065, w_075_066, w_075_067, w_075_068, w_075_069, w_075_070, w_075_071, w_075_072, w_075_073, w_075_074, w_075_075, w_075_076, w_075_077, w_075_078, w_075_079, w_075_080, w_075_081, w_075_082, w_075_083, w_075_084, w_075_085, w_075_086, w_075_087, w_075_088, w_075_089, w_075_090, w_075_091, w_075_092, w_075_093, w_075_094, w_075_095, w_075_096, w_075_097, w_075_098, w_075_099, w_075_100, w_075_101, w_075_102, w_075_103, w_075_104, w_075_105, w_075_106, w_075_107, w_075_108, w_075_109, w_075_110, w_075_111, w_075_112, w_075_113, w_075_114, w_075_115, w_075_116, w_075_117, w_075_118, w_075_119, w_075_120, w_075_121, w_075_122, w_075_123, w_075_124, w_075_125, w_075_126, w_075_127, w_075_128, w_075_129, w_075_130, w_075_131, w_075_132, w_075_133, w_075_134, w_075_135, w_075_136, w_075_137, w_075_138, w_075_139, w_075_140, w_075_141, w_075_142, w_075_143, w_075_144, w_075_145, w_075_146, w_075_147, w_075_148, w_075_149, w_075_150, w_075_151, w_075_152, w_075_153, w_075_154, w_075_155, w_075_156, w_075_157, w_075_158, w_075_159, w_075_160, w_075_161, w_075_162, w_075_163, w_075_164, w_075_165, w_075_166, w_075_167, w_075_168, w_075_169, w_075_170, w_075_171, w_075_172, w_075_173, w_075_174, w_075_175, w_075_176, w_075_177, w_075_178, w_075_179, w_075_180, w_075_181, w_075_182, w_075_183, w_075_184, w_075_185, w_075_186, w_075_187, w_075_188, w_075_189, w_075_190, w_075_191, w_075_192, w_075_193, w_075_194, w_075_195, w_075_196, w_075_197, w_075_198, w_075_199, w_075_200, w_075_201, w_075_202, w_075_203, w_075_204, w_075_205, w_075_206, w_075_207, w_075_208, w_075_209, w_075_210, w_075_211, w_075_212, w_075_213, w_075_214, w_075_215, w_075_216, w_075_217, w_075_218, w_075_219, w_075_220, w_075_221, w_075_222, w_075_223, w_075_224, w_075_225, w_075_226, w_075_227, w_075_228, w_075_229, w_075_230, w_075_231, w_075_232, w_075_233, w_075_234, w_075_235, w_075_236, w_075_237, w_075_238, w_075_239, w_075_240, w_075_241, w_075_242, w_075_243, w_075_244, w_075_245, w_075_246, w_075_247, w_075_248, w_075_249, w_075_250, w_075_251, w_075_252, w_075_253, w_075_254, w_075_255, w_075_256, w_075_257, w_075_258, w_075_259, w_075_260, w_075_261, w_075_262, w_075_263, w_075_264, w_075_265, w_075_266, w_075_267, w_075_268, w_075_269, w_075_270, w_075_271, w_075_272, w_075_273, w_075_274, w_075_275, w_075_276, w_075_277, w_075_278, w_075_279, w_075_280, w_075_281, w_075_282, w_075_283, w_075_284, w_075_285, w_075_286;
  wire w_076_000, w_076_001, w_076_002, w_076_003, w_076_004, w_076_005, w_076_006, w_076_007, w_076_008, w_076_009, w_076_010, w_076_011, w_076_012, w_076_013, w_076_014, w_076_015, w_076_016, w_076_017, w_076_018, w_076_019, w_076_020, w_076_021, w_076_022, w_076_023, w_076_024, w_076_025, w_076_026, w_076_027, w_076_029, w_076_031, w_076_032, w_076_033, w_076_034, w_076_035, w_076_036, w_076_037, w_076_038, w_076_039, w_076_040, w_076_041, w_076_042, w_076_043, w_076_044, w_076_045, w_076_046, w_076_047, w_076_048, w_076_049, w_076_050, w_076_051, w_076_052, w_076_053, w_076_054, w_076_055, w_076_057, w_076_058, w_076_059, w_076_060, w_076_061, w_076_062, w_076_063, w_076_064, w_076_065, w_076_066, w_076_067, w_076_068, w_076_069, w_076_070, w_076_071, w_076_072, w_076_073, w_076_074, w_076_075, w_076_076, w_076_077, w_076_078, w_076_079, w_076_080, w_076_081, w_076_082, w_076_083, w_076_084, w_076_085, w_076_086, w_076_087, w_076_088, w_076_089, w_076_090, w_076_091, w_076_092, w_076_093, w_076_094, w_076_095, w_076_096, w_076_097, w_076_098, w_076_099, w_076_100, w_076_101, w_076_102, w_076_103, w_076_104, w_076_105, w_076_106, w_076_107, w_076_108, w_076_109, w_076_110, w_076_111, w_076_112, w_076_113, w_076_114, w_076_115, w_076_116, w_076_117, w_076_118, w_076_119, w_076_120, w_076_121, w_076_122, w_076_123, w_076_124, w_076_125, w_076_126, w_076_127, w_076_128, w_076_129, w_076_130, w_076_131, w_076_132, w_076_133, w_076_134, w_076_135, w_076_136, w_076_137, w_076_138, w_076_139, w_076_140, w_076_141, w_076_142, w_076_143, w_076_144, w_076_147, w_076_148, w_076_149, w_076_150, w_076_151, w_076_152, w_076_153, w_076_154, w_076_155, w_076_156, w_076_157, w_076_158, w_076_159, w_076_160, w_076_161, w_076_162, w_076_163, w_076_164, w_076_165, w_076_166, w_076_167, w_076_168, w_076_169, w_076_170, w_076_171, w_076_172, w_076_173, w_076_174, w_076_175, w_076_176, w_076_177, w_076_178, w_076_179, w_076_180, w_076_181, w_076_182, w_076_183, w_076_185, w_076_186, w_076_187, w_076_188, w_076_189, w_076_190, w_076_191, w_076_192, w_076_194, w_076_195, w_076_196, w_076_197, w_076_198, w_076_199, w_076_200, w_076_201, w_076_202, w_076_203, w_076_204, w_076_205, w_076_206, w_076_207, w_076_208, w_076_209, w_076_210, w_076_211, w_076_212, w_076_213, w_076_214, w_076_215, w_076_216, w_076_217, w_076_218, w_076_219, w_076_220, w_076_221, w_076_222, w_076_223, w_076_224, w_076_225, w_076_226, w_076_227, w_076_228, w_076_229, w_076_230, w_076_231, w_076_232, w_076_233, w_076_234, w_076_235, w_076_236, w_076_237, w_076_238, w_076_239, w_076_240, w_076_241, w_076_242, w_076_243, w_076_244, w_076_245, w_076_246, w_076_247, w_076_248, w_076_249, w_076_250, w_076_251, w_076_252, w_076_253, w_076_254, w_076_255, w_076_256, w_076_257, w_076_258, w_076_259, w_076_260, w_076_261, w_076_262, w_076_263, w_076_265, w_076_266, w_076_267, w_076_268, w_076_270, w_076_271, w_076_272, w_076_273, w_076_274, w_076_275, w_076_276, w_076_277, w_076_278, w_076_279, w_076_280, w_076_281, w_076_282, w_076_284, w_076_285, w_076_286, w_076_287, w_076_288, w_076_289, w_076_290, w_076_291, w_076_292, w_076_293, w_076_294, w_076_295, w_076_296, w_076_297, w_076_298, w_076_299, w_076_300, w_076_301, w_076_302, w_076_303, w_076_304, w_076_305, w_076_306, w_076_307, w_076_308, w_076_309, w_076_310, w_076_311, w_076_312, w_076_314, w_076_315, w_076_316, w_076_317, w_076_318, w_076_319, w_076_320, w_076_321, w_076_322, w_076_323, w_076_324, w_076_325, w_076_326, w_076_327, w_076_328, w_076_329, w_076_330, w_076_331, w_076_332, w_076_333, w_076_334, w_076_335, w_076_336, w_076_337, w_076_338, w_076_339, w_076_340, w_076_341, w_076_342, w_076_343, w_076_344, w_076_345, w_076_346, w_076_347, w_076_348, w_076_349, w_076_350, w_076_351, w_076_352, w_076_353, w_076_354, w_076_355, w_076_356, w_076_357, w_076_358, w_076_359, w_076_360, w_076_361, w_076_362, w_076_363, w_076_364, w_076_365, w_076_366, w_076_367, w_076_368, w_076_369, w_076_370, w_076_371, w_076_372, w_076_373, w_076_374, w_076_375, w_076_376, w_076_377, w_076_378, w_076_379, w_076_380, w_076_381, w_076_382, w_076_383, w_076_384, w_076_385, w_076_386, w_076_387, w_076_388, w_076_389, w_076_390, w_076_391, w_076_392, w_076_393, w_076_394, w_076_395, w_076_396, w_076_397, w_076_399, w_076_400, w_076_401, w_076_402, w_076_403, w_076_404, w_076_405, w_076_406, w_076_407, w_076_408, w_076_409, w_076_410, w_076_411, w_076_412, w_076_413, w_076_414, w_076_415, w_076_416, w_076_417, w_076_418, w_076_419, w_076_420, w_076_421, w_076_422, w_076_423, w_076_424, w_076_425, w_076_426, w_076_427, w_076_428, w_076_429, w_076_430, w_076_431, w_076_432, w_076_433, w_076_435, w_076_436, w_076_437, w_076_438, w_076_439, w_076_440, w_076_441, w_076_442, w_076_443, w_076_444, w_076_445, w_076_446, w_076_447, w_076_448, w_076_449, w_076_450, w_076_451, w_076_452, w_076_454, w_076_455, w_076_456, w_076_457, w_076_458, w_076_459, w_076_460, w_076_461, w_076_462, w_076_463, w_076_464, w_076_465, w_076_466, w_076_467, w_076_468, w_076_469, w_076_470, w_076_471, w_076_472, w_076_473, w_076_474, w_076_475, w_076_476, w_076_477, w_076_478, w_076_479, w_076_480, w_076_481, w_076_482, w_076_483, w_076_484, w_076_485, w_076_487, w_076_488, w_076_489, w_076_491, w_076_492, w_076_493, w_076_494, w_076_495, w_076_496, w_076_497, w_076_498, w_076_499, w_076_500, w_076_501, w_076_502, w_076_503, w_076_504, w_076_505, w_076_506, w_076_507, w_076_508, w_076_509, w_076_510, w_076_511, w_076_512, w_076_513, w_076_514, w_076_515, w_076_516, w_076_517, w_076_518, w_076_519, w_076_520, w_076_521, w_076_522, w_076_523, w_076_524, w_076_525, w_076_526, w_076_527, w_076_528, w_076_529, w_076_530, w_076_531, w_076_532, w_076_534, w_076_535, w_076_536, w_076_537, w_076_538, w_076_539, w_076_540, w_076_541, w_076_542, w_076_543, w_076_544, w_076_545, w_076_546, w_076_547, w_076_548, w_076_549, w_076_550, w_076_551, w_076_552, w_076_553, w_076_554, w_076_555, w_076_556, w_076_557, w_076_558, w_076_559, w_076_560, w_076_561, w_076_562, w_076_563, w_076_564, w_076_565, w_076_566, w_076_568, w_076_570, w_076_571, w_076_572, w_076_574, w_076_575, w_076_576, w_076_577, w_076_578, w_076_579, w_076_580, w_076_581, w_076_582, w_076_583, w_076_584, w_076_585, w_076_586, w_076_587, w_076_588, w_076_589, w_076_590, w_076_591, w_076_592, w_076_593, w_076_594, w_076_595, w_076_596, w_076_597, w_076_598, w_076_599, w_076_601, w_076_602, w_076_603, w_076_604, w_076_605, w_076_606, w_076_607, w_076_608, w_076_609, w_076_611, w_076_612, w_076_613, w_076_616, w_076_617, w_076_618, w_076_619, w_076_620, w_076_621, w_076_622, w_076_623, w_076_624, w_076_625, w_076_626, w_076_627, w_076_628, w_076_629, w_076_631, w_076_632, w_076_633;
  wire w_077_000, w_077_002, w_077_003, w_077_005, w_077_009, w_077_011, w_077_012, w_077_014, w_077_017, w_077_018, w_077_019, w_077_022, w_077_023, w_077_025, w_077_027, w_077_028, w_077_029, w_077_031, w_077_032, w_077_034, w_077_035, w_077_038, w_077_040, w_077_041, w_077_042, w_077_045, w_077_050, w_077_051, w_077_052, w_077_053, w_077_058, w_077_059, w_077_062, w_077_066, w_077_067, w_077_068, w_077_071, w_077_072, w_077_074, w_077_075, w_077_077, w_077_078, w_077_079, w_077_080, w_077_081, w_077_083, w_077_085, w_077_087, w_077_090, w_077_092, w_077_094, w_077_095, w_077_097, w_077_100, w_077_101, w_077_103, w_077_105, w_077_107, w_077_109, w_077_111, w_077_112, w_077_114, w_077_115, w_077_116, w_077_117, w_077_118, w_077_119, w_077_120, w_077_123, w_077_124, w_077_125, w_077_126, w_077_127, w_077_128, w_077_129, w_077_130, w_077_132, w_077_134, w_077_136, w_077_137, w_077_138, w_077_139, w_077_141, w_077_145, w_077_149, w_077_153, w_077_155, w_077_160, w_077_162, w_077_163, w_077_164, w_077_165, w_077_167, w_077_171, w_077_174, w_077_176, w_077_177, w_077_178, w_077_180, w_077_182, w_077_185, w_077_187, w_077_188, w_077_190, w_077_192, w_077_194, w_077_197, w_077_203, w_077_204, w_077_206, w_077_208, w_077_211, w_077_212, w_077_214, w_077_216, w_077_220, w_077_223, w_077_224, w_077_225, w_077_226, w_077_227, w_077_228, w_077_229, w_077_232, w_077_233, w_077_236, w_077_237, w_077_238, w_077_241, w_077_242, w_077_244, w_077_245, w_077_246, w_077_249, w_077_250, w_077_251, w_077_252, w_077_254, w_077_255, w_077_256, w_077_258, w_077_260, w_077_263, w_077_264, w_077_270, w_077_271, w_077_273, w_077_274, w_077_275, w_077_277, w_077_279, w_077_280, w_077_281, w_077_283, w_077_284, w_077_289, w_077_290, w_077_292, w_077_294, w_077_296, w_077_299, w_077_301, w_077_304, w_077_306, w_077_309, w_077_311, w_077_312, w_077_313, w_077_314, w_077_316, w_077_317, w_077_319, w_077_321, w_077_322, w_077_323, w_077_324, w_077_325, w_077_326, w_077_327, w_077_328, w_077_329, w_077_330, w_077_335, w_077_336, w_077_337, w_077_338, w_077_339, w_077_341, w_077_343, w_077_345, w_077_346, w_077_347, w_077_348, w_077_352, w_077_354, w_077_355, w_077_359, w_077_361, w_077_365, w_077_372, w_077_374, w_077_375, w_077_378, w_077_381, w_077_385, w_077_387, w_077_389, w_077_391, w_077_394, w_077_395, w_077_401, w_077_403, w_077_404, w_077_405, w_077_406, w_077_407, w_077_411, w_077_412, w_077_414, w_077_415, w_077_416, w_077_417, w_077_418, w_077_419, w_077_421, w_077_422, w_077_423, w_077_425, w_077_426, w_077_428, w_077_429, w_077_432, w_077_433, w_077_438, w_077_439, w_077_441, w_077_442, w_077_444, w_077_446, w_077_450, w_077_452, w_077_453, w_077_454, w_077_455, w_077_456, w_077_464, w_077_465, w_077_466, w_077_467, w_077_468, w_077_471, w_077_475, w_077_476, w_077_477, w_077_478, w_077_479, w_077_480, w_077_483, w_077_485, w_077_488, w_077_489, w_077_492, w_077_493, w_077_494, w_077_496, w_077_497, w_077_499, w_077_501, w_077_503, w_077_505, w_077_507, w_077_512, w_077_513, w_077_514, w_077_515, w_077_516, w_077_517, w_077_518, w_077_519, w_077_520, w_077_521, w_077_522, w_077_523, w_077_524, w_077_525, w_077_526, w_077_527, w_077_529, w_077_531, w_077_532, w_077_533, w_077_537, w_077_538, w_077_539, w_077_540, w_077_544, w_077_546, w_077_551, w_077_552, w_077_553, w_077_554, w_077_555, w_077_556, w_077_559, w_077_560, w_077_562, w_077_563, w_077_566, w_077_567, w_077_568, w_077_569, w_077_570, w_077_571, w_077_572, w_077_573, w_077_577, w_077_579, w_077_582, w_077_583, w_077_584, w_077_586, w_077_587, w_077_589, w_077_590, w_077_591, w_077_592, w_077_593, w_077_594, w_077_595, w_077_596, w_077_597, w_077_598, w_077_603, w_077_604, w_077_605, w_077_607, w_077_609, w_077_610, w_077_612, w_077_613, w_077_614, w_077_615, w_077_617, w_077_618, w_077_619, w_077_620, w_077_624, w_077_626, w_077_627, w_077_628, w_077_629, w_077_630, w_077_631, w_077_632, w_077_633, w_077_634, w_077_635, w_077_636, w_077_637, w_077_638, w_077_640, w_077_641, w_077_642, w_077_643, w_077_644, w_077_645, w_077_646, w_077_647, w_077_648, w_077_649, w_077_650, w_077_651, w_077_652, w_077_653, w_077_654, w_077_655, w_077_656, w_077_657, w_077_660, w_077_661, w_077_662, w_077_663, w_077_664, w_077_665, w_077_666, w_077_668, w_077_670, w_077_673, w_077_675, w_077_677, w_077_678, w_077_679, w_077_683, w_077_684, w_077_685, w_077_687, w_077_688, w_077_690, w_077_693, w_077_694, w_077_697, w_077_699, w_077_700, w_077_705, w_077_707, w_077_708, w_077_709, w_077_712, w_077_714, w_077_716, w_077_718, w_077_719, w_077_720, w_077_721, w_077_723, w_077_725, w_077_726, w_077_727, w_077_729, w_077_732, w_077_733, w_077_735, w_077_741, w_077_742, w_077_743, w_077_745, w_077_746, w_077_747, w_077_750, w_077_751, w_077_752, w_077_753, w_077_756, w_077_757, w_077_759, w_077_760, w_077_761, w_077_762, w_077_763, w_077_764, w_077_765, w_077_766, w_077_768, w_077_769, w_077_772, w_077_773, w_077_775, w_077_779, w_077_780, w_077_784, w_077_788, w_077_789, w_077_790, w_077_792, w_077_793, w_077_796, w_077_797, w_077_800, w_077_802, w_077_805, w_077_807, w_077_808, w_077_810, w_077_812, w_077_815, w_077_816, w_077_817, w_077_823, w_077_826, w_077_827, w_077_828, w_077_829, w_077_831, w_077_835, w_077_839, w_077_841, w_077_843, w_077_847, w_077_848, w_077_849, w_077_851, w_077_852, w_077_854, w_077_856, w_077_859, w_077_861, w_077_862, w_077_863, w_077_864, w_077_865, w_077_866, w_077_870, w_077_873, w_077_874, w_077_875, w_077_877, w_077_878, w_077_880, w_077_881, w_077_882, w_077_884, w_077_885, w_077_887, w_077_888, w_077_889, w_077_890, w_077_892, w_077_893, w_077_895, w_077_896, w_077_897, w_077_901, w_077_902, w_077_903, w_077_904, w_077_905, w_077_906, w_077_907, w_077_909, w_077_910, w_077_913, w_077_914, w_077_915, w_077_920, w_077_921, w_077_927, w_077_928, w_077_930, w_077_931, w_077_934, w_077_935, w_077_936, w_077_940, w_077_941, w_077_943, w_077_945, w_077_946, w_077_947, w_077_951, w_077_953, w_077_956, w_077_957, w_077_958, w_077_960, w_077_961, w_077_964, w_077_965, w_077_967, w_077_968, w_077_969, w_077_971, w_077_972, w_077_974, w_077_976, w_077_977, w_077_978, w_077_979, w_077_981, w_077_983, w_077_984, w_077_986, w_077_989, w_077_991, w_077_993, w_077_994, w_077_995, w_077_999, w_077_1002, w_077_1006, w_077_1008, w_077_1009, w_077_1010, w_077_1012, w_077_1013, w_077_1014, w_077_1015, w_077_1016, w_077_1018, w_077_1019, w_077_1020, w_077_1021, w_077_1022, w_077_1023, w_077_1024, w_077_1025, w_077_1030, w_077_1031, w_077_1032, w_077_1033, w_077_1034, w_077_1035, w_077_1037, w_077_1040, w_077_1043, w_077_1044, w_077_1045, w_077_1048, w_077_1049, w_077_1052, w_077_1054, w_077_1057, w_077_1061, w_077_1063, w_077_1064, w_077_1065, w_077_1066, w_077_1067, w_077_1068, w_077_1070, w_077_1071, w_077_1072, w_077_1074, w_077_1077, w_077_1078, w_077_1079, w_077_1080, w_077_1082, w_077_1083, w_077_1084, w_077_1085, w_077_1087, w_077_1088, w_077_1089, w_077_1092, w_077_1095, w_077_1096, w_077_1097, w_077_1100, w_077_1101, w_077_1102, w_077_1105, w_077_1108, w_077_1109, w_077_1117, w_077_1118, w_077_1120, w_077_1121, w_077_1122, w_077_1123, w_077_1124, w_077_1125, w_077_1127, w_077_1129, w_077_1130, w_077_1131, w_077_1135, w_077_1136, w_077_1139, w_077_1141, w_077_1142, w_077_1143, w_077_1145, w_077_1147, w_077_1149, w_077_1150, w_077_1152, w_077_1155, w_077_1156, w_077_1158, w_077_1163, w_077_1164, w_077_1167, w_077_1168, w_077_1169, w_077_1170, w_077_1172, w_077_1176, w_077_1177, w_077_1178, w_077_1180, w_077_1183, w_077_1186, w_077_1188, w_077_1189, w_077_1191, w_077_1192, w_077_1194, w_077_1196, w_077_1204, w_077_1208, w_077_1210, w_077_1212, w_077_1213, w_077_1216, w_077_1219, w_077_1220, w_077_1223, w_077_1228, w_077_1231, w_077_1232, w_077_1235, w_077_1237, w_077_1238, w_077_1239, w_077_1242, w_077_1244, w_077_1245, w_077_1246, w_077_1247, w_077_1248, w_077_1251, w_077_1252, w_077_1255, w_077_1257, w_077_1258, w_077_1261, w_077_1263, w_077_1264, w_077_1266, w_077_1268, w_077_1270, w_077_1272, w_077_1274, w_077_1276, w_077_1279, w_077_1280, w_077_1281, w_077_1282, w_077_1283, w_077_1284, w_077_1285, w_077_1286, w_077_1287, w_077_1288, w_077_1289, w_077_1290, w_077_1291, w_077_1292, w_077_1294, w_077_1295, w_077_1296, w_077_1298, w_077_1299, w_077_1301, w_077_1303, w_077_1304, w_077_1305, w_077_1306, w_077_1307, w_077_1308, w_077_1309, w_077_1312, w_077_1315, w_077_1316, w_077_1317, w_077_1318, w_077_1319, w_077_1320, w_077_1321, w_077_1322, w_077_1324, w_077_1327, w_077_1328, w_077_1330, w_077_1331, w_077_1332, w_077_1335, w_077_1338, w_077_1340, w_077_1341, w_077_1343, w_077_1344, w_077_1345, w_077_1347, w_077_1348, w_077_1351, w_077_1353, w_077_1355, w_077_1356, w_077_1357, w_077_1359, w_077_1360, w_077_1362, w_077_1365, w_077_1366, w_077_1367, w_077_1369, w_077_1374, w_077_1375, w_077_1377, w_077_1378, w_077_1381, w_077_1382, w_077_1383, w_077_1384, w_077_1388, w_077_1389, w_077_1391, w_077_1392, w_077_1394, w_077_1396, w_077_1397, w_077_1399, w_077_1401, w_077_1402, w_077_1404, w_077_1405, w_077_1406, w_077_1409, w_077_1411, w_077_1414, w_077_1415, w_077_1417, w_077_1419, w_077_1421, w_077_1422, w_077_1424, w_077_1425, w_077_1431, w_077_1433, w_077_1435, w_077_1439, w_077_1440, w_077_1445, w_077_1447, w_077_1448, w_077_1449, w_077_1452, w_077_1454, w_077_1455, w_077_1456, w_077_1459, w_077_1460, w_077_1462, w_077_1463, w_077_1464, w_077_1467, w_077_1468, w_077_1472, w_077_1475, w_077_1476, w_077_1477, w_077_1480, w_077_1484, w_077_1487, w_077_1490, w_077_1492, w_077_1493, w_077_1497, w_077_1498, w_077_1499, w_077_1500, w_077_1504, w_077_1505, w_077_1506, w_077_1507, w_077_1509, w_077_1512, w_077_1514, w_077_1516, w_077_1517, w_077_1518, w_077_1519, w_077_1520, w_077_1521, w_077_1522, w_077_1527, w_077_1528, w_077_1529, w_077_1530, w_077_1532, w_077_1533, w_077_1534, w_077_1537, w_077_1538, w_077_1542, w_077_1543, w_077_1544, w_077_1546, w_077_1548, w_077_1550, w_077_1553, w_077_1554, w_077_1556, w_077_1558, w_077_1559, w_077_1560, w_077_1563, w_077_1568, w_077_1570, w_077_1571, w_077_1573, w_077_1574, w_077_1575, w_077_1576, w_077_1577, w_077_1578, w_077_1581, w_077_1582, w_077_1583, w_077_1585, w_077_1586, w_077_1587, w_077_1588, w_077_1591, w_077_1597, w_077_1600, w_077_1608, w_077_1610, w_077_1613, w_077_1615, w_077_1616, w_077_1617, w_077_1618, w_077_1621, w_077_1623, w_077_1624, w_077_1626, w_077_1627, w_077_1628, w_077_1629, w_077_1631, w_077_1632, w_077_1633, w_077_1635, w_077_1636, w_077_1638, w_077_1639, w_077_1640, w_077_1643, w_077_1645, w_077_1647, w_077_1650, w_077_1651, w_077_1652, w_077_1653, w_077_1655, w_077_1656, w_077_1658, w_077_1659, w_077_1661, w_077_1663, w_077_1664, w_077_1666, w_077_1667, w_077_1668, w_077_1669, w_077_1671, w_077_1672, w_077_1673, w_077_1675, w_077_1677, w_077_1678, w_077_1680, w_077_1681, w_077_1685, w_077_1686, w_077_1687, w_077_1688, w_077_1690, w_077_1691, w_077_1694, w_077_1695, w_077_1696, w_077_1697, w_077_1698, w_077_1699, w_077_1700, w_077_1701, w_077_1702, w_077_1703, w_077_1707, w_077_1708, w_077_1712, w_077_1713, w_077_1716, w_077_1718, w_077_1720, w_077_1721, w_077_1723, w_077_1724, w_077_1725, w_077_1726, w_077_1728, w_077_1730, w_077_1731, w_077_1732, w_077_1733, w_077_1734, w_077_1735, w_077_1736, w_077_1737, w_077_1738, w_077_1739, w_077_1740, w_077_1741, w_077_1742, w_077_1743, w_077_1744, w_077_1745, w_077_1748, w_077_1749, w_077_1751, w_077_1753, w_077_1756, w_077_1758, w_077_1760, w_077_1761, w_077_1763, w_077_1765, w_077_1768, w_077_1770, w_077_1772, w_077_1775, w_077_1779, w_077_1782, w_077_1784, w_077_1785, w_077_1786, w_077_1788, w_077_1789, w_077_1792, w_077_1793, w_077_1794, w_077_1795, w_077_1796, w_077_1799, w_077_1801, w_077_1802, w_077_1803, w_077_1804, w_077_1806, w_077_1807, w_077_1808, w_077_1809, w_077_1810, w_077_1812, w_077_1813, w_077_1814, w_077_1815, w_077_1816, w_077_1817, w_077_1819, w_077_1820, w_077_1824, w_077_1825, w_077_1826, w_077_1829, w_077_1830, w_077_1832, w_077_1834, w_077_1835, w_077_1836, w_077_1844, w_077_1847, w_077_1849, w_077_1852, w_077_1857, w_077_1859, w_077_1861, w_077_1862, w_077_1865, w_077_1871, w_077_1873, w_077_1875, w_077_1876, w_077_1886, w_077_1888, w_077_1890, w_077_1893, w_077_1898, w_077_1899, w_077_1900, w_077_1904, w_077_1905, w_077_1906, w_077_1907, w_077_1908, w_077_1909, w_077_1910, w_077_1912, w_077_1913, w_077_1915, w_077_1918, w_077_1920, w_077_1923, w_077_1924, w_077_1927, w_077_1933, w_077_1939, w_077_1944, w_077_1947, w_077_1949, w_077_1951, w_077_1952, w_077_1956, w_077_1959, w_077_1960, w_077_1961, w_077_1962, w_077_1966, w_077_1969, w_077_1970, w_077_1972, w_077_1979, w_077_1981, w_077_1984, w_077_1987, w_077_1992, w_077_1995, w_077_1997, w_077_1998, w_077_2000, w_077_2004, w_077_2005, w_077_2007, w_077_2010, w_077_2011, w_077_2012, w_077_2014, w_077_2017, w_077_2019, w_077_2026, w_077_2027, w_077_2029, w_077_2033, w_077_2038, w_077_2041, w_077_2043, w_077_2044, w_077_2045, w_077_2047, w_077_2049, w_077_2054, w_077_2060, w_077_2061, w_077_2064, w_077_2065, w_077_2067, w_077_2068, w_077_2070, w_077_2075, w_077_2080, w_077_2081, w_077_2085, w_077_2086, w_077_2095, w_077_2100, w_077_2101, w_077_2102, w_077_2107, w_077_2109, w_077_2112, w_077_2119, w_077_2121, w_077_2122, w_077_2125, w_077_2126, w_077_2127, w_077_2129, w_077_2134, w_077_2135, w_077_2143, w_077_2147, w_077_2151, w_077_2152, w_077_2157, w_077_2158, w_077_2159, w_077_2161, w_077_2163, w_077_2170, w_077_2171, w_077_2173, w_077_2175, w_077_2179, w_077_2182, w_077_2183, w_077_2185, w_077_2189, w_077_2191, w_077_2192, w_077_2195, w_077_2196, w_077_2198, w_077_2203, w_077_2205, w_077_2209, w_077_2210, w_077_2213, w_077_2216, w_077_2225, w_077_2228, w_077_2231, w_077_2237, w_077_2239, w_077_2243, w_077_2253, w_077_2254, w_077_2259, w_077_2262, w_077_2270, w_077_2273, w_077_2275, w_077_2277, w_077_2284, w_077_2291, w_077_2299, w_077_2302, w_077_2305, w_077_2309, w_077_2312, w_077_2316, w_077_2317, w_077_2318, w_077_2320, w_077_2321, w_077_2326, w_077_2327, w_077_2330, w_077_2334, w_077_2335, w_077_2346, w_077_2347, w_077_2351, w_077_2352, w_077_2358, w_077_2361, w_077_2362, w_077_2368, w_077_2369, w_077_2371, w_077_2372, w_077_2373, w_077_2380, w_077_2382, w_077_2385, w_077_2389, w_077_2390, w_077_2395, w_077_2396, w_077_2398, w_077_2400, w_077_2401, w_077_2402, w_077_2406, w_077_2410, w_077_2411, w_077_2416, w_077_2419, w_077_2420, w_077_2429, w_077_2431, w_077_2432, w_077_2433, w_077_2435, w_077_2436, w_077_2438, w_077_2439, w_077_2440, w_077_2444, w_077_2447, w_077_2448, w_077_2450, w_077_2455, w_077_2456, w_077_2457, w_077_2458, w_077_2459, w_077_2463, w_077_2467, w_077_2468, w_077_2470, w_077_2475, w_077_2476, w_077_2482, w_077_2487, w_077_2489, w_077_2494, w_077_2496, w_077_2497, w_077_2500, w_077_2506, w_077_2508, w_077_2513, w_077_2514, w_077_2515, w_077_2516, w_077_2517, w_077_2519, w_077_2527, w_077_2528, w_077_2530, w_077_2532, w_077_2537, w_077_2538, w_077_2543, w_077_2545, w_077_2547, w_077_2548, w_077_2555, w_077_2558, w_077_2563, w_077_2570, w_077_2571, w_077_2573, w_077_2575, w_077_2579, w_077_2581, w_077_2589, w_077_2593, w_077_2594, w_077_2596, w_077_2597, w_077_2602, w_077_2604, w_077_2605, w_077_2608, w_077_2609, w_077_2610, w_077_2614, w_077_2618, w_077_2619, w_077_2625, w_077_2627, w_077_2635, w_077_2643, w_077_2644, w_077_2651, w_077_2653, w_077_2655, w_077_2658, w_077_2659, w_077_2665, w_077_2678, w_077_2679, w_077_2681, w_077_2682, w_077_2683, w_077_2686, w_077_2688, w_077_2689, w_077_2691, w_077_2693, w_077_2698, w_077_2700, w_077_2701, w_077_2702, w_077_2704, w_077_2710, w_077_2711, w_077_2714, w_077_2715, w_077_2716, w_077_2719, w_077_2724, w_077_2726, w_077_2728, w_077_2730, w_077_2734, w_077_2737, w_077_2743, w_077_2745, w_077_2751, w_077_2756, w_077_2758, w_077_2759, w_077_2764, w_077_2765, w_077_2769, w_077_2770, w_077_2775, w_077_2778, w_077_2779, w_077_2781, w_077_2786, w_077_2794, w_077_2796, w_077_2797, w_077_2798, w_077_2799, w_077_2801, w_077_2804, w_077_2805, w_077_2819, w_077_2821, w_077_2825, w_077_2828, w_077_2831, w_077_2834, w_077_2835, w_077_2838, w_077_2842, w_077_2844, w_077_2846, w_077_2848, w_077_2854, w_077_2856, w_077_2858, w_077_2859, w_077_2862, w_077_2874, w_077_2877, w_077_2878, w_077_2881, w_077_2883, w_077_2884, w_077_2889, w_077_2891, w_077_2892, w_077_2893, w_077_2898, w_077_2902, w_077_2904, w_077_2905, w_077_2913, w_077_2914, w_077_2916, w_077_2924, w_077_2929, w_077_2931, w_077_2933, w_077_2937, w_077_2940, w_077_2947, w_077_2948, w_077_2949, w_077_2953, w_077_2955, w_077_2958, w_077_2965, w_077_2966, w_077_2968, w_077_2970, w_077_2975, w_077_2978, w_077_2981, w_077_2984, w_077_2987, w_077_2994, w_077_2995, w_077_3002, w_077_3005, w_077_3006, w_077_3009, w_077_3010, w_077_3013, w_077_3014, w_077_3016, w_077_3023, w_077_3024, w_077_3025, w_077_3026, w_077_3027, w_077_3033, w_077_3041, w_077_3045, w_077_3050, w_077_3052, w_077_3055, w_077_3058, w_077_3059, w_077_3062, w_077_3063, w_077_3070, w_077_3072, w_077_3074, w_077_3075, w_077_3076, w_077_3078, w_077_3079, w_077_3080, w_077_3085, w_077_3088, w_077_3089, w_077_3090, w_077_3092, w_077_3093, w_077_3094, w_077_3097, w_077_3098, w_077_3099, w_077_3102, w_077_3105, w_077_3107, w_077_3109, w_077_3111, w_077_3113, w_077_3114, w_077_3121, w_077_3123, w_077_3125, w_077_3127, w_077_3140, w_077_3141, w_077_3145, w_077_3148, w_077_3150, w_077_3152, w_077_3154, w_077_3155, w_077_3164, w_077_3167, w_077_3168, w_077_3172, w_077_3179, w_077_3180, w_077_3181, w_077_3182, w_077_3183, w_077_3184, w_077_3188, w_077_3189, w_077_3190, w_077_3191, w_077_3192, w_077_3194;
  wire w_078_000, w_078_001, w_078_002, w_078_003, w_078_004, w_078_005, w_078_006, w_078_007, w_078_008, w_078_009, w_078_010, w_078_011, w_078_012, w_078_013, w_078_014, w_078_015, w_078_016, w_078_017, w_078_018, w_078_019, w_078_020, w_078_021, w_078_022, w_078_023, w_078_024, w_078_025, w_078_026, w_078_027, w_078_028, w_078_029, w_078_030, w_078_031, w_078_032, w_078_033, w_078_034, w_078_035, w_078_036, w_078_037, w_078_038, w_078_039, w_078_040, w_078_041, w_078_042, w_078_043, w_078_044, w_078_045, w_078_046, w_078_047, w_078_048, w_078_049, w_078_050, w_078_052, w_078_053, w_078_054, w_078_055, w_078_056, w_078_057, w_078_058, w_078_059, w_078_060, w_078_061, w_078_062, w_078_063, w_078_064, w_078_065, w_078_066, w_078_067, w_078_068, w_078_069, w_078_070, w_078_071, w_078_072, w_078_073, w_078_074, w_078_075, w_078_076, w_078_077, w_078_078, w_078_079, w_078_080, w_078_081, w_078_082, w_078_083, w_078_084, w_078_085, w_078_086, w_078_087, w_078_088, w_078_089, w_078_090, w_078_091, w_078_092, w_078_093, w_078_094, w_078_095, w_078_096, w_078_097, w_078_098, w_078_099, w_078_100, w_078_101, w_078_102, w_078_103, w_078_104, w_078_105, w_078_106, w_078_107, w_078_108, w_078_109, w_078_110, w_078_111, w_078_112, w_078_113, w_078_114, w_078_116, w_078_117, w_078_118, w_078_119, w_078_120, w_078_121, w_078_122, w_078_123, w_078_124, w_078_125, w_078_126, w_078_127, w_078_128, w_078_129, w_078_130, w_078_131, w_078_132, w_078_133, w_078_134, w_078_135, w_078_136, w_078_137, w_078_138, w_078_139, w_078_140, w_078_141, w_078_142, w_078_143, w_078_144, w_078_145, w_078_146, w_078_147, w_078_148, w_078_149, w_078_150, w_078_151, w_078_152, w_078_153, w_078_154, w_078_155, w_078_156, w_078_157, w_078_158, w_078_159, w_078_160, w_078_161, w_078_162, w_078_163, w_078_164, w_078_165, w_078_166, w_078_167, w_078_168, w_078_169, w_078_170, w_078_171, w_078_172, w_078_173, w_078_174, w_078_175, w_078_176, w_078_177, w_078_178, w_078_179, w_078_180, w_078_181, w_078_182, w_078_183, w_078_184, w_078_185, w_078_186, w_078_187, w_078_188, w_078_189, w_078_190, w_078_191, w_078_192, w_078_193, w_078_194, w_078_195, w_078_196, w_078_197, w_078_198, w_078_199, w_078_200, w_078_201, w_078_202, w_078_203, w_078_204, w_078_205, w_078_206, w_078_207, w_078_208, w_078_209, w_078_210, w_078_211, w_078_212, w_078_213, w_078_214, w_078_215, w_078_216, w_078_217, w_078_218, w_078_219, w_078_220, w_078_221, w_078_222, w_078_223, w_078_224, w_078_225, w_078_226, w_078_227, w_078_228, w_078_229, w_078_230, w_078_231, w_078_232, w_078_233, w_078_234, w_078_235, w_078_236, w_078_237, w_078_238, w_078_239, w_078_240, w_078_241, w_078_242, w_078_243, w_078_244, w_078_245, w_078_246, w_078_247, w_078_248, w_078_249, w_078_250, w_078_251, w_078_252, w_078_253, w_078_254, w_078_255, w_078_256, w_078_257, w_078_258, w_078_259, w_078_260, w_078_261, w_078_262, w_078_263, w_078_264, w_078_265, w_078_266, w_078_267, w_078_268, w_078_269, w_078_270, w_078_271, w_078_272, w_078_273, w_078_274, w_078_275, w_078_276, w_078_277, w_078_278, w_078_279, w_078_280, w_078_281, w_078_282, w_078_283, w_078_284, w_078_285, w_078_286, w_078_287, w_078_288, w_078_289, w_078_290, w_078_291, w_078_292, w_078_293, w_078_294, w_078_295, w_078_296, w_078_297, w_078_298, w_078_299, w_078_300, w_078_301, w_078_302, w_078_303, w_078_304, w_078_305, w_078_306, w_078_307, w_078_308, w_078_309, w_078_310, w_078_311, w_078_312, w_078_313, w_078_314, w_078_315, w_078_316, w_078_317, w_078_318, w_078_319, w_078_320, w_078_321, w_078_322, w_078_323, w_078_324, w_078_325, w_078_326, w_078_327, w_078_328, w_078_329, w_078_330, w_078_331, w_078_332, w_078_333, w_078_334, w_078_335, w_078_336, w_078_337, w_078_338, w_078_339, w_078_340, w_078_341, w_078_342, w_078_343, w_078_344, w_078_345, w_078_346, w_078_347, w_078_348, w_078_349, w_078_350, w_078_351, w_078_352, w_078_353, w_078_354, w_078_355, w_078_356, w_078_357, w_078_358, w_078_359, w_078_360, w_078_361, w_078_362, w_078_363, w_078_364, w_078_365, w_078_366, w_078_367, w_078_368, w_078_369, w_078_370, w_078_371, w_078_372, w_078_373, w_078_374, w_078_375, w_078_376, w_078_377, w_078_378, w_078_379, w_078_380, w_078_381, w_078_382, w_078_383, w_078_384, w_078_385, w_078_386, w_078_387, w_078_388, w_078_389, w_078_390, w_078_391, w_078_392, w_078_393, w_078_394, w_078_395, w_078_396, w_078_397, w_078_398, w_078_399, w_078_400, w_078_401, w_078_402, w_078_403, w_078_404, w_078_405, w_078_406, w_078_407, w_078_408, w_078_409, w_078_410, w_078_411, w_078_412, w_078_413, w_078_414, w_078_415, w_078_416, w_078_417, w_078_418, w_078_419, w_078_420, w_078_421, w_078_422, w_078_423, w_078_424, w_078_425, w_078_426, w_078_427;
  wire w_079_000, w_079_002, w_079_003, w_079_006, w_079_007, w_079_008, w_079_009, w_079_011, w_079_014, w_079_015, w_079_017, w_079_019, w_079_020, w_079_022, w_079_027, w_079_030, w_079_031, w_079_033, w_079_034, w_079_035, w_079_036, w_079_037, w_079_038, w_079_039, w_079_042, w_079_043, w_079_044, w_079_045, w_079_046, w_079_047, w_079_049, w_079_051, w_079_052, w_079_053, w_079_054, w_079_055, w_079_057, w_079_058, w_079_059, w_079_061, w_079_066, w_079_072, w_079_073, w_079_075, w_079_077, w_079_078, w_079_079, w_079_081, w_079_082, w_079_083, w_079_086, w_079_089, w_079_090, w_079_091, w_079_092, w_079_096, w_079_097, w_079_098, w_079_104, w_079_111, w_079_112, w_079_116, w_079_121, w_079_123, w_079_124, w_079_125, w_079_127, w_079_131, w_079_132, w_079_137, w_079_138, w_079_140, w_079_143, w_079_144, w_079_150, w_079_152, w_079_153, w_079_155, w_079_158, w_079_160, w_079_161, w_079_163, w_079_164, w_079_165, w_079_167, w_079_168, w_079_169, w_079_170, w_079_171, w_079_172, w_079_173, w_079_174, w_079_175, w_079_177, w_079_178, w_079_179, w_079_183, w_079_185, w_079_187, w_079_188, w_079_191, w_079_192, w_079_193, w_079_198, w_079_200, w_079_201, w_079_207, w_079_208, w_079_209, w_079_210, w_079_211, w_079_212, w_079_214, w_079_215, w_079_217, w_079_218, w_079_219, w_079_220, w_079_222, w_079_223, w_079_224, w_079_225, w_079_227, w_079_229, w_079_231, w_079_232, w_079_234, w_079_235, w_079_236, w_079_239, w_079_241, w_079_242, w_079_244, w_079_245, w_079_246, w_079_247, w_079_249, w_079_250, w_079_251, w_079_253, w_079_254, w_079_258, w_079_259, w_079_267, w_079_268, w_079_269, w_079_270, w_079_272, w_079_273, w_079_274, w_079_275, w_079_278, w_079_281, w_079_282, w_079_284, w_079_285, w_079_292, w_079_294, w_079_298, w_079_299, w_079_300, w_079_301, w_079_302, w_079_303, w_079_306, w_079_307, w_079_308, w_079_309, w_079_313, w_079_315, w_079_317, w_079_321, w_079_323, w_079_326, w_079_328, w_079_331, w_079_332, w_079_333, w_079_335, w_079_337, w_079_338, w_079_340, w_079_345, w_079_346, w_079_348, w_079_349, w_079_350, w_079_351, w_079_352, w_079_353, w_079_354, w_079_355, w_079_363, w_079_364, w_079_365, w_079_366, w_079_367, w_079_369, w_079_372, w_079_373, w_079_375, w_079_376, w_079_377, w_079_378, w_079_380, w_079_381, w_079_382, w_079_384, w_079_386, w_079_388, w_079_389, w_079_390, w_079_392, w_079_393, w_079_394, w_079_395, w_079_396, w_079_397, w_079_398, w_079_400, w_079_403, w_079_404, w_079_408, w_079_409, w_079_410, w_079_415, w_079_417, w_079_418, w_079_419, w_079_422, w_079_423, w_079_424, w_079_425, w_079_427, w_079_428, w_079_429, w_079_430, w_079_431, w_079_432, w_079_433, w_079_434, w_079_435, w_079_437, w_079_441, w_079_445, w_079_446, w_079_450, w_079_451, w_079_452, w_079_454, w_079_455, w_079_460, w_079_466, w_079_470, w_079_473, w_079_475, w_079_476, w_079_478, w_079_479, w_079_481, w_079_482, w_079_483, w_079_485, w_079_486, w_079_487, w_079_488, w_079_489, w_079_491, w_079_492, w_079_493, w_079_494, w_079_497, w_079_500, w_079_501, w_079_503, w_079_506, w_079_508, w_079_509, w_079_510, w_079_511, w_079_512, w_079_513, w_079_514, w_079_515, w_079_519, w_079_523, w_079_524, w_079_525, w_079_526, w_079_527, w_079_528, w_079_530, w_079_531, w_079_534, w_079_535, w_079_536, w_079_539, w_079_540, w_079_543, w_079_550, w_079_552, w_079_555, w_079_557, w_079_558, w_079_559, w_079_560, w_079_564, w_079_565, w_079_569, w_079_570, w_079_571, w_079_572, w_079_573, w_079_574, w_079_575, w_079_576, w_079_579, w_079_582, w_079_584, w_079_585, w_079_588, w_079_589, w_079_591, w_079_592, w_079_593, w_079_595, w_079_597, w_079_598, w_079_599, w_079_601, w_079_603, w_079_604, w_079_606, w_079_607, w_079_609, w_079_611, w_079_612, w_079_613, w_079_614, w_079_617, w_079_618, w_079_619, w_079_620, w_079_621, w_079_623, w_079_626, w_079_627, w_079_628, w_079_629, w_079_631, w_079_636, w_079_637, w_079_639, w_079_640, w_079_641, w_079_642, w_079_644, w_079_645, w_079_646, w_079_647, w_079_648, w_079_649, w_079_650, w_079_651, w_079_653, w_079_657, w_079_658, w_079_659, w_079_660, w_079_664, w_079_665, w_079_666, w_079_668, w_079_669, w_079_674, w_079_675, w_079_677, w_079_679, w_079_681, w_079_683, w_079_686, w_079_692, w_079_695, w_079_698, w_079_699, w_079_701, w_079_705, w_079_708, w_079_709, w_079_710, w_079_711, w_079_714, w_079_717, w_079_721, w_079_722, w_079_724, w_079_725, w_079_729, w_079_731, w_079_732, w_079_735, w_079_737, w_079_739, w_079_740, w_079_741, w_079_742, w_079_743, w_079_745, w_079_748, w_079_750, w_079_752, w_079_754, w_079_757, w_079_761, w_079_763, w_079_767, w_079_768, w_079_769, w_079_772, w_079_773, w_079_776, w_079_778, w_079_779, w_079_782, w_079_783, w_079_786, w_079_787, w_079_788, w_079_790, w_079_793, w_079_794, w_079_795, w_079_796, w_079_797, w_079_798, w_079_799, w_079_801, w_079_802, w_079_804, w_079_807, w_079_808, w_079_809, w_079_810, w_079_811, w_079_812, w_079_815, w_079_816, w_079_817, w_079_818, w_079_822, w_079_823, w_079_824, w_079_825, w_079_827, w_079_828, w_079_830, w_079_831, w_079_832, w_079_833, w_079_835, w_079_836, w_079_838, w_079_839, w_079_840, w_079_841, w_079_843, w_079_846, w_079_848, w_079_849, w_079_850, w_079_851, w_079_852, w_079_854, w_079_855, w_079_856, w_079_857, w_079_860, w_079_861, w_079_864, w_079_865, w_079_866, w_079_868, w_079_870, w_079_872, w_079_873, w_079_874, w_079_877, w_079_878, w_079_879, w_079_880, w_079_881, w_079_882, w_079_883, w_079_885, w_079_886, w_079_887, w_079_888, w_079_890, w_079_891, w_079_894, w_079_895, w_079_897, w_079_898, w_079_900, w_079_902, w_079_903, w_079_905, w_079_908, w_079_909, w_079_911, w_079_912, w_079_913, w_079_914, w_079_915, w_079_921, w_079_922, w_079_924, w_079_925, w_079_926, w_079_929, w_079_930, w_079_932, w_079_934, w_079_935, w_079_936, w_079_939, w_079_940, w_079_941, w_079_944, w_079_945, w_079_946, w_079_947, w_079_949, w_079_950, w_079_951, w_079_952, w_079_958, w_079_959, w_079_960, w_079_962, w_079_963, w_079_964, w_079_965, w_079_966, w_079_967, w_079_968, w_079_969, w_079_972, w_079_973, w_079_974, w_079_976, w_079_978, w_079_979, w_079_980, w_079_981, w_079_983, w_079_984, w_079_986, w_079_987, w_079_988, w_079_990, w_079_991, w_079_992, w_079_994, w_079_997, w_079_998, w_079_999, w_079_1006, w_079_1007, w_079_1011, w_079_1012, w_079_1017, w_079_1018, w_079_1020, w_079_1022, w_079_1023, w_079_1025, w_079_1027, w_079_1028, w_079_1029, w_079_1031, w_079_1032, w_079_1033, w_079_1034, w_079_1035, w_079_1037, w_079_1038, w_079_1043, w_079_1044, w_079_1046, w_079_1048, w_079_1049, w_079_1050, w_079_1052, w_079_1053, w_079_1054, w_079_1055, w_079_1057, w_079_1058, w_079_1059, w_079_1060, w_079_1061, w_079_1063, w_079_1065, w_079_1068, w_079_1072, w_079_1073, w_079_1074, w_079_1075, w_079_1078, w_079_1082, w_079_1085, w_079_1086, w_079_1089, w_079_1091, w_079_1096, w_079_1097, w_079_1101, w_079_1102, w_079_1103, w_079_1105, w_079_1108, w_079_1109, w_079_1113, w_079_1120, w_079_1121, w_079_1127, w_079_1128, w_079_1130, w_079_1137, w_079_1138, w_079_1141, w_079_1142, w_079_1143, w_079_1144, w_079_1145, w_079_1147, w_079_1148, w_079_1150, w_079_1151, w_079_1154, w_079_1156, w_079_1158, w_079_1161, w_079_1162, w_079_1166, w_079_1169, w_079_1170, w_079_1172, w_079_1173, w_079_1175, w_079_1177, w_079_1178, w_079_1179, w_079_1182, w_079_1185, w_079_1186, w_079_1187, w_079_1188, w_079_1192, w_079_1196, w_079_1197, w_079_1198, w_079_1199, w_079_1200, w_079_1202, w_079_1205, w_079_1208, w_079_1210, w_079_1211, w_079_1212, w_079_1213, w_079_1214, w_079_1215, w_079_1216, w_079_1217, w_079_1218, w_079_1220, w_079_1221, w_079_1224, w_079_1226, w_079_1234, w_079_1236, w_079_1237, w_079_1239, w_079_1240, w_079_1241, w_079_1242, w_079_1246, w_079_1247, w_079_1248, w_079_1249, w_079_1251, w_079_1252, w_079_1253, w_079_1256, w_079_1262, w_079_1263, w_079_1264, w_079_1265, w_079_1271, w_079_1272, w_079_1273, w_079_1274, w_079_1276, w_079_1279, w_079_1281, w_079_1282, w_079_1283, w_079_1286, w_079_1287, w_079_1288, w_079_1290, w_079_1292, w_079_1293, w_079_1294, w_079_1295, w_079_1296, w_079_1299, w_079_1300, w_079_1301, w_079_1302, w_079_1303, w_079_1305, w_079_1306, w_079_1307, w_079_1308, w_079_1310, w_079_1311, w_079_1312, w_079_1313, w_079_1316, w_079_1317, w_079_1318, w_079_1320, w_079_1321, w_079_1325, w_079_1326, w_079_1327, w_079_1330, w_079_1331, w_079_1332, w_079_1335, w_079_1336, w_079_1338, w_079_1340, w_079_1342, w_079_1343, w_079_1344, w_079_1345, w_079_1352, w_079_1353, w_079_1354, w_079_1356, w_079_1357, w_079_1358, w_079_1359, w_079_1360, w_079_1364, w_079_1369, w_079_1370, w_079_1371, w_079_1373, w_079_1374, w_079_1375, w_079_1376, w_079_1377, w_079_1378, w_079_1379, w_079_1380, w_079_1382, w_079_1384, w_079_1385, w_079_1387, w_079_1391, w_079_1392, w_079_1393, w_079_1394, w_079_1395, w_079_1397, w_079_1398, w_079_1400, w_079_1402, w_079_1403, w_079_1404, w_079_1406, w_079_1410, w_079_1418, w_079_1419, w_079_1420, w_079_1425, w_079_1428, w_079_1430, w_079_1432, w_079_1434, w_079_1435, w_079_1436, w_079_1438, w_079_1439, w_079_1440, w_079_1441, w_079_1442, w_079_1444, w_079_1446, w_079_1448, w_079_1450, w_079_1451, w_079_1455, w_079_1459, w_079_1463, w_079_1465, w_079_1466, w_079_1467, w_079_1471, w_079_1473, w_079_1475, w_079_1478, w_079_1484, w_079_1485, w_079_1486, w_079_1487, w_079_1489, w_079_1491, w_079_1493, w_079_1494, w_079_1496, w_079_1497, w_079_1498, w_079_1500, w_079_1502, w_079_1503, w_079_1505, w_079_1507, w_079_1508, w_079_1511, w_079_1512, w_079_1513, w_079_1514, w_079_1515, w_079_1516, w_079_1517, w_079_1518, w_079_1519, w_079_1520, w_079_1521, w_079_1522, w_079_1526, w_079_1531, w_079_1534, w_079_1535, w_079_1536, w_079_1537, w_079_1539, w_079_1540, w_079_1543, w_079_1544, w_079_1545, w_079_1546, w_079_1548, w_079_1551, w_079_1553, w_079_1554, w_079_1555, w_079_1556, w_079_1557, w_079_1558, w_079_1561, w_079_1562, w_079_1564, w_079_1566, w_079_1567, w_079_1568, w_079_1569, w_079_1571, w_079_1574, w_079_1576, w_079_1580, w_079_1586, w_079_1593, w_079_1594, w_079_1595, w_079_1596, w_079_1597, w_079_1598, w_079_1600, w_079_1601, w_079_1602, w_079_1603, w_079_1604, w_079_1605, w_079_1608, w_079_1612, w_079_1613, w_079_1616, w_079_1617, w_079_1618, w_079_1619, w_079_1620, w_079_1621, w_079_1624, w_079_1625, w_079_1626, w_079_1632, w_079_1633, w_079_1634, w_079_1636, w_079_1637, w_079_1638, w_079_1640, w_079_1641, w_079_1642, w_079_1645, w_079_1647, w_079_1648, w_079_1649, w_079_1651, w_079_1653, w_079_1654, w_079_1655, w_079_1656, w_079_1657, w_079_1658, w_079_1659, w_079_1662, w_079_1666, w_079_1667, w_079_1668, w_079_1670, w_079_1674, w_079_1675, w_079_1676, w_079_1679, w_079_1683, w_079_1684, w_079_1685, w_079_1687, w_079_1690, w_079_1691, w_079_1692, w_079_1695, w_079_1696, w_079_1697, w_079_1699, w_079_1702, w_079_1706, w_079_1708, w_079_1711, w_079_1712, w_079_1713, w_079_1717, w_079_1718, w_079_1720, w_079_1721, w_079_1722, w_079_1725, w_079_1726, w_079_1729, w_079_1731, w_079_1733, w_079_1734, w_079_1735, w_079_1736, w_079_1737, w_079_1738, w_079_1740, w_079_1742, w_079_1746, w_079_1747, w_079_1749, w_079_1750, w_079_1751, w_079_1754, w_079_1756, w_079_1757, w_079_1758, w_079_1759, w_079_1760, w_079_1764, w_079_1766, w_079_1768, w_079_1769, w_079_1771, w_079_1775, w_079_1777, w_079_1779, w_079_1780, w_079_1781, w_079_1782, w_079_1785, w_079_1786, w_079_1790, w_079_1791, w_079_1793, w_079_1799, w_079_1801, w_079_1802, w_079_1804, w_079_1806, w_079_1807, w_079_1809, w_079_1811, w_079_1812, w_079_1813, w_079_1814, w_079_1815, w_079_1817, w_079_1818, w_079_1819, w_079_1820, w_079_1821, w_079_1822, w_079_1823, w_079_1824, w_079_1826, w_079_1827, w_079_1828, w_079_1830, w_079_1831, w_079_1832, w_079_1834, w_079_1837, w_079_1838, w_079_1839, w_079_1842, w_079_1844, w_079_1845, w_079_1846, w_079_1849, w_079_1850, w_079_1851, w_079_1855, w_079_1857, w_079_1859, w_079_1860, w_079_1861, w_079_1863, w_079_1865, w_079_1866, w_079_1869, w_079_1870, w_079_1871, w_079_1873, w_079_1875, w_079_1876, w_079_1878, w_079_1879, w_079_1880, w_079_1882, w_079_1883, w_079_1888, w_079_1889, w_079_1890, w_079_1891, w_079_1892, w_079_1893, w_079_1894, w_079_1896, w_079_1897, w_079_1898, w_079_1903, w_079_1904, w_079_1905, w_079_1907, w_079_1909, w_079_1910, w_079_1912, w_079_1914, w_079_1916, w_079_1917, w_079_1921, w_079_1922, w_079_1924, w_079_1925, w_079_1926, w_079_1927, w_079_1934, w_079_1935, w_079_1936, w_079_1938, w_079_1939, w_079_1940, w_079_1942, w_079_1943, w_079_1945, w_079_1946, w_079_1948, w_079_1950, w_079_1951, w_079_1952, w_079_1953, w_079_1954, w_079_1956, w_079_1957, w_079_1958, w_079_1959, w_079_1961, w_079_1962, w_079_1964, w_079_1965, w_079_1967, w_079_1968, w_079_1969, w_079_1971, w_079_1973, w_079_1974, w_079_1983, w_079_1984, w_079_1987, w_079_1989, w_079_1990, w_079_1997, w_079_1998, w_079_2000, w_079_2009, w_079_2010, w_079_2011, w_079_2015, w_079_2016, w_079_2017, w_079_2021, w_079_2022, w_079_2024, w_079_2026, w_079_2027, w_079_2028, w_079_2030, w_079_2032, w_079_2034, w_079_2035, w_079_2037, w_079_2038, w_079_2040, w_079_2041, w_079_2048, w_079_2050, w_079_2052, w_079_2060, w_079_2062, w_079_2068, w_079_2070, w_079_2072, w_079_2075, w_079_2077, w_079_2084, w_079_2087, w_079_2093, w_079_2095, w_079_2097, w_079_2105, w_079_2106, w_079_2108, w_079_2110, w_079_2111, w_079_2117, w_079_2121, w_079_2127, w_079_2130, w_079_2131, w_079_2132, w_079_2136, w_079_2137, w_079_2142, w_079_2147, w_079_2148, w_079_2152, w_079_2154, w_079_2163, w_079_2165, w_079_2166, w_079_2172, w_079_2181, w_079_2184, w_079_2185, w_079_2188, w_079_2189, w_079_2191, w_079_2193, w_079_2194, w_079_2197, w_079_2200, w_079_2203, w_079_2207, w_079_2210, w_079_2213, w_079_2215, w_079_2216, w_079_2218, w_079_2220, w_079_2223, w_079_2225, w_079_2226, w_079_2230, w_079_2234, w_079_2236, w_079_2247, w_079_2249, w_079_2259, w_079_2260, w_079_2266, w_079_2269, w_079_2270, w_079_2272, w_079_2275, w_079_2280, w_079_2281, w_079_2283, w_079_2284, w_079_2289, w_079_2291, w_079_2292, w_079_2294, w_079_2295, w_079_2297, w_079_2307, w_079_2311, w_079_2312, w_079_2323, w_079_2331, w_079_2332, w_079_2334, w_079_2335, w_079_2337, w_079_2338, w_079_2341, w_079_2342, w_079_2343, w_079_2346, w_079_2350, w_079_2353, w_079_2360, w_079_2370, w_079_2371, w_079_2373, w_079_2376, w_079_2384, w_079_2386, w_079_2387, w_079_2392, w_079_2393, w_079_2394, w_079_2395, w_079_2397, w_079_2401, w_079_2404, w_079_2406, w_079_2407, w_079_2408, w_079_2409, w_079_2412, w_079_2413, w_079_2421, w_079_2422, w_079_2423, w_079_2424, w_079_2433, w_079_2434, w_079_2439, w_079_2442, w_079_2447, w_079_2449, w_079_2453, w_079_2455, w_079_2458, w_079_2462, w_079_2464, w_079_2471, w_079_2472, w_079_2474, w_079_2479, w_079_2480, w_079_2481, w_079_2482, w_079_2484, w_079_2485, w_079_2488, w_079_2492, w_079_2499, w_079_2503, w_079_2509, w_079_2510, w_079_2511, w_079_2512, w_079_2519, w_079_2526, w_079_2530, w_079_2534, w_079_2535, w_079_2536, w_079_2540, w_079_2541, w_079_2548, w_079_2551, w_079_2552, w_079_2554, w_079_2556, w_079_2557, w_079_2558, w_079_2560, w_079_2568, w_079_2577, w_079_2580, w_079_2584, w_079_2585, w_079_2592, w_079_2594, w_079_2595, w_079_2596, w_079_2597, w_079_2598, w_079_2603, w_079_2604, w_079_2611, w_079_2613, w_079_2614, w_079_2616, w_079_2617, w_079_2619, w_079_2620, w_079_2625, w_079_2626, w_079_2630, w_079_2631, w_079_2633, w_079_2637, w_079_2638, w_079_2640, w_079_2641, w_079_2644, w_079_2645, w_079_2647, w_079_2653, w_079_2654, w_079_2656, w_079_2658, w_079_2664, w_079_2665, w_079_2666, w_079_2667, w_079_2670, w_079_2673, w_079_2674, w_079_2676, w_079_2678, w_079_2681, w_079_2682, w_079_2684, w_079_2689, w_079_2690, w_079_2696, w_079_2699, w_079_2703, w_079_2705, w_079_2710, w_079_2713, w_079_2717, w_079_2723, w_079_2724, w_079_2727, w_079_2731, w_079_2732, w_079_2734, w_079_2739, w_079_2741, w_079_2742, w_079_2747, w_079_2758, w_079_2760, w_079_2763, w_079_2765, w_079_2768, w_079_2772, w_079_2777, w_079_2778, w_079_2781, w_079_2782, w_079_2783, w_079_2784, w_079_2785, w_079_2786, w_079_2790, w_079_2792, w_079_2796, w_079_2802, w_079_2811, w_079_2816, w_079_2818, w_079_2822, w_079_2826, w_079_2827, w_079_2829, w_079_2830, w_079_2832, w_079_2834, w_079_2838, w_079_2839, w_079_2840, w_079_2851, w_079_2852, w_079_2855, w_079_2857, w_079_2860, w_079_2862, w_079_2866, w_079_2875, w_079_2876, w_079_2878, w_079_2881, w_079_2882, w_079_2884, w_079_2886, w_079_2888, w_079_2890, w_079_2891, w_079_2895, w_079_2902, w_079_2903, w_079_2909, w_079_2913, w_079_2917, w_079_2918, w_079_2920, w_079_2923, w_079_2924, w_079_2927, w_079_2928, w_079_2929, w_079_2930, w_079_2936, w_079_2941, w_079_2942, w_079_2948, w_079_2949, w_079_2952, w_079_2957, w_079_2959, w_079_2960, w_079_2961, w_079_2962, w_079_2965, w_079_2970, w_079_2972, w_079_2973, w_079_2976, w_079_2977, w_079_2984, w_079_2985, w_079_2986, w_079_2987, w_079_2988, w_079_2989, w_079_2992, w_079_2996, w_079_3001, w_079_3003, w_079_3005, w_079_3007, w_079_3009, w_079_3010, w_079_3011, w_079_3014;
  wire w_080_000, w_080_004, w_080_006, w_080_009, w_080_012, w_080_015, w_080_016, w_080_019, w_080_021, w_080_024, w_080_025, w_080_026, w_080_028, w_080_029, w_080_030, w_080_037, w_080_039, w_080_042, w_080_052, w_080_053, w_080_055, w_080_058, w_080_059, w_080_060, w_080_064, w_080_066, w_080_068, w_080_073, w_080_075, w_080_076, w_080_080, w_080_081, w_080_082, w_080_085, w_080_089, w_080_092, w_080_094, w_080_096, w_080_097, w_080_100, w_080_101, w_080_102, w_080_107, w_080_108, w_080_110, w_080_112, w_080_114, w_080_115, w_080_116, w_080_117, w_080_118, w_080_119, w_080_125, w_080_127, w_080_129, w_080_130, w_080_132, w_080_133, w_080_134, w_080_135, w_080_139, w_080_144, w_080_145, w_080_146, w_080_149, w_080_150, w_080_153, w_080_154, w_080_159, w_080_160, w_080_165, w_080_166, w_080_167, w_080_168, w_080_169, w_080_170, w_080_171, w_080_172, w_080_177, w_080_179, w_080_180, w_080_181, w_080_182, w_080_185, w_080_187, w_080_188, w_080_190, w_080_192, w_080_194, w_080_195, w_080_196, w_080_200, w_080_202, w_080_203, w_080_204, w_080_206, w_080_207, w_080_208, w_080_210, w_080_211, w_080_212, w_080_215, w_080_219, w_080_220, w_080_225, w_080_226, w_080_227, w_080_228, w_080_231, w_080_233, w_080_234, w_080_235, w_080_236, w_080_238, w_080_239, w_080_240, w_080_241, w_080_243, w_080_245, w_080_247, w_080_251, w_080_252, w_080_253, w_080_254, w_080_257, w_080_258, w_080_262, w_080_268, w_080_269, w_080_270, w_080_271, w_080_272, w_080_275, w_080_276, w_080_280, w_080_282, w_080_285, w_080_286, w_080_289, w_080_290, w_080_292, w_080_294, w_080_295, w_080_301, w_080_302, w_080_304, w_080_305, w_080_307, w_080_309, w_080_312, w_080_313, w_080_314, w_080_316, w_080_318, w_080_320, w_080_321, w_080_323, w_080_324, w_080_327, w_080_330, w_080_333, w_080_334, w_080_337, w_080_339, w_080_341, w_080_342, w_080_343, w_080_344, w_080_345, w_080_349, w_080_350, w_080_352, w_080_353, w_080_354, w_080_358, w_080_359, w_080_361, w_080_362, w_080_364, w_080_365, w_080_366, w_080_367, w_080_368, w_080_369, w_080_370, w_080_371, w_080_372, w_080_373, w_080_374, w_080_375, w_080_376, w_080_378, w_080_380, w_080_381, w_080_383, w_080_384, w_080_385, w_080_386, w_080_388, w_080_390, w_080_392, w_080_393, w_080_396, w_080_397, w_080_398, w_080_403, w_080_406, w_080_408, w_080_409, w_080_411, w_080_413, w_080_414, w_080_417, w_080_420, w_080_421, w_080_422, w_080_423, w_080_424, w_080_425, w_080_426, w_080_427, w_080_429, w_080_430, w_080_431, w_080_432, w_080_437, w_080_438, w_080_440, w_080_444, w_080_446, w_080_447, w_080_449, w_080_450, w_080_453, w_080_455, w_080_459, w_080_460, w_080_461, w_080_462, w_080_465, w_080_466, w_080_467, w_080_469, w_080_472, w_080_473, w_080_476, w_080_477, w_080_480, w_080_482, w_080_483, w_080_484, w_080_485, w_080_486, w_080_487, w_080_490, w_080_495, w_080_498, w_080_499, w_080_500, w_080_501, w_080_507, w_080_509, w_080_511, w_080_513, w_080_514, w_080_515, w_080_517, w_080_519, w_080_528, w_080_531, w_080_533, w_080_535, w_080_536, w_080_538, w_080_539, w_080_541, w_080_542, w_080_543, w_080_548, w_080_553, w_080_554, w_080_555, w_080_556, w_080_558, w_080_559, w_080_561, w_080_562, w_080_563, w_080_565, w_080_566, w_080_569, w_080_571, w_080_572, w_080_573, w_080_576, w_080_577, w_080_581, w_080_582, w_080_584, w_080_585, w_080_587, w_080_590, w_080_592, w_080_593, w_080_596, w_080_598, w_080_599, w_080_600, w_080_601, w_080_604, w_080_605, w_080_606, w_080_607, w_080_612, w_080_613, w_080_615, w_080_616, w_080_618, w_080_619, w_080_621, w_080_624, w_080_627, w_080_628, w_080_630, w_080_636, w_080_637, w_080_638, w_080_639, w_080_641, w_080_643, w_080_644, w_080_646, w_080_650, w_080_651, w_080_652, w_080_654, w_080_655, w_080_656, w_080_657, w_080_658, w_080_659, w_080_661, w_080_664, w_080_665, w_080_666, w_080_668, w_080_670, w_080_676, w_080_677, w_080_678, w_080_680, w_080_681, w_080_682, w_080_684, w_080_686, w_080_690, w_080_691, w_080_693, w_080_695, w_080_696, w_080_697, w_080_698, w_080_700, w_080_702, w_080_704, w_080_710, w_080_714, w_080_715, w_080_716, w_080_717, w_080_718, w_080_719, w_080_722, w_080_723, w_080_724, w_080_725, w_080_726, w_080_727, w_080_729, w_080_730, w_080_733, w_080_735, w_080_736, w_080_737, w_080_738, w_080_741, w_080_743, w_080_745, w_080_746, w_080_747, w_080_749, w_080_751, w_080_752, w_080_753, w_080_754, w_080_755, w_080_757, w_080_758, w_080_759, w_080_760, w_080_763, w_080_764, w_080_766, w_080_771, w_080_772, w_080_773, w_080_774, w_080_775, w_080_776, w_080_777, w_080_778, w_080_779, w_080_780, w_080_781, w_080_782, w_080_784, w_080_785, w_080_786, w_080_787, w_080_790, w_080_791, w_080_792, w_080_793, w_080_794, w_080_796, w_080_797, w_080_798, w_080_799, w_080_800, w_080_801, w_080_802, w_080_805, w_080_807, w_080_808, w_080_809, w_080_811, w_080_812, w_080_814, w_080_820, w_080_821, w_080_823, w_080_826, w_080_827, w_080_831, w_080_832, w_080_833, w_080_834, w_080_839, w_080_840, w_080_841, w_080_842, w_080_843, w_080_844, w_080_845, w_080_846, w_080_848, w_080_851, w_080_852, w_080_855, w_080_857, w_080_859, w_080_862, w_080_864, w_080_865, w_080_868, w_080_870, w_080_871, w_080_875, w_080_878, w_080_879, w_080_880, w_080_883, w_080_884, w_080_885, w_080_888, w_080_890, w_080_893, w_080_899, w_080_902, w_080_904, w_080_905, w_080_906, w_080_908, w_080_909, w_080_910, w_080_911, w_080_915, w_080_916, w_080_918, w_080_919, w_080_920, w_080_922, w_080_923, w_080_925, w_080_927, w_080_930, w_080_931, w_080_933, w_080_935, w_080_936, w_080_937, w_080_939, w_080_940, w_080_941, w_080_942, w_080_945, w_080_946, w_080_947, w_080_948, w_080_949, w_080_951, w_080_952, w_080_953, w_080_955, w_080_956, w_080_957, w_080_961, w_080_965, w_080_967, w_080_972, w_080_975, w_080_977, w_080_979, w_080_982, w_080_984, w_080_985, w_080_991, w_080_993, w_080_995, w_080_996, w_080_1001, w_080_1003, w_080_1006, w_080_1008, w_080_1011, w_080_1012, w_080_1013, w_080_1016, w_080_1017, w_080_1020, w_080_1021, w_080_1023, w_080_1024, w_080_1025, w_080_1026, w_080_1027, w_080_1029, w_080_1030, w_080_1031, w_080_1032, w_080_1033, w_080_1034, w_080_1036, w_080_1037, w_080_1040, w_080_1043, w_080_1044, w_080_1045, w_080_1046, w_080_1047, w_080_1048, w_080_1050, w_080_1051, w_080_1053, w_080_1055, w_080_1057, w_080_1061, w_080_1065, w_080_1066, w_080_1067, w_080_1069, w_080_1070, w_080_1071, w_080_1073, w_080_1074, w_080_1075, w_080_1077, w_080_1078, w_080_1079, w_080_1081, w_080_1082, w_080_1083, w_080_1084, w_080_1085, w_080_1086, w_080_1089, w_080_1091, w_080_1094, w_080_1096, w_080_1097, w_080_1098, w_080_1101, w_080_1102, w_080_1106, w_080_1107, w_080_1110, w_080_1113, w_080_1114, w_080_1115, w_080_1116, w_080_1118, w_080_1119, w_080_1121, w_080_1122, w_080_1123, w_080_1126, w_080_1127, w_080_1129, w_080_1131, w_080_1132, w_080_1134, w_080_1137, w_080_1138, w_080_1139, w_080_1140, w_080_1141, w_080_1142, w_080_1144, w_080_1146, w_080_1147, w_080_1149, w_080_1150, w_080_1151, w_080_1152, w_080_1153, w_080_1155, w_080_1156, w_080_1157, w_080_1160, w_080_1161, w_080_1162, w_080_1163, w_080_1166, w_080_1171, w_080_1172, w_080_1176, w_080_1177, w_080_1179, w_080_1180, w_080_1181, w_080_1182, w_080_1183, w_080_1185, w_080_1187, w_080_1188, w_080_1189, w_080_1190, w_080_1192, w_080_1193, w_080_1194, w_080_1197, w_080_1198, w_080_1199, w_080_1203, w_080_1205, w_080_1207, w_080_1209, w_080_1211, w_080_1212, w_080_1213, w_080_1215, w_080_1216, w_080_1217, w_080_1219, w_080_1221, w_080_1222, w_080_1224, w_080_1226, w_080_1228, w_080_1231, w_080_1233, w_080_1236, w_080_1237, w_080_1240, w_080_1241, w_080_1243, w_080_1244, w_080_1246, w_080_1247, w_080_1248, w_080_1254, w_080_1256, w_080_1259, w_080_1260, w_080_1261, w_080_1262, w_080_1263, w_080_1264, w_080_1265, w_080_1266, w_080_1270, w_080_1271, w_080_1272, w_080_1273, w_080_1274, w_080_1276, w_080_1277, w_080_1278, w_080_1279, w_080_1280, w_080_1282, w_080_1283, w_080_1284, w_080_1287, w_080_1288, w_080_1289, w_080_1290, w_080_1291, w_080_1294, w_080_1295, w_080_1297, w_080_1298, w_080_1299, w_080_1300, w_080_1302, w_080_1303, w_080_1307, w_080_1308, w_080_1309, w_080_1312, w_080_1314, w_080_1315, w_080_1319, w_080_1320, w_080_1322, w_080_1323, w_080_1324, w_080_1325, w_080_1327, w_080_1328, w_080_1330, w_080_1331, w_080_1333, w_080_1334, w_080_1337, w_080_1339, w_080_1341, w_080_1342, w_080_1343, w_080_1349, w_080_1350, w_080_1351, w_080_1353, w_080_1355, w_080_1356, w_080_1358, w_080_1359, w_080_1360, w_080_1362, w_080_1364, w_080_1365, w_080_1366, w_080_1367, w_080_1369, w_080_1371, w_080_1375, w_080_1376, w_080_1378, w_080_1379, w_080_1380, w_080_1382, w_080_1384, w_080_1386, w_080_1387, w_080_1388, w_080_1389, w_080_1392, w_080_1396, w_080_1397, w_080_1398, w_080_1399, w_080_1400, w_080_1401, w_080_1403, w_080_1404, w_080_1406, w_080_1408, w_080_1415, w_080_1416, w_080_1417, w_080_1418, w_080_1419, w_080_1421, w_080_1422, w_080_1427, w_080_1429, w_080_1430, w_080_1431, w_080_1433, w_080_1434, w_080_1435, w_080_1437, w_080_1439, w_080_1440, w_080_1441, w_080_1443, w_080_1444, w_080_1446, w_080_1447, w_080_1448, w_080_1449, w_080_1451, w_080_1458, w_080_1461, w_080_1462, w_080_1467, w_080_1470, w_080_1471, w_080_1472, w_080_1473, w_080_1474, w_080_1476, w_080_1479, w_080_1481, w_080_1488, w_080_1491, w_080_1493, w_080_1494, w_080_1504, w_080_1508, w_080_1509, w_080_1512, w_080_1516, w_080_1518, w_080_1521, w_080_1523, w_080_1525, w_080_1526, w_080_1538, w_080_1539, w_080_1543, w_080_1547, w_080_1551, w_080_1552, w_080_1555, w_080_1556, w_080_1559, w_080_1563, w_080_1566, w_080_1569, w_080_1571, w_080_1574, w_080_1580, w_080_1581, w_080_1585, w_080_1587, w_080_1596, w_080_1601, w_080_1603, w_080_1605, w_080_1607, w_080_1608, w_080_1610, w_080_1613, w_080_1617, w_080_1621, w_080_1622, w_080_1632, w_080_1640, w_080_1642, w_080_1643, w_080_1648, w_080_1651, w_080_1654, w_080_1659, w_080_1662, w_080_1664, w_080_1665, w_080_1669, w_080_1671, w_080_1672, w_080_1673, w_080_1675, w_080_1678, w_080_1685, w_080_1686, w_080_1688, w_080_1689, w_080_1699, w_080_1703, w_080_1706, w_080_1707, w_080_1711, w_080_1712, w_080_1714, w_080_1715, w_080_1717, w_080_1718, w_080_1720, w_080_1721, w_080_1727, w_080_1730, w_080_1732, w_080_1738, w_080_1739, w_080_1740, w_080_1743, w_080_1747, w_080_1751, w_080_1752, w_080_1757, w_080_1761, w_080_1763, w_080_1764, w_080_1765, w_080_1768, w_080_1771, w_080_1772, w_080_1775, w_080_1776, w_080_1778, w_080_1780, w_080_1783, w_080_1789, w_080_1791, w_080_1794, w_080_1796, w_080_1799, w_080_1803, w_080_1805, w_080_1806, w_080_1815, w_080_1817, w_080_1824, w_080_1825, w_080_1827, w_080_1828, w_080_1830, w_080_1835, w_080_1836, w_080_1837, w_080_1838, w_080_1846, w_080_1848, w_080_1860, w_080_1868, w_080_1874, w_080_1875, w_080_1877, w_080_1882, w_080_1889, w_080_1890, w_080_1892, w_080_1893, w_080_1894, w_080_1895, w_080_1896, w_080_1898, w_080_1899, w_080_1901, w_080_1903, w_080_1910, w_080_1912, w_080_1918, w_080_1922, w_080_1926, w_080_1930, w_080_1933, w_080_1936, w_080_1937, w_080_1940, w_080_1941, w_080_1942, w_080_1944, w_080_1945, w_080_1946, w_080_1948, w_080_1957, w_080_1958, w_080_1960, w_080_1966, w_080_1968, w_080_1969, w_080_1970, w_080_1971, w_080_1973, w_080_1974, w_080_1977, w_080_1979, w_080_1993, w_080_1994, w_080_1995, w_080_1996, w_080_1999, w_080_2000, w_080_2001, w_080_2003, w_080_2009, w_080_2010, w_080_2014, w_080_2018, w_080_2025, w_080_2030, w_080_2033, w_080_2034, w_080_2035, w_080_2041, w_080_2042, w_080_2045, w_080_2047, w_080_2051, w_080_2052, w_080_2059, w_080_2060, w_080_2062, w_080_2064, w_080_2066, w_080_2067, w_080_2068, w_080_2071, w_080_2072, w_080_2075, w_080_2078, w_080_2080, w_080_2091, w_080_2094, w_080_2095, w_080_2096, w_080_2102, w_080_2107, w_080_2110, w_080_2112, w_080_2115, w_080_2117, w_080_2120, w_080_2121, w_080_2126, w_080_2136, w_080_2137, w_080_2144, w_080_2145, w_080_2146, w_080_2149, w_080_2157, w_080_2162, w_080_2164, w_080_2167, w_080_2168, w_080_2172, w_080_2178, w_080_2180, w_080_2184, w_080_2189, w_080_2191, w_080_2193, w_080_2197, w_080_2204, w_080_2206, w_080_2207, w_080_2212, w_080_2213, w_080_2218, w_080_2220, w_080_2223, w_080_2227, w_080_2228, w_080_2229, w_080_2230, w_080_2235, w_080_2236, w_080_2237, w_080_2238, w_080_2240, w_080_2241, w_080_2250, w_080_2255, w_080_2257, w_080_2266, w_080_2268, w_080_2272, w_080_2274, w_080_2277, w_080_2278, w_080_2280, w_080_2283, w_080_2284, w_080_2289, w_080_2293, w_080_2297, w_080_2298, w_080_2302, w_080_2305, w_080_2307, w_080_2310, w_080_2312, w_080_2314, w_080_2316, w_080_2318, w_080_2320, w_080_2321, w_080_2327, w_080_2335, w_080_2336, w_080_2338, w_080_2341, w_080_2342, w_080_2344, w_080_2346, w_080_2352, w_080_2353, w_080_2355, w_080_2359, w_080_2360, w_080_2364, w_080_2365, w_080_2366, w_080_2369, w_080_2371, w_080_2372, w_080_2373, w_080_2379, w_080_2396, w_080_2398, w_080_2399, w_080_2401, w_080_2403, w_080_2404, w_080_2406, w_080_2411, w_080_2413, w_080_2415, w_080_2418, w_080_2419, w_080_2420, w_080_2424, w_080_2426, w_080_2428, w_080_2435, w_080_2436, w_080_2437, w_080_2438, w_080_2439, w_080_2442, w_080_2443, w_080_2450, w_080_2452, w_080_2457, w_080_2460, w_080_2466, w_080_2467, w_080_2470, w_080_2476, w_080_2479, w_080_2483, w_080_2485, w_080_2487, w_080_2488, w_080_2491, w_080_2492, w_080_2494, w_080_2495, w_080_2497, w_080_2501, w_080_2502, w_080_2507, w_080_2509, w_080_2511, w_080_2517, w_080_2518, w_080_2520, w_080_2522, w_080_2527, w_080_2534, w_080_2535, w_080_2536, w_080_2537, w_080_2552, w_080_2553, w_080_2554, w_080_2556, w_080_2560, w_080_2563, w_080_2567, w_080_2568, w_080_2569, w_080_2570, w_080_2574, w_080_2576, w_080_2578, w_080_2579, w_080_2580, w_080_2587, w_080_2591, w_080_2601, w_080_2605, w_080_2610, w_080_2611, w_080_2621, w_080_2622, w_080_2626, w_080_2627, w_080_2629, w_080_2631, w_080_2640, w_080_2642, w_080_2646, w_080_2648, w_080_2650, w_080_2651, w_080_2652, w_080_2654, w_080_2659, w_080_2662, w_080_2664, w_080_2668, w_080_2669, w_080_2672, w_080_2674, w_080_2675, w_080_2679, w_080_2681, w_080_2682, w_080_2687, w_080_2690, w_080_2691, w_080_2692, w_080_2696, w_080_2705, w_080_2706, w_080_2707, w_080_2708, w_080_2712, w_080_2719, w_080_2722, w_080_2724, w_080_2725, w_080_2727, w_080_2731, w_080_2732, w_080_2735, w_080_2738, w_080_2739, w_080_2740, w_080_2743, w_080_2750, w_080_2751, w_080_2754, w_080_2758, w_080_2759, w_080_2761, w_080_2764, w_080_2767, w_080_2770, w_080_2772, w_080_2777, w_080_2778, w_080_2779, w_080_2780, w_080_2782, w_080_2788, w_080_2795, w_080_2797, w_080_2799, w_080_2805, w_080_2810, w_080_2811, w_080_2814, w_080_2819, w_080_2827, w_080_2829, w_080_2830, w_080_2831, w_080_2833, w_080_2834, w_080_2837, w_080_2839, w_080_2843, w_080_2846, w_080_2850, w_080_2851, w_080_2853, w_080_2855, w_080_2857, w_080_2862, w_080_2864, w_080_2867, w_080_2870, w_080_2874, w_080_2875, w_080_2882, w_080_2886, w_080_2895, w_080_2896, w_080_2897, w_080_2898, w_080_2899, w_080_2905, w_080_2908, w_080_2915, w_080_2916, w_080_2920, w_080_2921, w_080_2926, w_080_2929, w_080_2932, w_080_2934, w_080_2936, w_080_2939, w_080_2943, w_080_2945, w_080_2946, w_080_2949, w_080_2952, w_080_2956, w_080_2962, w_080_2966, w_080_2969, w_080_2971, w_080_2975, w_080_2980, w_080_2981, w_080_2982, w_080_2985, w_080_2986, w_080_2995, w_080_2996, w_080_2999, w_080_3001, w_080_3003, w_080_3005, w_080_3007, w_080_3008, w_080_3010, w_080_3015, w_080_3017, w_080_3018, w_080_3022, w_080_3025, w_080_3026, w_080_3028, w_080_3031, w_080_3033, w_080_3034, w_080_3036, w_080_3038, w_080_3039, w_080_3041, w_080_3044, w_080_3045, w_080_3051, w_080_3052, w_080_3059, w_080_3061, w_080_3062, w_080_3065, w_080_3069, w_080_3073, w_080_3075, w_080_3080, w_080_3081, w_080_3083, w_080_3085, w_080_3088, w_080_3096, w_080_3102, w_080_3105, w_080_3107, w_080_3108, w_080_3110, w_080_3114, w_080_3115, w_080_3122, w_080_3123, w_080_3124, w_080_3125, w_080_3127, w_080_3134, w_080_3137, w_080_3145, w_080_3147, w_080_3148, w_080_3152, w_080_3161, w_080_3164, w_080_3166, w_080_3169, w_080_3182, w_080_3185, w_080_3187, w_080_3192, w_080_3202, w_080_3203, w_080_3207, w_080_3211, w_080_3213, w_080_3216, w_080_3218, w_080_3221, w_080_3225, w_080_3228, w_080_3229, w_080_3231, w_080_3232, w_080_3235, w_080_3238, w_080_3239, w_080_3242, w_080_3246, w_080_3250, w_080_3254, w_080_3255, w_080_3258, w_080_3279, w_080_3281, w_080_3283, w_080_3284, w_080_3287, w_080_3288, w_080_3290, w_080_3296, w_080_3300, w_080_3304, w_080_3307, w_080_3310, w_080_3311, w_080_3316, w_080_3318, w_080_3320, w_080_3332, w_080_3335, w_080_3336, w_080_3338, w_080_3339, w_080_3340, w_080_3343, w_080_3346, w_080_3348, w_080_3349, w_080_3350, w_080_3351, w_080_3352, w_080_3353, w_080_3355, w_080_3380, w_080_3382, w_080_3383, w_080_3384, w_080_3385, w_080_3386, w_080_3393, w_080_3396, w_080_3397, w_080_3398, w_080_3407, w_080_3418, w_080_3432, w_080_3433, w_080_3434, w_080_3436, w_080_3438, w_080_3439, w_080_3440, w_080_3441, w_080_3442, w_080_3443, w_080_3447, w_080_3448, w_080_3452, w_080_3457, w_080_3465, w_080_3467, w_080_3473, w_080_3476, w_080_3477, w_080_3483, w_080_3485, w_080_3490, w_080_3493, w_080_3500, w_080_3502, w_080_3503, w_080_3506, w_080_3507, w_080_3508, w_080_3512, w_080_3513, w_080_3514, w_080_3517, w_080_3518, w_080_3519, w_080_3520, w_080_3521, w_080_3522, w_080_3523, w_080_3525, w_080_3527, w_080_3528, w_080_3529, w_080_3530, w_080_3531, w_080_3532, w_080_3534;
  wire w_081_000, w_081_001, w_081_002, w_081_003, w_081_004, w_081_005, w_081_006, w_081_007, w_081_009, w_081_010, w_081_011, w_081_012, w_081_013, w_081_014, w_081_015, w_081_016, w_081_018, w_081_019, w_081_020, w_081_021, w_081_022, w_081_023, w_081_025, w_081_026, w_081_027, w_081_028, w_081_030, w_081_031, w_081_033, w_081_034, w_081_035, w_081_037, w_081_038, w_081_039, w_081_040, w_081_042, w_081_044, w_081_045, w_081_046, w_081_047, w_081_049, w_081_050, w_081_052, w_081_053, w_081_054, w_081_057, w_081_058, w_081_059, w_081_060, w_081_061, w_081_062, w_081_063, w_081_066, w_081_067, w_081_069, w_081_071, w_081_072, w_081_073, w_081_074, w_081_075, w_081_076, w_081_077, w_081_078, w_081_079, w_081_081, w_081_082, w_081_083, w_081_084, w_081_085, w_081_086, w_081_089, w_081_091, w_081_092, w_081_093, w_081_094, w_081_095, w_081_096, w_081_097, w_081_100, w_081_101, w_081_103, w_081_104, w_081_105, w_081_106, w_081_107, w_081_108, w_081_110, w_081_111, w_081_112, w_081_113, w_081_115, w_081_116, w_081_117, w_081_119, w_081_120, w_081_121, w_081_122, w_081_125, w_081_126, w_081_127, w_081_129, w_081_130, w_081_131, w_081_132, w_081_133, w_081_134, w_081_135, w_081_136, w_081_138, w_081_139, w_081_141, w_081_144, w_081_145, w_081_146, w_081_147, w_081_151, w_081_152, w_081_153, w_081_154, w_081_155, w_081_156, w_081_157, w_081_158, w_081_159, w_081_161, w_081_162, w_081_164, w_081_165, w_081_166, w_081_167, w_081_168, w_081_171, w_081_172, w_081_173, w_081_174, w_081_175, w_081_176, w_081_177, w_081_178, w_081_179, w_081_180, w_081_181, w_081_182, w_081_183, w_081_188, w_081_189, w_081_190, w_081_192, w_081_193, w_081_194, w_081_196, w_081_197, w_081_198, w_081_199, w_081_200, w_081_202, w_081_203, w_081_204, w_081_205, w_081_206, w_081_207, w_081_209, w_081_210, w_081_211, w_081_212, w_081_213, w_081_214, w_081_216, w_081_217, w_081_219, w_081_220, w_081_221, w_081_222, w_081_223, w_081_224, w_081_226, w_081_227, w_081_228, w_081_229, w_081_230, w_081_231, w_081_232, w_081_233, w_081_236, w_081_237, w_081_238, w_081_239, w_081_240, w_081_241, w_081_242, w_081_244, w_081_245, w_081_246, w_081_247, w_081_249, w_081_251, w_081_254, w_081_255, w_081_256, w_081_257, w_081_258, w_081_259, w_081_261, w_081_263, w_081_265, w_081_266, w_081_267, w_081_268, w_081_269, w_081_270, w_081_271, w_081_272, w_081_273, w_081_274, w_081_275, w_081_276, w_081_277, w_081_280, w_081_281, w_081_282, w_081_283, w_081_284, w_081_285, w_081_286, w_081_287, w_081_288, w_081_289, w_081_290, w_081_291, w_081_292, w_081_293, w_081_294, w_081_295, w_081_296, w_081_298, w_081_299, w_081_300, w_081_301, w_081_302, w_081_307, w_081_309, w_081_310, w_081_311, w_081_312, w_081_313, w_081_314, w_081_315, w_081_317, w_081_318, w_081_319, w_081_320, w_081_321, w_081_322, w_081_323, w_081_325, w_081_326, w_081_327, w_081_329, w_081_330, w_081_331, w_081_332, w_081_333, w_081_335, w_081_336, w_081_337, w_081_340, w_081_342, w_081_343, w_081_344, w_081_345, w_081_347, w_081_349, w_081_350, w_081_351, w_081_352, w_081_354, w_081_355, w_081_357, w_081_358, w_081_362, w_081_364, w_081_365, w_081_366, w_081_367, w_081_368, w_081_369, w_081_370, w_081_371, w_081_372, w_081_373, w_081_374, w_081_376, w_081_377, w_081_379, w_081_380, w_081_381, w_081_382, w_081_383, w_081_386, w_081_387, w_081_389, w_081_390, w_081_391, w_081_392, w_081_393, w_081_394, w_081_395, w_081_396, w_081_397, w_081_399, w_081_400, w_081_401, w_081_402, w_081_403, w_081_405, w_081_406, w_081_407, w_081_408, w_081_410, w_081_412, w_081_413, w_081_414, w_081_415, w_081_416, w_081_418, w_081_419, w_081_420, w_081_422, w_081_423, w_081_424, w_081_425, w_081_426, w_081_427, w_081_429, w_081_430, w_081_431, w_081_432, w_081_433, w_081_434, w_081_435, w_081_436, w_081_438, w_081_439, w_081_440, w_081_441, w_081_442, w_081_444, w_081_445, w_081_447, w_081_448, w_081_450, w_081_451, w_081_452, w_081_453, w_081_454, w_081_455, w_081_456, w_081_457, w_081_458, w_081_459, w_081_460, w_081_461, w_081_462, w_081_463, w_081_464, w_081_466, w_081_467, w_081_468, w_081_469, w_081_470, w_081_471, w_081_472, w_081_474, w_081_475, w_081_476, w_081_477, w_081_478, w_081_479, w_081_480, w_081_481, w_081_482, w_081_483, w_081_484, w_081_485, w_081_486, w_081_487, w_081_488, w_081_489, w_081_490, w_081_491, w_081_492, w_081_493, w_081_494, w_081_495, w_081_496, w_081_497, w_081_498, w_081_499, w_081_501, w_081_502, w_081_503, w_081_504, w_081_507, w_081_508, w_081_509, w_081_510, w_081_511, w_081_512, w_081_513, w_081_514, w_081_515, w_081_516, w_081_517, w_081_520, w_081_521, w_081_522, w_081_523, w_081_524, w_081_526, w_081_527, w_081_529, w_081_530, w_081_531, w_081_532, w_081_533, w_081_534, w_081_535, w_081_537, w_081_538, w_081_539, w_081_540, w_081_542, w_081_543, w_081_544, w_081_545, w_081_547, w_081_548, w_081_549, w_081_550, w_081_551, w_081_552, w_081_553, w_081_555, w_081_556, w_081_557, w_081_558, w_081_559, w_081_560, w_081_562, w_081_563, w_081_565, w_081_566, w_081_567, w_081_569, w_081_570, w_081_572, w_081_573, w_081_574, w_081_575, w_081_576, w_081_577, w_081_578, w_081_579, w_081_580, w_081_581, w_081_582, w_081_583, w_081_587, w_081_588, w_081_590, w_081_591, w_081_594, w_081_595, w_081_596, w_081_597, w_081_598, w_081_599, w_081_600, w_081_602, w_081_603, w_081_604, w_081_605, w_081_606, w_081_607, w_081_609, w_081_611, w_081_612, w_081_613, w_081_615, w_081_616, w_081_617, w_081_618, w_081_619, w_081_620, w_081_621, w_081_624, w_081_626, w_081_627, w_081_628, w_081_629, w_081_630, w_081_631, w_081_632, w_081_633, w_081_635, w_081_636, w_081_638, w_081_640, w_081_641, w_081_642, w_081_644, w_081_645, w_081_647, w_081_648, w_081_649, w_081_650, w_081_651, w_081_652, w_081_654, w_081_655, w_081_656, w_081_657, w_081_658, w_081_659, w_081_660, w_081_662, w_081_663, w_081_664, w_081_665, w_081_667, w_081_668, w_081_669, w_081_670, w_081_671, w_081_672, w_081_673, w_081_674, w_081_675, w_081_676, w_081_677, w_081_678, w_081_679, w_081_680, w_081_681, w_081_682, w_081_683, w_081_685, w_081_686, w_081_687, w_081_688, w_081_689, w_081_690, w_081_691, w_081_692, w_081_693, w_081_694, w_081_695, w_081_698, w_081_699, w_081_704, w_081_705, w_081_706, w_081_708, w_081_709, w_081_710, w_081_711, w_081_712, w_081_713, w_081_714, w_081_715, w_081_716, w_081_717, w_081_718, w_081_719, w_081_720, w_081_721, w_081_724, w_081_725, w_081_726, w_081_728, w_081_729, w_081_730, w_081_731, w_081_732, w_081_733, w_081_734, w_081_736, w_081_737, w_081_738, w_081_739, w_081_740, w_081_741, w_081_742, w_081_743, w_081_744, w_081_746, w_081_747, w_081_748, w_081_749, w_081_750, w_081_751, w_081_752, w_081_753, w_081_754, w_081_755, w_081_756, w_081_757, w_081_758, w_081_759, w_081_761, w_081_762, w_081_763, w_081_764, w_081_766, w_081_767, w_081_771, w_081_772, w_081_774, w_081_775, w_081_777, w_081_778, w_081_779, w_081_780, w_081_781, w_081_782, w_081_784, w_081_785, w_081_786, w_081_787, w_081_788, w_081_789, w_081_792, w_081_794, w_081_795, w_081_796, w_081_797, w_081_798, w_081_799, w_081_800, w_081_801, w_081_802, w_081_804, w_081_805, w_081_807, w_081_808, w_081_809, w_081_812, w_081_813, w_081_814, w_081_815, w_081_816, w_081_817, w_081_818, w_081_819, w_081_820, w_081_822, w_081_823, w_081_825, w_081_826, w_081_827, w_081_829, w_081_830, w_081_831, w_081_832, w_081_833, w_081_834, w_081_836, w_081_837, w_081_838, w_081_841, w_081_842, w_081_843, w_081_844, w_081_846, w_081_848, w_081_850, w_081_852, w_081_853, w_081_854, w_081_855, w_081_856, w_081_857, w_081_858, w_081_859, w_081_860, w_081_861, w_081_862, w_081_863, w_081_864, w_081_866, w_081_868, w_081_869, w_081_870, w_081_871, w_081_872, w_081_873, w_081_874, w_081_875, w_081_876, w_081_878, w_081_879, w_081_880, w_081_881, w_081_882, w_081_883, w_081_884, w_081_885, w_081_886, w_081_889, w_081_890, w_081_891, w_081_892, w_081_893, w_081_894, w_081_895, w_081_896, w_081_897, w_081_898, w_081_899, w_081_901, w_081_902, w_081_904, w_081_905, w_081_906, w_081_907, w_081_908, w_081_909, w_081_910, w_081_911, w_081_912, w_081_913, w_081_914, w_081_915, w_081_916, w_081_917, w_081_918, w_081_919, w_081_921, w_081_922, w_081_923, w_081_924, w_081_925, w_081_926, w_081_927, w_081_928, w_081_929, w_081_930, w_081_931, w_081_932, w_081_933, w_081_935, w_081_936, w_081_937, w_081_938, w_081_939, w_081_942, w_081_945, w_081_946, w_081_947, w_081_951, w_081_952, w_081_953, w_081_954, w_081_955, w_081_956, w_081_957, w_081_958, w_081_960, w_081_961, w_081_962, w_081_964, w_081_965, w_081_966, w_081_967, w_081_968, w_081_969, w_081_970, w_081_973, w_081_975, w_081_976, w_081_977, w_081_978, w_081_979, w_081_981, w_081_983, w_081_984, w_081_985, w_081_987, w_081_988, w_081_989, w_081_993, w_081_996, w_081_998, w_081_1000, w_081_1001, w_081_1003, w_081_1004, w_081_1005, w_081_1006, w_081_1007, w_081_1008, w_081_1009, w_081_1010, w_081_1011, w_081_1012, w_081_1014, w_081_1015, w_081_1017, w_081_1018, w_081_1021, w_081_1022, w_081_1026, w_081_1027, w_081_1029, w_081_1030, w_081_1031, w_081_1033, w_081_1034, w_081_1037, w_081_1038, w_081_1039, w_081_1040, w_081_1041, w_081_1043, w_081_1044, w_081_1045, w_081_1046, w_081_1047, w_081_1048, w_081_1049, w_081_1050, w_081_1051, w_081_1053, w_081_1054, w_081_1056, w_081_1057, w_081_1059, w_081_1061, w_081_1062, w_081_1063, w_081_1064, w_081_1065, w_081_1066, w_081_1068, w_081_1070, w_081_1072, w_081_1073, w_081_1074, w_081_1075, w_081_1077, w_081_1079, w_081_1081, w_081_1082, w_081_1083, w_081_1084, w_081_1085, w_081_1086, w_081_1088, w_081_1090, w_081_1091, w_081_1092, w_081_1094, w_081_1095, w_081_1096, w_081_1097, w_081_1100, w_081_1102, w_081_1103, w_081_1104, w_081_1106, w_081_1109, w_081_1110, w_081_1111, w_081_1112, w_081_1115, w_081_1116, w_081_1117, w_081_1118, w_081_1119, w_081_1120, w_081_1121, w_081_1122, w_081_1123, w_081_1124, w_081_1125, w_081_1126, w_081_1127, w_081_1129, w_081_1130, w_081_1131, w_081_1134, w_081_1135, w_081_1136, w_081_1137, w_081_1138, w_081_1139, w_081_1140, w_081_1142, w_081_1143, w_081_1146, w_081_1147, w_081_1148, w_081_1149, w_081_1150, w_081_1151, w_081_1152, w_081_1153, w_081_1154, w_081_1155, w_081_1158, w_081_1159, w_081_1164, w_081_1165, w_081_1167, w_081_1168, w_081_1169, w_081_1170, w_081_1171, w_081_1173, w_081_1174, w_081_1176, w_081_1177, w_081_1178, w_081_1179, w_081_1180, w_081_1181, w_081_1182, w_081_1183, w_081_1184, w_081_1185, w_081_1187, w_081_1189, w_081_1191, w_081_1193, w_081_1195, w_081_1197, w_081_1199, w_081_1201, w_081_1202, w_081_1203, w_081_1204, w_081_1208, w_081_1209, w_081_1210, w_081_1211, w_081_1212, w_081_1214, w_081_1215, w_081_1216, w_081_1218, w_081_1220, w_081_1222, w_081_1224, w_081_1226, w_081_1227, w_081_1228, w_081_1230, w_081_1231, w_081_1234, w_081_1236, w_081_1237, w_081_1240, w_081_1241, w_081_1246, w_081_1247, w_081_1248, w_081_1250, w_081_1251, w_081_1252, w_081_1253, w_081_1254, w_081_1255, w_081_1256, w_081_1257, w_081_1261, w_081_1263, w_081_1264, w_081_1265, w_081_1266, w_081_1267, w_081_1269, w_081_1271, w_081_1272, w_081_1276, w_081_1277, w_081_1278, w_081_1279, w_081_1283, w_081_1285, w_081_1287, w_081_1288, w_081_1289, w_081_1290, w_081_1291, w_081_1292, w_081_1295, w_081_1296, w_081_1297, w_081_1301, w_081_1302, w_081_1305, w_081_1306, w_081_1307, w_081_1308, w_081_1310, w_081_1311, w_081_1313, w_081_1314, w_081_1315, w_081_1316, w_081_1317, w_081_1318, w_081_1319, w_081_1322, w_081_1325, w_081_1326, w_081_1328, w_081_1329, w_081_1330, w_081_1332, w_081_1334, w_081_1335, w_081_1336, w_081_1337, w_081_1339, w_081_1340, w_081_1341, w_081_1342, w_081_1343;
  wire w_082_000, w_082_001, w_082_002, w_082_004, w_082_005, w_082_006, w_082_007, w_082_008, w_082_009, w_082_010, w_082_011, w_082_012, w_082_013, w_082_014, w_082_015, w_082_016, w_082_017, w_082_018, w_082_019, w_082_021, w_082_022, w_082_024, w_082_025, w_082_026, w_082_027, w_082_028, w_082_029, w_082_030, w_082_031, w_082_032, w_082_033, w_082_035, w_082_037, w_082_039, w_082_040, w_082_041, w_082_042, w_082_043, w_082_045, w_082_046, w_082_047, w_082_048, w_082_049, w_082_050, w_082_051, w_082_052, w_082_054, w_082_055, w_082_056, w_082_057, w_082_058, w_082_059, w_082_060, w_082_061, w_082_062, w_082_063, w_082_064, w_082_065, w_082_066, w_082_067, w_082_068, w_082_069, w_082_070, w_082_071, w_082_072, w_082_073, w_082_074, w_082_075, w_082_076, w_082_077, w_082_078, w_082_079, w_082_081, w_082_082, w_082_084, w_082_085, w_082_086, w_082_087, w_082_088, w_082_089, w_082_090, w_082_091, w_082_092, w_082_093, w_082_094, w_082_095, w_082_096, w_082_097, w_082_098, w_082_099, w_082_100, w_082_101, w_082_102, w_082_104, w_082_105, w_082_106, w_082_107, w_082_108, w_082_109, w_082_110, w_082_113, w_082_114, w_082_115, w_082_116, w_082_117, w_082_118, w_082_119, w_082_120, w_082_121, w_082_122, w_082_123, w_082_124, w_082_125, w_082_126, w_082_127, w_082_128, w_082_129, w_082_130, w_082_131, w_082_132, w_082_133, w_082_134, w_082_135, w_082_136, w_082_137, w_082_138, w_082_139, w_082_140, w_082_141, w_082_142, w_082_143, w_082_144, w_082_145, w_082_146, w_082_147, w_082_149, w_082_150, w_082_151, w_082_152, w_082_153, w_082_154, w_082_155, w_082_157, w_082_158, w_082_159, w_082_160, w_082_161, w_082_162, w_082_163, w_082_164, w_082_165, w_082_166, w_082_167, w_082_168, w_082_169, w_082_170, w_082_171, w_082_172, w_082_173, w_082_174, w_082_175, w_082_177, w_082_178, w_082_179, w_082_180, w_082_181, w_082_182, w_082_183, w_082_185, w_082_186, w_082_187, w_082_188, w_082_189, w_082_190, w_082_191, w_082_192, w_082_193, w_082_194, w_082_195, w_082_196, w_082_197, w_082_198, w_082_199, w_082_200, w_082_201, w_082_202, w_082_203, w_082_205, w_082_207, w_082_209, w_082_210, w_082_211, w_082_212, w_082_213, w_082_214, w_082_215, w_082_216, w_082_218, w_082_219, w_082_220, w_082_221, w_082_222, w_082_223, w_082_224, w_082_225, w_082_226, w_082_229, w_082_230, w_082_231, w_082_232, w_082_233, w_082_234, w_082_235, w_082_236, w_082_237, w_082_238, w_082_239, w_082_240, w_082_241, w_082_242, w_082_243, w_082_244, w_082_245, w_082_246, w_082_247, w_082_248, w_082_249, w_082_250, w_082_251, w_082_252, w_082_253, w_082_254, w_082_255, w_082_257, w_082_258, w_082_259, w_082_260, w_082_261, w_082_262, w_082_263, w_082_264, w_082_265, w_082_266, w_082_267, w_082_268, w_082_269, w_082_270, w_082_271, w_082_272, w_082_273, w_082_274, w_082_275, w_082_276, w_082_277, w_082_279, w_082_280, w_082_281, w_082_282, w_082_283, w_082_284, w_082_285, w_082_286, w_082_289, w_082_290, w_082_291, w_082_292, w_082_293, w_082_294, w_082_295, w_082_296, w_082_297, w_082_298, w_082_299, w_082_300, w_082_301, w_082_302, w_082_303, w_082_304, w_082_305, w_082_306, w_082_307, w_082_309, w_082_310, w_082_311, w_082_312, w_082_313, w_082_314, w_082_315, w_082_317, w_082_318, w_082_319, w_082_320, w_082_321, w_082_322, w_082_323, w_082_324, w_082_325, w_082_326, w_082_328, w_082_329, w_082_330, w_082_331, w_082_332, w_082_333, w_082_334, w_082_335, w_082_336, w_082_337, w_082_338, w_082_339, w_082_340, w_082_341, w_082_343, w_082_344, w_082_345, w_082_346, w_082_347, w_082_348, w_082_349, w_082_350, w_082_351, w_082_352, w_082_353, w_082_354, w_082_356, w_082_357, w_082_359, w_082_360, w_082_361, w_082_362, w_082_363, w_082_364, w_082_365, w_082_366, w_082_367, w_082_368, w_082_370, w_082_371, w_082_372, w_082_373, w_082_374, w_082_375, w_082_376, w_082_377, w_082_378, w_082_379, w_082_380, w_082_382, w_082_383, w_082_384, w_082_385, w_082_386, w_082_387, w_082_388, w_082_389, w_082_390, w_082_391, w_082_392, w_082_393, w_082_395, w_082_396, w_082_397, w_082_399, w_082_400, w_082_401, w_082_402, w_082_403, w_082_404, w_082_405, w_082_407, w_082_411, w_082_412, w_082_413, w_082_414, w_082_415, w_082_417, w_082_418, w_082_420, w_082_422, w_082_423, w_082_425, w_082_427, w_082_428, w_082_429, w_082_431, w_082_432, w_082_433, w_082_434, w_082_435, w_082_436, w_082_437, w_082_438, w_082_439, w_082_440, w_082_441, w_082_442, w_082_443, w_082_444, w_082_446, w_082_447, w_082_448, w_082_449, w_082_450, w_082_451, w_082_452, w_082_453, w_082_454, w_082_455, w_082_456, w_082_457, w_082_459, w_082_460, w_082_462, w_082_463, w_082_464, w_082_465, w_082_466, w_082_467, w_082_468, w_082_469, w_082_471, w_082_472, w_082_473, w_082_474, w_082_475, w_082_476, w_082_477, w_082_478, w_082_479, w_082_480, w_082_481, w_082_482, w_082_483, w_082_484, w_082_485, w_082_486, w_082_487, w_082_488, w_082_490, w_082_491, w_082_492, w_082_493, w_082_495, w_082_496, w_082_497, w_082_498, w_082_499, w_082_500, w_082_501, w_082_502, w_082_503, w_082_504, w_082_505, w_082_506, w_082_507, w_082_508, w_082_509, w_082_510, w_082_511, w_082_512, w_082_513, w_082_514, w_082_515, w_082_516, w_082_517, w_082_518, w_082_520, w_082_521, w_082_522, w_082_524, w_082_525, w_082_526, w_082_527, w_082_528, w_082_529, w_082_530, w_082_531, w_082_532, w_082_533, w_082_536, w_082_537, w_082_538, w_082_539, w_082_540, w_082_541, w_082_542, w_082_543, w_082_544, w_082_545, w_082_546, w_082_547, w_082_548, w_082_549, w_082_551, w_082_552, w_082_553, w_082_554, w_082_555, w_082_556, w_082_557, w_082_558, w_082_559, w_082_561, w_082_562, w_082_563, w_082_564, w_082_565, w_082_566, w_082_568, w_082_569, w_082_570, w_082_571, w_082_572, w_082_573, w_082_574, w_082_575, w_082_576, w_082_577, w_082_578, w_082_579, w_082_580, w_082_581, w_082_582, w_082_583, w_082_584, w_082_585, w_082_586, w_082_588, w_082_589, w_082_590, w_082_592, w_082_593, w_082_594, w_082_595, w_082_596, w_082_597, w_082_598, w_082_599, w_082_600, w_082_601, w_082_602, w_082_603, w_082_604, w_082_605, w_082_606, w_082_608, w_082_611, w_082_612, w_082_613, w_082_614, w_082_615, w_082_617, w_082_618, w_082_619, w_082_620, w_082_621, w_082_623, w_082_624, w_082_625, w_082_626, w_082_627, w_082_628, w_082_630, w_082_631, w_082_632, w_082_633, w_082_634, w_082_636, w_082_637, w_082_638, w_082_639, w_082_640, w_082_642, w_082_643, w_082_644, w_082_645, w_082_646, w_082_647, w_082_648, w_082_650, w_082_651, w_082_652, w_082_653, w_082_654, w_082_655, w_082_656, w_082_657, w_082_658, w_082_659, w_082_660, w_082_661, w_082_662, w_082_663, w_082_664, w_082_665, w_082_667, w_082_668, w_082_669, w_082_670, w_082_671, w_082_672, w_082_673, w_082_674, w_082_675, w_082_676, w_082_677, w_082_678, w_082_679, w_082_680, w_082_681, w_082_682, w_082_684, w_082_685, w_082_686, w_082_687, w_082_688, w_082_689, w_082_690, w_082_691, w_082_692, w_082_694, w_082_695, w_082_696, w_082_697, w_082_698, w_082_700, w_082_701, w_082_702, w_082_703, w_082_704, w_082_705, w_082_706, w_082_707, w_082_708, w_082_709, w_082_710, w_082_711, w_082_712, w_082_713, w_082_714, w_082_715, w_082_716, w_082_719, w_082_720, w_082_721, w_082_722, w_082_723, w_082_724, w_082_725, w_082_727, w_082_728, w_082_729, w_082_730, w_082_731, w_082_732, w_082_733, w_082_734, w_082_735, w_082_736, w_082_737, w_082_738, w_082_739, w_082_740, w_082_741, w_082_742, w_082_743, w_082_744, w_082_745, w_082_746, w_082_747, w_082_748, w_082_749, w_082_750, w_082_751, w_082_752, w_082_753, w_082_754, w_082_755, w_082_756, w_082_758, w_082_759, w_082_760, w_082_761, w_082_762, w_082_763, w_082_764, w_082_765, w_082_767, w_082_768, w_082_769, w_082_770, w_082_771, w_082_773, w_082_774, w_082_775, w_082_776, w_082_777, w_082_779, w_082_780, w_082_782, w_082_783, w_082_784, w_082_785, w_082_786, w_082_788, w_082_789, w_082_790, w_082_791, w_082_792, w_082_793, w_082_795, w_082_796, w_082_797, w_082_798, w_082_799, w_082_800, w_082_801, w_082_802, w_082_803, w_082_804, w_082_805, w_082_806, w_082_808, w_082_809, w_082_810, w_082_812, w_082_813, w_082_814, w_082_815, w_082_817, w_082_818, w_082_819, w_082_820, w_082_821, w_082_822, w_082_823, w_082_824, w_082_825, w_082_827, w_082_828, w_082_829, w_082_830, w_082_831, w_082_832, w_082_833, w_082_834, w_082_835, w_082_836, w_082_837, w_082_838, w_082_839, w_082_840, w_082_841, w_082_842, w_082_843, w_082_844, w_082_845, w_082_846, w_082_847, w_082_848, w_082_849, w_082_850, w_082_851, w_082_853, w_082_855, w_082_856, w_082_857, w_082_858, w_082_859, w_082_860, w_082_861, w_082_862, w_082_863, w_082_864, w_082_865, w_082_866, w_082_867, w_082_868, w_082_869, w_082_870, w_082_871, w_082_872, w_082_874, w_082_876, w_082_877, w_082_878, w_082_880, w_082_881, w_082_882, w_082_883, w_082_884, w_082_885, w_082_886, w_082_887, w_082_888, w_082_889, w_082_890, w_082_891, w_082_893, w_082_895, w_082_896, w_082_899, w_082_900, w_082_901, w_082_902, w_082_903, w_082_904, w_082_906, w_082_907, w_082_909, w_082_910, w_082_911, w_082_912, w_082_913, w_082_914, w_082_915, w_082_916, w_082_917, w_082_919, w_082_920, w_082_921, w_082_922, w_082_923, w_082_924, w_082_926, w_082_927, w_082_928, w_082_929, w_082_930, w_082_931, w_082_932, w_082_933, w_082_934, w_082_935, w_082_936, w_082_939, w_082_940, w_082_941;
  wire w_083_000, w_083_001, w_083_003, w_083_004, w_083_005, w_083_006, w_083_009, w_083_012, w_083_014, w_083_015, w_083_019, w_083_020, w_083_022, w_083_023, w_083_026, w_083_027, w_083_028, w_083_029, w_083_034, w_083_037, w_083_039, w_083_040, w_083_041, w_083_042, w_083_043, w_083_045, w_083_046, w_083_047, w_083_048, w_083_049, w_083_052, w_083_053, w_083_057, w_083_058, w_083_059, w_083_061, w_083_063, w_083_066, w_083_067, w_083_068, w_083_069, w_083_070, w_083_071, w_083_073, w_083_074, w_083_079, w_083_080, w_083_081, w_083_083, w_083_084, w_083_085, w_083_086, w_083_087, w_083_088, w_083_089, w_083_092, w_083_093, w_083_095, w_083_098, w_083_099, w_083_101, w_083_102, w_083_103, w_083_105, w_083_109, w_083_111, w_083_112, w_083_113, w_083_115, w_083_117, w_083_118, w_083_119, w_083_120, w_083_122, w_083_123, w_083_124, w_083_125, w_083_126, w_083_127, w_083_128, w_083_133, w_083_134, w_083_137, w_083_138, w_083_142, w_083_143, w_083_146, w_083_147, w_083_149, w_083_150, w_083_153, w_083_155, w_083_156, w_083_157, w_083_158, w_083_159, w_083_161, w_083_162, w_083_163, w_083_165, w_083_167, w_083_175, w_083_176, w_083_177, w_083_180, w_083_181, w_083_182, w_083_184, w_083_185, w_083_187, w_083_188, w_083_190, w_083_193, w_083_194, w_083_198, w_083_200, w_083_202, w_083_205, w_083_208, w_083_210, w_083_212, w_083_214, w_083_215, w_083_216, w_083_217, w_083_219, w_083_221, w_083_223, w_083_224, w_083_225, w_083_228, w_083_229, w_083_232, w_083_233, w_083_236, w_083_241, w_083_244, w_083_246, w_083_251, w_083_257, w_083_258, w_083_260, w_083_262, w_083_263, w_083_267, w_083_268, w_083_269, w_083_270, w_083_271, w_083_273, w_083_275, w_083_276, w_083_281, w_083_283, w_083_284, w_083_285, w_083_286, w_083_290, w_083_291, w_083_292, w_083_295, w_083_296, w_083_297, w_083_301, w_083_303, w_083_308, w_083_313, w_083_314, w_083_315, w_083_317, w_083_319, w_083_320, w_083_321, w_083_322, w_083_323, w_083_324, w_083_329, w_083_333, w_083_337, w_083_339, w_083_341, w_083_343, w_083_344, w_083_345, w_083_348, w_083_352, w_083_354, w_083_359, w_083_362, w_083_363, w_083_365, w_083_366, w_083_367, w_083_368, w_083_370, w_083_371, w_083_372, w_083_374, w_083_375, w_083_376, w_083_377, w_083_381, w_083_382, w_083_383, w_083_386, w_083_388, w_083_389, w_083_390, w_083_391, w_083_392, w_083_393, w_083_394, w_083_395, w_083_396, w_083_397, w_083_400, w_083_401, w_083_403, w_083_405, w_083_407, w_083_410, w_083_411, w_083_413, w_083_418, w_083_419, w_083_420, w_083_421, w_083_423, w_083_426, w_083_428, w_083_431, w_083_432, w_083_433, w_083_434, w_083_438, w_083_440, w_083_441, w_083_442, w_083_443, w_083_445, w_083_446, w_083_447, w_083_448, w_083_449, w_083_451, w_083_452, w_083_453, w_083_454, w_083_458, w_083_459, w_083_460, w_083_467, w_083_468, w_083_470, w_083_471, w_083_474, w_083_475, w_083_476, w_083_479, w_083_480, w_083_481, w_083_483, w_083_484, w_083_486, w_083_487, w_083_489, w_083_496, w_083_499, w_083_500, w_083_501, w_083_503, w_083_504, w_083_505, w_083_507, w_083_508, w_083_509, w_083_511, w_083_516, w_083_518, w_083_520, w_083_524, w_083_526, w_083_529, w_083_531, w_083_532, w_083_533, w_083_536, w_083_539, w_083_545, w_083_547, w_083_548, w_083_550, w_083_552, w_083_555, w_083_557, w_083_559, w_083_560, w_083_562, w_083_564, w_083_566, w_083_570, w_083_572, w_083_573, w_083_575, w_083_578, w_083_579, w_083_580, w_083_581, w_083_583, w_083_586, w_083_587, w_083_588, w_083_589, w_083_590, w_083_597, w_083_601, w_083_602, w_083_605, w_083_612, w_083_613, w_083_614, w_083_615, w_083_616, w_083_618, w_083_619, w_083_620, w_083_624, w_083_625, w_083_626, w_083_628, w_083_630, w_083_631, w_083_632, w_083_634, w_083_635, w_083_642, w_083_643, w_083_644, w_083_646, w_083_647, w_083_650, w_083_651, w_083_653, w_083_655, w_083_658, w_083_659, w_083_661, w_083_663, w_083_664, w_083_666, w_083_667, w_083_669, w_083_670, w_083_671, w_083_673, w_083_674, w_083_675, w_083_679, w_083_680, w_083_682, w_083_684, w_083_685, w_083_688, w_083_690, w_083_691, w_083_695, w_083_696, w_083_698, w_083_699, w_083_700, w_083_702, w_083_703, w_083_704, w_083_707, w_083_708, w_083_709, w_083_711, w_083_713, w_083_714, w_083_715, w_083_716, w_083_717, w_083_718, w_083_719, w_083_721, w_083_722, w_083_723, w_083_724, w_083_725, w_083_726, w_083_729, w_083_731, w_083_732, w_083_733, w_083_735, w_083_739, w_083_740, w_083_744, w_083_745, w_083_746, w_083_748, w_083_750, w_083_751, w_083_752, w_083_753, w_083_756, w_083_757, w_083_760, w_083_761, w_083_764, w_083_765, w_083_766, w_083_773, w_083_774, w_083_775, w_083_776, w_083_777, w_083_779, w_083_781, w_083_783, w_083_785, w_083_787, w_083_788, w_083_789, w_083_790, w_083_791, w_083_793, w_083_794, w_083_795, w_083_796, w_083_797, w_083_798, w_083_800, w_083_803, w_083_804, w_083_805, w_083_806, w_083_807, w_083_808, w_083_811, w_083_813, w_083_815, w_083_818, w_083_819, w_083_820, w_083_821, w_083_822, w_083_824, w_083_827, w_083_828, w_083_830, w_083_831, w_083_832, w_083_833, w_083_834, w_083_836, w_083_838, w_083_839, w_083_840, w_083_841, w_083_845, w_083_846, w_083_848, w_083_850, w_083_852, w_083_855, w_083_857, w_083_859, w_083_860, w_083_864, w_083_865, w_083_866, w_083_867, w_083_868, w_083_869, w_083_870, w_083_872, w_083_874, w_083_878, w_083_880, w_083_881, w_083_884, w_083_885, w_083_886, w_083_888, w_083_889, w_083_890, w_083_893, w_083_894, w_083_898, w_083_899, w_083_901, w_083_905, w_083_906, w_083_907, w_083_908, w_083_909, w_083_912, w_083_913, w_083_919, w_083_920, w_083_921, w_083_923, w_083_925, w_083_926, w_083_929, w_083_931, w_083_932, w_083_933, w_083_936, w_083_941, w_083_942, w_083_945, w_083_946, w_083_947, w_083_948, w_083_949, w_083_951, w_083_953, w_083_954, w_083_955, w_083_958, w_083_963, w_083_964, w_083_965, w_083_966, w_083_967, w_083_968, w_083_973, w_083_975, w_083_977, w_083_978, w_083_979, w_083_982, w_083_983, w_083_987, w_083_990, w_083_991, w_083_992, w_083_993, w_083_994, w_083_995, w_083_998, w_083_1004, w_083_1006, w_083_1009, w_083_1011, w_083_1012, w_083_1013, w_083_1016, w_083_1017, w_083_1019, w_083_1020, w_083_1023, w_083_1024, w_083_1025, w_083_1029, w_083_1031, w_083_1035, w_083_1038, w_083_1041, w_083_1042, w_083_1044, w_083_1046, w_083_1047, w_083_1049, w_083_1050, w_083_1051, w_083_1053, w_083_1054, w_083_1058, w_083_1060, w_083_1061, w_083_1062, w_083_1064, w_083_1065, w_083_1066, w_083_1067, w_083_1068, w_083_1070, w_083_1071, w_083_1072, w_083_1074, w_083_1080, w_083_1082, w_083_1085, w_083_1087, w_083_1088, w_083_1090, w_083_1091, w_083_1094, w_083_1096, w_083_1097, w_083_1098, w_083_1100, w_083_1102, w_083_1103, w_083_1106, w_083_1110, w_083_1114, w_083_1115, w_083_1116, w_083_1117, w_083_1118, w_083_1123, w_083_1125, w_083_1126, w_083_1128, w_083_1129, w_083_1132, w_083_1133, w_083_1137, w_083_1138, w_083_1140, w_083_1143, w_083_1145, w_083_1147, w_083_1152, w_083_1154, w_083_1161, w_083_1162, w_083_1164, w_083_1165, w_083_1170, w_083_1171, w_083_1172, w_083_1173, w_083_1174, w_083_1176, w_083_1179, w_083_1182, w_083_1183, w_083_1185, w_083_1186, w_083_1189, w_083_1190, w_083_1191, w_083_1192, w_083_1194, w_083_1196, w_083_1198, w_083_1202, w_083_1207, w_083_1209, w_083_1216, w_083_1218, w_083_1222, w_083_1227, w_083_1231, w_083_1232, w_083_1234, w_083_1235, w_083_1236, w_083_1241, w_083_1243, w_083_1244, w_083_1247, w_083_1248, w_083_1254, w_083_1257, w_083_1258, w_083_1261, w_083_1269, w_083_1270, w_083_1276, w_083_1279, w_083_1281, w_083_1283, w_083_1285, w_083_1286, w_083_1290, w_083_1297, w_083_1304, w_083_1305, w_083_1307, w_083_1309, w_083_1313, w_083_1317, w_083_1318, w_083_1330, w_083_1336, w_083_1337, w_083_1340, w_083_1344, w_083_1349, w_083_1353, w_083_1356, w_083_1357, w_083_1359, w_083_1360, w_083_1362, w_083_1364, w_083_1365, w_083_1369, w_083_1374, w_083_1382, w_083_1384, w_083_1388, w_083_1390, w_083_1394, w_083_1398, w_083_1402, w_083_1405, w_083_1410, w_083_1411, w_083_1417, w_083_1418, w_083_1419, w_083_1420, w_083_1424, w_083_1427, w_083_1428, w_083_1430, w_083_1431, w_083_1440, w_083_1443, w_083_1453, w_083_1455, w_083_1458, w_083_1463, w_083_1465, w_083_1469, w_083_1474, w_083_1478, w_083_1480, w_083_1481, w_083_1490, w_083_1493, w_083_1495, w_083_1496, w_083_1498, w_083_1499, w_083_1501, w_083_1505, w_083_1508, w_083_1509, w_083_1519, w_083_1520, w_083_1522, w_083_1524, w_083_1526, w_083_1535, w_083_1538, w_083_1539, w_083_1543, w_083_1544, w_083_1548, w_083_1549, w_083_1552, w_083_1555, w_083_1561, w_083_1563, w_083_1567, w_083_1568, w_083_1570, w_083_1573, w_083_1579, w_083_1581, w_083_1582, w_083_1594, w_083_1600, w_083_1607, w_083_1611, w_083_1612, w_083_1613, w_083_1619, w_083_1631, w_083_1632, w_083_1636, w_083_1638, w_083_1642, w_083_1643, w_083_1644, w_083_1647, w_083_1649, w_083_1654, w_083_1655, w_083_1667, w_083_1670, w_083_1671, w_083_1672, w_083_1673, w_083_1675, w_083_1676, w_083_1679, w_083_1687, w_083_1688, w_083_1691, w_083_1693, w_083_1695, w_083_1696, w_083_1704, w_083_1716, w_083_1717, w_083_1720, w_083_1722, w_083_1723, w_083_1724, w_083_1733, w_083_1734, w_083_1735, w_083_1737, w_083_1740, w_083_1745, w_083_1750, w_083_1751, w_083_1752, w_083_1759, w_083_1766, w_083_1767, w_083_1769, w_083_1773, w_083_1774, w_083_1775, w_083_1784, w_083_1785, w_083_1787, w_083_1790, w_083_1791, w_083_1792, w_083_1806, w_083_1807, w_083_1814, w_083_1815, w_083_1820, w_083_1825, w_083_1827, w_083_1828, w_083_1829, w_083_1830, w_083_1837, w_083_1838, w_083_1839, w_083_1842, w_083_1845, w_083_1847, w_083_1848, w_083_1855, w_083_1856, w_083_1868, w_083_1871, w_083_1872, w_083_1874, w_083_1875, w_083_1876, w_083_1877, w_083_1880, w_083_1882, w_083_1884, w_083_1885, w_083_1890, w_083_1892, w_083_1895, w_083_1897, w_083_1898, w_083_1901, w_083_1903, w_083_1906, w_083_1912, w_083_1916, w_083_1923, w_083_1926, w_083_1928, w_083_1930, w_083_1931, w_083_1932, w_083_1936, w_083_1941, w_083_1942, w_083_1943, w_083_1946, w_083_1949, w_083_1955, w_083_1957, w_083_1958, w_083_1962, w_083_1964, w_083_1970, w_083_1972, w_083_1975, w_083_1979, w_083_1980, w_083_1981, w_083_1984, w_083_1988, w_083_1992, w_083_1994, w_083_1995, w_083_1996, w_083_1997, w_083_1998, w_083_1999, w_083_2000, w_083_2001, w_083_2003, w_083_2005, w_083_2010, w_083_2015, w_083_2023, w_083_2030, w_083_2033, w_083_2034, w_083_2036, w_083_2043, w_083_2045, w_083_2050, w_083_2051, w_083_2055, w_083_2056, w_083_2059, w_083_2060, w_083_2077, w_083_2083, w_083_2087, w_083_2089, w_083_2093, w_083_2095, w_083_2096, w_083_2102, w_083_2105, w_083_2107, w_083_2108, w_083_2109, w_083_2111, w_083_2112, w_083_2113, w_083_2121, w_083_2122, w_083_2123, w_083_2125, w_083_2130, w_083_2131, w_083_2134, w_083_2136, w_083_2137, w_083_2143, w_083_2149, w_083_2151, w_083_2155, w_083_2158, w_083_2159, w_083_2160, w_083_2163, w_083_2168, w_083_2169, w_083_2173, w_083_2174, w_083_2180, w_083_2184, w_083_2187, w_083_2189, w_083_2193, w_083_2195, w_083_2196, w_083_2198, w_083_2201, w_083_2205, w_083_2206, w_083_2207, w_083_2208, w_083_2210, w_083_2212, w_083_2216, w_083_2217, w_083_2218, w_083_2224, w_083_2226, w_083_2228, w_083_2230, w_083_2231, w_083_2234, w_083_2240, w_083_2242, w_083_2243, w_083_2244, w_083_2248, w_083_2251, w_083_2256, w_083_2259, w_083_2272, w_083_2275, w_083_2277, w_083_2282, w_083_2285, w_083_2292, w_083_2293, w_083_2294, w_083_2295, w_083_2296, w_083_2297, w_083_2299, w_083_2300, w_083_2301, w_083_2303, w_083_2305, w_083_2309, w_083_2311, w_083_2314, w_083_2315, w_083_2320, w_083_2323, w_083_2325, w_083_2326, w_083_2327, w_083_2329, w_083_2330, w_083_2332, w_083_2333, w_083_2336, w_083_2338, w_083_2339, w_083_2340, w_083_2341, w_083_2343, w_083_2346, w_083_2349, w_083_2350, w_083_2351, w_083_2352, w_083_2354, w_083_2355, w_083_2362, w_083_2364, w_083_2365, w_083_2372, w_083_2376, w_083_2378, w_083_2389, w_083_2391, w_083_2392, w_083_2396, w_083_2399, w_083_2401, w_083_2406, w_083_2408, w_083_2410, w_083_2412, w_083_2417, w_083_2419, w_083_2421, w_083_2429, w_083_2430, w_083_2434, w_083_2437, w_083_2438, w_083_2439, w_083_2441, w_083_2446, w_083_2454, w_083_2458, w_083_2468, w_083_2476, w_083_2483, w_083_2485, w_083_2486, w_083_2487, w_083_2490, w_083_2491, w_083_2492, w_083_2493, w_083_2495, w_083_2496, w_083_2499, w_083_2502, w_083_2504, w_083_2506, w_083_2508, w_083_2518, w_083_2520, w_083_2525, w_083_2526, w_083_2530, w_083_2537, w_083_2538, w_083_2544, w_083_2545, w_083_2547, w_083_2557, w_083_2559, w_083_2562, w_083_2565, w_083_2568, w_083_2571, w_083_2576, w_083_2577, w_083_2581, w_083_2583, w_083_2586, w_083_2587, w_083_2591, w_083_2594, w_083_2601, w_083_2606, w_083_2607, w_083_2608, w_083_2609, w_083_2612, w_083_2615, w_083_2616, w_083_2625, w_083_2626, w_083_2627, w_083_2632, w_083_2639, w_083_2644, w_083_2645, w_083_2648, w_083_2649, w_083_2651, w_083_2654, w_083_2657, w_083_2659, w_083_2667, w_083_2672, w_083_2675, w_083_2679, w_083_2681, w_083_2685, w_083_2690, w_083_2694, w_083_2697, w_083_2698, w_083_2700, w_083_2711, w_083_2713, w_083_2719, w_083_2723, w_083_2725, w_083_2726, w_083_2729, w_083_2733, w_083_2739, w_083_2740, w_083_2745, w_083_2746, w_083_2752, w_083_2755, w_083_2763, w_083_2769, w_083_2771, w_083_2772, w_083_2775, w_083_2777, w_083_2780, w_083_2784, w_083_2786, w_083_2790, w_083_2791, w_083_2793, w_083_2796, w_083_2802, w_083_2807, w_083_2821, w_083_2824, w_083_2825, w_083_2827, w_083_2831, w_083_2839, w_083_2844, w_083_2845, w_083_2846, w_083_2850, w_083_2858, w_083_2861, w_083_2864, w_083_2865, w_083_2869, w_083_2877, w_083_2879, w_083_2883, w_083_2889, w_083_2891, w_083_2894, w_083_2898, w_083_2905, w_083_2907, w_083_2909, w_083_2913, w_083_2921, w_083_2922, w_083_2925, w_083_2927, w_083_2928, w_083_2929, w_083_2933, w_083_2936, w_083_2937, w_083_2939, w_083_2945, w_083_2949, w_083_2950, w_083_2956, w_083_2958, w_083_2961, w_083_2964, w_083_2965, w_083_2967, w_083_2968, w_083_2969, w_083_2971, w_083_2972, w_083_2976, w_083_2977, w_083_2982, w_083_2985, w_083_2987, w_083_2989, w_083_2993, w_083_2994, w_083_2998, w_083_3000, w_083_3001, w_083_3003, w_083_3006, w_083_3007, w_083_3010, w_083_3011, w_083_3016, w_083_3024, w_083_3026, w_083_3027, w_083_3028, w_083_3034, w_083_3045, w_083_3049, w_083_3054, w_083_3055, w_083_3056, w_083_3058, w_083_3061, w_083_3062, w_083_3063, w_083_3064, w_083_3067, w_083_3068, w_083_3069, w_083_3071, w_083_3080, w_083_3081, w_083_3086, w_083_3088, w_083_3094, w_083_3095, w_083_3100, w_083_3103, w_083_3109, w_083_3110, w_083_3112, w_083_3114, w_083_3115, w_083_3118, w_083_3119, w_083_3123, w_083_3125, w_083_3127, w_083_3134, w_083_3142, w_083_3143, w_083_3150, w_083_3151, w_083_3154, w_083_3157, w_083_3159, w_083_3163, w_083_3166, w_083_3167, w_083_3171, w_083_3172, w_083_3178, w_083_3179, w_083_3180, w_083_3181, w_083_3183, w_083_3184, w_083_3185, w_083_3189, w_083_3194, w_083_3196, w_083_3199, w_083_3206, w_083_3207, w_083_3208, w_083_3209, w_083_3210, w_083_3214, w_083_3215, w_083_3222, w_083_3223, w_083_3228, w_083_3229, w_083_3231, w_083_3232, w_083_3233, w_083_3234, w_083_3236, w_083_3238, w_083_3243, w_083_3244, w_083_3254, w_083_3257, w_083_3262, w_083_3263, w_083_3264, w_083_3266, w_083_3269, w_083_3271, w_083_3275, w_083_3279, w_083_3283, w_083_3284, w_083_3286, w_083_3289, w_083_3292, w_083_3298, w_083_3301, w_083_3306, w_083_3308, w_083_3311, w_083_3313, w_083_3315, w_083_3327, w_083_3331, w_083_3333, w_083_3334, w_083_3335, w_083_3338, w_083_3343, w_083_3344, w_083_3346, w_083_3347, w_083_3354, w_083_3355, w_083_3359, w_083_3363, w_083_3369, w_083_3376, w_083_3378, w_083_3380, w_083_3383, w_083_3387, w_083_3400, w_083_3402, w_083_3406, w_083_3408, w_083_3409, w_083_3411, w_083_3413, w_083_3417, w_083_3419, w_083_3423, w_083_3427, w_083_3428, w_083_3429, w_083_3431, w_083_3438, w_083_3442, w_083_3448, w_083_3451, w_083_3454, w_083_3455, w_083_3457, w_083_3461, w_083_3462, w_083_3466, w_083_3472, w_083_3474, w_083_3476, w_083_3479, w_083_3481, w_083_3483, w_083_3484, w_083_3486, w_083_3491, w_083_3493, w_083_3499, w_083_3500, w_083_3501, w_083_3503, w_083_3509, w_083_3510, w_083_3511, w_083_3513, w_083_3514, w_083_3516, w_083_3517, w_083_3518, w_083_3520, w_083_3521, w_083_3524, w_083_3526, w_083_3528, w_083_3535, w_083_3536, w_083_3538, w_083_3539, w_083_3541, w_083_3544, w_083_3546, w_083_3548, w_083_3551, w_083_3553, w_083_3554, w_083_3557, w_083_3562, w_083_3563, w_083_3567, w_083_3568, w_083_3569, w_083_3570, w_083_3572, w_083_3574, w_083_3577, w_083_3578, w_083_3580, w_083_3581, w_083_3582, w_083_3583, w_083_3584, w_083_3588, w_083_3589, w_083_3591, w_083_3596, w_083_3597, w_083_3598, w_083_3599, w_083_3600, w_083_3602, w_083_3604, w_083_3605, w_083_3609, w_083_3611, w_083_3613, w_083_3616, w_083_3618, w_083_3623, w_083_3625, w_083_3627, w_083_3628, w_083_3634, w_083_3635, w_083_3636, w_083_3637, w_083_3638, w_083_3640, w_083_3641, w_083_3648, w_083_3649, w_083_3650, w_083_3651, w_083_3656, w_083_3658, w_083_3660, w_083_3661, w_083_3664, w_083_3665, w_083_3670, w_083_3673, w_083_3679, w_083_3682, w_083_3683, w_083_3684, w_083_3686, w_083_3702, w_083_3708, w_083_3709, w_083_3710, w_083_3711, w_083_3713, w_083_3715, w_083_3718, w_083_3733, w_083_3737, w_083_3738, w_083_3742, w_083_3743, w_083_3744, w_083_3745, w_083_3748, w_083_3750, w_083_3752, w_083_3754, w_083_3755, w_083_3756, w_083_3758, w_083_3763, w_083_3769, w_083_3771, w_083_3775, w_083_3777, w_083_3780, w_083_3781, w_083_3786, w_083_3789, w_083_3796;
  wire w_084_000, w_084_001, w_084_003, w_084_007, w_084_009, w_084_010, w_084_011, w_084_012, w_084_014, w_084_015, w_084_016, w_084_019, w_084_022, w_084_023, w_084_024, w_084_025, w_084_027, w_084_030, w_084_033, w_084_035, w_084_037, w_084_041, w_084_044, w_084_045, w_084_046, w_084_047, w_084_049, w_084_054, w_084_057, w_084_058, w_084_059, w_084_060, w_084_061, w_084_064, w_084_066, w_084_069, w_084_071, w_084_074, w_084_075, w_084_076, w_084_077, w_084_080, w_084_081, w_084_082, w_084_083, w_084_084, w_084_086, w_084_087, w_084_088, w_084_089, w_084_090, w_084_093, w_084_097, w_084_098, w_084_099, w_084_100, w_084_102, w_084_103, w_084_104, w_084_107, w_084_108, w_084_111, w_084_117, w_084_119, w_084_126, w_084_127, w_084_129, w_084_131, w_084_133, w_084_137, w_084_139, w_084_140, w_084_142, w_084_146, w_084_151, w_084_152, w_084_153, w_084_155, w_084_156, w_084_157, w_084_162, w_084_163, w_084_164, w_084_166, w_084_170, w_084_175, w_084_179, w_084_180, w_084_181, w_084_185, w_084_186, w_084_187, w_084_189, w_084_190, w_084_192, w_084_195, w_084_197, w_084_199, w_084_201, w_084_205, w_084_206, w_084_210, w_084_212, w_084_214, w_084_217, w_084_220, w_084_222, w_084_226, w_084_227, w_084_228, w_084_229, w_084_230, w_084_231, w_084_233, w_084_235, w_084_236, w_084_241, w_084_243, w_084_247, w_084_256, w_084_257, w_084_258, w_084_260, w_084_261, w_084_262, w_084_263, w_084_265, w_084_266, w_084_267, w_084_269, w_084_270, w_084_271, w_084_272, w_084_276, w_084_277, w_084_279, w_084_281, w_084_284, w_084_286, w_084_287, w_084_288, w_084_289, w_084_293, w_084_294, w_084_295, w_084_297, w_084_298, w_084_299, w_084_306, w_084_308, w_084_309, w_084_310, w_084_315, w_084_316, w_084_320, w_084_323, w_084_324, w_084_325, w_084_327, w_084_328, w_084_329, w_084_332, w_084_333, w_084_334, w_084_337, w_084_338, w_084_343, w_084_344, w_084_345, w_084_347, w_084_348, w_084_349, w_084_351, w_084_354, w_084_355, w_084_358, w_084_360, w_084_361, w_084_363, w_084_366, w_084_369, w_084_370, w_084_374, w_084_375, w_084_376, w_084_377, w_084_379, w_084_380, w_084_381, w_084_382, w_084_383, w_084_384, w_084_385, w_084_386, w_084_389, w_084_390, w_084_391, w_084_392, w_084_394, w_084_395, w_084_396, w_084_398, w_084_399, w_084_400, w_084_401, w_084_403, w_084_404, w_084_406, w_084_407, w_084_408, w_084_409, w_084_412, w_084_413, w_084_414, w_084_416, w_084_417, w_084_419, w_084_422, w_084_425, w_084_428, w_084_432, w_084_433, w_084_434, w_084_435, w_084_436, w_084_437, w_084_438, w_084_440, w_084_441, w_084_442, w_084_444, w_084_445, w_084_447, w_084_448, w_084_449, w_084_454, w_084_455, w_084_458, w_084_459, w_084_460, w_084_463, w_084_464, w_084_466, w_084_467, w_084_468, w_084_469, w_084_470, w_084_471, w_084_473, w_084_476, w_084_477, w_084_478, w_084_483, w_084_484, w_084_487, w_084_490, w_084_497, w_084_498, w_084_499, w_084_510, w_084_511, w_084_512, w_084_513, w_084_514, w_084_515, w_084_518, w_084_523, w_084_525, w_084_528, w_084_531, w_084_537, w_084_538, w_084_541, w_084_550, w_084_552, w_084_553, w_084_558, w_084_559, w_084_561, w_084_566, w_084_567, w_084_568, w_084_577, w_084_581, w_084_582, w_084_588, w_084_594, w_084_598, w_084_599, w_084_603, w_084_604, w_084_609, w_084_612, w_084_613, w_084_624, w_084_625, w_084_626, w_084_627, w_084_631, w_084_634, w_084_635, w_084_636, w_084_637, w_084_638, w_084_640, w_084_641, w_084_642, w_084_648, w_084_651, w_084_652, w_084_653, w_084_657, w_084_660, w_084_662, w_084_663, w_084_664, w_084_670, w_084_672, w_084_673, w_084_674, w_084_676, w_084_683, w_084_688, w_084_689, w_084_691, w_084_693, w_084_696, w_084_699, w_084_701, w_084_707, w_084_709, w_084_710, w_084_717, w_084_718, w_084_719, w_084_722, w_084_726, w_084_730, w_084_735, w_084_743, w_084_744, w_084_748, w_084_752, w_084_755, w_084_757, w_084_762, w_084_763, w_084_766, w_084_769, w_084_770, w_084_779, w_084_783, w_084_788, w_084_789, w_084_795, w_084_797, w_084_798, w_084_800, w_084_801, w_084_803, w_084_806, w_084_807, w_084_810, w_084_811, w_084_812, w_084_814, w_084_817, w_084_822, w_084_828, w_084_837, w_084_838, w_084_845, w_084_862, w_084_865, w_084_869, w_084_871, w_084_872, w_084_873, w_084_874, w_084_875, w_084_882, w_084_883, w_084_886, w_084_887, w_084_891, w_084_893, w_084_894, w_084_896, w_084_901, w_084_903, w_084_911, w_084_916, w_084_920, w_084_921, w_084_922, w_084_923, w_084_924, w_084_925, w_084_926, w_084_930, w_084_932, w_084_936, w_084_939, w_084_940, w_084_942, w_084_943, w_084_946, w_084_948, w_084_950, w_084_954, w_084_956, w_084_965, w_084_967, w_084_968, w_084_969, w_084_972, w_084_976, w_084_978, w_084_981, w_084_983, w_084_984, w_084_986, w_084_988, w_084_990, w_084_993, w_084_996, w_084_997, w_084_1004, w_084_1006, w_084_1007, w_084_1011, w_084_1013, w_084_1014, w_084_1021, w_084_1035, w_084_1039, w_084_1040, w_084_1047, w_084_1049, w_084_1050, w_084_1051, w_084_1052, w_084_1053, w_084_1055, w_084_1058, w_084_1061, w_084_1063, w_084_1068, w_084_1072, w_084_1073, w_084_1076, w_084_1079, w_084_1081, w_084_1083, w_084_1084, w_084_1085, w_084_1087, w_084_1094, w_084_1095, w_084_1099, w_084_1100, w_084_1101, w_084_1114, w_084_1116, w_084_1117, w_084_1119, w_084_1121, w_084_1123, w_084_1124, w_084_1127, w_084_1129, w_084_1136, w_084_1138, w_084_1139, w_084_1140, w_084_1142, w_084_1152, w_084_1154, w_084_1155, w_084_1160, w_084_1161, w_084_1163, w_084_1165, w_084_1166, w_084_1170, w_084_1172, w_084_1173, w_084_1181, w_084_1184, w_084_1185, w_084_1194, w_084_1195, w_084_1198, w_084_1203, w_084_1207, w_084_1209, w_084_1210, w_084_1211, w_084_1212, w_084_1215, w_084_1216, w_084_1218, w_084_1220, w_084_1222, w_084_1227, w_084_1229, w_084_1232, w_084_1234, w_084_1237, w_084_1238, w_084_1244, w_084_1247, w_084_1251, w_084_1252, w_084_1253, w_084_1258, w_084_1263, w_084_1268, w_084_1269, w_084_1275, w_084_1276, w_084_1277, w_084_1279, w_084_1283, w_084_1285, w_084_1286, w_084_1287, w_084_1290, w_084_1296, w_084_1297, w_084_1299, w_084_1300, w_084_1301, w_084_1305, w_084_1306, w_084_1311, w_084_1312, w_084_1317, w_084_1319, w_084_1325, w_084_1329, w_084_1332, w_084_1333, w_084_1339, w_084_1340, w_084_1342, w_084_1344, w_084_1345, w_084_1349, w_084_1350, w_084_1351, w_084_1356, w_084_1358, w_084_1360, w_084_1365, w_084_1366, w_084_1367, w_084_1369, w_084_1372, w_084_1376, w_084_1377, w_084_1379, w_084_1384, w_084_1387, w_084_1388, w_084_1390, w_084_1397, w_084_1398, w_084_1401, w_084_1404, w_084_1411, w_084_1415, w_084_1419, w_084_1422, w_084_1427, w_084_1428, w_084_1439, w_084_1442, w_084_1444, w_084_1446, w_084_1454, w_084_1458, w_084_1461, w_084_1462, w_084_1463, w_084_1472, w_084_1473, w_084_1475, w_084_1476, w_084_1477, w_084_1479, w_084_1484, w_084_1490, w_084_1491, w_084_1492, w_084_1493, w_084_1505, w_084_1511, w_084_1513, w_084_1515, w_084_1520, w_084_1528, w_084_1530, w_084_1531, w_084_1535, w_084_1536, w_084_1538, w_084_1547, w_084_1549, w_084_1550, w_084_1551, w_084_1553, w_084_1554, w_084_1557, w_084_1558, w_084_1568, w_084_1569, w_084_1577, w_084_1583, w_084_1584, w_084_1586, w_084_1588, w_084_1589, w_084_1590, w_084_1592, w_084_1596, w_084_1597, w_084_1599, w_084_1600, w_084_1606, w_084_1610, w_084_1613, w_084_1617, w_084_1619, w_084_1627, w_084_1628, w_084_1630, w_084_1635, w_084_1636, w_084_1641, w_084_1642, w_084_1644, w_084_1645, w_084_1649, w_084_1650, w_084_1653, w_084_1657, w_084_1660, w_084_1661, w_084_1663, w_084_1664, w_084_1668, w_084_1671, w_084_1674, w_084_1678, w_084_1680, w_084_1681, w_084_1682, w_084_1684, w_084_1685, w_084_1686, w_084_1689, w_084_1692, w_084_1694, w_084_1699, w_084_1700, w_084_1703, w_084_1709, w_084_1710, w_084_1712, w_084_1713, w_084_1723, w_084_1724, w_084_1725, w_084_1726, w_084_1729, w_084_1730, w_084_1739, w_084_1744, w_084_1752, w_084_1754, w_084_1757, w_084_1758, w_084_1761, w_084_1763, w_084_1765, w_084_1770, w_084_1771, w_084_1773, w_084_1774, w_084_1776, w_084_1779, w_084_1781, w_084_1788, w_084_1795, w_084_1797, w_084_1798, w_084_1804, w_084_1805, w_084_1807, w_084_1809, w_084_1810, w_084_1811, w_084_1814, w_084_1815, w_084_1817, w_084_1819, w_084_1824, w_084_1825, w_084_1827, w_084_1828, w_084_1830, w_084_1834, w_084_1836, w_084_1839, w_084_1840, w_084_1841, w_084_1855, w_084_1858, w_084_1861, w_084_1863, w_084_1865, w_084_1866, w_084_1867, w_084_1872, w_084_1873, w_084_1876, w_084_1881, w_084_1883, w_084_1895, w_084_1897, w_084_1898, w_084_1903, w_084_1905, w_084_1906, w_084_1911, w_084_1915, w_084_1918, w_084_1923, w_084_1926, w_084_1930, w_084_1931, w_084_1936, w_084_1937, w_084_1938, w_084_1941, w_084_1945, w_084_1946, w_084_1953, w_084_1959, w_084_1967, w_084_1973, w_084_1974, w_084_1979, w_084_1980, w_084_1982, w_084_1985, w_084_1990, w_084_1995, w_084_1996, w_084_2001, w_084_2002, w_084_2004, w_084_2010, w_084_2014, w_084_2015, w_084_2020, w_084_2021, w_084_2024, w_084_2025, w_084_2028, w_084_2029, w_084_2032, w_084_2033, w_084_2035, w_084_2036, w_084_2037, w_084_2041, w_084_2048, w_084_2050, w_084_2053, w_084_2055, w_084_2059, w_084_2061, w_084_2066, w_084_2067, w_084_2072, w_084_2076, w_084_2080, w_084_2081, w_084_2082, w_084_2084, w_084_2089, w_084_2090, w_084_2091, w_084_2093, w_084_2094, w_084_2095, w_084_2098, w_084_2102, w_084_2106, w_084_2110, w_084_2112, w_084_2113, w_084_2120, w_084_2121, w_084_2123, w_084_2130, w_084_2133, w_084_2136, w_084_2137, w_084_2139, w_084_2140, w_084_2141, w_084_2144, w_084_2146, w_084_2147, w_084_2148, w_084_2150, w_084_2159, w_084_2161, w_084_2165, w_084_2167, w_084_2175, w_084_2178, w_084_2179, w_084_2183, w_084_2184, w_084_2196, w_084_2200, w_084_2206, w_084_2214, w_084_2217, w_084_2220, w_084_2221, w_084_2222, w_084_2224, w_084_2225, w_084_2228, w_084_2230, w_084_2239, w_084_2241, w_084_2242, w_084_2244, w_084_2245, w_084_2247, w_084_2249, w_084_2251, w_084_2254, w_084_2262, w_084_2268, w_084_2269, w_084_2271, w_084_2275, w_084_2277, w_084_2282, w_084_2283, w_084_2284, w_084_2288, w_084_2290, w_084_2291, w_084_2292, w_084_2294, w_084_2296, w_084_2304, w_084_2306, w_084_2307, w_084_2308, w_084_2310, w_084_2312, w_084_2314, w_084_2323, w_084_2324, w_084_2326, w_084_2334, w_084_2335, w_084_2337, w_084_2338, w_084_2341, w_084_2343, w_084_2349, w_084_2350, w_084_2353, w_084_2354, w_084_2359, w_084_2365, w_084_2366, w_084_2369, w_084_2370, w_084_2371, w_084_2379, w_084_2383, w_084_2386, w_084_2388, w_084_2390, w_084_2394, w_084_2397, w_084_2402, w_084_2403, w_084_2405, w_084_2406, w_084_2414, w_084_2415, w_084_2420, w_084_2423, w_084_2424, w_084_2426, w_084_2435, w_084_2436, w_084_2442, w_084_2443, w_084_2445, w_084_2446, w_084_2448, w_084_2451, w_084_2453, w_084_2459, w_084_2467, w_084_2480, w_084_2481, w_084_2482, w_084_2489, w_084_2491, w_084_2497, w_084_2498, w_084_2503, w_084_2505, w_084_2508, w_084_2509, w_084_2510, w_084_2512, w_084_2514, w_084_2517, w_084_2518, w_084_2520, w_084_2521, w_084_2524, w_084_2525, w_084_2526, w_084_2531, w_084_2535, w_084_2538, w_084_2539, w_084_2544, w_084_2546, w_084_2550, w_084_2552, w_084_2553, w_084_2557, w_084_2564, w_084_2566, w_084_2570, w_084_2573, w_084_2577, w_084_2581, w_084_2590, w_084_2592, w_084_2600, w_084_2601, w_084_2608, w_084_2612, w_084_2613, w_084_2619, w_084_2620, w_084_2623, w_084_2625, w_084_2626, w_084_2628, w_084_2630, w_084_2632, w_084_2634, w_084_2636, w_084_2637, w_084_2643, w_084_2645, w_084_2646, w_084_2647, w_084_2649, w_084_2660, w_084_2661, w_084_2662, w_084_2663, w_084_2667, w_084_2674, w_084_2676, w_084_2677, w_084_2678, w_084_2679, w_084_2680, w_084_2681, w_084_2685, w_084_2688, w_084_2692, w_084_2693, w_084_2694, w_084_2695, w_084_2696, w_084_2698, w_084_2703, w_084_2706, w_084_2709, w_084_2711, w_084_2713, w_084_2715, w_084_2718, w_084_2721, w_084_2723, w_084_2725, w_084_2726, w_084_2728, w_084_2730, w_084_2733, w_084_2734, w_084_2736, w_084_2739, w_084_2740, w_084_2741, w_084_2742, w_084_2746, w_084_2747, w_084_2748, w_084_2751, w_084_2754, w_084_2756, w_084_2762, w_084_2763, w_084_2765, w_084_2768, w_084_2769, w_084_2771, w_084_2772, w_084_2778, w_084_2785, w_084_2787, w_084_2789, w_084_2790, w_084_2791, w_084_2795, w_084_2797, w_084_2805, w_084_2807, w_084_2809, w_084_2810, w_084_2811, w_084_2812, w_084_2814, w_084_2820, w_084_2824, w_084_2832, w_084_2835, w_084_2840, w_084_2841, w_084_2844, w_084_2849, w_084_2852, w_084_2860, w_084_2861, w_084_2863, w_084_2868, w_084_2871, w_084_2873, w_084_2882, w_084_2887, w_084_2890, w_084_2891, w_084_2897, w_084_2898, w_084_2909, w_084_2913, w_084_2916, w_084_2918, w_084_2919, w_084_2925, w_084_2937, w_084_2939, w_084_2940, w_084_2942, w_084_2952, w_084_2956, w_084_2957, w_084_2958, w_084_2959, w_084_2965, w_084_2971, w_084_2972, w_084_2973, w_084_2975, w_084_2977, w_084_2987, w_084_2992, w_084_2994, w_084_2999, w_084_3000, w_084_3002, w_084_3004, w_084_3007, w_084_3009, w_084_3012, w_084_3014, w_084_3016, w_084_3019, w_084_3020, w_084_3022, w_084_3026, w_084_3027, w_084_3028, w_084_3039, w_084_3041, w_084_3042, w_084_3043, w_084_3044, w_084_3047, w_084_3048, w_084_3051, w_084_3054, w_084_3057, w_084_3066, w_084_3072, w_084_3074, w_084_3087, w_084_3089, w_084_3091, w_084_3092, w_084_3099, w_084_3102, w_084_3106, w_084_3109, w_084_3115, w_084_3117, w_084_3118, w_084_3119, w_084_3121, w_084_3122, w_084_3125, w_084_3136, w_084_3138, w_084_3140, w_084_3143, w_084_3154, w_084_3157, w_084_3166, w_084_3170, w_084_3175, w_084_3178, w_084_3181, w_084_3182, w_084_3183, w_084_3192, w_084_3197, w_084_3198, w_084_3202, w_084_3205, w_084_3208, w_084_3211, w_084_3212, w_084_3217, w_084_3221, w_084_3223, w_084_3224, w_084_3227, w_084_3230, w_084_3232, w_084_3233, w_084_3234, w_084_3235, w_084_3237, w_084_3242, w_084_3243, w_084_3248, w_084_3251, w_084_3256, w_084_3257, w_084_3258, w_084_3263, w_084_3266, w_084_3267, w_084_3268, w_084_3269, w_084_3274, w_084_3276, w_084_3280, w_084_3281, w_084_3282, w_084_3285, w_084_3286, w_084_3290, w_084_3292, w_084_3297, w_084_3299, w_084_3306, w_084_3308, w_084_3310, w_084_3311, w_084_3313, w_084_3320, w_084_3321, w_084_3325, w_084_3328, w_084_3329, w_084_3330, w_084_3332, w_084_3333, w_084_3339, w_084_3345, w_084_3349, w_084_3350, w_084_3351, w_084_3354, w_084_3357, w_084_3359, w_084_3362, w_084_3363, w_084_3367, w_084_3369, w_084_3372, w_084_3374, w_084_3375, w_084_3387, w_084_3393, w_084_3394, w_084_3399, w_084_3402, w_084_3405, w_084_3408, w_084_3413, w_084_3415, w_084_3416, w_084_3420, w_084_3422, w_084_3423, w_084_3425, w_084_3426, w_084_3427, w_084_3430, w_084_3431, w_084_3432, w_084_3437, w_084_3446, w_084_3452, w_084_3458, w_084_3468, w_084_3474, w_084_3475, w_084_3476, w_084_3477, w_084_3482, w_084_3486, w_084_3487, w_084_3489, w_084_3491, w_084_3496, w_084_3500, w_084_3501, w_084_3509, w_084_3515, w_084_3520, w_084_3522, w_084_3526, w_084_3531, w_084_3540, w_084_3541, w_084_3545, w_084_3548, w_084_3549, w_084_3550, w_084_3551, w_084_3552, w_084_3553, w_084_3556, w_084_3561, w_084_3563, w_084_3565, w_084_3573, w_084_3579, w_084_3582, w_084_3583, w_084_3587, w_084_3590, w_084_3591, w_084_3592, w_084_3594, w_084_3595, w_084_3596, w_084_3600, w_084_3604, w_084_3605, w_084_3612, w_084_3614, w_084_3615, w_084_3616, w_084_3617, w_084_3618, w_084_3620, w_084_3625, w_084_3626, w_084_3632, w_084_3633, w_084_3634, w_084_3646, w_084_3648, w_084_3649, w_084_3651, w_084_3654, w_084_3655, w_084_3660, w_084_3661, w_084_3662, w_084_3663, w_084_3665, w_084_3669, w_084_3678, w_084_3680, w_084_3682, w_084_3683, w_084_3684, w_084_3685, w_084_3687, w_084_3688, w_084_3691, w_084_3692, w_084_3696, w_084_3697, w_084_3703, w_084_3707, w_084_3711, w_084_3712, w_084_3713, w_084_3717, w_084_3726, w_084_3727, w_084_3738, w_084_3741, w_084_3747, w_084_3748, w_084_3750, w_084_3759, w_084_3761, w_084_3765, w_084_3766, w_084_3770, w_084_3771, w_084_3773, w_084_3774, w_084_3775, w_084_3779, w_084_3794, w_084_3795, w_084_3804, w_084_3810, w_084_3814, w_084_3815, w_084_3816, w_084_3817, w_084_3819, w_084_3820, w_084_3825, w_084_3831, w_084_3832, w_084_3833, w_084_3836, w_084_3839, w_084_3843, w_084_3847, w_084_3848, w_084_3849, w_084_3850, w_084_3852, w_084_3854, w_084_3855, w_084_3858, w_084_3862, w_084_3869, w_084_3870, w_084_3876, w_084_3877, w_084_3880, w_084_3882, w_084_3885, w_084_3888, w_084_3890, w_084_3891, w_084_3893, w_084_3897, w_084_3900, w_084_3901, w_084_3904, w_084_3908, w_084_3910, w_084_3912, w_084_3913, w_084_3916, w_084_3917, w_084_3921, w_084_3924, w_084_3928, w_084_3931, w_084_3934, w_084_3935, w_084_3936, w_084_3937, w_084_3940, w_084_3942, w_084_3943, w_084_3946, w_084_3949, w_084_3951, w_084_3953, w_084_3954, w_084_3955, w_084_3957, w_084_3959, w_084_3960, w_084_3963, w_084_3967, w_084_3968, w_084_3971, w_084_3972, w_084_3975, w_084_3976, w_084_3977, w_084_3982, w_084_3983, w_084_3985, w_084_3986, w_084_3988, w_084_3992, w_084_3997, w_084_3999, w_084_4002, w_084_4003, w_084_4004, w_084_4005, w_084_4011, w_084_4012, w_084_4020, w_084_4022, w_084_4024, w_084_4035, w_084_4036, w_084_4037, w_084_4040, w_084_4047, w_084_4049, w_084_4050, w_084_4052, w_084_4053, w_084_4060, w_084_4068, w_084_4069, w_084_4076, w_084_4078, w_084_4079, w_084_4085, w_084_4088, w_084_4091, w_084_4094, w_084_4096, w_084_4099, w_084_4103, w_084_4115, w_084_4131, w_084_4132, w_084_4141, w_084_4142, w_084_4147, w_084_4148, w_084_4149, w_084_4154, w_084_4155, w_084_4160, w_084_4162, w_084_4163, w_084_4164, w_084_4165, w_084_4170, w_084_4171, w_084_4188, w_084_4190, w_084_4191, w_084_4196, w_084_4197, w_084_4201, w_084_4203, w_084_4204, w_084_4205, w_084_4208, w_084_4210, w_084_4218, w_084_4219, w_084_4220, w_084_4222, w_084_4227, w_084_4232, w_084_4237, w_084_4238, w_084_4241, w_084_4242, w_084_4244, w_084_4249, w_084_4250, w_084_4252, w_084_4260, w_084_4264, w_084_4267, w_084_4270, w_084_4271, w_084_4272, w_084_4274, w_084_4282, w_084_4283, w_084_4284, w_084_4285, w_084_4287, w_084_4294, w_084_4298, w_084_4299, w_084_4303, w_084_4307, w_084_4311, w_084_4321, w_084_4324, w_084_4327, w_084_4328, w_084_4329, w_084_4330, w_084_4333, w_084_4334, w_084_4335, w_084_4346, w_084_4351, w_084_4352, w_084_4358, w_084_4361, w_084_4367, w_084_4371, w_084_4376, w_084_4378, w_084_4380, w_084_4383, w_084_4384, w_084_4385, w_084_4389, w_084_4390, w_084_4397, w_084_4400, w_084_4403, w_084_4405, w_084_4411, w_084_4412, w_084_4416, w_084_4422, w_084_4424, w_084_4426, w_084_4430, w_084_4433, w_084_4435, w_084_4442, w_084_4447, w_084_4453, w_084_4454, w_084_4458, w_084_4460, w_084_4461, w_084_4466, w_084_4467, w_084_4468, w_084_4469, w_084_4471, w_084_4472, w_084_4474, w_084_4483, w_084_4484, w_084_4490, w_084_4491, w_084_4494, w_084_4496, w_084_4498, w_084_4501, w_084_4503, w_084_4507, w_084_4511;
  wire w_085_000, w_085_001, w_085_003, w_085_004, w_085_005, w_085_006, w_085_007, w_085_008, w_085_009, w_085_010, w_085_011, w_085_012, w_085_013, w_085_014, w_085_015, w_085_016, w_085_017, w_085_019, w_085_020, w_085_021, w_085_022, w_085_023, w_085_024, w_085_025, w_085_026, w_085_027, w_085_028, w_085_029, w_085_030, w_085_031, w_085_032, w_085_033, w_085_034, w_085_035, w_085_036, w_085_037, w_085_038, w_085_039, w_085_040, w_085_042, w_085_043, w_085_044, w_085_045, w_085_046, w_085_047, w_085_048, w_085_049, w_085_050, w_085_051, w_085_052, w_085_053, w_085_054, w_085_055, w_085_056, w_085_057, w_085_058, w_085_061, w_085_062, w_085_064, w_085_065, w_085_067, w_085_068, w_085_069, w_085_070, w_085_071, w_085_072, w_085_073, w_085_074, w_085_075, w_085_076, w_085_077, w_085_078, w_085_079, w_085_080, w_085_082, w_085_083, w_085_085, w_085_087, w_085_088, w_085_089, w_085_090, w_085_091, w_085_092, w_085_093, w_085_094, w_085_096, w_085_097, w_085_098, w_085_099, w_085_100, w_085_101, w_085_102, w_085_103, w_085_104, w_085_105, w_085_106, w_085_107, w_085_109, w_085_110, w_085_111, w_085_112, w_085_113, w_085_114, w_085_115, w_085_116, w_085_117, w_085_118, w_085_120, w_085_121, w_085_122, w_085_123, w_085_124, w_085_126, w_085_127, w_085_128, w_085_129, w_085_130, w_085_131, w_085_132, w_085_133, w_085_135, w_085_138, w_085_139, w_085_140, w_085_142, w_085_144, w_085_145, w_085_146, w_085_147, w_085_148, w_085_149, w_085_150, w_085_151, w_085_152, w_085_153, w_085_154, w_085_155, w_085_156, w_085_157, w_085_158, w_085_160, w_085_161, w_085_162, w_085_163, w_085_164, w_085_165, w_085_166, w_085_167, w_085_168, w_085_169, w_085_170, w_085_171, w_085_172, w_085_173, w_085_174, w_085_175, w_085_176, w_085_177, w_085_178, w_085_179, w_085_180, w_085_181, w_085_182, w_085_183, w_085_184, w_085_185, w_085_186, w_085_187, w_085_189, w_085_190, w_085_191, w_085_194, w_085_195, w_085_196, w_085_197, w_085_198, w_085_199, w_085_200, w_085_201, w_085_202, w_085_203, w_085_204, w_085_205, w_085_206, w_085_208, w_085_210, w_085_211, w_085_213, w_085_214, w_085_215, w_085_216, w_085_217, w_085_218, w_085_219, w_085_220, w_085_221, w_085_222, w_085_223, w_085_224, w_085_225, w_085_227, w_085_228, w_085_229, w_085_230, w_085_231, w_085_232, w_085_233, w_085_234, w_085_235, w_085_236, w_085_237, w_085_238, w_085_239, w_085_241, w_085_242, w_085_243, w_085_245, w_085_246, w_085_247, w_085_248, w_085_249, w_085_251, w_085_252, w_085_253, w_085_255, w_085_256, w_085_257, w_085_258, w_085_259, w_085_260, w_085_262, w_085_263, w_085_264, w_085_265, w_085_266, w_085_267, w_085_268, w_085_269, w_085_270, w_085_271, w_085_272, w_085_273, w_085_275, w_085_277, w_085_278, w_085_279, w_085_280, w_085_283, w_085_284, w_085_285, w_085_286, w_085_287, w_085_289, w_085_290, w_085_291, w_085_292, w_085_293, w_085_294, w_085_295, w_085_296, w_085_297, w_085_298, w_085_300, w_085_301, w_085_302, w_085_303, w_085_304, w_085_305, w_085_306, w_085_307, w_085_309, w_085_310, w_085_311, w_085_312, w_085_313, w_085_314, w_085_315, w_085_316, w_085_317, w_085_318, w_085_319, w_085_320, w_085_321, w_085_322, w_085_323, w_085_324, w_085_325, w_085_326, w_085_327, w_085_328, w_085_329, w_085_330, w_085_331, w_085_332, w_085_333, w_085_334, w_085_335, w_085_336, w_085_337, w_085_338, w_085_339, w_085_341, w_085_342, w_085_343, w_085_344, w_085_345, w_085_346, w_085_347, w_085_348, w_085_349, w_085_350, w_085_351, w_085_352, w_085_353, w_085_354, w_085_355, w_085_356, w_085_357, w_085_358, w_085_359, w_085_360, w_085_361, w_085_362, w_085_363, w_085_364, w_085_365, w_085_366, w_085_368, w_085_369, w_085_370, w_085_371, w_085_372, w_085_373, w_085_374, w_085_376, w_085_377, w_085_378, w_085_379, w_085_380, w_085_382, w_085_383, w_085_384, w_085_385, w_085_386, w_085_387, w_085_389, w_085_390, w_085_391, w_085_392, w_085_393, w_085_394, w_085_395, w_085_396, w_085_397, w_085_398, w_085_399, w_085_400, w_085_401, w_085_402, w_085_403, w_085_404, w_085_405, w_085_406, w_085_407, w_085_408, w_085_409, w_085_410, w_085_411, w_085_412, w_085_413, w_085_414, w_085_415, w_085_416, w_085_417, w_085_418, w_085_419, w_085_420, w_085_421, w_085_422, w_085_423, w_085_425, w_085_426, w_085_427, w_085_428, w_085_429, w_085_430, w_085_431, w_085_432, w_085_433, w_085_435, w_085_436, w_085_438, w_085_439, w_085_440, w_085_441, w_085_442, w_085_444, w_085_445, w_085_446, w_085_447, w_085_449, w_085_450, w_085_451, w_085_452, w_085_453, w_085_454, w_085_455, w_085_456, w_085_457, w_085_458, w_085_461, w_085_462, w_085_463, w_085_464, w_085_466, w_085_468, w_085_469, w_085_470, w_085_471, w_085_472, w_085_473, w_085_476, w_085_477, w_085_478, w_085_479, w_085_480, w_085_481, w_085_483, w_085_485, w_085_486, w_085_488, w_085_489, w_085_490, w_085_491, w_085_492, w_085_493, w_085_494, w_085_495, w_085_497, w_085_498, w_085_499, w_085_500, w_085_501, w_085_502, w_085_503, w_085_504, w_085_505, w_085_506, w_085_507, w_085_509, w_085_510, w_085_511, w_085_512, w_085_513, w_085_514, w_085_515, w_085_516, w_085_517, w_085_518, w_085_520, w_085_522, w_085_524, w_085_525, w_085_526, w_085_527, w_085_528, w_085_531, w_085_532, w_085_533, w_085_535, w_085_536, w_085_537, w_085_538, w_085_539, w_085_541, w_085_542, w_085_543, w_085_544, w_085_546, w_085_547, w_085_548, w_085_549, w_085_550, w_085_551, w_085_552, w_085_553, w_085_554, w_085_555, w_085_556, w_085_557, w_085_560, w_085_561, w_085_562, w_085_563, w_085_564, w_085_565, w_085_566, w_085_567, w_085_568, w_085_569, w_085_570, w_085_571, w_085_573, w_085_574, w_085_575, w_085_576, w_085_577, w_085_578, w_085_579, w_085_580, w_085_581, w_085_583, w_085_584, w_085_585, w_085_586, w_085_587, w_085_588, w_085_589, w_085_590, w_085_591, w_085_592, w_085_593, w_085_594, w_085_595, w_085_597, w_085_599, w_085_600, w_085_602, w_085_603, w_085_604, w_085_605, w_085_606, w_085_607, w_085_608, w_085_609, w_085_610, w_085_611, w_085_612, w_085_614, w_085_615, w_085_616, w_085_617, w_085_618, w_085_619, w_085_620, w_085_621, w_085_622, w_085_623, w_085_624, w_085_625, w_085_626, w_085_627, w_085_628, w_085_629, w_085_630, w_085_631, w_085_632, w_085_633, w_085_634, w_085_635, w_085_636, w_085_637, w_085_638, w_085_640, w_085_642, w_085_643, w_085_644, w_085_645, w_085_646, w_085_647, w_085_648, w_085_649, w_085_650, w_085_651, w_085_652, w_085_655, w_085_656, w_085_657, w_085_658, w_085_661, w_085_662, w_085_663, w_085_664, w_085_665, w_085_666, w_085_667, w_085_668, w_085_669, w_085_670, w_085_672, w_085_673, w_085_674, w_085_675, w_085_676, w_085_677, w_085_678, w_085_680, w_085_681, w_085_682, w_085_683, w_085_684, w_085_685, w_085_686, w_085_687, w_085_688, w_085_689, w_085_692, w_085_693, w_085_694, w_085_695, w_085_696, w_085_697, w_085_698, w_085_699, w_085_700, w_085_701, w_085_703, w_085_704, w_085_705, w_085_706, w_085_707, w_085_708, w_085_709, w_085_710, w_085_711, w_085_712, w_085_714, w_085_716, w_085_717, w_085_718, w_085_719, w_085_720, w_085_722, w_085_723, w_085_724, w_085_727, w_085_728, w_085_729, w_085_730, w_085_731, w_085_732, w_085_733, w_085_734, w_085_735, w_085_736, w_085_737, w_085_738, w_085_739, w_085_740, w_085_741, w_085_743, w_085_744, w_085_745, w_085_746, w_085_747, w_085_748, w_085_750, w_085_751, w_085_754, w_085_755, w_085_756, w_085_757, w_085_758, w_085_760, w_085_761, w_085_762, w_085_764, w_085_765, w_085_766, w_085_767, w_085_768, w_085_769, w_085_770, w_085_771, w_085_772, w_085_773, w_085_774, w_085_775, w_085_777, w_085_778, w_085_779, w_085_780, w_085_781, w_085_782, w_085_783, w_085_784, w_085_785, w_085_786, w_085_787, w_085_788, w_085_789, w_085_790, w_085_791, w_085_792, w_085_793, w_085_795, w_085_797, w_085_798, w_085_799, w_085_800, w_085_801, w_085_802, w_085_803, w_085_804, w_085_805, w_085_807, w_085_808, w_085_809, w_085_810, w_085_814, w_085_815, w_085_817, w_085_818, w_085_819, w_085_820, w_085_822, w_085_823, w_085_824, w_085_825, w_085_826, w_085_827, w_085_829, w_085_830, w_085_831, w_085_833, w_085_834, w_085_835, w_085_836, w_085_837, w_085_838, w_085_839, w_085_841, w_085_842, w_085_843, w_085_844, w_085_846, w_085_847, w_085_848, w_085_849, w_085_850, w_085_851, w_085_852, w_085_853, w_085_854, w_085_855, w_085_857, w_085_858, w_085_859, w_085_860, w_085_862, w_085_863, w_085_864, w_085_865, w_085_866, w_085_867, w_085_869, w_085_870, w_085_871, w_085_872, w_085_873, w_085_874, w_085_875, w_085_876, w_085_877, w_085_878, w_085_879, w_085_880, w_085_881, w_085_882, w_085_883, w_085_884, w_085_885, w_085_886, w_085_887, w_085_888, w_085_889, w_085_890, w_085_891, w_085_892, w_085_893, w_085_894, w_085_895, w_085_896, w_085_898, w_085_899, w_085_900, w_085_901, w_085_902, w_085_903, w_085_904, w_085_905, w_085_906, w_085_907, w_085_908, w_085_909, w_085_910, w_085_911, w_085_913, w_085_914, w_085_916, w_085_917, w_085_918, w_085_919, w_085_920, w_085_921, w_085_922, w_085_923, w_085_924, w_085_925, w_085_926, w_085_927, w_085_928, w_085_929, w_085_930, w_085_931, w_085_932, w_085_934, w_085_935, w_085_936, w_085_937, w_085_938, w_085_939, w_085_940, w_085_941, w_085_943, w_085_944, w_085_945, w_085_947, w_085_948, w_085_949, w_085_950, w_085_951, w_085_952, w_085_953, w_085_954, w_085_955, w_085_957, w_085_958, w_085_959, w_085_960, w_085_961, w_085_963, w_085_964, w_085_966, w_085_967, w_085_968, w_085_970, w_085_972, w_085_973, w_085_974, w_085_975, w_085_976, w_085_977, w_085_978, w_085_979, w_085_980, w_085_981, w_085_982, w_085_983, w_085_984, w_085_985, w_085_986, w_085_987, w_085_988, w_085_989, w_085_990, w_085_991, w_085_992, w_085_993, w_085_994, w_085_995, w_085_996, w_085_997, w_085_998, w_085_999, w_085_1000;
  wire w_086_000, w_086_001, w_086_002, w_086_003, w_086_004, w_086_005, w_086_006, w_086_007, w_086_008, w_086_009, w_086_010, w_086_011, w_086_012, w_086_013, w_086_014, w_086_015, w_086_016, w_086_017, w_086_018, w_086_019, w_086_020, w_086_021, w_086_022, w_086_023, w_086_024, w_086_025, w_086_026, w_086_027, w_086_028, w_086_029, w_086_030, w_086_031, w_086_032, w_086_033, w_086_034, w_086_035, w_086_036, w_086_037, w_086_038, w_086_039, w_086_040, w_086_041, w_086_042, w_086_043, w_086_044, w_086_045, w_086_046, w_086_047, w_086_048, w_086_049, w_086_050, w_086_051, w_086_052, w_086_053, w_086_054, w_086_055, w_086_056, w_086_057, w_086_058, w_086_059, w_086_060, w_086_061, w_086_062, w_086_063, w_086_064, w_086_065, w_086_066, w_086_067, w_086_068, w_086_069, w_086_070, w_086_071, w_086_072, w_086_073, w_086_074, w_086_075, w_086_076, w_086_077, w_086_078, w_086_079, w_086_080, w_086_081, w_086_082, w_086_083, w_086_084, w_086_085, w_086_086, w_086_087, w_086_088, w_086_089, w_086_090, w_086_091, w_086_092, w_086_093, w_086_094, w_086_095, w_086_096, w_086_097, w_086_098, w_086_099, w_086_100, w_086_101, w_086_102, w_086_103, w_086_104, w_086_105, w_086_106, w_086_107, w_086_108, w_086_109, w_086_110, w_086_111, w_086_112, w_086_113, w_086_114, w_086_115, w_086_116, w_086_117, w_086_118, w_086_119, w_086_120, w_086_121, w_086_122, w_086_123, w_086_124, w_086_125, w_086_126, w_086_127, w_086_128, w_086_129, w_086_130, w_086_131, w_086_132, w_086_133, w_086_134, w_086_135, w_086_136, w_086_137, w_086_138, w_086_139, w_086_140, w_086_141, w_086_142, w_086_143, w_086_144, w_086_145, w_086_146, w_086_147, w_086_148, w_086_149, w_086_150, w_086_151, w_086_152, w_086_153, w_086_154, w_086_155, w_086_156, w_086_157, w_086_158, w_086_159, w_086_160, w_086_161, w_086_162, w_086_163, w_086_164, w_086_165, w_086_166, w_086_167, w_086_168, w_086_169, w_086_170, w_086_171, w_086_172, w_086_173, w_086_174, w_086_176, w_086_177, w_086_178, w_086_179, w_086_180, w_086_181, w_086_182, w_086_183, w_086_184, w_086_185, w_086_186, w_086_187, w_086_188, w_086_189, w_086_190, w_086_191, w_086_192, w_086_193, w_086_194, w_086_195, w_086_196, w_086_197, w_086_198, w_086_199, w_086_200, w_086_201, w_086_202, w_086_203, w_086_204, w_086_205, w_086_206, w_086_207, w_086_208, w_086_209, w_086_210, w_086_211, w_086_212, w_086_213, w_086_214, w_086_215, w_086_216, w_086_217, w_086_218, w_086_219, w_086_220, w_086_221, w_086_222, w_086_223, w_086_224, w_086_225, w_086_226, w_086_227, w_086_228, w_086_229, w_086_230, w_086_231, w_086_232, w_086_233, w_086_234, w_086_235, w_086_236, w_086_237, w_086_238, w_086_239, w_086_240, w_086_241, w_086_242, w_086_243, w_086_244, w_086_245, w_086_246, w_086_247, w_086_248, w_086_249, w_086_250, w_086_251, w_086_252, w_086_253, w_086_254, w_086_255, w_086_256, w_086_257, w_086_258, w_086_259, w_086_260, w_086_261, w_086_262, w_086_263, w_086_264, w_086_265, w_086_266, w_086_267, w_086_268, w_086_269, w_086_270, w_086_271, w_086_272, w_086_273, w_086_274, w_086_275, w_086_276, w_086_277, w_086_278, w_086_279, w_086_280, w_086_281, w_086_282, w_086_283, w_086_284, w_086_285, w_086_286, w_086_287, w_086_288, w_086_289, w_086_290, w_086_291, w_086_292, w_086_293;
  wire w_087_000, w_087_001, w_087_002, w_087_006, w_087_010, w_087_012, w_087_016, w_087_019, w_087_020, w_087_023, w_087_026, w_087_028, w_087_029, w_087_030, w_087_031, w_087_032, w_087_033, w_087_034, w_087_036, w_087_037, w_087_038, w_087_039, w_087_041, w_087_044, w_087_045, w_087_046, w_087_050, w_087_052, w_087_053, w_087_054, w_087_057, w_087_058, w_087_059, w_087_060, w_087_066, w_087_068, w_087_071, w_087_074, w_087_078, w_087_080, w_087_081, w_087_086, w_087_088, w_087_092, w_087_097, w_087_098, w_087_101, w_087_102, w_087_104, w_087_107, w_087_114, w_087_115, w_087_117, w_087_118, w_087_124, w_087_126, w_087_128, w_087_129, w_087_130, w_087_132, w_087_133, w_087_136, w_087_139, w_087_140, w_087_141, w_087_142, w_087_145, w_087_154, w_087_155, w_087_160, w_087_165, w_087_167, w_087_179, w_087_180, w_087_181, w_087_183, w_087_189, w_087_190, w_087_191, w_087_193, w_087_201, w_087_209, w_087_217, w_087_218, w_087_221, w_087_226, w_087_227, w_087_228, w_087_230, w_087_234, w_087_236, w_087_237, w_087_239, w_087_241, w_087_244, w_087_246, w_087_249, w_087_252, w_087_255, w_087_256, w_087_257, w_087_264, w_087_265, w_087_267, w_087_273, w_087_277, w_087_281, w_087_286, w_087_287, w_087_288, w_087_289, w_087_291, w_087_296, w_087_297, w_087_298, w_087_300, w_087_307, w_087_310, w_087_314, w_087_317, w_087_318, w_087_319, w_087_323, w_087_327, w_087_330, w_087_335, w_087_342, w_087_344, w_087_349, w_087_351, w_087_353, w_087_356, w_087_357, w_087_361, w_087_364, w_087_365, w_087_369, w_087_370, w_087_371, w_087_372, w_087_374, w_087_375, w_087_377, w_087_378, w_087_379, w_087_380, w_087_381, w_087_390, w_087_392, w_087_393, w_087_402, w_087_407, w_087_408, w_087_414, w_087_415, w_087_416, w_087_417, w_087_420, w_087_424, w_087_425, w_087_431, w_087_432, w_087_433, w_087_435, w_087_437, w_087_438, w_087_440, w_087_443, w_087_448, w_087_450, w_087_451, w_087_456, w_087_457, w_087_458, w_087_461, w_087_467, w_087_470, w_087_472, w_087_473, w_087_477, w_087_487, w_087_492, w_087_493, w_087_494, w_087_495, w_087_496, w_087_497, w_087_500, w_087_502, w_087_503, w_087_506, w_087_511, w_087_516, w_087_519, w_087_526, w_087_534, w_087_535, w_087_541, w_087_542, w_087_543, w_087_545, w_087_546, w_087_547, w_087_548, w_087_549, w_087_551, w_087_552, w_087_556, w_087_567, w_087_572, w_087_573, w_087_577, w_087_581, w_087_584, w_087_586, w_087_587, w_087_594, w_087_598, w_087_601, w_087_603, w_087_606, w_087_607, w_087_608, w_087_609, w_087_618, w_087_619, w_087_620, w_087_622, w_087_624, w_087_626, w_087_627, w_087_633, w_087_638, w_087_639, w_087_641, w_087_643, w_087_645, w_087_647, w_087_648, w_087_650, w_087_651, w_087_652, w_087_653, w_087_654, w_087_656, w_087_664, w_087_665, w_087_667, w_087_668, w_087_669, w_087_672, w_087_676, w_087_677, w_087_678, w_087_683, w_087_699, w_087_700, w_087_704, w_087_706, w_087_710, w_087_713, w_087_716, w_087_717, w_087_723, w_087_724, w_087_725, w_087_730, w_087_731, w_087_739, w_087_743, w_087_745, w_087_746, w_087_752, w_087_753, w_087_754, w_087_756, w_087_760, w_087_761, w_087_764, w_087_765, w_087_767, w_087_770, w_087_771, w_087_782, w_087_785, w_087_789, w_087_791, w_087_796, w_087_797, w_087_798, w_087_799, w_087_800, w_087_801, w_087_804, w_087_805, w_087_814, w_087_817, w_087_818, w_087_826, w_087_831, w_087_832, w_087_846, w_087_847, w_087_848, w_087_850, w_087_854, w_087_856, w_087_858, w_087_863, w_087_866, w_087_875, w_087_878, w_087_880, w_087_881, w_087_882, w_087_884, w_087_888, w_087_891, w_087_892, w_087_900, w_087_902, w_087_903, w_087_904, w_087_905, w_087_909, w_087_916, w_087_917, w_087_922, w_087_924, w_087_931, w_087_932, w_087_933, w_087_934, w_087_938, w_087_943, w_087_946, w_087_948, w_087_951, w_087_956, w_087_957, w_087_959, w_087_963, w_087_967, w_087_970, w_087_971, w_087_972, w_087_976, w_087_977, w_087_989, w_087_993, w_087_998, w_087_999, w_087_1000, w_087_1005, w_087_1008, w_087_1013, w_087_1014, w_087_1022, w_087_1023, w_087_1026, w_087_1029, w_087_1030, w_087_1034, w_087_1036, w_087_1038, w_087_1039, w_087_1043, w_087_1045, w_087_1049, w_087_1052, w_087_1054, w_087_1059, w_087_1061, w_087_1066, w_087_1069, w_087_1074, w_087_1085, w_087_1086, w_087_1087, w_087_1096, w_087_1097, w_087_1100, w_087_1104, w_087_1105, w_087_1107, w_087_1115, w_087_1116, w_087_1118, w_087_1121, w_087_1124, w_087_1131, w_087_1132, w_087_1135, w_087_1136, w_087_1140, w_087_1143, w_087_1146, w_087_1147, w_087_1152, w_087_1153, w_087_1154, w_087_1158, w_087_1159, w_087_1166, w_087_1168, w_087_1169, w_087_1170, w_087_1171, w_087_1177, w_087_1182, w_087_1183, w_087_1188, w_087_1190, w_087_1192, w_087_1195, w_087_1196, w_087_1198, w_087_1199, w_087_1201, w_087_1204, w_087_1206, w_087_1208, w_087_1210, w_087_1215, w_087_1219, w_087_1220, w_087_1221, w_087_1228, w_087_1229, w_087_1230, w_087_1233, w_087_1236, w_087_1239, w_087_1240, w_087_1242, w_087_1246, w_087_1252, w_087_1255, w_087_1256, w_087_1257, w_087_1263, w_087_1267, w_087_1268, w_087_1274, w_087_1275, w_087_1276, w_087_1278, w_087_1281, w_087_1282, w_087_1287, w_087_1292, w_087_1298, w_087_1301, w_087_1304, w_087_1307, w_087_1309, w_087_1311, w_087_1312, w_087_1316, w_087_1318, w_087_1319, w_087_1324, w_087_1326, w_087_1327, w_087_1329, w_087_1331, w_087_1334, w_087_1337, w_087_1339, w_087_1346, w_087_1347, w_087_1351, w_087_1353, w_087_1354, w_087_1360, w_087_1362, w_087_1366, w_087_1370, w_087_1373, w_087_1376, w_087_1380, w_087_1388, w_087_1390, w_087_1391, w_087_1392, w_087_1395, w_087_1399, w_087_1401, w_087_1403, w_087_1404, w_087_1408, w_087_1418, w_087_1421, w_087_1422, w_087_1425, w_087_1426, w_087_1428, w_087_1434, w_087_1436, w_087_1440, w_087_1445, w_087_1448, w_087_1449, w_087_1451, w_087_1456, w_087_1460, w_087_1467, w_087_1468, w_087_1469, w_087_1472, w_087_1473, w_087_1475, w_087_1477, w_087_1478, w_087_1482, w_087_1484, w_087_1491, w_087_1495, w_087_1496, w_087_1498, w_087_1500, w_087_1501, w_087_1502, w_087_1504, w_087_1507, w_087_1510, w_087_1517, w_087_1520, w_087_1529, w_087_1530, w_087_1540, w_087_1541, w_087_1544, w_087_1547, w_087_1548, w_087_1549, w_087_1557, w_087_1565, w_087_1566, w_087_1567, w_087_1573, w_087_1574, w_087_1576, w_087_1581, w_087_1585, w_087_1589, w_087_1596, w_087_1597, w_087_1604, w_087_1605, w_087_1606, w_087_1607, w_087_1609, w_087_1611, w_087_1612, w_087_1616, w_087_1620, w_087_1622, w_087_1633, w_087_1635, w_087_1636, w_087_1637, w_087_1641, w_087_1642, w_087_1645, w_087_1647, w_087_1649, w_087_1653, w_087_1656, w_087_1662, w_087_1673, w_087_1675, w_087_1676, w_087_1678, w_087_1679, w_087_1685, w_087_1692, w_087_1693, w_087_1695, w_087_1697, w_087_1700, w_087_1702, w_087_1703, w_087_1705, w_087_1706, w_087_1711, w_087_1714, w_087_1716, w_087_1721, w_087_1722, w_087_1727, w_087_1728, w_087_1729, w_087_1731, w_087_1733, w_087_1737, w_087_1739, w_087_1745, w_087_1746, w_087_1748, w_087_1753, w_087_1759, w_087_1767, w_087_1769, w_087_1774, w_087_1777, w_087_1780, w_087_1781, w_087_1784, w_087_1787, w_087_1790, w_087_1793, w_087_1797, w_087_1798, w_087_1802, w_087_1804, w_087_1807, w_087_1808, w_087_1811, w_087_1814, w_087_1815, w_087_1816, w_087_1817, w_087_1818, w_087_1819, w_087_1820, w_087_1827, w_087_1830, w_087_1831, w_087_1834, w_087_1838, w_087_1841, w_087_1846, w_087_1849, w_087_1854, w_087_1857, w_087_1858, w_087_1859, w_087_1861, w_087_1862, w_087_1863, w_087_1868, w_087_1870, w_087_1873, w_087_1882, w_087_1887, w_087_1888, w_087_1901, w_087_1902, w_087_1907, w_087_1909, w_087_1910, w_087_1912, w_087_1914, w_087_1917, w_087_1922, w_087_1930, w_087_1932, w_087_1933, w_087_1938, w_087_1946, w_087_1947, w_087_1948, w_087_1949, w_087_1950, w_087_1951, w_087_1952, w_087_1953, w_087_1954, w_087_1956, w_087_1957, w_087_1961, w_087_1962, w_087_1963, w_087_1964, w_087_1965, w_087_1966, w_087_1967, w_087_1968, w_087_1970, w_087_1974, w_087_1978, w_087_1979, w_087_1980, w_087_1981, w_087_1982, w_087_1984, w_087_1986, w_087_1987, w_087_1989, w_087_1999, w_087_2001, w_087_2004, w_087_2006, w_087_2011, w_087_2013, w_087_2014, w_087_2015, w_087_2016, w_087_2020, w_087_2022, w_087_2027, w_087_2028, w_087_2032, w_087_2034, w_087_2040, w_087_2041, w_087_2045, w_087_2046, w_087_2047, w_087_2052, w_087_2054, w_087_2057, w_087_2060, w_087_2062, w_087_2064, w_087_2065, w_087_2068, w_087_2069, w_087_2072, w_087_2074, w_087_2076, w_087_2077, w_087_2078, w_087_2082, w_087_2084, w_087_2091, w_087_2092, w_087_2096, w_087_2097, w_087_2106, w_087_2111, w_087_2114, w_087_2115, w_087_2117, w_087_2118, w_087_2127, w_087_2133, w_087_2135, w_087_2138, w_087_2141, w_087_2147, w_087_2149, w_087_2153, w_087_2154, w_087_2161, w_087_2162, w_087_2166, w_087_2167, w_087_2168, w_087_2170, w_087_2172, w_087_2179, w_087_2181, w_087_2183, w_087_2184, w_087_2185, w_087_2192, w_087_2193, w_087_2195, w_087_2197, w_087_2199, w_087_2204, w_087_2207, w_087_2212, w_087_2213, w_087_2214, w_087_2215, w_087_2216, w_087_2219, w_087_2220, w_087_2229, w_087_2235, w_087_2237, w_087_2238, w_087_2239, w_087_2243, w_087_2244, w_087_2248, w_087_2250, w_087_2251, w_087_2255, w_087_2259, w_087_2261, w_087_2265, w_087_2268, w_087_2269, w_087_2272, w_087_2274, w_087_2278, w_087_2281, w_087_2282, w_087_2283, w_087_2289, w_087_2290, w_087_2291, w_087_2294, w_087_2295, w_087_2298, w_087_2305, w_087_2308, w_087_2309, w_087_2313, w_087_2321, w_087_2325, w_087_2326, w_087_2328, w_087_2329, w_087_2330, w_087_2331, w_087_2335, w_087_2337, w_087_2348, w_087_2355, w_087_2356, w_087_2357, w_087_2362, w_087_2363, w_087_2365, w_087_2370, w_087_2373, w_087_2378, w_087_2382, w_087_2387, w_087_2388, w_087_2389, w_087_2390, w_087_2396, w_087_2400, w_087_2401, w_087_2410, w_087_2413, w_087_2415, w_087_2418, w_087_2419, w_087_2424, w_087_2425, w_087_2430, w_087_2431, w_087_2432, w_087_2435, w_087_2438, w_087_2439, w_087_2441, w_087_2442, w_087_2443, w_087_2447, w_087_2448, w_087_2450, w_087_2452, w_087_2456, w_087_2457, w_087_2461, w_087_2463, w_087_2464, w_087_2466, w_087_2468, w_087_2469, w_087_2471, w_087_2475, w_087_2477, w_087_2482, w_087_2489, w_087_2492, w_087_2495, w_087_2499, w_087_2500, w_087_2513, w_087_2515, w_087_2516, w_087_2517, w_087_2519, w_087_2529, w_087_2531, w_087_2535, w_087_2536, w_087_2540, w_087_2542, w_087_2546, w_087_2551, w_087_2555, w_087_2558, w_087_2566, w_087_2570, w_087_2572, w_087_2573, w_087_2574, w_087_2579, w_087_2597, w_087_2598, w_087_2599, w_087_2602, w_087_2606, w_087_2611, w_087_2613, w_087_2615, w_087_2632, w_087_2642, w_087_2644, w_087_2648, w_087_2649, w_087_2651, w_087_2654, w_087_2656, w_087_2664, w_087_2665, w_087_2667, w_087_2672, w_087_2674, w_087_2685, w_087_2687, w_087_2699, w_087_2700, w_087_2702, w_087_2703, w_087_2706, w_087_2711, w_087_2714, w_087_2715, w_087_2724, w_087_2728, w_087_2733, w_087_2737, w_087_2740, w_087_2741, w_087_2748, w_087_2753, w_087_2757, w_087_2758, w_087_2763, w_087_2764, w_087_2765, w_087_2767, w_087_2773, w_087_2776, w_087_2778, w_087_2780, w_087_2787, w_087_2797, w_087_2799, w_087_2801, w_087_2804, w_087_2807, w_087_2810, w_087_2818, w_087_2828, w_087_2829, w_087_2831, w_087_2834, w_087_2835, w_087_2838, w_087_2840, w_087_2841, w_087_2842, w_087_2848, w_087_2850, w_087_2861, w_087_2862, w_087_2865, w_087_2866, w_087_2867, w_087_2868, w_087_2869, w_087_2875, w_087_2876, w_087_2877, w_087_2882, w_087_2884, w_087_2888, w_087_2889, w_087_2890, w_087_2894, w_087_2896, w_087_2899, w_087_2904, w_087_2915, w_087_2916, w_087_2917, w_087_2919, w_087_2920, w_087_2921, w_087_2923, w_087_2926, w_087_2930, w_087_2932, w_087_2935, w_087_2937, w_087_2940, w_087_2945, w_087_2947, w_087_2948, w_087_2958, w_087_2960, w_087_2963, w_087_2975, w_087_2976, w_087_2983, w_087_2985, w_087_2987, w_087_2991, w_087_2993, w_087_2995, w_087_2996, w_087_2999, w_087_3003, w_087_3004, w_087_3005, w_087_3010, w_087_3014, w_087_3016, w_087_3019, w_087_3032, w_087_3035, w_087_3036, w_087_3040, w_087_3041, w_087_3049, w_087_3050, w_087_3055, w_087_3056, w_087_3058, w_087_3060, w_087_3063, w_087_3068, w_087_3069, w_087_3070, w_087_3072, w_087_3073, w_087_3078, w_087_3079, w_087_3081, w_087_3082, w_087_3083, w_087_3086, w_087_3088, w_087_3089, w_087_3090, w_087_3095, w_087_3097, w_087_3098, w_087_3100, w_087_3102, w_087_3104, w_087_3108, w_087_3113, w_087_3116, w_087_3117, w_087_3119, w_087_3126, w_087_3127, w_087_3132, w_087_3133, w_087_3136, w_087_3143, w_087_3147, w_087_3156, w_087_3158, w_087_3167, w_087_3170, w_087_3176, w_087_3177, w_087_3181, w_087_3182, w_087_3183, w_087_3186, w_087_3187, w_087_3189, w_087_3198, w_087_3205, w_087_3207, w_087_3208, w_087_3216, w_087_3223, w_087_3227, w_087_3228, w_087_3229, w_087_3230, w_087_3233, w_087_3234, w_087_3236, w_087_3238, w_087_3239, w_087_3241, w_087_3243, w_087_3245, w_087_3247, w_087_3248, w_087_3250, w_087_3252, w_087_3253, w_087_3257, w_087_3259, w_087_3263, w_087_3271, w_087_3273, w_087_3274, w_087_3277, w_087_3278, w_087_3281, w_087_3288, w_087_3295, w_087_3296, w_087_3299, w_087_3304, w_087_3305, w_087_3309, w_087_3310, w_087_3314, w_087_3321, w_087_3322, w_087_3323, w_087_3324, w_087_3326, w_087_3329, w_087_3332, w_087_3333, w_087_3336, w_087_3337, w_087_3340, w_087_3342, w_087_3343, w_087_3344, w_087_3346, w_087_3347, w_087_3351, w_087_3356, w_087_3360, w_087_3365, w_087_3372, w_087_3375, w_087_3376, w_087_3383, w_087_3390, w_087_3392, w_087_3395, w_087_3396, w_087_3398, w_087_3400, w_087_3402, w_087_3406, w_087_3411, w_087_3417, w_087_3423, w_087_3427, w_087_3431, w_087_3433, w_087_3438, w_087_3445, w_087_3446, w_087_3448, w_087_3449, w_087_3450, w_087_3452, w_087_3458, w_087_3459, w_087_3471, w_087_3472, w_087_3474, w_087_3476, w_087_3477, w_087_3478, w_087_3484, w_087_3492, w_087_3494, w_087_3495, w_087_3497, w_087_3502, w_087_3503, w_087_3505, w_087_3506, w_087_3508, w_087_3512, w_087_3518, w_087_3520, w_087_3521, w_087_3523, w_087_3524, w_087_3530, w_087_3531, w_087_3537, w_087_3540, w_087_3541, w_087_3544, w_087_3545, w_087_3546, w_087_3551, w_087_3553, w_087_3554, w_087_3557, w_087_3560, w_087_3561, w_087_3562, w_087_3564, w_087_3565, w_087_3570, w_087_3574, w_087_3576, w_087_3577, w_087_3580, w_087_3583, w_087_3585, w_087_3588, w_087_3589, w_087_3590, w_087_3591, w_087_3598, w_087_3601, w_087_3608, w_087_3614, w_087_3620, w_087_3622, w_087_3623, w_087_3640, w_087_3643, w_087_3648, w_087_3649, w_087_3650, w_087_3651, w_087_3654, w_087_3660, w_087_3663, w_087_3666, w_087_3667, w_087_3668, w_087_3669, w_087_3681, w_087_3685, w_087_3690, w_087_3691, w_087_3694, w_087_3697, w_087_3701, w_087_3703, w_087_3705, w_087_3706, w_087_3707, w_087_3709, w_087_3713, w_087_3718, w_087_3728, w_087_3732, w_087_3735, w_087_3737, w_087_3739, w_087_3743, w_087_3744, w_087_3748, w_087_3753, w_087_3755, w_087_3759, w_087_3761, w_087_3762, w_087_3763, w_087_3765, w_087_3773, w_087_3779, w_087_3781, w_087_3782, w_087_3786, w_087_3789, w_087_3790, w_087_3792, w_087_3795, w_087_3799, w_087_3803, w_087_3807, w_087_3816, w_087_3818, w_087_3819, w_087_3822, w_087_3826, w_087_3827, w_087_3832, w_087_3835, w_087_3854, w_087_3855, w_087_3856, w_087_3858, w_087_3866, w_087_3868, w_087_3878, w_087_3882, w_087_3888, w_087_3892, w_087_3895, w_087_3896, w_087_3897, w_087_3903, w_087_3904, w_087_3906, w_087_3910, w_087_3914, w_087_3916, w_087_3917, w_087_3923, w_087_3926, w_087_3927, w_087_3929, w_087_3930, w_087_3931, w_087_3932, w_087_3934, w_087_3938, w_087_3942, w_087_3943, w_087_3946, w_087_3950, w_087_3955, w_087_3958, w_087_3959, w_087_3960, w_087_3963, w_087_3964, w_087_3972, w_087_3974, w_087_3977, w_087_3979, w_087_3983, w_087_3984, w_087_3989, w_087_3992, w_087_3993, w_087_3994, w_087_3997, w_087_4001, w_087_4002, w_087_4003, w_087_4005, w_087_4008, w_087_4017, w_087_4019, w_087_4022, w_087_4026, w_087_4027, w_087_4030, w_087_4031, w_087_4040, w_087_4041, w_087_4045, w_087_4052, w_087_4053, w_087_4055, w_087_4056, w_087_4057, w_087_4059, w_087_4061, w_087_4062, w_087_4064, w_087_4066, w_087_4069, w_087_4073, w_087_4075, w_087_4076, w_087_4077, w_087_4080, w_087_4082, w_087_4086, w_087_4091, w_087_4092, w_087_4093, w_087_4097, w_087_4101, w_087_4102, w_087_4105, w_087_4106, w_087_4108, w_087_4109, w_087_4110, w_087_4111, w_087_4112, w_087_4113, w_087_4115, w_087_4116, w_087_4117, w_087_4119, w_087_4121, w_087_4127, w_087_4129, w_087_4130, w_087_4132, w_087_4135, w_087_4136, w_087_4145, w_087_4149, w_087_4152, w_087_4159, w_087_4161, w_087_4163, w_087_4166, w_087_4171, w_087_4177, w_087_4179, w_087_4188, w_087_4189, w_087_4196, w_087_4202, w_087_4205, w_087_4210, w_087_4211, w_087_4220, w_087_4226, w_087_4227, w_087_4228, w_087_4231, w_087_4232, w_087_4234, w_087_4235, w_087_4241, w_087_4242, w_087_4246, w_087_4247, w_087_4248, w_087_4250, w_087_4260, w_087_4268, w_087_4269, w_087_4270, w_087_4273, w_087_4274, w_087_4277, w_087_4278, w_087_4284, w_087_4291, w_087_4296, w_087_4303, w_087_4305, w_087_4306, w_087_4311, w_087_4312, w_087_4316, w_087_4317, w_087_4329, w_087_4330, w_087_4332, w_087_4334, w_087_4335, w_087_4339, w_087_4340, w_087_4342, w_087_4344, w_087_4345, w_087_4359, w_087_4361, w_087_4362, w_087_4364, w_087_4367, w_087_4375, w_087_4378, w_087_4379, w_087_4395, w_087_4397, w_087_4398, w_087_4399, w_087_4415, w_087_4416, w_087_4419, w_087_4420, w_087_4421, w_087_4422, w_087_4427, w_087_4430, w_087_4431, w_087_4432, w_087_4437, w_087_4441, w_087_4442, w_087_4445, w_087_4448, w_087_4452, w_087_4453, w_087_4456, w_087_4459, w_087_4462, w_087_4463, w_087_4465, w_087_4466, w_087_4471, w_087_4473, w_087_4479, w_087_4484, w_087_4486, w_087_4489, w_087_4492, w_087_4501, w_087_4503, w_087_4504, w_087_4505, w_087_4510, w_087_4512, w_087_4514, w_087_4516, w_087_4518, w_087_4524, w_087_4525, w_087_4526, w_087_4527, w_087_4529, w_087_4531, w_087_4532, w_087_4534, w_087_4538, w_087_4545, w_087_4546, w_087_4553, w_087_4556, w_087_4558, w_087_4561, w_087_4562, w_087_4568, w_087_4571, w_087_4574, w_087_4575, w_087_4586, w_087_4589, w_087_4590, w_087_4593, w_087_4595, w_087_4596, w_087_4597, w_087_4602, w_087_4603, w_087_4605, w_087_4607, w_087_4611, w_087_4612, w_087_4613, w_087_4619, w_087_4629, w_087_4630, w_087_4634, w_087_4637, w_087_4640, w_087_4642, w_087_4644, w_087_4652, w_087_4659, w_087_4660, w_087_4661, w_087_4665, w_087_4669, w_087_4670, w_087_4674, w_087_4680, w_087_4683, w_087_4689, w_087_4690, w_087_4692, w_087_4695, w_087_4698, w_087_4699, w_087_4702, w_087_4705, w_087_4706, w_087_4707, w_087_4710, w_087_4723, w_087_4726, w_087_4730, w_087_4731, w_087_4735, w_087_4736, w_087_4737, w_087_4740, w_087_4742, w_087_4744, w_087_4745, w_087_4753, w_087_4755, w_087_4762, w_087_4764, w_087_4766, w_087_4767, w_087_4768, w_087_4774, w_087_4777, w_087_4778, w_087_4780, w_087_4781, w_087_4783, w_087_4785, w_087_4794, w_087_4796, w_087_4806, w_087_4811, w_087_4813, w_087_4815, w_087_4816, w_087_4819, w_087_4820, w_087_4824, w_087_4825, w_087_4827, w_087_4830, w_087_4833, w_087_4837, w_087_4843, w_087_4844, w_087_4847, w_087_4848, w_087_4853, w_087_4858, w_087_4860, w_087_4863, w_087_4871, w_087_4873, w_087_4877, w_087_4878, w_087_4880, w_087_4881, w_087_4884, w_087_4888, w_087_4890, w_087_4892, w_087_4899, w_087_4901, w_087_4904, w_087_4906, w_087_4908, w_087_4912, w_087_4922, w_087_4924, w_087_4925, w_087_4927, w_087_4934, w_087_4938, w_087_4940, w_087_4942, w_087_4945, w_087_4947, w_087_4948, w_087_4949, w_087_4950, w_087_4951, w_087_4953, w_087_4955, w_087_4956, w_087_4957, w_087_4958, w_087_4959, w_087_4960, w_087_4961, w_087_4962, w_087_4963, w_087_4964, w_087_4965, w_087_4967;
  wire w_088_001, w_088_003, w_088_004, w_088_005, w_088_008, w_088_009, w_088_011, w_088_013, w_088_016, w_088_017, w_088_018, w_088_019, w_088_020, w_088_022, w_088_023, w_088_026, w_088_027, w_088_028, w_088_029, w_088_030, w_088_031, w_088_033, w_088_034, w_088_036, w_088_039, w_088_040, w_088_041, w_088_042, w_088_046, w_088_047, w_088_048, w_088_051, w_088_053, w_088_056, w_088_059, w_088_062, w_088_063, w_088_064, w_088_065, w_088_066, w_088_067, w_088_072, w_088_074, w_088_077, w_088_079, w_088_081, w_088_082, w_088_083, w_088_084, w_088_090, w_088_093, w_088_094, w_088_095, w_088_096, w_088_097, w_088_098, w_088_099, w_088_100, w_088_103, w_088_104, w_088_105, w_088_106, w_088_111, w_088_115, w_088_117, w_088_118, w_088_120, w_088_123, w_088_127, w_088_128, w_088_130, w_088_131, w_088_132, w_088_133, w_088_137, w_088_142, w_088_143, w_088_144, w_088_147, w_088_149, w_088_151, w_088_154, w_088_155, w_088_158, w_088_161, w_088_165, w_088_166, w_088_167, w_088_169, w_088_170, w_088_171, w_088_173, w_088_175, w_088_176, w_088_177, w_088_179, w_088_180, w_088_184, w_088_185, w_088_188, w_088_189, w_088_190, w_088_191, w_088_192, w_088_193, w_088_199, w_088_200, w_088_201, w_088_204, w_088_205, w_088_206, w_088_207, w_088_208, w_088_210, w_088_211, w_088_212, w_088_215, w_088_218, w_088_219, w_088_222, w_088_224, w_088_226, w_088_227, w_088_231, w_088_232, w_088_234, w_088_235, w_088_236, w_088_238, w_088_240, w_088_241, w_088_242, w_088_245, w_088_246, w_088_247, w_088_250, w_088_251, w_088_253, w_088_254, w_088_256, w_088_265, w_088_268, w_088_271, w_088_272, w_088_273, w_088_275, w_088_276, w_088_277, w_088_279, w_088_280, w_088_281, w_088_283, w_088_285, w_088_287, w_088_288, w_088_291, w_088_292, w_088_293, w_088_295, w_088_296, w_088_297, w_088_298, w_088_301, w_088_302, w_088_304, w_088_306, w_088_308, w_088_310, w_088_319, w_088_321, w_088_327, w_088_328, w_088_334, w_088_335, w_088_337, w_088_338, w_088_340, w_088_341, w_088_343, w_088_345, w_088_348, w_088_350, w_088_351, w_088_352, w_088_354, w_088_355, w_088_356, w_088_360, w_088_362, w_088_363, w_088_364, w_088_369, w_088_372, w_088_374, w_088_375, w_088_377, w_088_379, w_088_380, w_088_382, w_088_390, w_088_391, w_088_392, w_088_394, w_088_395, w_088_396, w_088_397, w_088_398, w_088_403, w_088_404, w_088_405, w_088_409, w_088_411, w_088_412, w_088_415, w_088_416, w_088_417, w_088_418, w_088_421, w_088_423, w_088_424, w_088_426, w_088_427, w_088_428, w_088_429, w_088_430, w_088_432, w_088_433, w_088_434, w_088_436, w_088_437, w_088_438, w_088_439, w_088_440, w_088_443, w_088_445, w_088_446, w_088_447, w_088_448, w_088_449, w_088_450, w_088_452, w_088_453, w_088_455, w_088_456, w_088_458, w_088_464, w_088_466, w_088_467, w_088_469, w_088_471, w_088_472, w_088_474, w_088_480, w_088_481, w_088_483, w_088_484, w_088_489, w_088_490, w_088_493, w_088_495, w_088_497, w_088_499, w_088_500, w_088_501, w_088_502, w_088_503, w_088_504, w_088_505, w_088_507, w_088_509, w_088_512, w_088_513, w_088_514, w_088_520, w_088_522, w_088_524, w_088_525, w_088_528, w_088_530, w_088_531, w_088_533, w_088_535, w_088_536, w_088_537, w_088_538, w_088_539, w_088_540, w_088_541, w_088_543, w_088_546, w_088_547, w_088_549, w_088_551, w_088_552, w_088_553, w_088_555, w_088_556, w_088_557, w_088_558, w_088_560, w_088_561, w_088_562, w_088_563, w_088_567, w_088_569, w_088_570, w_088_571, w_088_572, w_088_573, w_088_579, w_088_580, w_088_581, w_088_583, w_088_584, w_088_585, w_088_586, w_088_587, w_088_588, w_088_589, w_088_591, w_088_592, w_088_593, w_088_598, w_088_600, w_088_601, w_088_603, w_088_604, w_088_605, w_088_606, w_088_609, w_088_614, w_088_615, w_088_616, w_088_620, w_088_623, w_088_625, w_088_626, w_088_627, w_088_628, w_088_629, w_088_631, w_088_632, w_088_633, w_088_636, w_088_637, w_088_640, w_088_641, w_088_644, w_088_645, w_088_647, w_088_648, w_088_649, w_088_650, w_088_651, w_088_652, w_088_653, w_088_654, w_088_655, w_088_658, w_088_660, w_088_662, w_088_663, w_088_664, w_088_668, w_088_669, w_088_670, w_088_676, w_088_677, w_088_678, w_088_680, w_088_682, w_088_684, w_088_686, w_088_688, w_088_689, w_088_691, w_088_697, w_088_699, w_088_700, w_088_702, w_088_704, w_088_705, w_088_706, w_088_707, w_088_709, w_088_710, w_088_711, w_088_712, w_088_713, w_088_714, w_088_715, w_088_719, w_088_720, w_088_721, w_088_722, w_088_724, w_088_726, w_088_727, w_088_729, w_088_733, w_088_738, w_088_739, w_088_741, w_088_746, w_088_748, w_088_749, w_088_750, w_088_753, w_088_754, w_088_756, w_088_758, w_088_761, w_088_764, w_088_765, w_088_766, w_088_768, w_088_772, w_088_774, w_088_776, w_088_778, w_088_783, w_088_784, w_088_786, w_088_788, w_088_791, w_088_792, w_088_793, w_088_794, w_088_797, w_088_800, w_088_801, w_088_802, w_088_804, w_088_806, w_088_808, w_088_809, w_088_810, w_088_811, w_088_814, w_088_818, w_088_819, w_088_820, w_088_821, w_088_823, w_088_824, w_088_826, w_088_827, w_088_828, w_088_831, w_088_832, w_088_834, w_088_837, w_088_838, w_088_840, w_088_841, w_088_843, w_088_844, w_088_845, w_088_846, w_088_850, w_088_853, w_088_854, w_088_855, w_088_858, w_088_859, w_088_864, w_088_866, w_088_869, w_088_871, w_088_875, w_088_876, w_088_878, w_088_881, w_088_882, w_088_883, w_088_884, w_088_886, w_088_887, w_088_888, w_088_890, w_088_892, w_088_893, w_088_895, w_088_896, w_088_897, w_088_898, w_088_900, w_088_902, w_088_905, w_088_906, w_088_907, w_088_909, w_088_913, w_088_917, w_088_918, w_088_920, w_088_922, w_088_923, w_088_929, w_088_933, w_088_934, w_088_935, w_088_936, w_088_937, w_088_942, w_088_943, w_088_947, w_088_948, w_088_950, w_088_951, w_088_952, w_088_953, w_088_956, w_088_957, w_088_958, w_088_959, w_088_962, w_088_964, w_088_967, w_088_969, w_088_970, w_088_971, w_088_975, w_088_976, w_088_978, w_088_983, w_088_985, w_088_986, w_088_989, w_088_991, w_088_994, w_088_995, w_088_998, w_088_999, w_088_1000, w_088_1001, w_088_1003, w_088_1004, w_088_1005, w_088_1006, w_088_1007, w_088_1011, w_088_1012, w_088_1014, w_088_1017, w_088_1021, w_088_1024, w_088_1027, w_088_1029, w_088_1030, w_088_1031, w_088_1034, w_088_1035, w_088_1040, w_088_1041, w_088_1044, w_088_1046, w_088_1047, w_088_1048, w_088_1049, w_088_1050, w_088_1053, w_088_1055, w_088_1056, w_088_1057, w_088_1058, w_088_1061, w_088_1062, w_088_1063, w_088_1064, w_088_1065, w_088_1066, w_088_1075, w_088_1077, w_088_1079, w_088_1080, w_088_1087, w_088_1091, w_088_1094, w_088_1095, w_088_1097, w_088_1102, w_088_1104, w_088_1108, w_088_1111, w_088_1113, w_088_1114, w_088_1115, w_088_1120, w_088_1121, w_088_1128, w_088_1132, w_088_1133, w_088_1137, w_088_1140, w_088_1141, w_088_1149, w_088_1156, w_088_1160, w_088_1161, w_088_1171, w_088_1173, w_088_1175, w_088_1179, w_088_1182, w_088_1184, w_088_1185, w_088_1187, w_088_1191, w_088_1196, w_088_1197, w_088_1198, w_088_1206, w_088_1207, w_088_1209, w_088_1216, w_088_1218, w_088_1221, w_088_1222, w_088_1226, w_088_1229, w_088_1231, w_088_1232, w_088_1238, w_088_1242, w_088_1243, w_088_1244, w_088_1247, w_088_1250, w_088_1254, w_088_1257, w_088_1259, w_088_1271, w_088_1274, w_088_1277, w_088_1278, w_088_1283, w_088_1284, w_088_1285, w_088_1287, w_088_1289, w_088_1292, w_088_1295, w_088_1301, w_088_1302, w_088_1307, w_088_1310, w_088_1311, w_088_1318, w_088_1319, w_088_1324, w_088_1325, w_088_1326, w_088_1329, w_088_1332, w_088_1335, w_088_1336, w_088_1340, w_088_1343, w_088_1345, w_088_1348, w_088_1350, w_088_1353, w_088_1368, w_088_1370, w_088_1372, w_088_1374, w_088_1375, w_088_1377, w_088_1378, w_088_1383, w_088_1384, w_088_1386, w_088_1397, w_088_1401, w_088_1405, w_088_1409, w_088_1413, w_088_1416, w_088_1417, w_088_1423, w_088_1424, w_088_1427, w_088_1428, w_088_1431, w_088_1433, w_088_1441, w_088_1444, w_088_1447, w_088_1448, w_088_1452, w_088_1457, w_088_1459, w_088_1460, w_088_1464, w_088_1471, w_088_1476, w_088_1479, w_088_1481, w_088_1484, w_088_1488, w_088_1489, w_088_1494, w_088_1495, w_088_1496, w_088_1497, w_088_1498, w_088_1501, w_088_1502, w_088_1509, w_088_1510, w_088_1518, w_088_1522, w_088_1526, w_088_1527, w_088_1529, w_088_1538, w_088_1541, w_088_1545, w_088_1552, w_088_1556, w_088_1562, w_088_1571, w_088_1572, w_088_1577, w_088_1581, w_088_1584, w_088_1587, w_088_1589, w_088_1593, w_088_1595, w_088_1596, w_088_1598, w_088_1599, w_088_1600, w_088_1608, w_088_1612, w_088_1616, w_088_1617, w_088_1618, w_088_1619, w_088_1620, w_088_1634, w_088_1635, w_088_1638, w_088_1640, w_088_1641, w_088_1642, w_088_1645, w_088_1646, w_088_1647, w_088_1648, w_088_1650, w_088_1656, w_088_1657, w_088_1660, w_088_1662, w_088_1663, w_088_1665, w_088_1667, w_088_1669, w_088_1670, w_088_1672, w_088_1675, w_088_1679, w_088_1680, w_088_1681, w_088_1686, w_088_1690, w_088_1692, w_088_1694, w_088_1703, w_088_1704, w_088_1706, w_088_1707, w_088_1714, w_088_1717, w_088_1722, w_088_1724, w_088_1730, w_088_1731, w_088_1734, w_088_1735, w_088_1737, w_088_1738, w_088_1741, w_088_1746, w_088_1750, w_088_1752, w_088_1763, w_088_1765, w_088_1768, w_088_1773, w_088_1775, w_088_1776, w_088_1777, w_088_1784, w_088_1792, w_088_1796, w_088_1803, w_088_1805, w_088_1806, w_088_1809, w_088_1810, w_088_1811, w_088_1813, w_088_1814, w_088_1818, w_088_1823, w_088_1826, w_088_1828, w_088_1830, w_088_1832, w_088_1833, w_088_1834, w_088_1835, w_088_1837, w_088_1838, w_088_1843, w_088_1845, w_088_1846, w_088_1847, w_088_1852, w_088_1855, w_088_1856, w_088_1860, w_088_1868, w_088_1873, w_088_1874, w_088_1876, w_088_1879, w_088_1880, w_088_1883, w_088_1887, w_088_1891, w_088_1894, w_088_1896, w_088_1897, w_088_1899, w_088_1900, w_088_1903, w_088_1904, w_088_1905, w_088_1906, w_088_1909, w_088_1911, w_088_1913, w_088_1921, w_088_1923, w_088_1925, w_088_1926, w_088_1927, w_088_1929, w_088_1931, w_088_1933, w_088_1934, w_088_1938, w_088_1939, w_088_1942, w_088_1944, w_088_1946, w_088_1951, w_088_1952, w_088_1953, w_088_1956, w_088_1958, w_088_1962, w_088_1969, w_088_1971, w_088_1977, w_088_1979, w_088_1994, w_088_1998, w_088_2000, w_088_2001, w_088_2005, w_088_2011, w_088_2017, w_088_2019, w_088_2020, w_088_2022, w_088_2026, w_088_2027, w_088_2032, w_088_2038, w_088_2045, w_088_2046, w_088_2049, w_088_2053, w_088_2054, w_088_2058, w_088_2060, w_088_2063, w_088_2064, w_088_2066, w_088_2072, w_088_2081, w_088_2083, w_088_2088, w_088_2089, w_088_2090, w_088_2100, w_088_2102, w_088_2107, w_088_2109, w_088_2111, w_088_2117, w_088_2118, w_088_2120, w_088_2124, w_088_2128, w_088_2131, w_088_2133, w_088_2136, w_088_2138, w_088_2139, w_088_2143, w_088_2147, w_088_2149, w_088_2154, w_088_2157, w_088_2159, w_088_2161, w_088_2163, w_088_2164, w_088_2167, w_088_2169, w_088_2172, w_088_2179, w_088_2180, w_088_2182, w_088_2194, w_088_2196, w_088_2198, w_088_2202, w_088_2204, w_088_2209, w_088_2214, w_088_2217, w_088_2218, w_088_2219, w_088_2221, w_088_2230, w_088_2234, w_088_2236, w_088_2238, w_088_2240, w_088_2241, w_088_2243, w_088_2244, w_088_2247, w_088_2248, w_088_2256, w_088_2257, w_088_2258, w_088_2259, w_088_2261, w_088_2262, w_088_2264, w_088_2278, w_088_2280, w_088_2284, w_088_2285, w_088_2288, w_088_2290, w_088_2292, w_088_2293, w_088_2298, w_088_2299, w_088_2304, w_088_2306, w_088_2310, w_088_2311, w_088_2314, w_088_2317, w_088_2321, w_088_2322, w_088_2329, w_088_2330, w_088_2332, w_088_2334, w_088_2335, w_088_2337, w_088_2342, w_088_2344, w_088_2349, w_088_2350, w_088_2353, w_088_2354, w_088_2355, w_088_2356, w_088_2358, w_088_2359, w_088_2360, w_088_2361, w_088_2362, w_088_2365, w_088_2369, w_088_2371, w_088_2372, w_088_2376, w_088_2378, w_088_2384, w_088_2396, w_088_2397, w_088_2399, w_088_2401, w_088_2403, w_088_2404, w_088_2407, w_088_2409, w_088_2412, w_088_2416, w_088_2419, w_088_2420, w_088_2421, w_088_2426, w_088_2431, w_088_2432, w_088_2445, w_088_2452, w_088_2453, w_088_2456, w_088_2463, w_088_2464, w_088_2465, w_088_2467, w_088_2469, w_088_2470, w_088_2472, w_088_2477, w_088_2479, w_088_2482, w_088_2483, w_088_2488, w_088_2490, w_088_2493, w_088_2494, w_088_2497, w_088_2498, w_088_2499, w_088_2500, w_088_2501, w_088_2512, w_088_2513, w_088_2515, w_088_2525, w_088_2530, w_088_2539, w_088_2541, w_088_2545, w_088_2547, w_088_2553, w_088_2557, w_088_2558, w_088_2560, w_088_2565, w_088_2572, w_088_2577, w_088_2579, w_088_2584, w_088_2590, w_088_2591, w_088_2594, w_088_2598, w_088_2607, w_088_2613, w_088_2617, w_088_2620, w_088_2621, w_088_2632, w_088_2635, w_088_2639, w_088_2644, w_088_2645, w_088_2662, w_088_2668, w_088_2669, w_088_2683, w_088_2688, w_088_2690, w_088_2691, w_088_2696, w_088_2703, w_088_2706, w_088_2708, w_088_2721, w_088_2722, w_088_2726, w_088_2733, w_088_2736, w_088_2737, w_088_2738, w_088_2743, w_088_2744, w_088_2749, w_088_2750, w_088_2754, w_088_2756, w_088_2759, w_088_2760, w_088_2762, w_088_2764, w_088_2767, w_088_2770, w_088_2778, w_088_2779, w_088_2780, w_088_2782, w_088_2786, w_088_2789, w_088_2792, w_088_2793, w_088_2795, w_088_2797, w_088_2798, w_088_2806, w_088_2811, w_088_2821, w_088_2822, w_088_2823, w_088_2825, w_088_2826, w_088_2828, w_088_2830, w_088_2835, w_088_2836, w_088_2839, w_088_2843, w_088_2844, w_088_2846, w_088_2847, w_088_2848, w_088_2851, w_088_2852, w_088_2854, w_088_2855, w_088_2862, w_088_2864, w_088_2865, w_088_2869, w_088_2872, w_088_2873, w_088_2879, w_088_2888, w_088_2893, w_088_2902, w_088_2915, w_088_2916, w_088_2919, w_088_2922, w_088_2925, w_088_2927, w_088_2935, w_088_2936, w_088_2943, w_088_2945, w_088_2946, w_088_2947, w_088_2948, w_088_2949, w_088_2953, w_088_2958, w_088_2960, w_088_2962, w_088_2973, w_088_2981, w_088_2991, w_088_2997, w_088_3001, w_088_3002, w_088_3004, w_088_3006, w_088_3007, w_088_3008, w_088_3010, w_088_3011, w_088_3013, w_088_3018, w_088_3021, w_088_3022, w_088_3026, w_088_3027, w_088_3030, w_088_3034, w_088_3036, w_088_3041, w_088_3042, w_088_3046, w_088_3048, w_088_3049, w_088_3054, w_088_3057, w_088_3061, w_088_3063, w_088_3065, w_088_3068, w_088_3070, w_088_3071, w_088_3072, w_088_3073, w_088_3075, w_088_3077, w_088_3080, w_088_3081, w_088_3085, w_088_3088, w_088_3089, w_088_3091, w_088_3095, w_088_3097, w_088_3099, w_088_3100, w_088_3106, w_088_3107, w_088_3109, w_088_3110, w_088_3113, w_088_3117, w_088_3120, w_088_3122, w_088_3124, w_088_3125, w_088_3126, w_088_3132, w_088_3137, w_088_3141, w_088_3148, w_088_3151, w_088_3159, w_088_3161, w_088_3162, w_088_3164, w_088_3165, w_088_3166, w_088_3167, w_088_3168, w_088_3170, w_088_3171, w_088_3174, w_088_3184, w_088_3186, w_088_3187, w_088_3188, w_088_3190, w_088_3193, w_088_3197, w_088_3203, w_088_3211, w_088_3214, w_088_3216, w_088_3220, w_088_3224, w_088_3230, w_088_3233, w_088_3234, w_088_3235, w_088_3237, w_088_3239, w_088_3243, w_088_3246, w_088_3253, w_088_3255, w_088_3260, w_088_3262, w_088_3275, w_088_3276, w_088_3277, w_088_3278, w_088_3283, w_088_3284, w_088_3285, w_088_3287, w_088_3294, w_088_3298, w_088_3299, w_088_3307, w_088_3313, w_088_3314, w_088_3318, w_088_3319, w_088_3328, w_088_3329, w_088_3331, w_088_3334, w_088_3338, w_088_3340, w_088_3342, w_088_3349, w_088_3350, w_088_3351, w_088_3357, w_088_3359, w_088_3360, w_088_3364, w_088_3367, w_088_3375, w_088_3377, w_088_3387, w_088_3391, w_088_3392, w_088_3395, w_088_3396, w_088_3398, w_088_3400, w_088_3401, w_088_3402, w_088_3405, w_088_3406, w_088_3410, w_088_3411, w_088_3438, w_088_3442, w_088_3444, w_088_3445, w_088_3446, w_088_3448, w_088_3451, w_088_3455, w_088_3457, w_088_3464, w_088_3465, w_088_3466, w_088_3471, w_088_3474, w_088_3475, w_088_3481, w_088_3486, w_088_3491, w_088_3499, w_088_3500, w_088_3504, w_088_3507, w_088_3510, w_088_3511, w_088_3513, w_088_3517, w_088_3518, w_088_3523, w_088_3525, w_088_3527, w_088_3529, w_088_3530, w_088_3531, w_088_3538, w_088_3541, w_088_3548, w_088_3553, w_088_3555, w_088_3556, w_088_3557, w_088_3559, w_088_3561, w_088_3565, w_088_3571, w_088_3572, w_088_3574, w_088_3580, w_088_3581, w_088_3583, w_088_3584, w_088_3585, w_088_3587, w_088_3590, w_088_3593, w_088_3595, w_088_3596, w_088_3600, w_088_3608, w_088_3609, w_088_3610, w_088_3617, w_088_3619, w_088_3624, w_088_3625, w_088_3627, w_088_3631, w_088_3632, w_088_3635, w_088_3639, w_088_3640, w_088_3642, w_088_3643, w_088_3646, w_088_3647, w_088_3648, w_088_3649, w_088_3653, w_088_3654, w_088_3668, w_088_3671, w_088_3674, w_088_3681, w_088_3683, w_088_3690, w_088_3695, w_088_3696, w_088_3702, w_088_3709, w_088_3710, w_088_3712, w_088_3716, w_088_3718, w_088_3719, w_088_3721, w_088_3722, w_088_3725, w_088_3726, w_088_3733, w_088_3735, w_088_3736, w_088_3750, w_088_3754, w_088_3758, w_088_3760, w_088_3772, w_088_3777, w_088_3781, w_088_3782, w_088_3786, w_088_3787, w_088_3794, w_088_3802, w_088_3803, w_088_3815, w_088_3816, w_088_3818, w_088_3819, w_088_3822, w_088_3826, w_088_3827, w_088_3841, w_088_3842, w_088_3843, w_088_3846, w_088_3849, w_088_3853, w_088_3855, w_088_3857, w_088_3858, w_088_3859, w_088_3864, w_088_3865, w_088_3873, w_088_3874, w_088_3876, w_088_3884, w_088_3885, w_088_3888, w_088_3890, w_088_3891, w_088_3894, w_088_3895, w_088_3896, w_088_3900, w_088_3904, w_088_3905, w_088_3906, w_088_3917, w_088_3919, w_088_3921, w_088_3924, w_088_3927, w_088_3928, w_088_3929;
  wire w_089_000, w_089_001, w_089_003, w_089_004, w_089_005, w_089_006, w_089_007, w_089_008, w_089_009, w_089_011, w_089_012, w_089_013, w_089_014, w_089_015, w_089_017, w_089_018, w_089_019, w_089_020, w_089_022, w_089_023, w_089_024, w_089_026, w_089_027, w_089_028, w_089_029, w_089_030, w_089_032, w_089_033, w_089_034, w_089_035, w_089_036, w_089_037, w_089_038, w_089_039, w_089_040, w_089_042, w_089_043, w_089_044, w_089_045, w_089_046, w_089_047, w_089_048, w_089_049, w_089_050, w_089_051, w_089_054, w_089_055, w_089_056, w_089_057, w_089_059, w_089_060, w_089_061, w_089_062, w_089_063, w_089_064, w_089_066, w_089_067, w_089_069, w_089_070, w_089_071, w_089_072, w_089_073, w_089_074, w_089_075, w_089_078, w_089_079, w_089_080, w_089_081, w_089_082, w_089_084, w_089_085, w_089_086, w_089_087, w_089_088, w_089_089, w_089_090, w_089_091, w_089_092, w_089_093, w_089_094, w_089_095, w_089_096, w_089_097, w_089_098, w_089_099, w_089_100, w_089_101, w_089_102, w_089_103, w_089_104, w_089_105, w_089_106, w_089_107, w_089_108, w_089_109, w_089_110, w_089_111, w_089_112, w_089_115, w_089_116, w_089_117, w_089_118, w_089_119, w_089_120, w_089_121, w_089_122, w_089_123, w_089_124, w_089_125, w_089_126, w_089_127, w_089_130, w_089_131, w_089_132, w_089_133, w_089_134, w_089_137, w_089_138, w_089_139, w_089_140, w_089_141, w_089_142, w_089_143, w_089_146, w_089_147, w_089_149, w_089_150, w_089_151, w_089_152, w_089_153, w_089_154, w_089_155, w_089_156, w_089_157, w_089_158, w_089_159, w_089_160, w_089_162, w_089_163, w_089_164, w_089_165, w_089_167, w_089_168, w_089_169, w_089_170, w_089_171, w_089_172, w_089_173, w_089_175, w_089_176, w_089_177, w_089_178, w_089_179, w_089_180, w_089_181, w_089_182, w_089_185, w_089_186, w_089_187, w_089_188, w_089_189, w_089_190, w_089_191, w_089_192, w_089_193, w_089_194, w_089_195, w_089_196, w_089_197, w_089_198, w_089_199, w_089_201, w_089_202, w_089_204, w_089_205, w_089_206, w_089_207, w_089_208, w_089_209, w_089_210, w_089_212, w_089_214, w_089_215, w_089_216, w_089_217, w_089_218, w_089_219, w_089_220, w_089_221, w_089_222, w_089_223, w_089_224, w_089_225, w_089_226, w_089_228, w_089_230, w_089_231, w_089_232, w_089_234, w_089_235, w_089_236, w_089_238, w_089_239, w_089_240, w_089_241, w_089_243, w_089_246, w_089_247, w_089_248, w_089_249, w_089_251, w_089_254, w_089_255, w_089_256, w_089_257, w_089_258, w_089_260, w_089_262, w_089_263, w_089_264, w_089_265, w_089_266, w_089_267, w_089_268, w_089_269, w_089_270, w_089_271, w_089_272, w_089_273, w_089_274, w_089_276, w_089_278, w_089_280, w_089_281, w_089_282, w_089_283, w_089_285, w_089_286, w_089_287, w_089_288, w_089_289, w_089_290, w_089_291, w_089_292, w_089_294, w_089_295, w_089_298, w_089_299, w_089_300, w_089_301, w_089_302, w_089_304, w_089_305, w_089_306, w_089_307, w_089_309, w_089_310, w_089_311, w_089_312, w_089_314, w_089_316, w_089_317, w_089_318, w_089_319, w_089_320, w_089_321, w_089_322, w_089_323, w_089_324, w_089_326, w_089_327, w_089_328, w_089_330, w_089_331, w_089_334, w_089_335, w_089_336, w_089_337, w_089_338, w_089_340, w_089_342, w_089_343, w_089_345, w_089_346, w_089_347, w_089_348, w_089_350, w_089_352, w_089_354, w_089_355, w_089_357, w_089_358, w_089_360, w_089_362, w_089_365, w_089_366, w_089_367, w_089_368, w_089_369, w_089_371, w_089_372, w_089_373, w_089_374, w_089_375, w_089_376, w_089_377, w_089_379, w_089_380, w_089_381, w_089_382, w_089_384, w_089_385, w_089_387, w_089_389, w_089_390, w_089_391, w_089_392, w_089_393, w_089_398, w_089_399, w_089_400, w_089_401, w_089_403, w_089_404, w_089_409, w_089_410, w_089_411, w_089_412, w_089_413, w_089_415, w_089_416, w_089_417, w_089_418, w_089_419, w_089_421, w_089_422, w_089_423, w_089_424, w_089_425, w_089_426, w_089_427, w_089_428, w_089_429, w_089_430, w_089_432, w_089_435, w_089_436, w_089_437, w_089_438, w_089_439, w_089_440, w_089_441, w_089_442, w_089_443, w_089_444, w_089_445, w_089_446, w_089_447, w_089_448, w_089_449, w_089_450, w_089_453, w_089_454, w_089_455, w_089_457, w_089_458, w_089_461, w_089_462, w_089_464, w_089_466, w_089_467, w_089_469, w_089_470, w_089_471, w_089_472, w_089_473, w_089_474, w_089_476, w_089_478, w_089_479, w_089_480, w_089_481, w_089_482, w_089_484, w_089_486, w_089_488, w_089_489, w_089_490, w_089_491, w_089_492, w_089_493, w_089_496, w_089_497, w_089_500, w_089_502, w_089_503, w_089_504, w_089_505, w_089_506, w_089_507, w_089_508, w_089_509, w_089_511, w_089_512, w_089_514, w_089_515, w_089_516, w_089_518, w_089_519, w_089_521, w_089_522, w_089_523, w_089_524, w_089_526, w_089_527, w_089_528, w_089_529, w_089_530, w_089_531, w_089_533, w_089_535, w_089_536, w_089_537, w_089_538, w_089_539, w_089_541, w_089_542, w_089_543, w_089_544, w_089_548, w_089_551, w_089_552, w_089_553, w_089_554, w_089_556, w_089_557, w_089_560, w_089_562, w_089_563, w_089_564, w_089_565, w_089_567, w_089_569, w_089_570, w_089_572, w_089_573, w_089_575, w_089_576, w_089_577, w_089_578, w_089_579, w_089_580, w_089_581, w_089_582, w_089_583, w_089_584, w_089_586, w_089_587, w_089_588, w_089_589, w_089_590, w_089_591, w_089_592, w_089_594, w_089_595, w_089_596, w_089_599, w_089_600, w_089_602, w_089_603, w_089_604, w_089_605, w_089_606, w_089_607, w_089_608, w_089_610, w_089_611, w_089_613, w_089_616, w_089_617, w_089_618, w_089_619, w_089_620, w_089_621, w_089_622, w_089_624, w_089_625, w_089_626, w_089_630, w_089_632, w_089_633, w_089_635, w_089_636, w_089_637, w_089_639, w_089_640, w_089_641, w_089_642, w_089_643, w_089_645, w_089_646, w_089_647, w_089_648, w_089_649, w_089_653, w_089_656, w_089_657, w_089_658, w_089_659, w_089_660, w_089_661, w_089_662, w_089_664, w_089_665, w_089_666, w_089_667, w_089_668, w_089_669, w_089_670, w_089_672, w_089_673, w_089_675, w_089_676, w_089_678, w_089_679, w_089_680, w_089_681, w_089_682, w_089_683, w_089_684, w_089_685, w_089_687, w_089_688, w_089_690, w_089_692, w_089_693, w_089_694, w_089_695, w_089_696, w_089_697, w_089_698, w_089_699, w_089_700, w_089_701, w_089_702, w_089_703, w_089_704, w_089_705, w_089_706, w_089_707, w_089_708, w_089_709, w_089_710, w_089_712, w_089_713, w_089_714, w_089_716, w_089_717, w_089_718, w_089_719, w_089_720, w_089_722, w_089_723, w_089_724, w_089_725, w_089_727, w_089_729, w_089_730, w_089_731, w_089_732, w_089_734, w_089_737, w_089_738, w_089_739, w_089_740, w_089_741, w_089_743, w_089_744, w_089_745, w_089_746, w_089_747, w_089_748, w_089_749, w_089_750, w_089_751, w_089_752, w_089_755, w_089_756, w_089_757, w_089_758, w_089_759, w_089_761, w_089_762, w_089_764, w_089_765, w_089_766, w_089_767, w_089_768, w_089_770, w_089_771, w_089_772, w_089_774, w_089_775, w_089_776, w_089_780, w_089_781, w_089_783, w_089_785, w_089_787, w_089_788, w_089_789, w_089_790, w_089_791, w_089_792, w_089_793, w_089_795, w_089_796, w_089_799, w_089_800, w_089_802, w_089_804, w_089_805, w_089_806, w_089_807, w_089_808, w_089_809, w_089_810, w_089_812, w_089_813, w_089_814, w_089_815, w_089_816, w_089_817, w_089_818, w_089_819, w_089_820, w_089_821, w_089_825, w_089_826, w_089_828, w_089_830, w_089_831, w_089_832, w_089_833, w_089_834, w_089_835, w_089_836, w_089_837, w_089_838, w_089_840, w_089_841, w_089_843, w_089_844, w_089_846, w_089_847, w_089_848, w_089_849, w_089_850, w_089_851, w_089_852, w_089_853, w_089_854, w_089_856, w_089_857, w_089_858, w_089_859, w_089_860, w_089_861, w_089_862, w_089_863, w_089_865, w_089_866, w_089_867, w_089_868, w_089_869, w_089_870, w_089_871, w_089_872, w_089_873, w_089_874, w_089_876, w_089_877, w_089_878, w_089_884, w_089_885, w_089_887, w_089_888, w_089_889, w_089_890, w_089_891, w_089_892, w_089_893, w_089_894, w_089_895, w_089_896, w_089_897, w_089_898, w_089_899, w_089_901, w_089_902, w_089_903, w_089_905, w_089_906, w_089_908, w_089_909, w_089_912, w_089_913, w_089_914, w_089_916, w_089_918, w_089_919, w_089_920, w_089_921, w_089_922, w_089_924, w_089_925, w_089_926, w_089_927, w_089_928, w_089_929, w_089_930, w_089_932, w_089_933, w_089_934, w_089_935, w_089_936, w_089_938, w_089_939, w_089_940, w_089_942, w_089_943, w_089_944, w_089_945, w_089_946, w_089_947, w_089_950, w_089_951, w_089_953, w_089_954, w_089_955, w_089_957, w_089_958, w_089_959, w_089_961, w_089_963, w_089_965, w_089_967, w_089_968, w_089_969, w_089_970, w_089_971, w_089_972, w_089_973, w_089_974, w_089_975, w_089_976, w_089_977, w_089_979, w_089_980, w_089_981, w_089_982, w_089_983, w_089_985, w_089_986, w_089_987, w_089_990, w_089_991, w_089_992, w_089_994, w_089_995, w_089_996, w_089_998, w_089_999, w_089_1000, w_089_1001, w_089_1002, w_089_1003, w_089_1004, w_089_1005, w_089_1006, w_089_1007, w_089_1008, w_089_1009, w_089_1010, w_089_1011, w_089_1012, w_089_1014, w_089_1015, w_089_1016, w_089_1019, w_089_1020, w_089_1022, w_089_1023, w_089_1024, w_089_1025, w_089_1030, w_089_1031, w_089_1032, w_089_1033, w_089_1034, w_089_1035, w_089_1037, w_089_1039, w_089_1040, w_089_1041, w_089_1042, w_089_1044, w_089_1046, w_089_1047, w_089_1048, w_089_1049, w_089_1050, w_089_1051, w_089_1052, w_089_1053, w_089_1054, w_089_1055, w_089_1056, w_089_1057, w_089_1058, w_089_1059, w_089_1061, w_089_1063, w_089_1065, w_089_1066, w_089_1067, w_089_1068, w_089_1069, w_089_1070, w_089_1071, w_089_1073, w_089_1077, w_089_1079, w_089_1080, w_089_1081, w_089_1082, w_089_1083, w_089_1084, w_089_1085, w_089_1086, w_089_1087, w_089_1088, w_089_1089, w_089_1091, w_089_1093, w_089_1095, w_089_1098, w_089_1100, w_089_1101, w_089_1102, w_089_1103, w_089_1105, w_089_1106, w_089_1107, w_089_1108, w_089_1109, w_089_1110, w_089_1111, w_089_1112, w_089_1114, w_089_1115, w_089_1116, w_089_1117, w_089_1118, w_089_1119, w_089_1120, w_089_1121, w_089_1122, w_089_1123, w_089_1125, w_089_1127, w_089_1128, w_089_1129, w_089_1130, w_089_1133, w_089_1134, w_089_1135, w_089_1137, w_089_1138, w_089_1139, w_089_1140, w_089_1141, w_089_1142, w_089_1145, w_089_1146, w_089_1147, w_089_1148, w_089_1149, w_089_1153, w_089_1154, w_089_1156, w_089_1157, w_089_1158, w_089_1159, w_089_1160, w_089_1161, w_089_1162, w_089_1166, w_089_1167, w_089_1168, w_089_1169, w_089_1171, w_089_1172, w_089_1173, w_089_1174, w_089_1175, w_089_1176, w_089_1178, w_089_1179, w_089_1180, w_089_1181, w_089_1182, w_089_1183, w_089_1184, w_089_1185, w_089_1186, w_089_1187;
  wire w_090_001, w_090_002, w_090_004, w_090_006, w_090_009, w_090_010, w_090_015, w_090_016, w_090_018, w_090_019, w_090_020, w_090_021, w_090_022, w_090_024, w_090_025, w_090_026, w_090_028, w_090_029, w_090_031, w_090_033, w_090_034, w_090_036, w_090_037, w_090_038, w_090_039, w_090_040, w_090_042, w_090_043, w_090_044, w_090_045, w_090_046, w_090_047, w_090_048, w_090_051, w_090_052, w_090_053, w_090_054, w_090_055, w_090_056, w_090_061, w_090_063, w_090_064, w_090_065, w_090_066, w_090_068, w_090_072, w_090_073, w_090_074, w_090_076, w_090_077, w_090_080, w_090_082, w_090_084, w_090_085, w_090_086, w_090_087, w_090_088, w_090_089, w_090_090, w_090_091, w_090_092, w_090_093, w_090_094, w_090_095, w_090_098, w_090_100, w_090_102, w_090_103, w_090_104, w_090_105, w_090_106, w_090_107, w_090_108, w_090_109, w_090_110, w_090_111, w_090_112, w_090_113, w_090_114, w_090_115, w_090_117, w_090_118, w_090_121, w_090_123, w_090_125, w_090_126, w_090_128, w_090_132, w_090_134, w_090_136, w_090_137, w_090_138, w_090_139, w_090_142, w_090_143, w_090_144, w_090_147, w_090_148, w_090_149, w_090_151, w_090_153, w_090_154, w_090_155, w_090_156, w_090_157, w_090_159, w_090_161, w_090_162, w_090_163, w_090_164, w_090_166, w_090_169, w_090_170, w_090_171, w_090_172, w_090_173, w_090_176, w_090_177, w_090_179, w_090_180, w_090_184, w_090_186, w_090_188, w_090_189, w_090_191, w_090_195, w_090_197, w_090_198, w_090_200, w_090_201, w_090_202, w_090_203, w_090_207, w_090_208, w_090_209, w_090_210, w_090_211, w_090_212, w_090_213, w_090_214, w_090_215, w_090_216, w_090_219, w_090_220, w_090_221, w_090_222, w_090_223, w_090_225, w_090_226, w_090_227, w_090_229, w_090_231, w_090_232, w_090_234, w_090_235, w_090_236, w_090_238, w_090_239, w_090_240, w_090_241, w_090_242, w_090_244, w_090_245, w_090_246, w_090_247, w_090_248, w_090_250, w_090_254, w_090_255, w_090_256, w_090_258, w_090_260, w_090_262, w_090_263, w_090_265, w_090_266, w_090_269, w_090_270, w_090_272, w_090_277, w_090_278, w_090_279, w_090_282, w_090_285, w_090_286, w_090_287, w_090_288, w_090_290, w_090_293, w_090_294, w_090_296, w_090_297, w_090_298, w_090_299, w_090_300, w_090_302, w_090_303, w_090_306, w_090_310, w_090_311, w_090_312, w_090_313, w_090_316, w_090_317, w_090_318, w_090_319, w_090_320, w_090_321, w_090_323, w_090_326, w_090_329, w_090_330, w_090_331, w_090_333, w_090_334, w_090_335, w_090_337, w_090_338, w_090_339, w_090_342, w_090_343, w_090_344, w_090_345, w_090_346, w_090_351, w_090_352, w_090_354, w_090_356, w_090_357, w_090_358, w_090_359, w_090_360, w_090_361, w_090_362, w_090_364, w_090_366, w_090_367, w_090_373, w_090_374, w_090_375, w_090_378, w_090_379, w_090_380, w_090_381, w_090_383, w_090_384, w_090_385, w_090_388, w_090_389, w_090_390, w_090_391, w_090_392, w_090_395, w_090_396, w_090_398, w_090_400, w_090_401, w_090_402, w_090_403, w_090_405, w_090_407, w_090_409, w_090_410, w_090_414, w_090_415, w_090_416, w_090_418, w_090_419, w_090_420, w_090_421, w_090_422, w_090_423, w_090_425, w_090_427, w_090_429, w_090_431, w_090_433, w_090_434, w_090_435, w_090_437, w_090_438, w_090_439, w_090_441, w_090_443, w_090_446, w_090_447, w_090_448, w_090_449, w_090_450, w_090_451, w_090_452, w_090_454, w_090_457, w_090_460, w_090_461, w_090_462, w_090_464, w_090_465, w_090_466, w_090_467, w_090_468, w_090_470, w_090_471, w_090_472, w_090_473, w_090_474, w_090_476, w_090_478, w_090_480, w_090_481, w_090_482, w_090_483, w_090_485, w_090_486, w_090_487, w_090_489, w_090_492, w_090_493, w_090_494, w_090_495, w_090_496, w_090_497, w_090_498, w_090_499, w_090_500, w_090_501, w_090_502, w_090_503, w_090_509, w_090_511, w_090_512, w_090_513, w_090_515, w_090_517, w_090_518, w_090_519, w_090_520, w_090_521, w_090_525, w_090_526, w_090_527, w_090_528, w_090_529, w_090_530, w_090_532, w_090_533, w_090_535, w_090_536, w_090_538, w_090_539, w_090_540, w_090_541, w_090_543, w_090_544, w_090_545, w_090_546, w_090_547, w_090_548, w_090_549, w_090_550, w_090_551, w_090_553, w_090_554, w_090_555, w_090_556, w_090_557, w_090_560, w_090_561, w_090_562, w_090_563, w_090_565, w_090_568, w_090_569, w_090_570, w_090_571, w_090_574, w_090_575, w_090_576, w_090_577, w_090_578, w_090_579, w_090_580, w_090_581, w_090_582, w_090_583, w_090_584, w_090_585, w_090_586, w_090_587, w_090_588, w_090_594, w_090_596, w_090_597, w_090_598, w_090_599, w_090_600, w_090_602, w_090_603, w_090_606, w_090_607, w_090_608, w_090_610, w_090_612, w_090_613, w_090_616, w_090_617, w_090_618, w_090_619, w_090_620, w_090_621, w_090_623, w_090_624, w_090_626, w_090_629, w_090_630, w_090_635, w_090_636, w_090_637, w_090_641, w_090_643, w_090_644, w_090_645, w_090_646, w_090_647, w_090_648, w_090_650, w_090_651, w_090_654, w_090_655, w_090_656, w_090_657, w_090_659, w_090_660, w_090_662, w_090_663, w_090_665, w_090_667, w_090_670, w_090_671, w_090_672, w_090_674, w_090_676, w_090_677, w_090_678, w_090_680, w_090_681, w_090_682, w_090_683, w_090_684, w_090_686, w_090_687, w_090_688, w_090_689, w_090_691, w_090_692, w_090_693, w_090_694, w_090_697, w_090_701, w_090_703, w_090_704, w_090_705, w_090_706, w_090_707, w_090_708, w_090_709, w_090_712, w_090_714, w_090_715, w_090_718, w_090_719, w_090_723, w_090_728, w_090_729, w_090_732, w_090_740, w_090_742, w_090_743, w_090_744, w_090_745, w_090_747, w_090_752, w_090_758, w_090_759, w_090_760, w_090_762, w_090_763, w_090_764, w_090_772, w_090_773, w_090_774, w_090_777, w_090_778, w_090_782, w_090_786, w_090_787, w_090_789, w_090_791, w_090_796, w_090_797, w_090_799, w_090_801, w_090_804, w_090_805, w_090_806, w_090_807, w_090_809, w_090_810, w_090_811, w_090_813, w_090_814, w_090_815, w_090_817, w_090_818, w_090_819, w_090_820, w_090_821, w_090_822, w_090_823, w_090_829, w_090_831, w_090_834, w_090_835, w_090_837, w_090_838, w_090_839, w_090_840, w_090_843, w_090_845, w_090_846, w_090_847, w_090_848, w_090_849, w_090_851, w_090_852, w_090_857, w_090_859, w_090_862, w_090_864, w_090_865, w_090_867, w_090_871, w_090_872, w_090_875, w_090_878, w_090_879, w_090_880, w_090_881, w_090_882, w_090_883, w_090_884, w_090_885, w_090_886, w_090_887, w_090_889, w_090_890, w_090_891, w_090_892, w_090_893, w_090_895, w_090_897, w_090_898, w_090_900, w_090_903, w_090_904, w_090_907, w_090_909, w_090_911, w_090_914, w_090_916, w_090_919, w_090_921, w_090_924, w_090_930, w_090_931, w_090_932, w_090_935, w_090_936, w_090_937, w_090_938, w_090_940, w_090_942, w_090_944, w_090_945, w_090_946, w_090_947, w_090_948, w_090_950, w_090_953, w_090_956, w_090_957, w_090_959, w_090_960, w_090_961, w_090_962, w_090_964, w_090_966, w_090_968, w_090_969, w_090_970, w_090_972, w_090_973, w_090_974, w_090_977, w_090_978, w_090_980, w_090_981, w_090_982, w_090_983, w_090_985, w_090_986, w_090_989, w_090_991, w_090_993, w_090_995, w_090_999, w_090_1000, w_090_1001, w_090_1005, w_090_1009, w_090_1010, w_090_1012, w_090_1014, w_090_1016, w_090_1018, w_090_1019, w_090_1020, w_090_1021, w_090_1022, w_090_1025, w_090_1029, w_090_1030, w_090_1032, w_090_1036, w_090_1037, w_090_1038, w_090_1040, w_090_1041, w_090_1042, w_090_1043, w_090_1046, w_090_1047, w_090_1048, w_090_1057, w_090_1058, w_090_1060, w_090_1062, w_090_1066, w_090_1067, w_090_1069, w_090_1070, w_090_1072, w_090_1073, w_090_1075, w_090_1077, w_090_1080, w_090_1081, w_090_1084, w_090_1086, w_090_1088, w_090_1090, w_090_1091, w_090_1093, w_090_1095, w_090_1097, w_090_1098, w_090_1101, w_090_1103, w_090_1107, w_090_1108, w_090_1109, w_090_1112, w_090_1113, w_090_1116, w_090_1117, w_090_1118, w_090_1119, w_090_1120, w_090_1121, w_090_1122, w_090_1126, w_090_1127, w_090_1128, w_090_1129, w_090_1130, w_090_1132, w_090_1138, w_090_1141, w_090_1144, w_090_1145, w_090_1146, w_090_1147, w_090_1148, w_090_1150, w_090_1151, w_090_1152, w_090_1153, w_090_1154, w_090_1155, w_090_1156, w_090_1158, w_090_1159, w_090_1160, w_090_1161, w_090_1162, w_090_1163, w_090_1164, w_090_1165, w_090_1166, w_090_1167, w_090_1168, w_090_1171, w_090_1176, w_090_1178, w_090_1180, w_090_1181, w_090_1182, w_090_1184, w_090_1192, w_090_1195, w_090_1197, w_090_1198, w_090_1199, w_090_1200, w_090_1202, w_090_1206, w_090_1210, w_090_1211, w_090_1213, w_090_1214, w_090_1215, w_090_1217, w_090_1223, w_090_1224, w_090_1226, w_090_1230, w_090_1231, w_090_1232, w_090_1233, w_090_1240, w_090_1244, w_090_1245, w_090_1246, w_090_1247, w_090_1249, w_090_1250, w_090_1252, w_090_1253, w_090_1255, w_090_1256, w_090_1259, w_090_1261, w_090_1263, w_090_1264, w_090_1266, w_090_1267, w_090_1268, w_090_1269, w_090_1271, w_090_1272, w_090_1274, w_090_1276, w_090_1277, w_090_1278, w_090_1280, w_090_1281, w_090_1285, w_090_1286, w_090_1288, w_090_1291, w_090_1292, w_090_1295, w_090_1297, w_090_1299, w_090_1301, w_090_1303, w_090_1305, w_090_1307, w_090_1308, w_090_1310, w_090_1311, w_090_1314, w_090_1315, w_090_1316, w_090_1317, w_090_1319, w_090_1320, w_090_1323, w_090_1325, w_090_1327, w_090_1329, w_090_1330, w_090_1331, w_090_1334, w_090_1339, w_090_1341, w_090_1342, w_090_1344, w_090_1345, w_090_1347, w_090_1348, w_090_1358, w_090_1360, w_090_1361, w_090_1363, w_090_1366, w_090_1368, w_090_1372, w_090_1376, w_090_1378, w_090_1383, w_090_1384, w_090_1387, w_090_1389, w_090_1392, w_090_1397, w_090_1398, w_090_1401, w_090_1402, w_090_1403, w_090_1405, w_090_1406, w_090_1408, w_090_1410, w_090_1411, w_090_1412, w_090_1413, w_090_1415, w_090_1418, w_090_1422, w_090_1424, w_090_1425, w_090_1432, w_090_1433, w_090_1434, w_090_1435, w_090_1437, w_090_1438, w_090_1441, w_090_1442, w_090_1444, w_090_1447, w_090_1450, w_090_1453, w_090_1456, w_090_1457, w_090_1459, w_090_1460, w_090_1461, w_090_1463, w_090_1468, w_090_1471, w_090_1477, w_090_1478, w_090_1480, w_090_1481, w_090_1491, w_090_1492, w_090_1494, w_090_1496, w_090_1499, w_090_1505, w_090_1506, w_090_1507, w_090_1510, w_090_1511, w_090_1512, w_090_1513, w_090_1516, w_090_1517, w_090_1518, w_090_1519, w_090_1523, w_090_1524, w_090_1526, w_090_1527, w_090_1528, w_090_1529, w_090_1532, w_090_1533, w_090_1536, w_090_1537, w_090_1538, w_090_1539, w_090_1541, w_090_1543, w_090_1544, w_090_1545, w_090_1546, w_090_1548, w_090_1553, w_090_1555, w_090_1558, w_090_1560, w_090_1562, w_090_1563, w_090_1564, w_090_1566, w_090_1567, w_090_1568, w_090_1575, w_090_1576, w_090_1577, w_090_1578, w_090_1582, w_090_1583, w_090_1586, w_090_1589, w_090_1590, w_090_1591, w_090_1592, w_090_1594, w_090_1597, w_090_1606, w_090_1607, w_090_1609, w_090_1613, w_090_1615, w_090_1617, w_090_1619, w_090_1620, w_090_1622, w_090_1623, w_090_1627, w_090_1631, w_090_1634, w_090_1636, w_090_1641, w_090_1642, w_090_1643, w_090_1645, w_090_1646, w_090_1647, w_090_1648, w_090_1651, w_090_1653, w_090_1656, w_090_1657, w_090_1658, w_090_1659, w_090_1661, w_090_1662, w_090_1664, w_090_1665, w_090_1666, w_090_1672, w_090_1673, w_090_1674, w_090_1676, w_090_1678, w_090_1680, w_090_1681, w_090_1682, w_090_1691, w_090_1692, w_090_1694, w_090_1696, w_090_1697, w_090_1700, w_090_1702, w_090_1703, w_090_1709, w_090_1711, w_090_1712, w_090_1716, w_090_1717, w_090_1718, w_090_1719, w_090_1721, w_090_1722, w_090_1723, w_090_1726, w_090_1728, w_090_1729, w_090_1730, w_090_1732, w_090_1734, w_090_1736, w_090_1739, w_090_1740, w_090_1741, w_090_1742, w_090_1743, w_090_1745, w_090_1747, w_090_1748, w_090_1756, w_090_1759, w_090_1763, w_090_1764, w_090_1765, w_090_1766, w_090_1767, w_090_1768, w_090_1773, w_090_1774, w_090_1775, w_090_1776, w_090_1778, w_090_1780, w_090_1781, w_090_1782, w_090_1783, w_090_1785, w_090_1786, w_090_1788, w_090_1791, w_090_1792, w_090_1793, w_090_1795, w_090_1799, w_090_1800, w_090_1802, w_090_1804, w_090_1807, w_090_1808, w_090_1811, w_090_1812, w_090_1813, w_090_1816, w_090_1819, w_090_1822, w_090_1824, w_090_1825, w_090_1826, w_090_1827, w_090_1828, w_090_1830, w_090_1833, w_090_1834, w_090_1836, w_090_1837, w_090_1839, w_090_1840, w_090_1841, w_090_1842, w_090_1843, w_090_1852, w_090_1855, w_090_1856, w_090_1860, w_090_1862, w_090_1863, w_090_1864, w_090_1866, w_090_1869, w_090_1870, w_090_1872, w_090_1873, w_090_1877, w_090_1878, w_090_1879, w_090_1880, w_090_1881, w_090_1886, w_090_1889, w_090_1891, w_090_1892, w_090_1895, w_090_1897, w_090_1899, w_090_1900, w_090_1902, w_090_1906, w_090_1908, w_090_1909, w_090_1911, w_090_1916, w_090_1920, w_090_1921, w_090_1922, w_090_1923, w_090_1926, w_090_1929, w_090_1930, w_090_1931, w_090_1938, w_090_1940, w_090_1943, w_090_1944, w_090_1945, w_090_1946, w_090_1950, w_090_1951, w_090_1952, w_090_1953, w_090_1960, w_090_1961, w_090_1964, w_090_1969, w_090_1970, w_090_1972, w_090_1973, w_090_1976, w_090_1979, w_090_1980, w_090_1982, w_090_1983, w_090_1985, w_090_1987, w_090_1988, w_090_1990, w_090_1992, w_090_1993, w_090_1994, w_090_1995, w_090_1996, w_090_1997, w_090_1999, w_090_2000, w_090_2005, w_090_2007, w_090_2011, w_090_2012, w_090_2013, w_090_2015, w_090_2016, w_090_2018, w_090_2019, w_090_2021, w_090_2022, w_090_2023, w_090_2025, w_090_2029, w_090_2030, w_090_2031, w_090_2032, w_090_2033, w_090_2034, w_090_2041, w_090_2042, w_090_2043, w_090_2044, w_090_2045, w_090_2046, w_090_2048, w_090_2051, w_090_2052, w_090_2054, w_090_2055, w_090_2059, w_090_2061, w_090_2064, w_090_2067, w_090_2068, w_090_2069, w_090_2070, w_090_2072, w_090_2077, w_090_2078, w_090_2083, w_090_2084, w_090_2086, w_090_2092, w_090_2093, w_090_2094, w_090_2095, w_090_2097, w_090_2099, w_090_2100, w_090_2103, w_090_2104, w_090_2105, w_090_2107, w_090_2108, w_090_2112, w_090_2113, w_090_2114, w_090_2115, w_090_2116, w_090_2119, w_090_2122, w_090_2125, w_090_2126, w_090_2128, w_090_2131, w_090_2132, w_090_2133, w_090_2134, w_090_2136, w_090_2138, w_090_2139, w_090_2141, w_090_2143, w_090_2146, w_090_2147, w_090_2149, w_090_2150, w_090_2151, w_090_2152, w_090_2153, w_090_2154, w_090_2155, w_090_2161, w_090_2162, w_090_2166, w_090_2167, w_090_2169, w_090_2170, w_090_2171, w_090_2172;
  wire w_091_001, w_091_003, w_091_004, w_091_010, w_091_011, w_091_013, w_091_014, w_091_015, w_091_016, w_091_017, w_091_018, w_091_019, w_091_022, w_091_023, w_091_024, w_091_025, w_091_026, w_091_027, w_091_034, w_091_035, w_091_036, w_091_038, w_091_039, w_091_042, w_091_044, w_091_047, w_091_050, w_091_051, w_091_052, w_091_054, w_091_058, w_091_059, w_091_060, w_091_062, w_091_066, w_091_067, w_091_068, w_091_069, w_091_070, w_091_071, w_091_072, w_091_074, w_091_075, w_091_076, w_091_077, w_091_081, w_091_083, w_091_084, w_091_085, w_091_088, w_091_089, w_091_090, w_091_092, w_091_094, w_091_097, w_091_098, w_091_099, w_091_101, w_091_105, w_091_106, w_091_108, w_091_110, w_091_112, w_091_113, w_091_114, w_091_115, w_091_119, w_091_120, w_091_122, w_091_123, w_091_126, w_091_127, w_091_128, w_091_129, w_091_131, w_091_132, w_091_135, w_091_136, w_091_137, w_091_142, w_091_143, w_091_146, w_091_148, w_091_152, w_091_153, w_091_154, w_091_155, w_091_156, w_091_160, w_091_161, w_091_165, w_091_167, w_091_168, w_091_171, w_091_172, w_091_173, w_091_175, w_091_176, w_091_179, w_091_186, w_091_190, w_091_192, w_091_193, w_091_205, w_091_207, w_091_209, w_091_213, w_091_214, w_091_216, w_091_221, w_091_225, w_091_226, w_091_229, w_091_233, w_091_235, w_091_236, w_091_237, w_091_239, w_091_241, w_091_242, w_091_243, w_091_249, w_091_250, w_091_253, w_091_255, w_091_257, w_091_258, w_091_259, w_091_262, w_091_263, w_091_265, w_091_266, w_091_267, w_091_270, w_091_271, w_091_272, w_091_274, w_091_275, w_091_278, w_091_280, w_091_281, w_091_282, w_091_283, w_091_286, w_091_288, w_091_289, w_091_291, w_091_293, w_091_294, w_091_295, w_091_296, w_091_297, w_091_299, w_091_300, w_091_302, w_091_304, w_091_305, w_091_307, w_091_308, w_091_311, w_091_313, w_091_314, w_091_316, w_091_320, w_091_321, w_091_322, w_091_324, w_091_325, w_091_326, w_091_327, w_091_330, w_091_331, w_091_334, w_091_335, w_091_337, w_091_338, w_091_339, w_091_342, w_091_343, w_091_345, w_091_346, w_091_351, w_091_352, w_091_354, w_091_357, w_091_362, w_091_363, w_091_364, w_091_365, w_091_366, w_091_368, w_091_369, w_091_370, w_091_377, w_091_380, w_091_384, w_091_385, w_091_388, w_091_394, w_091_395, w_091_396, w_091_397, w_091_400, w_091_402, w_091_403, w_091_405, w_091_407, w_091_408, w_091_410, w_091_411, w_091_413, w_091_414, w_091_417, w_091_419, w_091_421, w_091_422, w_091_423, w_091_424, w_091_425, w_091_426, w_091_432, w_091_433, w_091_436, w_091_438, w_091_441, w_091_444, w_091_447, w_091_448, w_091_451, w_091_454, w_091_455, w_091_456, w_091_457, w_091_458, w_091_461, w_091_466, w_091_467, w_091_468, w_091_470, w_091_471, w_091_476, w_091_478, w_091_479, w_091_480, w_091_481, w_091_482, w_091_486, w_091_488, w_091_490, w_091_491, w_091_492, w_091_493, w_091_497, w_091_498, w_091_500, w_091_501, w_091_502, w_091_510, w_091_513, w_091_514, w_091_518, w_091_521, w_091_523, w_091_526, w_091_527, w_091_528, w_091_531, w_091_533, w_091_534, w_091_535, w_091_536, w_091_537, w_091_538, w_091_539, w_091_541, w_091_544, w_091_548, w_091_549, w_091_550, w_091_551, w_091_552, w_091_553, w_091_555, w_091_556, w_091_558, w_091_559, w_091_560, w_091_562, w_091_565, w_091_567, w_091_569, w_091_570, w_091_572, w_091_573, w_091_576, w_091_578, w_091_582, w_091_583, w_091_589, w_091_590, w_091_591, w_091_592, w_091_593, w_091_595, w_091_596, w_091_598, w_091_599, w_091_604, w_091_605, w_091_606, w_091_607, w_091_610, w_091_618, w_091_619, w_091_624, w_091_626, w_091_629, w_091_630, w_091_631, w_091_632, w_091_635, w_091_636, w_091_637, w_091_640, w_091_641, w_091_642, w_091_643, w_091_646, w_091_647, w_091_651, w_091_653, w_091_656, w_091_658, w_091_660, w_091_661, w_091_662, w_091_668, w_091_674, w_091_675, w_091_681, w_091_682, w_091_686, w_091_690, w_091_691, w_091_693, w_091_694, w_091_695, w_091_705, w_091_706, w_091_708, w_091_709, w_091_712, w_091_717, w_091_719, w_091_720, w_091_722, w_091_723, w_091_725, w_091_726, w_091_727, w_091_728, w_091_730, w_091_731, w_091_734, w_091_735, w_091_736, w_091_737, w_091_738, w_091_740, w_091_741, w_091_742, w_091_743, w_091_744, w_091_747, w_091_748, w_091_749, w_091_750, w_091_755, w_091_760, w_091_762, w_091_764, w_091_766, w_091_767, w_091_768, w_091_769, w_091_771, w_091_772, w_091_777, w_091_778, w_091_779, w_091_780, w_091_781, w_091_782, w_091_786, w_091_789, w_091_792, w_091_793, w_091_794, w_091_795, w_091_797, w_091_798, w_091_799, w_091_801, w_091_804, w_091_805, w_091_806, w_091_808, w_091_809, w_091_811, w_091_816, w_091_818, w_091_821, w_091_822, w_091_823, w_091_827, w_091_828, w_091_829, w_091_830, w_091_831, w_091_832, w_091_834, w_091_840, w_091_841, w_091_842, w_091_845, w_091_846, w_091_847, w_091_849, w_091_850, w_091_851, w_091_853, w_091_863, w_091_866, w_091_867, w_091_869, w_091_870, w_091_874, w_091_875, w_091_876, w_091_877, w_091_878, w_091_879, w_091_881, w_091_882, w_091_883, w_091_885, w_091_886, w_091_887, w_091_889, w_091_890, w_091_892, w_091_893, w_091_897, w_091_898, w_091_901, w_091_903, w_091_904, w_091_907, w_091_908, w_091_913, w_091_918, w_091_919, w_091_920, w_091_922, w_091_923, w_091_924, w_091_925, w_091_926, w_091_927, w_091_928, w_091_929, w_091_930, w_091_931, w_091_932, w_091_933, w_091_935, w_091_936, w_091_938, w_091_940, w_091_941, w_091_943, w_091_944, w_091_945, w_091_946, w_091_947, w_091_948, w_091_949, w_091_950, w_091_952, w_091_954, w_091_956, w_091_957, w_091_959, w_091_960, w_091_964, w_091_965, w_091_966, w_091_967, w_091_970, w_091_971, w_091_973, w_091_974, w_091_977, w_091_979, w_091_980, w_091_982, w_091_984, w_091_985, w_091_986, w_091_987, w_091_990, w_091_994, w_091_998, w_091_999, w_091_1005, w_091_1006, w_091_1010, w_091_1011, w_091_1012, w_091_1015, w_091_1017, w_091_1019, w_091_1020, w_091_1021, w_091_1025, w_091_1026, w_091_1032, w_091_1033, w_091_1034, w_091_1035, w_091_1037, w_091_1038, w_091_1039, w_091_1040, w_091_1046, w_091_1047, w_091_1051, w_091_1053, w_091_1057, w_091_1058, w_091_1059, w_091_1061, w_091_1062, w_091_1066, w_091_1070, w_091_1071, w_091_1072, w_091_1073, w_091_1075, w_091_1081, w_091_1082, w_091_1084, w_091_1087, w_091_1090, w_091_1091, w_091_1094, w_091_1096, w_091_1097, w_091_1098, w_091_1099, w_091_1102, w_091_1103, w_091_1105, w_091_1106, w_091_1107, w_091_1108, w_091_1112, w_091_1113, w_091_1114, w_091_1115, w_091_1116, w_091_1117, w_091_1118, w_091_1123, w_091_1128, w_091_1130, w_091_1131, w_091_1133, w_091_1134, w_091_1137, w_091_1138, w_091_1139, w_091_1140, w_091_1143, w_091_1144, w_091_1145, w_091_1146, w_091_1147, w_091_1148, w_091_1152, w_091_1155, w_091_1156, w_091_1161, w_091_1162, w_091_1165, w_091_1166, w_091_1168, w_091_1174, w_091_1175, w_091_1178, w_091_1179, w_091_1181, w_091_1182, w_091_1184, w_091_1185, w_091_1187, w_091_1189, w_091_1192, w_091_1193, w_091_1194, w_091_1198, w_091_1199, w_091_1201, w_091_1207, w_091_1209, w_091_1212, w_091_1213, w_091_1215, w_091_1216, w_091_1219, w_091_1220, w_091_1221, w_091_1222, w_091_1223, w_091_1225, w_091_1227, w_091_1228, w_091_1229, w_091_1230, w_091_1233, w_091_1234, w_091_1237, w_091_1242, w_091_1244, w_091_1245, w_091_1246, w_091_1247, w_091_1249, w_091_1252, w_091_1253, w_091_1254, w_091_1255, w_091_1256, w_091_1257, w_091_1259, w_091_1260, w_091_1263, w_091_1264, w_091_1268, w_091_1269, w_091_1270, w_091_1271, w_091_1272, w_091_1277, w_091_1279, w_091_1280, w_091_1284, w_091_1286, w_091_1287, w_091_1288, w_091_1290, w_091_1292, w_091_1293, w_091_1294, w_091_1295, w_091_1296, w_091_1297, w_091_1298, w_091_1300, w_091_1302, w_091_1303, w_091_1305, w_091_1307, w_091_1308, w_091_1309, w_091_1310, w_091_1315, w_091_1317, w_091_1318, w_091_1324, w_091_1325, w_091_1327, w_091_1328, w_091_1329, w_091_1330, w_091_1331, w_091_1334, w_091_1341, w_091_1342, w_091_1346, w_091_1347, w_091_1348, w_091_1349, w_091_1350, w_091_1352, w_091_1353, w_091_1354, w_091_1355, w_091_1357, w_091_1361, w_091_1365, w_091_1367, w_091_1370, w_091_1371, w_091_1373, w_091_1374, w_091_1376, w_091_1382, w_091_1383, w_091_1384, w_091_1386, w_091_1387, w_091_1389, w_091_1392, w_091_1394, w_091_1396, w_091_1397, w_091_1402, w_091_1403, w_091_1404, w_091_1405, w_091_1406, w_091_1407, w_091_1409, w_091_1410, w_091_1412, w_091_1418, w_091_1420, w_091_1421, w_091_1422, w_091_1423, w_091_1425, w_091_1427, w_091_1428, w_091_1430, w_091_1432, w_091_1433, w_091_1434, w_091_1435, w_091_1437, w_091_1440, w_091_1443, w_091_1444, w_091_1445, w_091_1447, w_091_1453, w_091_1456, w_091_1459, w_091_1460, w_091_1461, w_091_1462, w_091_1463, w_091_1465, w_091_1466, w_091_1467, w_091_1473, w_091_1474, w_091_1475, w_091_1476, w_091_1477, w_091_1478, w_091_1480, w_091_1486, w_091_1487, w_091_1491, w_091_1498, w_091_1499, w_091_1503, w_091_1507, w_091_1508, w_091_1510, w_091_1511, w_091_1512, w_091_1517, w_091_1518, w_091_1520, w_091_1525, w_091_1526, w_091_1527, w_091_1528, w_091_1529, w_091_1531, w_091_1533, w_091_1534, w_091_1535, w_091_1536, w_091_1537, w_091_1540, w_091_1543, w_091_1544, w_091_1545, w_091_1546, w_091_1549, w_091_1551, w_091_1552, w_091_1553, w_091_1557, w_091_1559, w_091_1560, w_091_1561, w_091_1564, w_091_1565, w_091_1566, w_091_1568, w_091_1569, w_091_1570, w_091_1571, w_091_1572, w_091_1574, w_091_1577, w_091_1581, w_091_1582, w_091_1584, w_091_1586, w_091_1588, w_091_1589, w_091_1590, w_091_1591, w_091_1594, w_091_1597, w_091_1598, w_091_1600, w_091_1602, w_091_1604, w_091_1608, w_091_1610, w_091_1611, w_091_1612, w_091_1613, w_091_1615, w_091_1616, w_091_1620, w_091_1622, w_091_1623, w_091_1624, w_091_1627, w_091_1629, w_091_1630, w_091_1632, w_091_1633, w_091_1634, w_091_1640, w_091_1644, w_091_1646, w_091_1647, w_091_1650, w_091_1651, w_091_1653, w_091_1654, w_091_1655, w_091_1658, w_091_1660, w_091_1661, w_091_1662, w_091_1663, w_091_1664, w_091_1665, w_091_1666, w_091_1667, w_091_1668, w_091_1669, w_091_1672, w_091_1673, w_091_1674, w_091_1676, w_091_1677, w_091_1679, w_091_1682, w_091_1683, w_091_1685, w_091_1686, w_091_1688, w_091_1689, w_091_1690, w_091_1694, w_091_1696, w_091_1698, w_091_1700, w_091_1701, w_091_1702, w_091_1703, w_091_1705, w_091_1708, w_091_1711, w_091_1714, w_091_1715, w_091_1723, w_091_1725, w_091_1726, w_091_1728, w_091_1732, w_091_1733, w_091_1736, w_091_1738, w_091_1739, w_091_1742, w_091_1744, w_091_1745, w_091_1747, w_091_1748, w_091_1750, w_091_1752, w_091_1754, w_091_1755, w_091_1758, w_091_1759, w_091_1761, w_091_1763, w_091_1764, w_091_1766, w_091_1769, w_091_1770, w_091_1771, w_091_1772, w_091_1776, w_091_1777, w_091_1779, w_091_1781, w_091_1783, w_091_1786, w_091_1787, w_091_1788, w_091_1789, w_091_1791, w_091_1792, w_091_1793, w_091_1795, w_091_1798, w_091_1799, w_091_1802, w_091_1803, w_091_1805, w_091_1806, w_091_1808, w_091_1809, w_091_1813, w_091_1815, w_091_1816, w_091_1817, w_091_1818, w_091_1819, w_091_1821, w_091_1825, w_091_1826, w_091_1827, w_091_1828, w_091_1829, w_091_1831, w_091_1832, w_091_1833, w_091_1836, w_091_1837, w_091_1840, w_091_1841, w_091_1847, w_091_1848, w_091_1849, w_091_1851, w_091_1853, w_091_1854, w_091_1855, w_091_1856, w_091_1861, w_091_1865, w_091_1866, w_091_1868, w_091_1869, w_091_1871, w_091_1874, w_091_1875, w_091_1876, w_091_1877, w_091_1878, w_091_1879, w_091_1881, w_091_1883, w_091_1884, w_091_1886, w_091_1887, w_091_1888, w_091_1891, w_091_1892, w_091_1895, w_091_1896, w_091_1897, w_091_1898, w_091_1901, w_091_1902, w_091_1904, w_091_1908, w_091_1909, w_091_1911, w_091_1912, w_091_1915, w_091_1916, w_091_1917, w_091_1918, w_091_1919, w_091_1920, w_091_1923, w_091_1924, w_091_1925, w_091_1927, w_091_1928, w_091_1930, w_091_1932, w_091_1933, w_091_1934, w_091_1936, w_091_1938, w_091_1940, w_091_1943, w_091_1944, w_091_1950, w_091_1956, w_091_1963, w_091_1964, w_091_1966, w_091_1972, w_091_1973, w_091_1974, w_091_1978, w_091_1979, w_091_1982, w_091_1985, w_091_1986, w_091_1988, w_091_1989, w_091_1991, w_091_1993, w_091_1996, w_091_1998, w_091_2010, w_091_2011, w_091_2013, w_091_2017, w_091_2024, w_091_2025, w_091_2026, w_091_2028, w_091_2029, w_091_2030, w_091_2032, w_091_2033, w_091_2034, w_091_2035, w_091_2039, w_091_2040, w_091_2041, w_091_2042, w_091_2044, w_091_2051, w_091_2055, w_091_2062, w_091_2083, w_091_2084, w_091_2085, w_091_2086, w_091_2097, w_091_2098, w_091_2115, w_091_2121, w_091_2122, w_091_2123, w_091_2125, w_091_2126, w_091_2141, w_091_2151, w_091_2155, w_091_2172, w_091_2173, w_091_2179, w_091_2188, w_091_2192, w_091_2193, w_091_2195, w_091_2196, w_091_2198, w_091_2202, w_091_2203, w_091_2208, w_091_2214, w_091_2218, w_091_2219, w_091_2221, w_091_2223, w_091_2229, w_091_2234, w_091_2235, w_091_2236, w_091_2238, w_091_2241, w_091_2248, w_091_2255, w_091_2256, w_091_2257, w_091_2258, w_091_2264, w_091_2267, w_091_2270, w_091_2273, w_091_2278, w_091_2280, w_091_2284, w_091_2287, w_091_2292, w_091_2301, w_091_2304, w_091_2309, w_091_2312, w_091_2313, w_091_2317, w_091_2319, w_091_2321, w_091_2322, w_091_2327, w_091_2329, w_091_2339, w_091_2341, w_091_2342, w_091_2343, w_091_2344, w_091_2345, w_091_2353, w_091_2354, w_091_2360, w_091_2365, w_091_2371, w_091_2373, w_091_2376, w_091_2382, w_091_2383, w_091_2385, w_091_2386, w_091_2391, w_091_2398, w_091_2403, w_091_2404, w_091_2409, w_091_2411, w_091_2415, w_091_2416, w_091_2419, w_091_2421, w_091_2426, w_091_2429, w_091_2434, w_091_2437, w_091_2438, w_091_2440, w_091_2446, w_091_2449, w_091_2452, w_091_2454, w_091_2467, w_091_2468, w_091_2473, w_091_2477, w_091_2478, w_091_2483, w_091_2487, w_091_2492, w_091_2494, w_091_2495, w_091_2496, w_091_2499, w_091_2502, w_091_2503, w_091_2504, w_091_2505, w_091_2506, w_091_2508, w_091_2510, w_091_2512, w_091_2515, w_091_2520, w_091_2526, w_091_2528, w_091_2531, w_091_2532, w_091_2533, w_091_2540, w_091_2546, w_091_2549, w_091_2550, w_091_2557, w_091_2559, w_091_2564, w_091_2568, w_091_2569, w_091_2570, w_091_2571, w_091_2573, w_091_2578, w_091_2581, w_091_2588, w_091_2589, w_091_2590, w_091_2593, w_091_2598, w_091_2605, w_091_2612, w_091_2618, w_091_2620, w_091_2622, w_091_2623, w_091_2625, w_091_2628, w_091_2630, w_091_2632, w_091_2639, w_091_2640, w_091_2642, w_091_2647, w_091_2653, w_091_2654, w_091_2664, w_091_2666, w_091_2670, w_091_2671, w_091_2674, w_091_2678, w_091_2679, w_091_2681, w_091_2685, w_091_2687, w_091_2691, w_091_2692, w_091_2693, w_091_2694, w_091_2695, w_091_2696, w_091_2697, w_091_2698, w_091_2701, w_091_2707, w_091_2710, w_091_2713, w_091_2714, w_091_2716, w_091_2717, w_091_2718, w_091_2719, w_091_2723, w_091_2729, w_091_2733, w_091_2734, w_091_2735, w_091_2737, w_091_2744, w_091_2750, w_091_2753, w_091_2758, w_091_2762, w_091_2767, w_091_2769, w_091_2775, w_091_2784, w_091_2785, w_091_2786, w_091_2789, w_091_2794, w_091_2796, w_091_2801, w_091_2803, w_091_2807, w_091_2808, w_091_2809, w_091_2812, w_091_2818, w_091_2824, w_091_2830, w_091_2831, w_091_2833, w_091_2838, w_091_2839, w_091_2844, w_091_2845, w_091_2850, w_091_2856, w_091_2857, w_091_2859, w_091_2863, w_091_2864, w_091_2868, w_091_2869, w_091_2870, w_091_2875, w_091_2877, w_091_2883, w_091_2884, w_091_2885, w_091_2886, w_091_2887, w_091_2888, w_091_2891, w_091_2892, w_091_2898, w_091_2902, w_091_2906, w_091_2909, w_091_2917, w_091_2921, w_091_2922, w_091_2924, w_091_2925, w_091_2928, w_091_2929, w_091_2932, w_091_2940, w_091_2941, w_091_2943, w_091_2949, w_091_2950, w_091_2952, w_091_2953, w_091_2954, w_091_2957, w_091_2966, w_091_2967, w_091_2969, w_091_2972, w_091_2973, w_091_2974, w_091_2975, w_091_2980, w_091_2983, w_091_2987, w_091_2990, w_091_2991, w_091_2994, w_091_2996, w_091_2998, w_091_3002, w_091_3003, w_091_3007, w_091_3009, w_091_3025, w_091_3029, w_091_3030, w_091_3032, w_091_3035, w_091_3037, w_091_3041, w_091_3042, w_091_3045, w_091_3046, w_091_3049, w_091_3053, w_091_3056, w_091_3057, w_091_3058, w_091_3059, w_091_3060, w_091_3064, w_091_3065, w_091_3066, w_091_3068;
  wire w_092_001, w_092_004, w_092_008, w_092_010, w_092_015, w_092_019, w_092_020, w_092_024, w_092_026, w_092_030, w_092_031, w_092_032, w_092_035, w_092_038, w_092_040, w_092_044, w_092_045, w_092_047, w_092_048, w_092_055, w_092_058, w_092_059, w_092_061, w_092_062, w_092_063, w_092_066, w_092_067, w_092_069, w_092_071, w_092_072, w_092_073, w_092_074, w_092_075, w_092_076, w_092_080, w_092_081, w_092_082, w_092_083, w_092_088, w_092_091, w_092_093, w_092_095, w_092_096, w_092_097, w_092_098, w_092_100, w_092_102, w_092_104, w_092_107, w_092_109, w_092_110, w_092_111, w_092_113, w_092_114, w_092_115, w_092_118, w_092_119, w_092_120, w_092_122, w_092_123, w_092_124, w_092_125, w_092_126, w_092_127, w_092_128, w_092_129, w_092_130, w_092_131, w_092_133, w_092_135, w_092_136, w_092_138, w_092_140, w_092_142, w_092_143, w_092_144, w_092_145, w_092_146, w_092_148, w_092_153, w_092_155, w_092_156, w_092_157, w_092_162, w_092_163, w_092_164, w_092_166, w_092_167, w_092_170, w_092_175, w_092_179, w_092_180, w_092_181, w_092_183, w_092_187, w_092_189, w_092_190, w_092_191, w_092_192, w_092_195, w_092_197, w_092_199, w_092_200, w_092_201, w_092_216, w_092_222, w_092_223, w_092_225, w_092_227, w_092_231, w_092_234, w_092_236, w_092_238, w_092_246, w_092_248, w_092_250, w_092_251, w_092_255, w_092_257, w_092_260, w_092_261, w_092_262, w_092_263, w_092_264, w_092_267, w_092_270, w_092_274, w_092_275, w_092_279, w_092_283, w_092_286, w_092_288, w_092_292, w_092_294, w_092_297, w_092_298, w_092_299, w_092_305, w_092_311, w_092_313, w_092_321, w_092_331, w_092_333, w_092_334, w_092_344, w_092_345, w_092_348, w_092_364, w_092_365, w_092_372, w_092_374, w_092_375, w_092_379, w_092_380, w_092_381, w_092_383, w_092_385, w_092_387, w_092_388, w_092_394, w_092_398, w_092_401, w_092_403, w_092_411, w_092_413, w_092_417, w_092_421, w_092_424, w_092_432, w_092_433, w_092_435, w_092_443, w_092_449, w_092_459, w_092_460, w_092_464, w_092_466, w_092_467, w_092_470, w_092_471, w_092_475, w_092_482, w_092_484, w_092_488, w_092_492, w_092_496, w_092_498, w_092_500, w_092_509, w_092_512, w_092_514, w_092_518, w_092_530, w_092_533, w_092_535, w_092_537, w_092_539, w_092_542, w_092_550, w_092_551, w_092_561, w_092_564, w_092_570, w_092_573, w_092_579, w_092_583, w_092_584, w_092_586, w_092_587, w_092_590, w_092_593, w_092_595, w_092_596, w_092_603, w_092_605, w_092_607, w_092_608, w_092_609, w_092_615, w_092_626, w_092_631, w_092_632, w_092_633, w_092_636, w_092_637, w_092_642, w_092_646, w_092_653, w_092_656, w_092_657, w_092_659, w_092_665, w_092_668, w_092_676, w_092_690, w_092_691, w_092_700, w_092_701, w_092_707, w_092_712, w_092_715, w_092_716, w_092_720, w_092_722, w_092_725, w_092_728, w_092_729, w_092_737, w_092_744, w_092_745, w_092_746, w_092_748, w_092_751, w_092_757, w_092_760, w_092_762, w_092_768, w_092_769, w_092_771, w_092_772, w_092_773, w_092_775, w_092_778, w_092_781, w_092_787, w_092_790, w_092_792, w_092_794, w_092_798, w_092_801, w_092_808, w_092_811, w_092_813, w_092_816, w_092_819, w_092_822, w_092_823, w_092_825, w_092_826, w_092_828, w_092_835, w_092_839, w_092_840, w_092_842, w_092_843, w_092_846, w_092_848, w_092_849, w_092_851, w_092_854, w_092_855, w_092_861, w_092_866, w_092_870, w_092_874, w_092_875, w_092_876, w_092_879, w_092_881, w_092_887, w_092_888, w_092_894, w_092_896, w_092_898, w_092_900, w_092_902, w_092_920, w_092_932, w_092_935, w_092_936, w_092_941, w_092_946, w_092_948, w_092_952, w_092_956, w_092_958, w_092_959, w_092_960, w_092_962, w_092_963, w_092_964, w_092_971, w_092_972, w_092_974, w_092_982, w_092_983, w_092_984, w_092_985, w_092_986, w_092_989, w_092_990, w_092_992, w_092_995, w_092_1000, w_092_1002, w_092_1012, w_092_1015, w_092_1018, w_092_1022, w_092_1023, w_092_1026, w_092_1027, w_092_1030, w_092_1033, w_092_1036, w_092_1037, w_092_1038, w_092_1039, w_092_1041, w_092_1042, w_092_1052, w_092_1053, w_092_1058, w_092_1060, w_092_1065, w_092_1068, w_092_1072, w_092_1074, w_092_1075, w_092_1076, w_092_1078, w_092_1081, w_092_1082, w_092_1083, w_092_1086, w_092_1089, w_092_1094, w_092_1097, w_092_1099, w_092_1102, w_092_1103, w_092_1110, w_092_1118, w_092_1120, w_092_1133, w_092_1140, w_092_1143, w_092_1145, w_092_1148, w_092_1149, w_092_1151, w_092_1152, w_092_1153, w_092_1154, w_092_1159, w_092_1164, w_092_1165, w_092_1174, w_092_1180, w_092_1184, w_092_1192, w_092_1196, w_092_1200, w_092_1201, w_092_1207, w_092_1208, w_092_1210, w_092_1213, w_092_1215, w_092_1218, w_092_1219, w_092_1221, w_092_1226, w_092_1229, w_092_1230, w_092_1239, w_092_1241, w_092_1246, w_092_1247, w_092_1250, w_092_1253, w_092_1255, w_092_1259, w_092_1262, w_092_1264, w_092_1266, w_092_1267, w_092_1269, w_092_1277, w_092_1281, w_092_1283, w_092_1286, w_092_1287, w_092_1294, w_092_1300, w_092_1301, w_092_1308, w_092_1309, w_092_1313, w_092_1320, w_092_1327, w_092_1330, w_092_1334, w_092_1336, w_092_1337, w_092_1338, w_092_1340, w_092_1341, w_092_1350, w_092_1351, w_092_1352, w_092_1353, w_092_1358, w_092_1362, w_092_1366, w_092_1367, w_092_1370, w_092_1371, w_092_1374, w_092_1381, w_092_1382, w_092_1385, w_092_1386, w_092_1400, w_092_1401, w_092_1402, w_092_1404, w_092_1406, w_092_1414, w_092_1415, w_092_1417, w_092_1418, w_092_1422, w_092_1424, w_092_1426, w_092_1429, w_092_1432, w_092_1434, w_092_1437, w_092_1440, w_092_1441, w_092_1445, w_092_1446, w_092_1449, w_092_1456, w_092_1457, w_092_1458, w_092_1466, w_092_1468, w_092_1474, w_092_1475, w_092_1481, w_092_1484, w_092_1486, w_092_1490, w_092_1491, w_092_1494, w_092_1502, w_092_1506, w_092_1507, w_092_1510, w_092_1512, w_092_1516, w_092_1517, w_092_1519, w_092_1521, w_092_1522, w_092_1525, w_092_1530, w_092_1535, w_092_1538, w_092_1539, w_092_1541, w_092_1542, w_092_1545, w_092_1550, w_092_1551, w_092_1555, w_092_1564, w_092_1572, w_092_1576, w_092_1579, w_092_1580, w_092_1581, w_092_1592, w_092_1594, w_092_1604, w_092_1614, w_092_1617, w_092_1618, w_092_1629, w_092_1630, w_092_1631, w_092_1637, w_092_1638, w_092_1641, w_092_1643, w_092_1644, w_092_1649, w_092_1650, w_092_1655, w_092_1664, w_092_1665, w_092_1666, w_092_1678, w_092_1680, w_092_1683, w_092_1684, w_092_1685, w_092_1688, w_092_1689, w_092_1693, w_092_1698, w_092_1699, w_092_1708, w_092_1712, w_092_1715, w_092_1723, w_092_1724, w_092_1727, w_092_1728, w_092_1731, w_092_1735, w_092_1738, w_092_1739, w_092_1741, w_092_1742, w_092_1746, w_092_1751, w_092_1763, w_092_1766, w_092_1771, w_092_1772, w_092_1775, w_092_1777, w_092_1779, w_092_1780, w_092_1787, w_092_1795, w_092_1798, w_092_1802, w_092_1805, w_092_1807, w_092_1810, w_092_1813, w_092_1825, w_092_1826, w_092_1829, w_092_1830, w_092_1835, w_092_1840, w_092_1847, w_092_1849, w_092_1855, w_092_1859, w_092_1863, w_092_1865, w_092_1868, w_092_1875, w_092_1878, w_092_1880, w_092_1882, w_092_1889, w_092_1891, w_092_1897, w_092_1900, w_092_1906, w_092_1909, w_092_1911, w_092_1913, w_092_1915, w_092_1916, w_092_1925, w_092_1933, w_092_1934, w_092_1936, w_092_1937, w_092_1942, w_092_1943, w_092_1952, w_092_1954, w_092_1960, w_092_1963, w_092_1966, w_092_1971, w_092_1974, w_092_1976, w_092_1979, w_092_1982, w_092_1985, w_092_1987, w_092_1990, w_092_1991, w_092_1992, w_092_1993, w_092_1994, w_092_1996, w_092_1998, w_092_2003, w_092_2006, w_092_2008, w_092_2014, w_092_2019, w_092_2022, w_092_2026, w_092_2031, w_092_2032, w_092_2034, w_092_2044, w_092_2050, w_092_2052, w_092_2053, w_092_2055, w_092_2059, w_092_2060, w_092_2061, w_092_2066, w_092_2068, w_092_2069, w_092_2070, w_092_2072, w_092_2079, w_092_2080, w_092_2084, w_092_2093, w_092_2096, w_092_2098, w_092_2102, w_092_2104, w_092_2110, w_092_2115, w_092_2120, w_092_2129, w_092_2130, w_092_2132, w_092_2136, w_092_2138, w_092_2149, w_092_2150, w_092_2152, w_092_2153, w_092_2160, w_092_2163, w_092_2164, w_092_2167, w_092_2168, w_092_2171, w_092_2173, w_092_2174, w_092_2177, w_092_2182, w_092_2183, w_092_2184, w_092_2185, w_092_2188, w_092_2189, w_092_2193, w_092_2198, w_092_2200, w_092_2201, w_092_2204, w_092_2205, w_092_2209, w_092_2211, w_092_2213, w_092_2215, w_092_2219, w_092_2220, w_092_2223, w_092_2226, w_092_2233, w_092_2238, w_092_2241, w_092_2242, w_092_2246, w_092_2249, w_092_2258, w_092_2259, w_092_2267, w_092_2270, w_092_2271, w_092_2273, w_092_2274, w_092_2275, w_092_2278, w_092_2279, w_092_2280, w_092_2281, w_092_2289, w_092_2292, w_092_2297, w_092_2298, w_092_2302, w_092_2304, w_092_2310, w_092_2324, w_092_2326, w_092_2335, w_092_2339, w_092_2345, w_092_2347, w_092_2352, w_092_2355, w_092_2356, w_092_2364, w_092_2369, w_092_2370, w_092_2374, w_092_2379, w_092_2383, w_092_2386, w_092_2387, w_092_2392, w_092_2394, w_092_2398, w_092_2400, w_092_2405, w_092_2406, w_092_2415, w_092_2418, w_092_2420, w_092_2423, w_092_2425, w_092_2426, w_092_2429, w_092_2431, w_092_2435, w_092_2438, w_092_2439, w_092_2447, w_092_2448, w_092_2453, w_092_2461, w_092_2462, w_092_2463, w_092_2465, w_092_2473, w_092_2481, w_092_2483, w_092_2489, w_092_2491, w_092_2497, w_092_2503, w_092_2509, w_092_2510, w_092_2511, w_092_2514, w_092_2515, w_092_2516, w_092_2518, w_092_2527, w_092_2533, w_092_2537, w_092_2540, w_092_2542, w_092_2546, w_092_2549, w_092_2550, w_092_2554, w_092_2555, w_092_2559, w_092_2560, w_092_2561, w_092_2565, w_092_2568, w_092_2571, w_092_2573, w_092_2578, w_092_2581, w_092_2582, w_092_2586, w_092_2587, w_092_2590, w_092_2591, w_092_2592, w_092_2594, w_092_2598, w_092_2601, w_092_2611, w_092_2614, w_092_2618, w_092_2621, w_092_2625, w_092_2630, w_092_2634, w_092_2636, w_092_2637, w_092_2638, w_092_2640, w_092_2642, w_092_2646, w_092_2649, w_092_2650, w_092_2658, w_092_2659, w_092_2661, w_092_2663, w_092_2666, w_092_2668, w_092_2669, w_092_2670, w_092_2672, w_092_2675, w_092_2676, w_092_2682, w_092_2686, w_092_2687, w_092_2694, w_092_2695, w_092_2700, w_092_2708, w_092_2711, w_092_2716, w_092_2719, w_092_2722, w_092_2724, w_092_2726, w_092_2729, w_092_2730, w_092_2731, w_092_2734, w_092_2735, w_092_2742, w_092_2746, w_092_2748, w_092_2759, w_092_2762, w_092_2765, w_092_2766, w_092_2772, w_092_2775, w_092_2776, w_092_2778, w_092_2782, w_092_2783, w_092_2785, w_092_2786, w_092_2792, w_092_2796, w_092_2801, w_092_2808, w_092_2813, w_092_2816, w_092_2818, w_092_2819, w_092_2824, w_092_2827, w_092_2830, w_092_2831, w_092_2833, w_092_2838, w_092_2846, w_092_2848, w_092_2849, w_092_2851, w_092_2857, w_092_2859, w_092_2860, w_092_2865, w_092_2868, w_092_2869, w_092_2871, w_092_2872, w_092_2873, w_092_2878, w_092_2884, w_092_2889, w_092_2890, w_092_2894, w_092_2896, w_092_2897, w_092_2902, w_092_2904, w_092_2906, w_092_2909, w_092_2912, w_092_2917, w_092_2924, w_092_2927, w_092_2932, w_092_2937, w_092_2945, w_092_2950, w_092_2952, w_092_2956, w_092_2960, w_092_2963, w_092_2966, w_092_2968, w_092_2970, w_092_2971, w_092_2975, w_092_2978, w_092_2979, w_092_2988, w_092_2989, w_092_2992, w_092_2997, w_092_2998, w_092_3000, w_092_3006, w_092_3007, w_092_3008, w_092_3015, w_092_3022, w_092_3025, w_092_3027, w_092_3029, w_092_3030, w_092_3035, w_092_3037, w_092_3045, w_092_3046, w_092_3051, w_092_3055, w_092_3057, w_092_3058, w_092_3060, w_092_3070, w_092_3072, w_092_3074, w_092_3078, w_092_3084, w_092_3089, w_092_3093, w_092_3098, w_092_3101, w_092_3105, w_092_3107, w_092_3109, w_092_3111, w_092_3112, w_092_3117, w_092_3118, w_092_3122, w_092_3128, w_092_3130, w_092_3131, w_092_3147, w_092_3152, w_092_3163, w_092_3171, w_092_3174, w_092_3175, w_092_3177, w_092_3182, w_092_3183, w_092_3184, w_092_3186, w_092_3189, w_092_3194, w_092_3200, w_092_3209, w_092_3210, w_092_3212, w_092_3215, w_092_3216, w_092_3217, w_092_3220, w_092_3221, w_092_3222, w_092_3224, w_092_3229, w_092_3231, w_092_3235, w_092_3237, w_092_3240, w_092_3243, w_092_3245, w_092_3248, w_092_3256, w_092_3260, w_092_3263, w_092_3264, w_092_3265, w_092_3269, w_092_3271, w_092_3273, w_092_3274, w_092_3275, w_092_3276, w_092_3277, w_092_3278, w_092_3285, w_092_3293, w_092_3295, w_092_3296, w_092_3298, w_092_3301, w_092_3302, w_092_3307, w_092_3308, w_092_3310, w_092_3314, w_092_3315, w_092_3321, w_092_3324, w_092_3326, w_092_3327, w_092_3331, w_092_3334, w_092_3335, w_092_3336, w_092_3338, w_092_3340, w_092_3349, w_092_3351, w_092_3352, w_092_3357, w_092_3364, w_092_3365, w_092_3366, w_092_3369, w_092_3376, w_092_3377, w_092_3378, w_092_3381, w_092_3382, w_092_3383, w_092_3387, w_092_3395, w_092_3397, w_092_3399, w_092_3400, w_092_3402, w_092_3404, w_092_3405, w_092_3408, w_092_3409, w_092_3421, w_092_3422, w_092_3424, w_092_3427, w_092_3429, w_092_3431, w_092_3432, w_092_3439, w_092_3447, w_092_3449, w_092_3455, w_092_3456, w_092_3458, w_092_3460, w_092_3461, w_092_3464, w_092_3469, w_092_3470, w_092_3480, w_092_3484, w_092_3485, w_092_3488, w_092_3489, w_092_3490, w_092_3492, w_092_3493, w_092_3505, w_092_3508, w_092_3514, w_092_3520, w_092_3529, w_092_3532, w_092_3537, w_092_3543, w_092_3546, w_092_3547, w_092_3550, w_092_3551, w_092_3553, w_092_3557, w_092_3559, w_092_3563, w_092_3566, w_092_3568, w_092_3573, w_092_3577, w_092_3583, w_092_3584, w_092_3587, w_092_3590, w_092_3591, w_092_3592, w_092_3593, w_092_3595, w_092_3597, w_092_3598, w_092_3599, w_092_3601, w_092_3602, w_092_3611, w_092_3612, w_092_3615, w_092_3616, w_092_3617, w_092_3623, w_092_3629, w_092_3639, w_092_3644, w_092_3647, w_092_3652, w_092_3659, w_092_3661, w_092_3662, w_092_3663, w_092_3665, w_092_3672, w_092_3673, w_092_3674, w_092_3681, w_092_3682, w_092_3684, w_092_3688, w_092_3689, w_092_3690, w_092_3693, w_092_3705, w_092_3711, w_092_3716, w_092_3725, w_092_3727, w_092_3728, w_092_3730, w_092_3731, w_092_3736, w_092_3738, w_092_3753, w_092_3756, w_092_3757, w_092_3763, w_092_3764, w_092_3765, w_092_3769, w_092_3770, w_092_3774, w_092_3776, w_092_3779, w_092_3780, w_092_3782, w_092_3783, w_092_3785, w_092_3788, w_092_3790, w_092_3793, w_092_3798, w_092_3801, w_092_3805, w_092_3806, w_092_3808, w_092_3811, w_092_3814, w_092_3816, w_092_3817, w_092_3826, w_092_3827, w_092_3835, w_092_3836, w_092_3839, w_092_3841, w_092_3843, w_092_3844, w_092_3851, w_092_3852, w_092_3853, w_092_3855, w_092_3858, w_092_3864, w_092_3869, w_092_3875, w_092_3876, w_092_3880, w_092_3883, w_092_3884, w_092_3885, w_092_3886, w_092_3887, w_092_3890, w_092_3898, w_092_3899, w_092_3901, w_092_3911, w_092_3913, w_092_3914, w_092_3923, w_092_3928, w_092_3929, w_092_3934, w_092_3935, w_092_3956, w_092_3958, w_092_3960, w_092_3961, w_092_3962, w_092_3964, w_092_3966, w_092_3968, w_092_3970, w_092_3971, w_092_3972, w_092_3975, w_092_3977, w_092_3981, w_092_3983, w_092_3984, w_092_3985, w_092_3988, w_092_3994, w_092_3997, w_092_4002, w_092_4004, w_092_4005, w_092_4006, w_092_4012, w_092_4013, w_092_4020, w_092_4022, w_092_4028, w_092_4030, w_092_4032, w_092_4038, w_092_4043, w_092_4048, w_092_4050, w_092_4052, w_092_4053, w_092_4054, w_092_4057, w_092_4059, w_092_4060, w_092_4062, w_092_4064, w_092_4073, w_092_4075, w_092_4086, w_092_4088, w_092_4090, w_092_4098, w_092_4101, w_092_4104, w_092_4105, w_092_4107, w_092_4109, w_092_4110, w_092_4113, w_092_4119, w_092_4120, w_092_4122, w_092_4130, w_092_4143, w_092_4144, w_092_4145, w_092_4146, w_092_4147, w_092_4149, w_092_4150, w_092_4152, w_092_4153, w_092_4157, w_092_4159, w_092_4163, w_092_4165, w_092_4172, w_092_4186, w_092_4194, w_092_4198, w_092_4199, w_092_4201, w_092_4203, w_092_4205, w_092_4207, w_092_4210, w_092_4215, w_092_4219, w_092_4220, w_092_4225, w_092_4227, w_092_4229, w_092_4234, w_092_4243, w_092_4244, w_092_4247, w_092_4249, w_092_4250, w_092_4251, w_092_4253, w_092_4254, w_092_4255, w_092_4258, w_092_4262, w_092_4265, w_092_4268, w_092_4269, w_092_4270, w_092_4271, w_092_4276, w_092_4278, w_092_4286, w_092_4289, w_092_4290, w_092_4299, w_092_4300, w_092_4303, w_092_4305, w_092_4308, w_092_4309, w_092_4310, w_092_4311, w_092_4312, w_092_4318, w_092_4319, w_092_4324, w_092_4327, w_092_4329, w_092_4331, w_092_4334, w_092_4335, w_092_4338, w_092_4342, w_092_4344, w_092_4350, w_092_4352, w_092_4357, w_092_4358, w_092_4376, w_092_4380, w_092_4381, w_092_4383, w_092_4384, w_092_4395, w_092_4396, w_092_4399, w_092_4401, w_092_4406, w_092_4407, w_092_4410, w_092_4411, w_092_4414, w_092_4415, w_092_4420, w_092_4421, w_092_4422, w_092_4424, w_092_4426, w_092_4428, w_092_4440, w_092_4448, w_092_4452, w_092_4453, w_092_4455, w_092_4456, w_092_4461, w_092_4465, w_092_4466, w_092_4467, w_092_4469, w_092_4470, w_092_4480, w_092_4481, w_092_4492, w_092_4494, w_092_4500, w_092_4509, w_092_4521, w_092_4522, w_092_4529, w_092_4533, w_092_4534, w_092_4543, w_092_4545, w_092_4546, w_092_4548, w_092_4550, w_092_4557, w_092_4560, w_092_4562, w_092_4567, w_092_4571, w_092_4572, w_092_4573, w_092_4581, w_092_4584, w_092_4588, w_092_4591, w_092_4593, w_092_4596, w_092_4599, w_092_4602, w_092_4605, w_092_4609, w_092_4616, w_092_4630, w_092_4634, w_092_4635, w_092_4639, w_092_4641, w_092_4642, w_092_4645, w_092_4646, w_092_4649, w_092_4652, w_092_4654, w_092_4663, w_092_4667, w_092_4668, w_092_4669, w_092_4672, w_092_4677, w_092_4683, w_092_4685, w_092_4689, w_092_4690, w_092_4704, w_092_4706, w_092_4707, w_092_4713, w_092_4714, w_092_4717, w_092_4725, w_092_4726, w_092_4733, w_092_4734, w_092_4735, w_092_4736, w_092_4737, w_092_4742, w_092_4744, w_092_4748, w_092_4757, w_092_4761, w_092_4762, w_092_4764, w_092_4765, w_092_4771, w_092_4774, w_092_4775, w_092_4776, w_092_4777, w_092_4782, w_092_4784, w_092_4785, w_092_4787, w_092_4788, w_092_4789, w_092_4790, w_092_4791, w_092_4794, w_092_4800, w_092_4801, w_092_4802, w_092_4803, w_092_4804, w_092_4805, w_092_4807, w_092_4809, w_092_4810, w_092_4811, w_092_4812, w_092_4813, w_092_4814, w_092_4815, w_092_4816, w_092_4817, w_092_4818, w_092_4819, w_092_4820, w_092_4822;
  wire w_093_000, w_093_001, w_093_002, w_093_003, w_093_004, w_093_005, w_093_006, w_093_007, w_093_008, w_093_009, w_093_010, w_093_011, w_093_013, w_093_015, w_093_016, w_093_017, w_093_018, w_093_021, w_093_023, w_093_024, w_093_026, w_093_027, w_093_031, w_093_033, w_093_035, w_093_036, w_093_038, w_093_039, w_093_040, w_093_042, w_093_043, w_093_044, w_093_046, w_093_050, w_093_051, w_093_053, w_093_056, w_093_057, w_093_058, w_093_059, w_093_060, w_093_061, w_093_062, w_093_063, w_093_066, w_093_068, w_093_069, w_093_070, w_093_071, w_093_072, w_093_073, w_093_075, w_093_076, w_093_077, w_093_078, w_093_081, w_093_082, w_093_085, w_093_086, w_093_087, w_093_089, w_093_091, w_093_093, w_093_096, w_093_098, w_093_102, w_093_104, w_093_105, w_093_106, w_093_109, w_093_111, w_093_112, w_093_113, w_093_115, w_093_116, w_093_117, w_093_118, w_093_119, w_093_120, w_093_121, w_093_122, w_093_127, w_093_130, w_093_132, w_093_133, w_093_134, w_093_136, w_093_138, w_093_139, w_093_140, w_093_143, w_093_144, w_093_146, w_093_147, w_093_151, w_093_152, w_093_155, w_093_156, w_093_157, w_093_159, w_093_160, w_093_165, w_093_166, w_093_167, w_093_168, w_093_169, w_093_170, w_093_173, w_093_174, w_093_175, w_093_179, w_093_180, w_093_183, w_093_184, w_093_185, w_093_186, w_093_187, w_093_190, w_093_191, w_093_192, w_093_193, w_093_194, w_093_195, w_093_197, w_093_199, w_093_200, w_093_201, w_093_202, w_093_203, w_093_204, w_093_205, w_093_206, w_093_207, w_093_208, w_093_209, w_093_210, w_093_211, w_093_212, w_093_213, w_093_214, w_093_215, w_093_216, w_093_217, w_093_220, w_093_222, w_093_224, w_093_226, w_093_227, w_093_228, w_093_229, w_093_230, w_093_232, w_093_233, w_093_235, w_093_236, w_093_237, w_093_238, w_093_239, w_093_240, w_093_241, w_093_242, w_093_243, w_093_244, w_093_246, w_093_248, w_093_249, w_093_250, w_093_251, w_093_254, w_093_255, w_093_257, w_093_259, w_093_260, w_093_261, w_093_262, w_093_263, w_093_264, w_093_267, w_093_268, w_093_269, w_093_270, w_093_271, w_093_272, w_093_274, w_093_276, w_093_279, w_093_280, w_093_281, w_093_282, w_093_283, w_093_284, w_093_285, w_093_287, w_093_289, w_093_291, w_093_292, w_093_293, w_093_296, w_093_297, w_093_299, w_093_300, w_093_301, w_093_304, w_093_305, w_093_307, w_093_308, w_093_309, w_093_311, w_093_312, w_093_313, w_093_314, w_093_316, w_093_318, w_093_319, w_093_320, w_093_323, w_093_325, w_093_326, w_093_328, w_093_330, w_093_331, w_093_332, w_093_333, w_093_334, w_093_335, w_093_336, w_093_337, w_093_338, w_093_339, w_093_340, w_093_341, w_093_342, w_093_343, w_093_344, w_093_345, w_093_347, w_093_348, w_093_349, w_093_350, w_093_352, w_093_353, w_093_354, w_093_355, w_093_356, w_093_357, w_093_358, w_093_359, w_093_362, w_093_367, w_093_368, w_093_371, w_093_372, w_093_373, w_093_374, w_093_376, w_093_378, w_093_379, w_093_380, w_093_381, w_093_382, w_093_387, w_093_389, w_093_390, w_093_392, w_093_395, w_093_396, w_093_397, w_093_399, w_093_400, w_093_401, w_093_403, w_093_405, w_093_406, w_093_407, w_093_408, w_093_410, w_093_412, w_093_413, w_093_417, w_093_421, w_093_423, w_093_424, w_093_426, w_093_427, w_093_429, w_093_430, w_093_433, w_093_434, w_093_437, w_093_438, w_093_441, w_093_442, w_093_445, w_093_448, w_093_450, w_093_455, w_093_459, w_093_460, w_093_462, w_093_464, w_093_465, w_093_467, w_093_468, w_093_471, w_093_475, w_093_478, w_093_480, w_093_483, w_093_487, w_093_488, w_093_490, w_093_493, w_093_496, w_093_497, w_093_498, w_093_500, w_093_504, w_093_507, w_093_508, w_093_510, w_093_511, w_093_512, w_093_513, w_093_514, w_093_515, w_093_516, w_093_517, w_093_519, w_093_520, w_093_521, w_093_525, w_093_526, w_093_529, w_093_530, w_093_533, w_093_534, w_093_538, w_093_540, w_093_544, w_093_548, w_093_549, w_093_550, w_093_556, w_093_559, w_093_561, w_093_562, w_093_566, w_093_570, w_093_571, w_093_572, w_093_574, w_093_577, w_093_578, w_093_579, w_093_581, w_093_582, w_093_585, w_093_589, w_093_590, w_093_591, w_093_592, w_093_599, w_093_600, w_093_602, w_093_603, w_093_605, w_093_606, w_093_608, w_093_609, w_093_611, w_093_615, w_093_616, w_093_618, w_093_619, w_093_620, w_093_621, w_093_623, w_093_626, w_093_627, w_093_628, w_093_629, w_093_630, w_093_632, w_093_633, w_093_635, w_093_637, w_093_641, w_093_643, w_093_646, w_093_649, w_093_650, w_093_651, w_093_652, w_093_655, w_093_661, w_093_662, w_093_663, w_093_667, w_093_670, w_093_676, w_093_677, w_093_678, w_093_682, w_093_683, w_093_684, w_093_686, w_093_690, w_093_691, w_093_694, w_093_696, w_093_697, w_093_698, w_093_706, w_093_708, w_093_709, w_093_710, w_093_713, w_093_717, w_093_722, w_093_726, w_093_729, w_093_730, w_093_732, w_093_735, w_093_736, w_093_738, w_093_740, w_093_741, w_093_742, w_093_743, w_093_744, w_093_746, w_093_747, w_093_750, w_093_751, w_093_753, w_093_756, w_093_757, w_093_761, w_093_768, w_093_771, w_093_774, w_093_775, w_093_776, w_093_778, w_093_779, w_093_780, w_093_781, w_093_782, w_093_784, w_093_785, w_093_786, w_093_789, w_093_792, w_093_795, w_093_796, w_093_797, w_093_798, w_093_804, w_093_806, w_093_812, w_093_819, w_093_820, w_093_821, w_093_822, w_093_823, w_093_825, w_093_826, w_093_827, w_093_829, w_093_832, w_093_833, w_093_835, w_093_836, w_093_837, w_093_838, w_093_839, w_093_842, w_093_843, w_093_844, w_093_853, w_093_854, w_093_858, w_093_859, w_093_860, w_093_861, w_093_863, w_093_867, w_093_869, w_093_873, w_093_875, w_093_880, w_093_882, w_093_884, w_093_885, w_093_887, w_093_890, w_093_892, w_093_893, w_093_896, w_093_897, w_093_899, w_093_901, w_093_902, w_093_904, w_093_905, w_093_906, w_093_907, w_093_908, w_093_909, w_093_910, w_093_912, w_093_913, w_093_915, w_093_916, w_093_924, w_093_925, w_093_926, w_093_927, w_093_929, w_093_930, w_093_934, w_093_935, w_093_936, w_093_937, w_093_940, w_093_941, w_093_942, w_093_944, w_093_945, w_093_947, w_093_948, w_093_949, w_093_950, w_093_953, w_093_954, w_093_956, w_093_957, w_093_958, w_093_959, w_093_963, w_093_965, w_093_966, w_093_968, w_093_969, w_093_971, w_093_973, w_093_977, w_093_980, w_093_984, w_093_985, w_093_988, w_093_989, w_093_998, w_093_1001, w_093_1005, w_093_1007, w_093_1008, w_093_1010, w_093_1011, w_093_1012, w_093_1015, w_093_1017, w_093_1018, w_093_1019, w_093_1024, w_093_1025, w_093_1026, w_093_1028, w_093_1031, w_093_1032, w_093_1036, w_093_1040, w_093_1041, w_093_1042, w_093_1044, w_093_1045, w_093_1047, w_093_1049, w_093_1052, w_093_1056, w_093_1058, w_093_1061, w_093_1062, w_093_1065, w_093_1066, w_093_1067, w_093_1069, w_093_1070, w_093_1071, w_093_1072, w_093_1073, w_093_1075, w_093_1078, w_093_1083, w_093_1084, w_093_1089, w_093_1092, w_093_1094, w_093_1095, w_093_1098, w_093_1099, w_093_1101, w_093_1102, w_093_1103, w_093_1104, w_093_1106, w_093_1113, w_093_1114, w_093_1116, w_093_1118, w_093_1121, w_093_1123, w_093_1124, w_093_1130, w_093_1131, w_093_1132, w_093_1135, w_093_1136, w_093_1137, w_093_1138, w_093_1141, w_093_1142, w_093_1143, w_093_1148, w_093_1149, w_093_1150, w_093_1151, w_093_1153, w_093_1154, w_093_1155, w_093_1157, w_093_1158, w_093_1160, w_093_1165, w_093_1166, w_093_1167, w_093_1168, w_093_1169, w_093_1172, w_093_1173, w_093_1175, w_093_1178, w_093_1182, w_093_1183, w_093_1184, w_093_1185, w_093_1193, w_093_1194, w_093_1195, w_093_1196, w_093_1202, w_093_1204, w_093_1206, w_093_1209, w_093_1210, w_093_1212, w_093_1214, w_093_1215, w_093_1216, w_093_1217, w_093_1219, w_093_1221, w_093_1222, w_093_1223, w_093_1224, w_093_1226, w_093_1229, w_093_1231, w_093_1233, w_093_1235, w_093_1236, w_093_1237, w_093_1238, w_093_1239, w_093_1242, w_093_1243, w_093_1245, w_093_1246, w_093_1247, w_093_1251, w_093_1253, w_093_1254, w_093_1255, w_093_1256, w_093_1258, w_093_1260, w_093_1261, w_093_1265, w_093_1266, w_093_1267, w_093_1268, w_093_1277, w_093_1279, w_093_1281, w_093_1284, w_093_1288, w_093_1290, w_093_1296, w_093_1297, w_093_1299, w_093_1304, w_093_1307, w_093_1310, w_093_1311, w_093_1312, w_093_1313, w_093_1316, w_093_1318, w_093_1319, w_093_1320, w_093_1321, w_093_1322, w_093_1325, w_093_1327, w_093_1328, w_093_1329, w_093_1330, w_093_1332, w_093_1333, w_093_1336, w_093_1337, w_093_1338, w_093_1339, w_093_1340, w_093_1343, w_093_1345, w_093_1347, w_093_1348, w_093_1350, w_093_1353, w_093_1355, w_093_1357, w_093_1358, w_093_1359, w_093_1364, w_093_1366, w_093_1368, w_093_1370, w_093_1373, w_093_1374, w_093_1376, w_093_1377, w_093_1378, w_093_1380, w_093_1383, w_093_1384, w_093_1385, w_093_1387, w_093_1390, w_093_1391, w_093_1394, w_093_1395, w_093_1397, w_093_1398, w_093_1400, w_093_1403, w_093_1405, w_093_1406, w_093_1407, w_093_1410, w_093_1411, w_093_1419, w_093_1421, w_093_1422, w_093_1423, w_093_1424, w_093_1427, w_093_1430, w_093_1432, w_093_1433, w_093_1434, w_093_1436, w_093_1437, w_093_1438, w_093_1439, w_093_1441, w_093_1442, w_093_1443, w_093_1445, w_093_1446, w_093_1447, w_093_1448, w_093_1449, w_093_1451, w_093_1452, w_093_1453, w_093_1457, w_093_1461, w_093_1463, w_093_1466, w_093_1469, w_093_1470, w_093_1471, w_093_1472, w_093_1473, w_093_1475, w_093_1478, w_093_1479, w_093_1481, w_093_1484, w_093_1485, w_093_1486, w_093_1488, w_093_1490, w_093_1498, w_093_1499, w_093_1501, w_093_1503, w_093_1504, w_093_1505, w_093_1506, w_093_1507, w_093_1510, w_093_1511, w_093_1512, w_093_1514, w_093_1517, w_093_1519, w_093_1520, w_093_1521, w_093_1522, w_093_1524, w_093_1525, w_093_1526, w_093_1527, w_093_1528, w_093_1532, w_093_1533, w_093_1537, w_093_1538, w_093_1540, w_093_1541, w_093_1542, w_093_1548, w_093_1549, w_093_1551, w_093_1552, w_093_1553, w_093_1554, w_093_1556, w_093_1557, w_093_1561, w_093_1563, w_093_1564, w_093_1566, w_093_1567, w_093_1568, w_093_1574, w_093_1576, w_093_1577, w_093_1579, w_093_1581, w_093_1582, w_093_1583, w_093_1584, w_093_1586, w_093_1587, w_093_1589, w_093_1594, w_093_1596, w_093_1597, w_093_1598, w_093_1600, w_093_1601, w_093_1603, w_093_1604, w_093_1607, w_093_1610, w_093_1611, w_093_1613, w_093_1617, w_093_1619, w_093_1620, w_093_1624, w_093_1626, w_093_1627, w_093_1631, w_093_1633, w_093_1635, w_093_1638, w_093_1639, w_093_1643, w_093_1645, w_093_1646, w_093_1647, w_093_1653, w_093_1655, w_093_1656, w_093_1659, w_093_1660, w_093_1661, w_093_1663, w_093_1673, w_093_1674, w_093_1676, w_093_1678, w_093_1680, w_093_1682, w_093_1683, w_093_1684, w_093_1687, w_093_1688, w_093_1691, w_093_1693, w_093_1694, w_093_1695, w_093_1699, w_093_1701, w_093_1702, w_093_1704, w_093_1705, w_093_1706, w_093_1709, w_093_1710, w_093_1711, w_093_1713, w_093_1715, w_093_1719, w_093_1720, w_093_1722, w_093_1724, w_093_1725, w_093_1726, w_093_1728, w_093_1731, w_093_1733, w_093_1736, w_093_1741, w_093_1742, w_093_1744, w_093_1745, w_093_1746, w_093_1748, w_093_1750, w_093_1752, w_093_1754, w_093_1755, w_093_1756, w_093_1757, w_093_1759, w_093_1760, w_093_1764, w_093_1765, w_093_1766, w_093_1767, w_093_1770, w_093_1771, w_093_1772, w_093_1777, w_093_1781, w_093_1783, w_093_1784, w_093_1787, w_093_1788, w_093_1789, w_093_1790, w_093_1795, w_093_1796, w_093_1798, w_093_1799, w_093_1800, w_093_1801, w_093_1803, w_093_1804, w_093_1806, w_093_1812, w_093_1813, w_093_1815, w_093_1820, w_093_1823, w_093_1825, w_093_1826, w_093_1827, w_093_1829, w_093_1830, w_093_1831, w_093_1832, w_093_1833, w_093_1835, w_093_1838, w_093_1839, w_093_1841, w_093_1842, w_093_1844, w_093_1847, w_093_1848, w_093_1851, w_093_1853, w_093_1854, w_093_1857, w_093_1860, w_093_1862, w_093_1863, w_093_1865, w_093_1866, w_093_1871, w_093_1875, w_093_1877, w_093_1878, w_093_1881, w_093_1882, w_093_1886, w_093_1887, w_093_1888, w_093_1889, w_093_1892, w_093_1894, w_093_1898, w_093_1904, w_093_1905, w_093_1906, w_093_1911, w_093_1912, w_093_1913, w_093_1914, w_093_1916, w_093_1920, w_093_1921, w_093_1922, w_093_1924, w_093_1926, w_093_1927, w_093_1932, w_093_1933, w_093_1935, w_093_1942, w_093_1944, w_093_1945, w_093_1946, w_093_1947, w_093_1948, w_093_1951, w_093_1952, w_093_1953, w_093_1954, w_093_1958, w_093_1961, w_093_1963, w_093_1965, w_093_1966, w_093_1968, w_093_1969, w_093_1972, w_093_1973, w_093_1974, w_093_1978, w_093_1980, w_093_1981, w_093_1982, w_093_1985, w_093_1986, w_093_1987, w_093_1988, w_093_1990, w_093_1991, w_093_1994, w_093_1996, w_093_1999, w_093_2000, w_093_2001, w_093_2002, w_093_2003, w_093_2006, w_093_2007, w_093_2008, w_093_2014, w_093_2017, w_093_2018, w_093_2019, w_093_2021, w_093_2025, w_093_2028, w_093_2029, w_093_2032, w_093_2035, w_093_2036, w_093_2038, w_093_2039, w_093_2040, w_093_2043, w_093_2045, w_093_2046, w_093_2048, w_093_2049, w_093_2051, w_093_2052, w_093_2055, w_093_2056, w_093_2058, w_093_2062, w_093_2063, w_093_2074, w_093_2077, w_093_2079, w_093_2080, w_093_2081, w_093_2089, w_093_2090, w_093_2091, w_093_2093, w_093_2094, w_093_2096, w_093_2098, w_093_2099, w_093_2100, w_093_2101, w_093_2104, w_093_2107, w_093_2108, w_093_2109, w_093_2110, w_093_2111, w_093_2113, w_093_2115, w_093_2119, w_093_2121, w_093_2127, w_093_2128, w_093_2131, w_093_2134, w_093_2139, w_093_2140, w_093_2141, w_093_2142, w_093_2145, w_093_2146, w_093_2147, w_093_2148, w_093_2150, w_093_2152, w_093_2153, w_093_2154, w_093_2157, w_093_2160, w_093_2161, w_093_2163, w_093_2165, w_093_2167, w_093_2168, w_093_2169, w_093_2172, w_093_2174, w_093_2175, w_093_2176, w_093_2178, w_093_2180, w_093_2181, w_093_2182, w_093_2184, w_093_2185, w_093_2187, w_093_2188, w_093_2190, w_093_2191, w_093_2194, w_093_2196, w_093_2197, w_093_2198, w_093_2200, w_093_2201, w_093_2202, w_093_2203, w_093_2204, w_093_2206, w_093_2207, w_093_2209, w_093_2210, w_093_2212, w_093_2213, w_093_2215, w_093_2217, w_093_2218, w_093_2219, w_093_2220, w_093_2223, w_093_2228, w_093_2230, w_093_2232, w_093_2234, w_093_2236, w_093_2237, w_093_2238, w_093_2241, w_093_2242, w_093_2244, w_093_2245, w_093_2248, w_093_2249, w_093_2250, w_093_2251, w_093_2252, w_093_2253, w_093_2254, w_093_2257, w_093_2259, w_093_2264, w_093_2265, w_093_2266, w_093_2267, w_093_2268, w_093_2269, w_093_2275, w_093_2278, w_093_2281, w_093_2283, w_093_2284, w_093_2285, w_093_2287, w_093_2288, w_093_2289, w_093_2292, w_093_2295, w_093_2297, w_093_2299, w_093_2300, w_093_2302, w_093_2303, w_093_2305, w_093_2306, w_093_2308;
  wire w_094_000, w_094_002, w_094_003, w_094_004, w_094_005, w_094_006, w_094_008, w_094_009, w_094_011, w_094_012, w_094_014, w_094_017, w_094_018, w_094_019, w_094_023, w_094_024, w_094_025, w_094_026, w_094_027, w_094_028, w_094_030, w_094_032, w_094_033, w_094_034, w_094_037, w_094_040, w_094_041, w_094_042, w_094_043, w_094_045, w_094_046, w_094_050, w_094_051, w_094_054, w_094_055, w_094_056, w_094_058, w_094_059, w_094_060, w_094_064, w_094_065, w_094_066, w_094_067, w_094_068, w_094_069, w_094_071, w_094_072, w_094_075, w_094_076, w_094_077, w_094_078, w_094_080, w_094_082, w_094_084, w_094_086, w_094_088, w_094_091, w_094_093, w_094_094, w_094_097, w_094_099, w_094_100, w_094_101, w_094_102, w_094_103, w_094_104, w_094_106, w_094_108, w_094_109, w_094_110, w_094_111, w_094_113, w_094_116, w_094_117, w_094_119, w_094_120, w_094_121, w_094_123, w_094_124, w_094_126, w_094_128, w_094_131, w_094_132, w_094_133, w_094_134, w_094_141, w_094_146, w_094_147, w_094_148, w_094_150, w_094_151, w_094_155, w_094_157, w_094_158, w_094_160, w_094_161, w_094_162, w_094_163, w_094_166, w_094_167, w_094_168, w_094_169, w_094_170, w_094_173, w_094_174, w_094_177, w_094_178, w_094_179, w_094_183, w_094_186, w_094_192, w_094_193, w_094_201, w_094_203, w_094_204, w_094_209, w_094_211, w_094_212, w_094_215, w_094_216, w_094_217, w_094_218, w_094_219, w_094_220, w_094_221, w_094_222, w_094_223, w_094_224, w_094_225, w_094_228, w_094_231, w_094_232, w_094_234, w_094_235, w_094_237, w_094_239, w_094_240, w_094_243, w_094_244, w_094_245, w_094_246, w_094_248, w_094_249, w_094_251, w_094_252, w_094_253, w_094_256, w_094_257, w_094_262, w_094_263, w_094_265, w_094_266, w_094_267, w_094_269, w_094_270, w_094_272, w_094_274, w_094_276, w_094_277, w_094_278, w_094_280, w_094_285, w_094_289, w_094_290, w_094_291, w_094_292, w_094_293, w_094_294, w_094_297, w_094_299, w_094_303, w_094_309, w_094_310, w_094_313, w_094_314, w_094_315, w_094_317, w_094_319, w_094_320, w_094_324, w_094_326, w_094_327, w_094_328, w_094_329, w_094_330, w_094_332, w_094_333, w_094_335, w_094_336, w_094_339, w_094_340, w_094_342, w_094_343, w_094_344, w_094_350, w_094_351, w_094_352, w_094_354, w_094_355, w_094_359, w_094_361, w_094_362, w_094_363, w_094_364, w_094_368, w_094_372, w_094_373, w_094_376, w_094_377, w_094_381, w_094_383, w_094_384, w_094_385, w_094_386, w_094_388, w_094_390, w_094_392, w_094_393, w_094_395, w_094_404, w_094_405, w_094_406, w_094_407, w_094_408, w_094_412, w_094_413, w_094_414, w_094_415, w_094_416, w_094_417, w_094_420, w_094_421, w_094_422, w_094_424, w_094_426, w_094_428, w_094_429, w_094_433, w_094_436, w_094_437, w_094_438, w_094_439, w_094_442, w_094_448, w_094_450, w_094_451, w_094_452, w_094_453, w_094_454, w_094_455, w_094_456, w_094_457, w_094_458, w_094_460, w_094_461, w_094_462, w_094_464, w_094_466, w_094_467, w_094_469, w_094_471, w_094_474, w_094_476, w_094_481, w_094_482, w_094_485, w_094_486, w_094_487, w_094_489, w_094_490, w_094_491, w_094_492, w_094_493, w_094_496, w_094_497, w_094_498, w_094_499, w_094_500, w_094_501, w_094_502, w_094_504, w_094_506, w_094_508, w_094_517, w_094_520, w_094_523, w_094_525, w_094_529, w_094_531, w_094_533, w_094_535, w_094_539, w_094_540, w_094_542, w_094_543, w_094_544, w_094_546, w_094_547, w_094_550, w_094_551, w_094_552, w_094_555, w_094_557, w_094_558, w_094_562, w_094_565, w_094_568, w_094_571, w_094_572, w_094_573, w_094_575, w_094_578, w_094_580, w_094_581, w_094_583, w_094_584, w_094_585, w_094_587, w_094_588, w_094_592, w_094_593, w_094_596, w_094_598, w_094_599, w_094_600, w_094_602, w_094_603, w_094_605, w_094_607, w_094_608, w_094_610, w_094_613, w_094_615, w_094_616, w_094_618, w_094_619, w_094_621, w_094_626, w_094_629, w_094_630, w_094_633, w_094_636, w_094_639, w_094_640, w_094_641, w_094_644, w_094_649, w_094_651, w_094_652, w_094_656, w_094_658, w_094_659, w_094_661, w_094_663, w_094_664, w_094_666, w_094_674, w_094_675, w_094_677, w_094_683, w_094_686, w_094_687, w_094_690, w_094_694, w_094_699, w_094_701, w_094_702, w_094_706, w_094_710, w_094_712, w_094_719, w_094_724, w_094_725, w_094_726, w_094_727, w_094_730, w_094_732, w_094_736, w_094_737, w_094_739, w_094_740, w_094_741, w_094_742, w_094_743, w_094_744, w_094_745, w_094_747, w_094_749, w_094_751, w_094_752, w_094_753, w_094_754, w_094_756, w_094_758, w_094_759, w_094_774, w_094_775, w_094_776, w_094_779, w_094_782, w_094_784, w_094_794, w_094_797, w_094_799, w_094_805, w_094_808, w_094_809, w_094_811, w_094_818, w_094_823, w_094_826, w_094_836, w_094_840, w_094_851, w_094_867, w_094_870, w_094_873, w_094_876, w_094_877, w_094_879, w_094_880, w_094_882, w_094_883, w_094_886, w_094_888, w_094_892, w_094_897, w_094_899, w_094_903, w_094_905, w_094_906, w_094_908, w_094_913, w_094_914, w_094_917, w_094_918, w_094_928, w_094_936, w_094_944, w_094_947, w_094_949, w_094_951, w_094_952, w_094_962, w_094_969, w_094_970, w_094_975, w_094_976, w_094_980, w_094_985, w_094_986, w_094_995, w_094_1006, w_094_1009, w_094_1010, w_094_1012, w_094_1019, w_094_1027, w_094_1032, w_094_1034, w_094_1038, w_094_1044, w_094_1045, w_094_1046, w_094_1047, w_094_1050, w_094_1053, w_094_1054, w_094_1057, w_094_1058, w_094_1059, w_094_1061, w_094_1064, w_094_1067, w_094_1068, w_094_1070, w_094_1083, w_094_1084, w_094_1092, w_094_1101, w_094_1102, w_094_1107, w_094_1109, w_094_1111, w_094_1118, w_094_1120, w_094_1121, w_094_1123, w_094_1126, w_094_1129, w_094_1132, w_094_1136, w_094_1138, w_094_1144, w_094_1145, w_094_1146, w_094_1149, w_094_1151, w_094_1152, w_094_1155, w_094_1156, w_094_1157, w_094_1162, w_094_1163, w_094_1170, w_094_1177, w_094_1182, w_094_1184, w_094_1192, w_094_1194, w_094_1197, w_094_1203, w_094_1207, w_094_1208, w_094_1212, w_094_1221, w_094_1224, w_094_1230, w_094_1232, w_094_1237, w_094_1238, w_094_1239, w_094_1248, w_094_1252, w_094_1254, w_094_1271, w_094_1273, w_094_1275, w_094_1276, w_094_1283, w_094_1284, w_094_1288, w_094_1290, w_094_1293, w_094_1294, w_094_1296, w_094_1300, w_094_1301, w_094_1322, w_094_1325, w_094_1327, w_094_1330, w_094_1332, w_094_1336, w_094_1338, w_094_1341, w_094_1346, w_094_1347, w_094_1350, w_094_1354, w_094_1356, w_094_1357, w_094_1359, w_094_1362, w_094_1368, w_094_1372, w_094_1374, w_094_1376, w_094_1381, w_094_1382, w_094_1390, w_094_1393, w_094_1396, w_094_1403, w_094_1410, w_094_1411, w_094_1413, w_094_1414, w_094_1415, w_094_1416, w_094_1419, w_094_1421, w_094_1423, w_094_1430, w_094_1435, w_094_1438, w_094_1440, w_094_1445, w_094_1452, w_094_1453, w_094_1456, w_094_1459, w_094_1461, w_094_1464, w_094_1466, w_094_1467, w_094_1470, w_094_1471, w_094_1473, w_094_1474, w_094_1475, w_094_1476, w_094_1477, w_094_1483, w_094_1486, w_094_1490, w_094_1498, w_094_1500, w_094_1504, w_094_1509, w_094_1510, w_094_1512, w_094_1521, w_094_1522, w_094_1523, w_094_1525, w_094_1528, w_094_1530, w_094_1531, w_094_1532, w_094_1534, w_094_1535, w_094_1539, w_094_1540, w_094_1547, w_094_1552, w_094_1553, w_094_1556, w_094_1558, w_094_1560, w_094_1561, w_094_1562, w_094_1563, w_094_1566, w_094_1567, w_094_1572, w_094_1573, w_094_1574, w_094_1575, w_094_1579, w_094_1580, w_094_1582, w_094_1583, w_094_1585, w_094_1587, w_094_1588, w_094_1592, w_094_1607, w_094_1616, w_094_1617, w_094_1626, w_094_1629, w_094_1632, w_094_1637, w_094_1642, w_094_1648, w_094_1649, w_094_1651, w_094_1654, w_094_1660, w_094_1664, w_094_1671, w_094_1672, w_094_1675, w_094_1682, w_094_1684, w_094_1686, w_094_1690, w_094_1692, w_094_1698, w_094_1703, w_094_1705, w_094_1706, w_094_1707, w_094_1713, w_094_1714, w_094_1718, w_094_1721, w_094_1723, w_094_1728, w_094_1729, w_094_1731, w_094_1732, w_094_1736, w_094_1739, w_094_1742, w_094_1747, w_094_1748, w_094_1752, w_094_1753, w_094_1757, w_094_1758, w_094_1759, w_094_1761, w_094_1762, w_094_1765, w_094_1766, w_094_1767, w_094_1769, w_094_1776, w_094_1778, w_094_1779, w_094_1780, w_094_1792, w_094_1793, w_094_1795, w_094_1797, w_094_1799, w_094_1801, w_094_1802, w_094_1803, w_094_1806, w_094_1813, w_094_1814, w_094_1816, w_094_1821, w_094_1822, w_094_1824, w_094_1825, w_094_1826, w_094_1827, w_094_1830, w_094_1831, w_094_1838, w_094_1843, w_094_1844, w_094_1847, w_094_1859, w_094_1870, w_094_1873, w_094_1876, w_094_1878, w_094_1880, w_094_1881, w_094_1883, w_094_1884, w_094_1889, w_094_1894, w_094_1896, w_094_1900, w_094_1902, w_094_1905, w_094_1907, w_094_1915, w_094_1920, w_094_1922, w_094_1926, w_094_1930, w_094_1931, w_094_1934, w_094_1937, w_094_1940, w_094_1944, w_094_1947, w_094_1949, w_094_1953, w_094_1956, w_094_1960, w_094_1962, w_094_1968, w_094_1969, w_094_1970, w_094_1981, w_094_1982, w_094_1984, w_094_1986, w_094_1987, w_094_1989, w_094_1994, w_094_1998, w_094_2000, w_094_2002, w_094_2012, w_094_2013, w_094_2015, w_094_2018, w_094_2019, w_094_2024, w_094_2026, w_094_2029, w_094_2033, w_094_2036, w_094_2037, w_094_2043, w_094_2045, w_094_2049, w_094_2054, w_094_2060, w_094_2073, w_094_2079, w_094_2083, w_094_2087, w_094_2088, w_094_2090, w_094_2096, w_094_2100, w_094_2104, w_094_2105, w_094_2106, w_094_2112, w_094_2116, w_094_2119, w_094_2121, w_094_2131, w_094_2133, w_094_2140, w_094_2142, w_094_2145, w_094_2151, w_094_2153, w_094_2154, w_094_2155, w_094_2156, w_094_2158, w_094_2168, w_094_2174, w_094_2178, w_094_2186, w_094_2190, w_094_2193, w_094_2194, w_094_2196, w_094_2201, w_094_2212, w_094_2221, w_094_2222, w_094_2224, w_094_2225, w_094_2227, w_094_2229, w_094_2230, w_094_2233, w_094_2235, w_094_2242, w_094_2248, w_094_2250, w_094_2252, w_094_2253, w_094_2254, w_094_2256, w_094_2257, w_094_2262, w_094_2267, w_094_2271, w_094_2273, w_094_2277, w_094_2281, w_094_2284, w_094_2289, w_094_2298, w_094_2299, w_094_2300, w_094_2305, w_094_2306, w_094_2308, w_094_2316, w_094_2323, w_094_2325, w_094_2326, w_094_2327, w_094_2335, w_094_2339, w_094_2340, w_094_2344, w_094_2346, w_094_2348, w_094_2350, w_094_2351, w_094_2353, w_094_2355, w_094_2357, w_094_2359, w_094_2361, w_094_2363, w_094_2371, w_094_2374, w_094_2376, w_094_2378, w_094_2379, w_094_2381, w_094_2395, w_094_2396, w_094_2403, w_094_2404, w_094_2405, w_094_2406, w_094_2412, w_094_2413, w_094_2416, w_094_2424, w_094_2425, w_094_2428, w_094_2437, w_094_2442, w_094_2449, w_094_2456, w_094_2457, w_094_2458, w_094_2462, w_094_2465, w_094_2468, w_094_2471, w_094_2475, w_094_2477, w_094_2480, w_094_2485, w_094_2486, w_094_2488, w_094_2497, w_094_2509, w_094_2512, w_094_2515, w_094_2517, w_094_2522, w_094_2526, w_094_2528, w_094_2533, w_094_2537, w_094_2539, w_094_2545, w_094_2546, w_094_2559, w_094_2563, w_094_2568, w_094_2577, w_094_2582, w_094_2585, w_094_2586, w_094_2594, w_094_2600, w_094_2601, w_094_2602, w_094_2604, w_094_2605, w_094_2607, w_094_2615, w_094_2619, w_094_2620, w_094_2634, w_094_2641, w_094_2644, w_094_2645, w_094_2646, w_094_2648, w_094_2651, w_094_2654, w_094_2659, w_094_2666, w_094_2667, w_094_2669, w_094_2673, w_094_2679, w_094_2680, w_094_2682, w_094_2685, w_094_2688, w_094_2692, w_094_2693, w_094_2697, w_094_2698, w_094_2700, w_094_2706, w_094_2711, w_094_2714, w_094_2716, w_094_2719, w_094_2723, w_094_2729, w_094_2731, w_094_2733, w_094_2734, w_094_2735, w_094_2737, w_094_2738, w_094_2740, w_094_2741, w_094_2742, w_094_2743, w_094_2750, w_094_2761, w_094_2767, w_094_2769, w_094_2770, w_094_2771, w_094_2772, w_094_2774, w_094_2778, w_094_2779, w_094_2780, w_094_2786, w_094_2787, w_094_2789, w_094_2791, w_094_2794, w_094_2796, w_094_2797, w_094_2800, w_094_2803, w_094_2804, w_094_2808, w_094_2810, w_094_2813, w_094_2818, w_094_2824, w_094_2825, w_094_2829, w_094_2833, w_094_2835, w_094_2842, w_094_2843, w_094_2846, w_094_2856, w_094_2859, w_094_2860, w_094_2869, w_094_2872, w_094_2873, w_094_2875, w_094_2876, w_094_2878, w_094_2883, w_094_2884, w_094_2885, w_094_2888, w_094_2889, w_094_2895, w_094_2896, w_094_2898, w_094_2901, w_094_2902, w_094_2905, w_094_2909, w_094_2910, w_094_2912, w_094_2913, w_094_2916, w_094_2919, w_094_2928, w_094_2931, w_094_2937, w_094_2945, w_094_2952, w_094_2953, w_094_2954, w_094_2955, w_094_2960, w_094_2964, w_094_2968, w_094_2975, w_094_2977, w_094_2979, w_094_2980, w_094_2985, w_094_2987, w_094_2995, w_094_2996, w_094_3006, w_094_3007, w_094_3008, w_094_3011, w_094_3017, w_094_3019, w_094_3021, w_094_3027, w_094_3031, w_094_3034, w_094_3035, w_094_3050, w_094_3051, w_094_3055, w_094_3057, w_094_3058, w_094_3062, w_094_3065, w_094_3068, w_094_3072, w_094_3075, w_094_3076, w_094_3077, w_094_3078, w_094_3079, w_094_3081, w_094_3090, w_094_3095, w_094_3097, w_094_3098, w_094_3099, w_094_3100, w_094_3102, w_094_3105, w_094_3106, w_094_3110, w_094_3111, w_094_3113, w_094_3119, w_094_3126, w_094_3127, w_094_3130, w_094_3131, w_094_3133, w_094_3134, w_094_3135, w_094_3138, w_094_3140, w_094_3141, w_094_3142, w_094_3144, w_094_3152, w_094_3153, w_094_3154, w_094_3157, w_094_3159, w_094_3166, w_094_3167, w_094_3168, w_094_3172, w_094_3180, w_094_3185, w_094_3187, w_094_3189, w_094_3198, w_094_3201, w_094_3203, w_094_3206, w_094_3207, w_094_3208, w_094_3211, w_094_3212, w_094_3213, w_094_3214, w_094_3219, w_094_3227, w_094_3228, w_094_3230, w_094_3238, w_094_3243, w_094_3244, w_094_3245, w_094_3246, w_094_3252, w_094_3253, w_094_3254, w_094_3259, w_094_3260, w_094_3264, w_094_3270, w_094_3274, w_094_3281, w_094_3282, w_094_3288, w_094_3291, w_094_3292, w_094_3294, w_094_3295, w_094_3299, w_094_3303, w_094_3306, w_094_3307, w_094_3310, w_094_3311, w_094_3312, w_094_3313, w_094_3316, w_094_3319, w_094_3320, w_094_3327, w_094_3336, w_094_3337, w_094_3341, w_094_3343, w_094_3344, w_094_3347, w_094_3357, w_094_3364, w_094_3371, w_094_3376, w_094_3379, w_094_3385, w_094_3386, w_094_3389, w_094_3394, w_094_3397, w_094_3398, w_094_3402, w_094_3411, w_094_3414, w_094_3418, w_094_3420, w_094_3422, w_094_3423, w_094_3425, w_094_3427, w_094_3428, w_094_3429, w_094_3438, w_094_3452, w_094_3453, w_094_3455, w_094_3458, w_094_3464, w_094_3470, w_094_3472, w_094_3476, w_094_3477, w_094_3480, w_094_3486, w_094_3487, w_094_3490, w_094_3491, w_094_3492, w_094_3505, w_094_3508, w_094_3509, w_094_3512, w_094_3514, w_094_3516, w_094_3519, w_094_3528, w_094_3529, w_094_3532, w_094_3534, w_094_3535, w_094_3543, w_094_3545, w_094_3547, w_094_3554, w_094_3559, w_094_3563, w_094_3574, w_094_3577, w_094_3582, w_094_3583, w_094_3587, w_094_3588, w_094_3589, w_094_3593, w_094_3598, w_094_3602, w_094_3607, w_094_3609, w_094_3616, w_094_3621, w_094_3623, w_094_3624, w_094_3625, w_094_3630, w_094_3632, w_094_3635, w_094_3640, w_094_3642, w_094_3649, w_094_3654, w_094_3655, w_094_3658, w_094_3665, w_094_3666, w_094_3670, w_094_3671, w_094_3672, w_094_3676, w_094_3679, w_094_3682, w_094_3687, w_094_3689, w_094_3691, w_094_3692, w_094_3693, w_094_3695, w_094_3698, w_094_3699, w_094_3702, w_094_3704, w_094_3707, w_094_3710, w_094_3712, w_094_3726, w_094_3739, w_094_3740, w_094_3743, w_094_3745, w_094_3746, w_094_3747, w_094_3752, w_094_3757, w_094_3761, w_094_3768, w_094_3769, w_094_3772, w_094_3778, w_094_3781, w_094_3784, w_094_3790, w_094_3791, w_094_3794, w_094_3796, w_094_3799, w_094_3800, w_094_3802, w_094_3805, w_094_3806, w_094_3807, w_094_3808, w_094_3809, w_094_3811, w_094_3819, w_094_3824, w_094_3827, w_094_3828, w_094_3829, w_094_3837, w_094_3839, w_094_3841, w_094_3842, w_094_3845, w_094_3850, w_094_3852, w_094_3854, w_094_3855, w_094_3857, w_094_3860, w_094_3861, w_094_3862, w_094_3863, w_094_3868, w_094_3871, w_094_3876, w_094_3880, w_094_3882, w_094_3886, w_094_3892, w_094_3894, w_094_3897, w_094_3901, w_094_3907, w_094_3912, w_094_3918, w_094_3920, w_094_3921, w_094_3925, w_094_3927, w_094_3928, w_094_3929, w_094_3932, w_094_3938, w_094_3946, w_094_3947, w_094_3948, w_094_3953, w_094_3957, w_094_3965, w_094_3969, w_094_3972, w_094_3973, w_094_3974, w_094_3975, w_094_3978, w_094_3980, w_094_3981, w_094_3985, w_094_3986, w_094_3989, w_094_3991, w_094_3992, w_094_3993, w_094_3997, w_094_3998, w_094_4004, w_094_4008, w_094_4009, w_094_4010, w_094_4011, w_094_4015, w_094_4017, w_094_4018, w_094_4019, w_094_4020, w_094_4028, w_094_4030, w_094_4031, w_094_4032, w_094_4033, w_094_4037, w_094_4054, w_094_4057, w_094_4060, w_094_4062, w_094_4063, w_094_4065, w_094_4073, w_094_4077, w_094_4082, w_094_4085, w_094_4086, w_094_4094, w_094_4115, w_094_4116, w_094_4119, w_094_4120, w_094_4122, w_094_4124, w_094_4127, w_094_4129, w_094_4130, w_094_4135, w_094_4137, w_094_4143, w_094_4144, w_094_4160, w_094_4161, w_094_4164, w_094_4167, w_094_4168, w_094_4175, w_094_4177, w_094_4185, w_094_4191, w_094_4192, w_094_4197, w_094_4198, w_094_4204, w_094_4210, w_094_4212, w_094_4217, w_094_4219, w_094_4226, w_094_4228, w_094_4231, w_094_4234, w_094_4236, w_094_4238, w_094_4239, w_094_4241, w_094_4242, w_094_4243, w_094_4244, w_094_4245, w_094_4246, w_094_4247, w_094_4248, w_094_4249, w_094_4250;
  wire w_095_000, w_095_003, w_095_004, w_095_005, w_095_007, w_095_010, w_095_011, w_095_012, w_095_014, w_095_016, w_095_017, w_095_019, w_095_020, w_095_023, w_095_024, w_095_028, w_095_030, w_095_031, w_095_034, w_095_035, w_095_038, w_095_040, w_095_041, w_095_042, w_095_045, w_095_046, w_095_047, w_095_048, w_095_051, w_095_054, w_095_055, w_095_056, w_095_057, w_095_060, w_095_064, w_095_065, w_095_066, w_095_067, w_095_072, w_095_073, w_095_077, w_095_078, w_095_080, w_095_082, w_095_085, w_095_086, w_095_087, w_095_088, w_095_091, w_095_094, w_095_095, w_095_099, w_095_100, w_095_101, w_095_102, w_095_109, w_095_112, w_095_114, w_095_115, w_095_117, w_095_119, w_095_120, w_095_121, w_095_123, w_095_126, w_095_127, w_095_128, w_095_130, w_095_131, w_095_132, w_095_133, w_095_134, w_095_139, w_095_140, w_095_141, w_095_142, w_095_144, w_095_145, w_095_146, w_095_148, w_095_149, w_095_156, w_095_157, w_095_161, w_095_164, w_095_165, w_095_166, w_095_168, w_095_170, w_095_171, w_095_175, w_095_178, w_095_179, w_095_181, w_095_182, w_095_183, w_095_186, w_095_187, w_095_189, w_095_190, w_095_193, w_095_195, w_095_197, w_095_198, w_095_199, w_095_202, w_095_205, w_095_206, w_095_208, w_095_211, w_095_214, w_095_217, w_095_218, w_095_220, w_095_221, w_095_223, w_095_225, w_095_226, w_095_232, w_095_233, w_095_236, w_095_237, w_095_238, w_095_239, w_095_241, w_095_243, w_095_244, w_095_245, w_095_246, w_095_248, w_095_249, w_095_251, w_095_252, w_095_253, w_095_258, w_095_259, w_095_260, w_095_261, w_095_262, w_095_263, w_095_266, w_095_267, w_095_268, w_095_271, w_095_272, w_095_274, w_095_275, w_095_278, w_095_281, w_095_284, w_095_288, w_095_291, w_095_294, w_095_296, w_095_298, w_095_300, w_095_305, w_095_306, w_095_307, w_095_308, w_095_309, w_095_312, w_095_313, w_095_314, w_095_315, w_095_318, w_095_319, w_095_322, w_095_323, w_095_324, w_095_325, w_095_326, w_095_328, w_095_329, w_095_330, w_095_336, w_095_337, w_095_338, w_095_341, w_095_343, w_095_344, w_095_347, w_095_348, w_095_349, w_095_351, w_095_352, w_095_355, w_095_357, w_095_358, w_095_359, w_095_361, w_095_363, w_095_364, w_095_366, w_095_367, w_095_368, w_095_370, w_095_372, w_095_373, w_095_374, w_095_375, w_095_376, w_095_378, w_095_379, w_095_383, w_095_386, w_095_389, w_095_391, w_095_392, w_095_395, w_095_397, w_095_402, w_095_406, w_095_410, w_095_411, w_095_412, w_095_414, w_095_416, w_095_418, w_095_419, w_095_422, w_095_425, w_095_429, w_095_433, w_095_434, w_095_436, w_095_437, w_095_438, w_095_439, w_095_440, w_095_441, w_095_442, w_095_443, w_095_444, w_095_445, w_095_446, w_095_447, w_095_451, w_095_453, w_095_454, w_095_455, w_095_458, w_095_459, w_095_461, w_095_462, w_095_463, w_095_464, w_095_466, w_095_467, w_095_468, w_095_469, w_095_472, w_095_473, w_095_475, w_095_477, w_095_478, w_095_479, w_095_484, w_095_489, w_095_493, w_095_498, w_095_502, w_095_505, w_095_506, w_095_508, w_095_514, w_095_516, w_095_517, w_095_518, w_095_519, w_095_521, w_095_522, w_095_524, w_095_526, w_095_527, w_095_529, w_095_530, w_095_532, w_095_535, w_095_536, w_095_537, w_095_543, w_095_548, w_095_551, w_095_552, w_095_553, w_095_555, w_095_556, w_095_559, w_095_561, w_095_562, w_095_563, w_095_566, w_095_567, w_095_569, w_095_570, w_095_572, w_095_573, w_095_575, w_095_576, w_095_578, w_095_580, w_095_583, w_095_585, w_095_589, w_095_595, w_095_598, w_095_599, w_095_602, w_095_604, w_095_605, w_095_607, w_095_608, w_095_609, w_095_612, w_095_613, w_095_614, w_095_616, w_095_618, w_095_623, w_095_624, w_095_627, w_095_630, w_095_631, w_095_633, w_095_636, w_095_637, w_095_638, w_095_639, w_095_644, w_095_647, w_095_651, w_095_652, w_095_655, w_095_656, w_095_659, w_095_660, w_095_663, w_095_664, w_095_665, w_095_666, w_095_669, w_095_670, w_095_672, w_095_674, w_095_675, w_095_678, w_095_682, w_095_683, w_095_684, w_095_687, w_095_688, w_095_691, w_095_692, w_095_693, w_095_694, w_095_697, w_095_701, w_095_705, w_095_707, w_095_711, w_095_713, w_095_714, w_095_716, w_095_717, w_095_718, w_095_719, w_095_720, w_095_722, w_095_725, w_095_728, w_095_732, w_095_733, w_095_735, w_095_739, w_095_740, w_095_741, w_095_743, w_095_744, w_095_746, w_095_747, w_095_748, w_095_752, w_095_753, w_095_754, w_095_757, w_095_758, w_095_760, w_095_762, w_095_764, w_095_765, w_095_766, w_095_768, w_095_769, w_095_772, w_095_774, w_095_776, w_095_779, w_095_780, w_095_782, w_095_787, w_095_788, w_095_791, w_095_792, w_095_793, w_095_794, w_095_796, w_095_799, w_095_800, w_095_805, w_095_806, w_095_807, w_095_808, w_095_809, w_095_810, w_095_811, w_095_815, w_095_817, w_095_820, w_095_822, w_095_823, w_095_826, w_095_832, w_095_833, w_095_836, w_095_837, w_095_838, w_095_840, w_095_843, w_095_844, w_095_845, w_095_847, w_095_848, w_095_849, w_095_851, w_095_853, w_095_854, w_095_860, w_095_863, w_095_864, w_095_865, w_095_866, w_095_867, w_095_869, w_095_870, w_095_871, w_095_872, w_095_873, w_095_875, w_095_879, w_095_885, w_095_886, w_095_887, w_095_890, w_095_894, w_095_897, w_095_901, w_095_906, w_095_907, w_095_911, w_095_913, w_095_915, w_095_916, w_095_923, w_095_925, w_095_926, w_095_928, w_095_930, w_095_931, w_095_933, w_095_935, w_095_937, w_095_938, w_095_939, w_095_940, w_095_941, w_095_946, w_095_947, w_095_961, w_095_968, w_095_970, w_095_973, w_095_974, w_095_975, w_095_976, w_095_984, w_095_989, w_095_992, w_095_996, w_095_998, w_095_999, w_095_1001, w_095_1006, w_095_1011, w_095_1012, w_095_1018, w_095_1021, w_095_1022, w_095_1025, w_095_1026, w_095_1034, w_095_1040, w_095_1046, w_095_1048, w_095_1055, w_095_1058, w_095_1060, w_095_1071, w_095_1072, w_095_1075, w_095_1078, w_095_1087, w_095_1088, w_095_1092, w_095_1095, w_095_1096, w_095_1100, w_095_1105, w_095_1110, w_095_1112, w_095_1116, w_095_1119, w_095_1123, w_095_1127, w_095_1132, w_095_1140, w_095_1145, w_095_1148, w_095_1151, w_095_1159, w_095_1160, w_095_1161, w_095_1168, w_095_1173, w_095_1174, w_095_1178, w_095_1188, w_095_1190, w_095_1191, w_095_1202, w_095_1205, w_095_1207, w_095_1210, w_095_1211, w_095_1212, w_095_1214, w_095_1215, w_095_1221, w_095_1222, w_095_1223, w_095_1225, w_095_1227, w_095_1228, w_095_1229, w_095_1230, w_095_1246, w_095_1250, w_095_1253, w_095_1264, w_095_1265, w_095_1271, w_095_1272, w_095_1276, w_095_1284, w_095_1290, w_095_1292, w_095_1294, w_095_1300, w_095_1302, w_095_1306, w_095_1311, w_095_1312, w_095_1314, w_095_1315, w_095_1319, w_095_1321, w_095_1325, w_095_1328, w_095_1329, w_095_1332, w_095_1338, w_095_1340, w_095_1341, w_095_1357, w_095_1362, w_095_1366, w_095_1368, w_095_1369, w_095_1373, w_095_1376, w_095_1380, w_095_1381, w_095_1384, w_095_1389, w_095_1390, w_095_1394, w_095_1399, w_095_1402, w_095_1404, w_095_1412, w_095_1415, w_095_1416, w_095_1417, w_095_1419, w_095_1420, w_095_1424, w_095_1428, w_095_1429, w_095_1434, w_095_1442, w_095_1443, w_095_1450, w_095_1453, w_095_1454, w_095_1455, w_095_1457, w_095_1462, w_095_1463, w_095_1466, w_095_1467, w_095_1469, w_095_1474, w_095_1475, w_095_1477, w_095_1490, w_095_1495, w_095_1497, w_095_1503, w_095_1504, w_095_1507, w_095_1508, w_095_1509, w_095_1516, w_095_1518, w_095_1521, w_095_1522, w_095_1523, w_095_1525, w_095_1527, w_095_1545, w_095_1546, w_095_1547, w_095_1551, w_095_1554, w_095_1557, w_095_1558, w_095_1559, w_095_1561, w_095_1562, w_095_1566, w_095_1569, w_095_1570, w_095_1578, w_095_1583, w_095_1587, w_095_1592, w_095_1597, w_095_1598, w_095_1603, w_095_1606, w_095_1610, w_095_1613, w_095_1614, w_095_1618, w_095_1619, w_095_1622, w_095_1627, w_095_1629, w_095_1635, w_095_1636, w_095_1642, w_095_1643, w_095_1646, w_095_1653, w_095_1654, w_095_1656, w_095_1670, w_095_1676, w_095_1677, w_095_1682, w_095_1687, w_095_1695, w_095_1706, w_095_1707, w_095_1709, w_095_1713, w_095_1717, w_095_1718, w_095_1724, w_095_1727, w_095_1731, w_095_1736, w_095_1740, w_095_1741, w_095_1743, w_095_1745, w_095_1746, w_095_1754, w_095_1756, w_095_1759, w_095_1760, w_095_1762, w_095_1768, w_095_1769, w_095_1771, w_095_1773, w_095_1774, w_095_1775, w_095_1780, w_095_1782, w_095_1788, w_095_1798, w_095_1803, w_095_1807, w_095_1809, w_095_1810, w_095_1812, w_095_1815, w_095_1818, w_095_1819, w_095_1821, w_095_1832, w_095_1835, w_095_1838, w_095_1841, w_095_1843, w_095_1848, w_095_1852, w_095_1858, w_095_1866, w_095_1871, w_095_1873, w_095_1874, w_095_1876, w_095_1878, w_095_1879, w_095_1888, w_095_1890, w_095_1893, w_095_1894, w_095_1900, w_095_1906, w_095_1908, w_095_1911, w_095_1912, w_095_1913, w_095_1923, w_095_1924, w_095_1926, w_095_1928, w_095_1940, w_095_1941, w_095_1944, w_095_1949, w_095_1950, w_095_1953, w_095_1961, w_095_1962, w_095_1967, w_095_1971, w_095_1972, w_095_1973, w_095_1974, w_095_1977, w_095_1979, w_095_1980, w_095_1992, w_095_2008, w_095_2009, w_095_2012, w_095_2013, w_095_2014, w_095_2017, w_095_2020, w_095_2028, w_095_2029, w_095_2031, w_095_2032, w_095_2040, w_095_2041, w_095_2046, w_095_2047, w_095_2049, w_095_2051, w_095_2053, w_095_2054, w_095_2055, w_095_2060, w_095_2061, w_095_2066, w_095_2068, w_095_2071, w_095_2074, w_095_2076, w_095_2084, w_095_2094, w_095_2095, w_095_2109, w_095_2113, w_095_2114, w_095_2118, w_095_2121, w_095_2124, w_095_2128, w_095_2129, w_095_2130, w_095_2132, w_095_2139, w_095_2142, w_095_2143, w_095_2145, w_095_2149, w_095_2155, w_095_2157, w_095_2159, w_095_2163, w_095_2164, w_095_2167, w_095_2171, w_095_2175, w_095_2177, w_095_2179, w_095_2181, w_095_2185, w_095_2191, w_095_2196, w_095_2201, w_095_2205, w_095_2208, w_095_2211, w_095_2212, w_095_2213, w_095_2215, w_095_2221, w_095_2222, w_095_2223, w_095_2225, w_095_2226, w_095_2227, w_095_2231, w_095_2232, w_095_2233, w_095_2237, w_095_2243, w_095_2248, w_095_2250, w_095_2256, w_095_2257, w_095_2258, w_095_2260, w_095_2269, w_095_2273, w_095_2277, w_095_2291, w_095_2296, w_095_2298, w_095_2299, w_095_2301, w_095_2306, w_095_2313, w_095_2314, w_095_2318, w_095_2320, w_095_2324, w_095_2331, w_095_2334, w_095_2336, w_095_2340, w_095_2343, w_095_2345, w_095_2346, w_095_2347, w_095_2350, w_095_2352, w_095_2353, w_095_2360, w_095_2363, w_095_2368, w_095_2378, w_095_2380, w_095_2385, w_095_2388, w_095_2394, w_095_2396, w_095_2399, w_095_2403, w_095_2404, w_095_2409, w_095_2412, w_095_2418, w_095_2420, w_095_2427, w_095_2430, w_095_2437, w_095_2438, w_095_2441, w_095_2449, w_095_2451, w_095_2452, w_095_2456, w_095_2460, w_095_2466, w_095_2468, w_095_2472, w_095_2473, w_095_2475, w_095_2480, w_095_2485, w_095_2487, w_095_2488, w_095_2489, w_095_2490, w_095_2492, w_095_2493, w_095_2502, w_095_2505, w_095_2512, w_095_2524, w_095_2526, w_095_2527, w_095_2528, w_095_2529, w_095_2534, w_095_2535, w_095_2537, w_095_2540, w_095_2546, w_095_2551, w_095_2552, w_095_2555, w_095_2569, w_095_2570, w_095_2572, w_095_2579, w_095_2580, w_095_2584, w_095_2589, w_095_2593, w_095_2598, w_095_2599, w_095_2607, w_095_2609, w_095_2611, w_095_2613, w_095_2616, w_095_2619, w_095_2620, w_095_2623, w_095_2625, w_095_2628, w_095_2629, w_095_2636, w_095_2638, w_095_2639, w_095_2645, w_095_2653, w_095_2654, w_095_2655, w_095_2658, w_095_2667, w_095_2676, w_095_2684, w_095_2688, w_095_2694, w_095_2699, w_095_2700, w_095_2701, w_095_2702, w_095_2706, w_095_2714, w_095_2718, w_095_2725, w_095_2727, w_095_2729, w_095_2738, w_095_2749, w_095_2750, w_095_2754, w_095_2755, w_095_2756, w_095_2758, w_095_2759, w_095_2762, w_095_2771, w_095_2775, w_095_2776, w_095_2779, w_095_2780, w_095_2783, w_095_2784, w_095_2786, w_095_2788, w_095_2790, w_095_2794, w_095_2798, w_095_2811, w_095_2814, w_095_2816, w_095_2821, w_095_2822, w_095_2823, w_095_2824, w_095_2830, w_095_2839, w_095_2842, w_095_2843, w_095_2844, w_095_2847, w_095_2855, w_095_2856, w_095_2857, w_095_2862, w_095_2864, w_095_2870, w_095_2872, w_095_2873, w_095_2875, w_095_2883, w_095_2885, w_095_2887, w_095_2888, w_095_2891, w_095_2893, w_095_2895, w_095_2901, w_095_2902, w_095_2904, w_095_2913, w_095_2914, w_095_2918, w_095_2919, w_095_2920, w_095_2927, w_095_2930, w_095_2931, w_095_2935, w_095_2936, w_095_2940, w_095_2941, w_095_2942, w_095_2944, w_095_2947, w_095_2948, w_095_2955, w_095_2964, w_095_2975, w_095_2978, w_095_2993, w_095_2997, w_095_3002, w_095_3003, w_095_3007, w_095_3008, w_095_3010, w_095_3013, w_095_3014, w_095_3017, w_095_3019, w_095_3021, w_095_3023, w_095_3024, w_095_3025, w_095_3026, w_095_3043, w_095_3045, w_095_3047, w_095_3048, w_095_3050, w_095_3052, w_095_3054, w_095_3059, w_095_3061, w_095_3069, w_095_3071, w_095_3079, w_095_3083, w_095_3093, w_095_3097, w_095_3098, w_095_3103, w_095_3108, w_095_3110, w_095_3111, w_095_3112, w_095_3116, w_095_3119, w_095_3126, w_095_3128, w_095_3135, w_095_3136, w_095_3139, w_095_3149, w_095_3152, w_095_3155, w_095_3157, w_095_3158, w_095_3164, w_095_3176, w_095_3178, w_095_3184, w_095_3192, w_095_3194, w_095_3195, w_095_3200, w_095_3203, w_095_3204, w_095_3207, w_095_3208, w_095_3209, w_095_3217, w_095_3219, w_095_3220, w_095_3222, w_095_3225, w_095_3230, w_095_3231, w_095_3232, w_095_3234, w_095_3235, w_095_3236, w_095_3241, w_095_3243, w_095_3248, w_095_3254, w_095_3255, w_095_3256, w_095_3257, w_095_3259, w_095_3263, w_095_3264, w_095_3269, w_095_3273, w_095_3274, w_095_3279, w_095_3280, w_095_3281, w_095_3285, w_095_3286, w_095_3295, w_095_3297, w_095_3298, w_095_3300, w_095_3301, w_095_3304, w_095_3305, w_095_3310, w_095_3311, w_095_3316, w_095_3317, w_095_3320, w_095_3323, w_095_3324, w_095_3328, w_095_3333, w_095_3335, w_095_3340, w_095_3343, w_095_3346, w_095_3349, w_095_3350, w_095_3353, w_095_3354, w_095_3357, w_095_3360, w_095_3372, w_095_3373, w_095_3381, w_095_3383, w_095_3392, w_095_3396, w_095_3401, w_095_3411, w_095_3412, w_095_3414, w_095_3415, w_095_3420, w_095_3421, w_095_3422, w_095_3432, w_095_3437, w_095_3443, w_095_3446, w_095_3453, w_095_3454, w_095_3457, w_095_3458, w_095_3459, w_095_3460, w_095_3464, w_095_3466, w_095_3468, w_095_3469, w_095_3470, w_095_3480, w_095_3481, w_095_3482, w_095_3485, w_095_3486, w_095_3493, w_095_3495, w_095_3500, w_095_3501, w_095_3502, w_095_3509, w_095_3510, w_095_3512, w_095_3515, w_095_3519, w_095_3520, w_095_3521, w_095_3522, w_095_3526, w_095_3528, w_095_3530, w_095_3534, w_095_3537, w_095_3538, w_095_3540, w_095_3542, w_095_3546, w_095_3557, w_095_3558, w_095_3565, w_095_3567, w_095_3571, w_095_3574, w_095_3579, w_095_3582, w_095_3586, w_095_3587, w_095_3590, w_095_3591, w_095_3602, w_095_3604, w_095_3613, w_095_3615, w_095_3616, w_095_3620, w_095_3622, w_095_3624, w_095_3628, w_095_3630, w_095_3638, w_095_3641, w_095_3651, w_095_3652, w_095_3657, w_095_3658, w_095_3659, w_095_3660, w_095_3662, w_095_3664, w_095_3667, w_095_3674, w_095_3676, w_095_3679, w_095_3683, w_095_3688, w_095_3689, w_095_3691, w_095_3695, w_095_3706, w_095_3713, w_095_3719, w_095_3722, w_095_3723, w_095_3728, w_095_3730, w_095_3731, w_095_3738, w_095_3751, w_095_3753, w_095_3757, w_095_3763, w_095_3765, w_095_3769, w_095_3777, w_095_3779, w_095_3780, w_095_3782, w_095_3785, w_095_3786, w_095_3787, w_095_3788, w_095_3790, w_095_3791, w_095_3797, w_095_3800, w_095_3804, w_095_3805, w_095_3806, w_095_3807, w_095_3811, w_095_3813, w_095_3814, w_095_3825, w_095_3826, w_095_3827, w_095_3828, w_095_3831, w_095_3833, w_095_3838, w_095_3839, w_095_3847, w_095_3848, w_095_3850, w_095_3851, w_095_3852, w_095_3854, w_095_3868, w_095_3872, w_095_3883, w_095_3884, w_095_3885, w_095_3896, w_095_3897, w_095_3900, w_095_3902, w_095_3904, w_095_3909, w_095_3911, w_095_3912, w_095_3915, w_095_3917, w_095_3926, w_095_3928, w_095_3934, w_095_3937, w_095_3938, w_095_3939, w_095_3940, w_095_3950, w_095_3958, w_095_3959, w_095_3961, w_095_3963, w_095_3966, w_095_3967, w_095_3971, w_095_3976, w_095_3977, w_095_3979, w_095_3984, w_095_3994, w_095_3997, w_095_4000, w_095_4001, w_095_4003, w_095_4004, w_095_4005, w_095_4006, w_095_4009, w_095_4011, w_095_4015, w_095_4016, w_095_4019, w_095_4025, w_095_4027, w_095_4039, w_095_4040, w_095_4044, w_095_4047, w_095_4048;
  wire w_096_000, w_096_001, w_096_002, w_096_003, w_096_004, w_096_005, w_096_006, w_096_007, w_096_008, w_096_010, w_096_011, w_096_012, w_096_013, w_096_014, w_096_016, w_096_017, w_096_018, w_096_019, w_096_020, w_096_021, w_096_022, w_096_023, w_096_024, w_096_025, w_096_026, w_096_027, w_096_028, w_096_029, w_096_030, w_096_031, w_096_032, w_096_033, w_096_034, w_096_035, w_096_036, w_096_037, w_096_038, w_096_039, w_096_040, w_096_041, w_096_042, w_096_043, w_096_044, w_096_046, w_096_047, w_096_048, w_096_049, w_096_050, w_096_051, w_096_052, w_096_053, w_096_054, w_096_055, w_096_056, w_096_057, w_096_058, w_096_059, w_096_060, w_096_061, w_096_062, w_096_063, w_096_064, w_096_065, w_096_066, w_096_067, w_096_068, w_096_069, w_096_070, w_096_071, w_096_072, w_096_073, w_096_074, w_096_075, w_096_076, w_096_077, w_096_078, w_096_079, w_096_080, w_096_081, w_096_082, w_096_083, w_096_084, w_096_085, w_096_086, w_096_087, w_096_088, w_096_089, w_096_091, w_096_092, w_096_093, w_096_094, w_096_095, w_096_096, w_096_097, w_096_098, w_096_099, w_096_100, w_096_101, w_096_102, w_096_103, w_096_104, w_096_105, w_096_106, w_096_107, w_096_108, w_096_109, w_096_110, w_096_111, w_096_112, w_096_113, w_096_114, w_096_115, w_096_116, w_096_117, w_096_118, w_096_119, w_096_120, w_096_121, w_096_122, w_096_123, w_096_124, w_096_125, w_096_126, w_096_127, w_096_128, w_096_129, w_096_130, w_096_131, w_096_132, w_096_133, w_096_134, w_096_135, w_096_136, w_096_137, w_096_138, w_096_139, w_096_140, w_096_141, w_096_142, w_096_143, w_096_144, w_096_145, w_096_146, w_096_147, w_096_148, w_096_149, w_096_150, w_096_151, w_096_152, w_096_154, w_096_155, w_096_156, w_096_157, w_096_158, w_096_159, w_096_160, w_096_161, w_096_162, w_096_163, w_096_164, w_096_165, w_096_166, w_096_167, w_096_168, w_096_169, w_096_170, w_096_171, w_096_172, w_096_173, w_096_174, w_096_175, w_096_176, w_096_177, w_096_178, w_096_179, w_096_180, w_096_181, w_096_182, w_096_183, w_096_184, w_096_185, w_096_186, w_096_188, w_096_189, w_096_190, w_096_191, w_096_192, w_096_193, w_096_194, w_096_195, w_096_196, w_096_197, w_096_198, w_096_199, w_096_200, w_096_201, w_096_202, w_096_203, w_096_204, w_096_205, w_096_206, w_096_207, w_096_208, w_096_209, w_096_210, w_096_211, w_096_212, w_096_213, w_096_214, w_096_215, w_096_216, w_096_217, w_096_218, w_096_219, w_096_220, w_096_221, w_096_222, w_096_223, w_096_224, w_096_225, w_096_226, w_096_227, w_096_228, w_096_229, w_096_230, w_096_231, w_096_232, w_096_233, w_096_234, w_096_235, w_096_236, w_096_237, w_096_238, w_096_239, w_096_240, w_096_241, w_096_242, w_096_243, w_096_244, w_096_245, w_096_246, w_096_247, w_096_248, w_096_249, w_096_250, w_096_251, w_096_252, w_096_253, w_096_254, w_096_255, w_096_256, w_096_257, w_096_258, w_096_259, w_096_260, w_096_261, w_096_262, w_096_263, w_096_264, w_096_265, w_096_266, w_096_267, w_096_268, w_096_269, w_096_270, w_096_271, w_096_272, w_096_273, w_096_274, w_096_275, w_096_276, w_096_277, w_096_278, w_096_279, w_096_280, w_096_281, w_096_282, w_096_283, w_096_284, w_096_285, w_096_286, w_096_287, w_096_288, w_096_290, w_096_291, w_096_292, w_096_293, w_096_294, w_096_295, w_096_296, w_096_297, w_096_298, w_096_299, w_096_300, w_096_301, w_096_302, w_096_303, w_096_304, w_096_305, w_096_306, w_096_307, w_096_308, w_096_309, w_096_310, w_096_311, w_096_312, w_096_313, w_096_314, w_096_315, w_096_316, w_096_317, w_096_318, w_096_319, w_096_320, w_096_321, w_096_322, w_096_323, w_096_324, w_096_325, w_096_326, w_096_327, w_096_328, w_096_329, w_096_330, w_096_331, w_096_332, w_096_333, w_096_334, w_096_335, w_096_336, w_096_337, w_096_338, w_096_339, w_096_340, w_096_341, w_096_342, w_096_343, w_096_344, w_096_345, w_096_346, w_096_347, w_096_348, w_096_349, w_096_350, w_096_351, w_096_352, w_096_353, w_096_354, w_096_355, w_096_356, w_096_357, w_096_358, w_096_359, w_096_360, w_096_361, w_096_362, w_096_363, w_096_364, w_096_365, w_096_366, w_096_367, w_096_368, w_096_369, w_096_370, w_096_371, w_096_372, w_096_373, w_096_374, w_096_375, w_096_376, w_096_377, w_096_378, w_096_379, w_096_380, w_096_381, w_096_383, w_096_384, w_096_385, w_096_386, w_096_387, w_096_388, w_096_389, w_096_390, w_096_391, w_096_392, w_096_393, w_096_394, w_096_395, w_096_396, w_096_397, w_096_398, w_096_399, w_096_400, w_096_401, w_096_402, w_096_403, w_096_404, w_096_405, w_096_406, w_096_407, w_096_408, w_096_409, w_096_410, w_096_411, w_096_412, w_096_413, w_096_414, w_096_416, w_096_417, w_096_418, w_096_419, w_096_420, w_096_421, w_096_422, w_096_423, w_096_424, w_096_425, w_096_426, w_096_427, w_096_428, w_096_429, w_096_430, w_096_431, w_096_432, w_096_433, w_096_435, w_096_436, w_096_437, w_096_438, w_096_439, w_096_440, w_096_441, w_096_442, w_096_443, w_096_445, w_096_446, w_096_447, w_096_448, w_096_449, w_096_450, w_096_451, w_096_452, w_096_453, w_096_454, w_096_455, w_096_456, w_096_457, w_096_458, w_096_459, w_096_460, w_096_461, w_096_462, w_096_463, w_096_464, w_096_465, w_096_466, w_096_467, w_096_468, w_096_469, w_096_470, w_096_471, w_096_472, w_096_473, w_096_474, w_096_475, w_096_476, w_096_477, w_096_478, w_096_479, w_096_480, w_096_481, w_096_482, w_096_483, w_096_484, w_096_485, w_096_486, w_096_487, w_096_488, w_096_489, w_096_490, w_096_491, w_096_492, w_096_493, w_096_494, w_096_495, w_096_496, w_096_497, w_096_498, w_096_499, w_096_500, w_096_502, w_096_503, w_096_504, w_096_505, w_096_509, w_096_510, w_096_511, w_096_512, w_096_513, w_096_514, w_096_515, w_096_516, w_096_517, w_096_518, w_096_520;
  wire w_097_001, w_097_002, w_097_004, w_097_005, w_097_007, w_097_008, w_097_009, w_097_012, w_097_014, w_097_015, w_097_016, w_097_017, w_097_018, w_097_019, w_097_020, w_097_021, w_097_024, w_097_026, w_097_027, w_097_028, w_097_030, w_097_031, w_097_032, w_097_036, w_097_038, w_097_040, w_097_041, w_097_042, w_097_044, w_097_045, w_097_046, w_097_047, w_097_049, w_097_050, w_097_051, w_097_052, w_097_054, w_097_055, w_097_057, w_097_058, w_097_059, w_097_060, w_097_062, w_097_063, w_097_064, w_097_065, w_097_066, w_097_068, w_097_071, w_097_073, w_097_074, w_097_075, w_097_076, w_097_078, w_097_081, w_097_083, w_097_084, w_097_085, w_097_086, w_097_087, w_097_088, w_097_089, w_097_092, w_097_093, w_097_095, w_097_096, w_097_097, w_097_098, w_097_099, w_097_100, w_097_101, w_097_102, w_097_103, w_097_104, w_097_105, w_097_106, w_097_107, w_097_108, w_097_109, w_097_111, w_097_112, w_097_113, w_097_114, w_097_115, w_097_120, w_097_124, w_097_126, w_097_128, w_097_129, w_097_130, w_097_131, w_097_132, w_097_133, w_097_134, w_097_135, w_097_137, w_097_138, w_097_139, w_097_140, w_097_142, w_097_144, w_097_146, w_097_147, w_097_148, w_097_149, w_097_150, w_097_152, w_097_153, w_097_155, w_097_156, w_097_158, w_097_160, w_097_161, w_097_162, w_097_163, w_097_164, w_097_165, w_097_167, w_097_170, w_097_171, w_097_173, w_097_175, w_097_176, w_097_179, w_097_181, w_097_185, w_097_186, w_097_187, w_097_190, w_097_193, w_097_195, w_097_196, w_097_198, w_097_200, w_097_201, w_097_202, w_097_205, w_097_207, w_097_208, w_097_209, w_097_210, w_097_211, w_097_213, w_097_215, w_097_217, w_097_219, w_097_220, w_097_221, w_097_224, w_097_225, w_097_227, w_097_229, w_097_230, w_097_231, w_097_232, w_097_233, w_097_234, w_097_236, w_097_237, w_097_238, w_097_240, w_097_241, w_097_243, w_097_244, w_097_245, w_097_248, w_097_249, w_097_250, w_097_252, w_097_253, w_097_255, w_097_256, w_097_257, w_097_258, w_097_260, w_097_263, w_097_264, w_097_266, w_097_267, w_097_268, w_097_271, w_097_272, w_097_273, w_097_274, w_097_275, w_097_279, w_097_280, w_097_281, w_097_282, w_097_286, w_097_289, w_097_290, w_097_292, w_097_293, w_097_294, w_097_295, w_097_296, w_097_297, w_097_298, w_097_300, w_097_301, w_097_304, w_097_305, w_097_309, w_097_312, w_097_314, w_097_315, w_097_316, w_097_317, w_097_319, w_097_320, w_097_321, w_097_322, w_097_323, w_097_324, w_097_326, w_097_327, w_097_328, w_097_329, w_097_330, w_097_331, w_097_333, w_097_334, w_097_335, w_097_337, w_097_339, w_097_340, w_097_341, w_097_342, w_097_343, w_097_345, w_097_346, w_097_350, w_097_352, w_097_355, w_097_356, w_097_357, w_097_358, w_097_360, w_097_362, w_097_363, w_097_364, w_097_365, w_097_366, w_097_367, w_097_369, w_097_370, w_097_371, w_097_372, w_097_373, w_097_375, w_097_376, w_097_377, w_097_378, w_097_379, w_097_380, w_097_381, w_097_382, w_097_383, w_097_384, w_097_385, w_097_389, w_097_392, w_097_393, w_097_394, w_097_395, w_097_396, w_097_397, w_097_398, w_097_399, w_097_400, w_097_401, w_097_402, w_097_404, w_097_406, w_097_407, w_097_408, w_097_409, w_097_410, w_097_411, w_097_414, w_097_415, w_097_416, w_097_418, w_097_420, w_097_421, w_097_423, w_097_425, w_097_426, w_097_427, w_097_428, w_097_432, w_097_433, w_097_434, w_097_435, w_097_436, w_097_437, w_097_438, w_097_440, w_097_441, w_097_442, w_097_443, w_097_444, w_097_445, w_097_446, w_097_447, w_097_449, w_097_451, w_097_452, w_097_454, w_097_456, w_097_457, w_097_459, w_097_460, w_097_462, w_097_463, w_097_464, w_097_465, w_097_466, w_097_475, w_097_479, w_097_480, w_097_481, w_097_482, w_097_483, w_097_485, w_097_487, w_097_491, w_097_493, w_097_494, w_097_495, w_097_496, w_097_498, w_097_504, w_097_505, w_097_506, w_097_508, w_097_510, w_097_512, w_097_513, w_097_516, w_097_517, w_097_518, w_097_519, w_097_520, w_097_523, w_097_524, w_097_525, w_097_526, w_097_527, w_097_528, w_097_529, w_097_530, w_097_532, w_097_533, w_097_536, w_097_537, w_097_539, w_097_542, w_097_544, w_097_547, w_097_548, w_097_550, w_097_553, w_097_554, w_097_555, w_097_557, w_097_559, w_097_561, w_097_563, w_097_564, w_097_565, w_097_567, w_097_568, w_097_569, w_097_570, w_097_571, w_097_572, w_097_573, w_097_574, w_097_578, w_097_580, w_097_582, w_097_586, w_097_588, w_097_589, w_097_590, w_097_593, w_097_595, w_097_596, w_097_598, w_097_600, w_097_601, w_097_603, w_097_605, w_097_607, w_097_610, w_097_611, w_097_612, w_097_613, w_097_619, w_097_620, w_097_624, w_097_626, w_097_627, w_097_628, w_097_629, w_097_630, w_097_632, w_097_633, w_097_635, w_097_638, w_097_639, w_097_641, w_097_643, w_097_644, w_097_645, w_097_647, w_097_649, w_097_650, w_097_651, w_097_652, w_097_653, w_097_654, w_097_655, w_097_656, w_097_658, w_097_660, w_097_662, w_097_665, w_097_666, w_097_668, w_097_674, w_097_675, w_097_676, w_097_677, w_097_679, w_097_680, w_097_681, w_097_683, w_097_685, w_097_686, w_097_689, w_097_690, w_097_692, w_097_693, w_097_695, w_097_696, w_097_697, w_097_698, w_097_702, w_097_704, w_097_706, w_097_708, w_097_710, w_097_712, w_097_713, w_097_714, w_097_715, w_097_716, w_097_717, w_097_719, w_097_720, w_097_721, w_097_723, w_097_726, w_097_727, w_097_728, w_097_729, w_097_730, w_097_731, w_097_732, w_097_733, w_097_734, w_097_735, w_097_736, w_097_737, w_097_739, w_097_740, w_097_742, w_097_744, w_097_747, w_097_750, w_097_751, w_097_753, w_097_757, w_097_759, w_097_760, w_097_761, w_097_762, w_097_763, w_097_765, w_097_767, w_097_768, w_097_769, w_097_770, w_097_771, w_097_772, w_097_773, w_097_778, w_097_781, w_097_782, w_097_787, w_097_790, w_097_791, w_097_793, w_097_795, w_097_796, w_097_797, w_097_798, w_097_799, w_097_800, w_097_802, w_097_804, w_097_805, w_097_806, w_097_807, w_097_808, w_097_810, w_097_811, w_097_813, w_097_814, w_097_815, w_097_820, w_097_822, w_097_823, w_097_825, w_097_826, w_097_827, w_097_829, w_097_831, w_097_833, w_097_834, w_097_835, w_097_837, w_097_838, w_097_839, w_097_840, w_097_842, w_097_843, w_097_844, w_097_845, w_097_846, w_097_848, w_097_849, w_097_851, w_097_853, w_097_855, w_097_856, w_097_857, w_097_858, w_097_859, w_097_860, w_097_862, w_097_864, w_097_865, w_097_866, w_097_867, w_097_869, w_097_870, w_097_871, w_097_874, w_097_875, w_097_876, w_097_877, w_097_878, w_097_879, w_097_880, w_097_881, w_097_882, w_097_883, w_097_884, w_097_885, w_097_886, w_097_887, w_097_890, w_097_891, w_097_893, w_097_894, w_097_895, w_097_899, w_097_900, w_097_901, w_097_902, w_097_903, w_097_904, w_097_905, w_097_906, w_097_907, w_097_908, w_097_909, w_097_912, w_097_913, w_097_916, w_097_918, w_097_919, w_097_920, w_097_921, w_097_924, w_097_925, w_097_926, w_097_929, w_097_930, w_097_931, w_097_933, w_097_934, w_097_935, w_097_937, w_097_938, w_097_939, w_097_940, w_097_941, w_097_942, w_097_943, w_097_944, w_097_945, w_097_946, w_097_948, w_097_949, w_097_951, w_097_952, w_097_953, w_097_955, w_097_956, w_097_957, w_097_961, w_097_962, w_097_963, w_097_964, w_097_965, w_097_966, w_097_968, w_097_970, w_097_972, w_097_973, w_097_977, w_097_978, w_097_979, w_097_980, w_097_981, w_097_982, w_097_984, w_097_985, w_097_987, w_097_988, w_097_989, w_097_990, w_097_991, w_097_992, w_097_993, w_097_994, w_097_995, w_097_996, w_097_997, w_097_999, w_097_1001, w_097_1003, w_097_1006, w_097_1008, w_097_1011, w_097_1012, w_097_1014, w_097_1017, w_097_1020, w_097_1021, w_097_1022, w_097_1023, w_097_1024, w_097_1026, w_097_1027, w_097_1028, w_097_1030, w_097_1031, w_097_1034, w_097_1035, w_097_1036, w_097_1037, w_097_1039, w_097_1040, w_097_1041, w_097_1043, w_097_1044, w_097_1046, w_097_1047, w_097_1048, w_097_1050, w_097_1052, w_097_1053, w_097_1054, w_097_1055, w_097_1058, w_097_1059, w_097_1060, w_097_1063, w_097_1064, w_097_1065, w_097_1066, w_097_1068, w_097_1069, w_097_1070, w_097_1072, w_097_1075, w_097_1076, w_097_1078, w_097_1079, w_097_1081, w_097_1084, w_097_1087, w_097_1088, w_097_1089, w_097_1090, w_097_1091, w_097_1092, w_097_1093, w_097_1094, w_097_1095, w_097_1096, w_097_1097, w_097_1098, w_097_1100, w_097_1101, w_097_1102, w_097_1104, w_097_1106, w_097_1108, w_097_1110, w_097_1111, w_097_1112, w_097_1113, w_097_1114, w_097_1115, w_097_1118, w_097_1119, w_097_1120, w_097_1121, w_097_1122, w_097_1123, w_097_1125, w_097_1128, w_097_1129, w_097_1131, w_097_1133, w_097_1134, w_097_1136, w_097_1139, w_097_1140, w_097_1142, w_097_1143, w_097_1148, w_097_1149, w_097_1150, w_097_1151, w_097_1153, w_097_1154, w_097_1156, w_097_1158, w_097_1159, w_097_1160, w_097_1163, w_097_1164, w_097_1166, w_097_1167, w_097_1168, w_097_1169, w_097_1170, w_097_1174, w_097_1176, w_097_1177, w_097_1179, w_097_1181, w_097_1182, w_097_1184, w_097_1185, w_097_1187, w_097_1189, w_097_1190, w_097_1191, w_097_1193, w_097_1194, w_097_1195, w_097_1196, w_097_1198, w_097_1199, w_097_1202, w_097_1203, w_097_1206, w_097_1207, w_097_1208, w_097_1209, w_097_1210, w_097_1211, w_097_1213, w_097_1214, w_097_1216, w_097_1217, w_097_1218, w_097_1219, w_097_1220, w_097_1221, w_097_1227, w_097_1228, w_097_1229, w_097_1230, w_097_1232, w_097_1233, w_097_1234, w_097_1235, w_097_1236, w_097_1237, w_097_1239, w_097_1241, w_097_1242, w_097_1243, w_097_1244, w_097_1248, w_097_1250, w_097_1251, w_097_1253, w_097_1257, w_097_1258, w_097_1259, w_097_1260, w_097_1262, w_097_1265, w_097_1266, w_097_1267, w_097_1269, w_097_1270, w_097_1272, w_097_1275, w_097_1277, w_097_1278, w_097_1279, w_097_1280, w_097_1281, w_097_1282, w_097_1283, w_097_1287, w_097_1288, w_097_1289, w_097_1292, w_097_1293, w_097_1295, w_097_1296, w_097_1297, w_097_1300, w_097_1301, w_097_1302, w_097_1303, w_097_1304, w_097_1305, w_097_1306, w_097_1309, w_097_1310, w_097_1314, w_097_1315, w_097_1316, w_097_1317, w_097_1319, w_097_1320, w_097_1321, w_097_1322, w_097_1325, w_097_1328, w_097_1329, w_097_1330, w_097_1332, w_097_1333, w_097_1334, w_097_1335, w_097_1339, w_097_1341, w_097_1343, w_097_1344, w_097_1346, w_097_1348, w_097_1350, w_097_1352, w_097_1353, w_097_1354, w_097_1356, w_097_1358, w_097_1359, w_097_1360, w_097_1361, w_097_1363, w_097_1365, w_097_1366, w_097_1367, w_097_1368, w_097_1370, w_097_1372, w_097_1373, w_097_1374, w_097_1375, w_097_1378, w_097_1379, w_097_1380, w_097_1381, w_097_1383, w_097_1384, w_097_1386, w_097_1387, w_097_1388, w_097_1389, w_097_1390, w_097_1391, w_097_1392, w_097_1394, w_097_1395, w_097_1402, w_097_1403, w_097_1404, w_097_1405, w_097_1406, w_097_1407, w_097_1408, w_097_1410, w_097_1412, w_097_1413, w_097_1415, w_097_1416, w_097_1417, w_097_1419, w_097_1420, w_097_1421, w_097_1423, w_097_1424, w_097_1425, w_097_1426, w_097_1427, w_097_1428, w_097_1429, w_097_1430, w_097_1435, w_097_1436, w_097_1437, w_097_1438, w_097_1439, w_097_1440, w_097_1441, w_097_1442, w_097_1443, w_097_1446, w_097_1447, w_097_1448, w_097_1449, w_097_1451, w_097_1452, w_097_1453, w_097_1454, w_097_1455, w_097_1456, w_097_1460, w_097_1461, w_097_1462, w_097_1464, w_097_1467, w_097_1469, w_097_1472, w_097_1475, w_097_1476, w_097_1477, w_097_1480, w_097_1481, w_097_1483, w_097_1484, w_097_1485, w_097_1486, w_097_1489, w_097_1490, w_097_1493, w_097_1495, w_097_1496, w_097_1497, w_097_1502, w_097_1505, w_097_1507, w_097_1508, w_097_1510, w_097_1511, w_097_1513, w_097_1517, w_097_1519, w_097_1520, w_097_1523, w_097_1524, w_097_1525, w_097_1526, w_097_1527, w_097_1528, w_097_1529, w_097_1530, w_097_1532, w_097_1533, w_097_1534, w_097_1535, w_097_1536, w_097_1537, w_097_1540, w_097_1541, w_097_1542, w_097_1543, w_097_1544, w_097_1545, w_097_1546, w_097_1548, w_097_1549, w_097_1551, w_097_1552, w_097_1553, w_097_1554, w_097_1555, w_097_1556, w_097_1557, w_097_1559, w_097_1560, w_097_1561, w_097_1562, w_097_1563, w_097_1564, w_097_1565, w_097_1569, w_097_1570, w_097_1571, w_097_1572, w_097_1573, w_097_1574, w_097_1575, w_097_1577, w_097_1579, w_097_1581, w_097_1582, w_097_1583, w_097_1585, w_097_1588, w_097_1589, w_097_1592, w_097_1594, w_097_1595, w_097_1596, w_097_1598, w_097_1599, w_097_1601, w_097_1603, w_097_1604, w_097_1605, w_097_1606, w_097_1607, w_097_1608, w_097_1610, w_097_1612, w_097_1613, w_097_1616, w_097_1617, w_097_1618, w_097_1619, w_097_1622, w_097_1623, w_097_1625, w_097_1626, w_097_1627, w_097_1628, w_097_1629, w_097_1630, w_097_1631, w_097_1632, w_097_1633, w_097_1636, w_097_1637, w_097_1639, w_097_1640, w_097_1641, w_097_1642, w_097_1644, w_097_1645, w_097_1647, w_097_1648;
  wire w_098_000, w_098_001, w_098_002, w_098_004, w_098_005, w_098_006, w_098_007, w_098_008, w_098_009, w_098_010, w_098_011, w_098_012, w_098_013, w_098_014, w_098_015, w_098_016, w_098_017, w_098_018, w_098_019, w_098_022, w_098_023, w_098_024, w_098_026, w_098_027, w_098_029, w_098_030, w_098_031, w_098_032, w_098_033, w_098_034, w_098_035, w_098_036, w_098_037, w_098_038, w_098_039, w_098_040, w_098_041, w_098_042, w_098_044, w_098_045, w_098_048, w_098_050, w_098_051, w_098_052, w_098_053, w_098_054, w_098_056, w_098_057, w_098_058, w_098_059, w_098_060, w_098_062, w_098_063, w_098_065, w_098_066, w_098_067, w_098_069, w_098_070, w_098_071, w_098_074, w_098_075, w_098_076, w_098_077, w_098_078, w_098_079, w_098_080, w_098_081, w_098_082, w_098_086, w_098_087, w_098_088, w_098_089, w_098_093, w_098_095, w_098_096, w_098_097, w_098_099, w_098_101, w_098_102, w_098_104, w_098_105, w_098_106, w_098_107, w_098_111, w_098_112, w_098_113, w_098_115, w_098_117, w_098_121, w_098_122, w_098_123, w_098_124, w_098_128, w_098_130, w_098_131, w_098_135, w_098_137, w_098_141, w_098_142, w_098_143, w_098_144, w_098_145, w_098_147, w_098_149, w_098_152, w_098_154, w_098_155, w_098_156, w_098_157, w_098_158, w_098_159, w_098_160, w_098_165, w_098_166, w_098_167, w_098_168, w_098_169, w_098_173, w_098_174, w_098_176, w_098_177, w_098_180, w_098_182, w_098_183, w_098_185, w_098_186, w_098_187, w_098_188, w_098_189, w_098_190, w_098_192, w_098_195, w_098_196, w_098_198, w_098_199, w_098_200, w_098_203, w_098_204, w_098_207, w_098_208, w_098_209, w_098_210, w_098_213, w_098_217, w_098_219, w_098_220, w_098_221, w_098_223, w_098_224, w_098_229, w_098_231, w_098_235, w_098_237, w_098_238, w_098_239, w_098_245, w_098_247, w_098_248, w_098_249, w_098_250, w_098_251, w_098_252, w_098_254, w_098_255, w_098_256, w_098_257, w_098_259, w_098_261, w_098_263, w_098_264, w_098_265, w_098_266, w_098_267, w_098_268, w_098_269, w_098_272, w_098_273, w_098_275, w_098_278, w_098_280, w_098_281, w_098_282, w_098_283, w_098_284, w_098_285, w_098_287, w_098_288, w_098_290, w_098_293, w_098_294, w_098_295, w_098_296, w_098_297, w_098_299, w_098_301, w_098_304, w_098_305, w_098_306, w_098_308, w_098_309, w_098_310, w_098_311, w_098_312, w_098_313, w_098_314, w_098_315, w_098_317, w_098_318, w_098_320, w_098_321, w_098_322, w_098_327, w_098_328, w_098_331, w_098_338, w_098_339, w_098_340, w_098_342, w_098_348, w_098_349, w_098_351, w_098_352, w_098_356, w_098_358, w_098_359, w_098_363, w_098_364, w_098_365, w_098_366, w_098_367, w_098_368, w_098_369, w_098_370, w_098_373, w_098_374, w_098_376, w_098_378, w_098_379, w_098_381, w_098_382, w_098_383, w_098_384, w_098_386, w_098_387, w_098_388, w_098_389, w_098_390, w_098_391, w_098_392, w_098_393, w_098_394, w_098_395, w_098_398, w_098_399, w_098_400, w_098_401, w_098_402, w_098_404, w_098_405, w_098_406, w_098_408, w_098_410, w_098_411, w_098_412, w_098_413, w_098_414, w_098_416, w_098_418, w_098_419, w_098_420, w_098_421, w_098_422, w_098_423, w_098_424, w_098_426, w_098_428, w_098_429, w_098_430, w_098_432, w_098_434, w_098_435, w_098_437, w_098_439, w_098_440, w_098_442, w_098_443, w_098_445, w_098_449, w_098_450, w_098_451, w_098_452, w_098_453, w_098_454, w_098_456, w_098_457, w_098_459, w_098_463, w_098_464, w_098_468, w_098_469, w_098_472, w_098_473, w_098_474, w_098_475, w_098_476, w_098_477, w_098_481, w_098_482, w_098_483, w_098_484, w_098_486, w_098_488, w_098_489, w_098_490, w_098_491, w_098_492, w_098_493, w_098_494, w_098_496, w_098_497, w_098_498, w_098_500, w_098_503, w_098_506, w_098_508, w_098_509, w_098_510, w_098_511, w_098_512, w_098_513, w_098_514, w_098_517, w_098_518, w_098_521, w_098_525, w_098_527, w_098_528, w_098_530, w_098_531, w_098_533, w_098_534, w_098_536, w_098_538, w_098_540, w_098_543, w_098_544, w_098_545, w_098_546, w_098_547, w_098_549, w_098_550, w_098_553, w_098_554, w_098_555, w_098_557, w_098_558, w_098_559, w_098_560, w_098_562, w_098_563, w_098_565, w_098_566, w_098_567, w_098_568, w_098_571, w_098_572, w_098_573, w_098_576, w_098_578, w_098_579, w_098_580, w_098_584, w_098_585, w_098_589, w_098_590, w_098_591, w_098_592, w_098_593, w_098_595, w_098_596, w_098_598, w_098_599, w_098_600, w_098_602, w_098_603, w_098_608, w_098_609, w_098_615, w_098_616, w_098_617, w_098_619, w_098_620, w_098_621, w_098_623, w_098_624, w_098_625, w_098_627, w_098_629, w_098_630, w_098_631, w_098_632, w_098_633, w_098_637, w_098_638, w_098_639, w_098_640, w_098_641, w_098_642, w_098_646, w_098_647, w_098_648, w_098_650, w_098_652, w_098_653, w_098_654, w_098_657, w_098_659, w_098_660, w_098_661, w_098_662, w_098_663, w_098_664, w_098_666, w_098_672, w_098_673, w_098_675, w_098_676, w_098_678, w_098_681, w_098_682, w_098_683, w_098_684, w_098_686, w_098_687, w_098_688, w_098_692, w_098_693, w_098_695, w_098_696, w_098_697, w_098_699, w_098_706, w_098_707, w_098_709, w_098_710, w_098_714, w_098_715, w_098_716, w_098_717, w_098_719, w_098_720, w_098_721, w_098_723, w_098_724, w_098_725, w_098_726, w_098_728, w_098_729, w_098_730, w_098_734, w_098_735, w_098_736, w_098_737, w_098_739, w_098_741, w_098_742, w_098_743, w_098_744, w_098_745, w_098_746, w_098_747, w_098_748, w_098_750, w_098_751, w_098_752, w_098_755, w_098_757, w_098_759, w_098_760, w_098_761, w_098_762, w_098_763, w_098_765, w_098_767, w_098_768, w_098_770, w_098_771, w_098_773, w_098_774, w_098_776, w_098_779, w_098_780, w_098_781, w_098_782, w_098_783, w_098_784, w_098_785, w_098_789, w_098_791, w_098_792, w_098_793, w_098_794, w_098_796, w_098_799, w_098_800, w_098_801, w_098_802, w_098_803, w_098_804, w_098_806, w_098_807, w_098_808, w_098_809, w_098_810, w_098_811, w_098_812, w_098_814, w_098_817, w_098_819, w_098_820, w_098_821, w_098_822, w_098_826, w_098_827, w_098_829, w_098_833, w_098_834, w_098_838, w_098_839, w_098_840, w_098_841, w_098_843, w_098_844, w_098_845, w_098_847, w_098_848, w_098_849, w_098_851, w_098_853, w_098_854, w_098_857, w_098_858, w_098_860, w_098_861, w_098_862, w_098_863, w_098_864, w_098_865, w_098_868, w_098_871, w_098_873, w_098_876, w_098_877, w_098_880, w_098_881, w_098_882, w_098_886, w_098_887, w_098_888, w_098_889, w_098_890, w_098_892, w_098_894, w_098_896, w_098_898, w_098_899, w_098_900, w_098_901, w_098_902, w_098_903, w_098_904, w_098_905, w_098_909, w_098_910, w_098_911, w_098_912, w_098_913, w_098_914, w_098_915, w_098_916, w_098_919, w_098_920, w_098_922, w_098_924, w_098_925, w_098_926, w_098_928, w_098_929, w_098_930, w_098_931, w_098_932, w_098_933, w_098_934, w_098_935, w_098_936, w_098_937, w_098_938, w_098_939, w_098_940, w_098_945, w_098_947, w_098_948, w_098_949, w_098_950, w_098_951, w_098_953, w_098_954, w_098_958, w_098_960, w_098_961, w_098_962, w_098_963, w_098_965, w_098_971, w_098_973, w_098_975, w_098_976, w_098_981, w_098_982, w_098_984, w_098_986, w_098_987, w_098_991, w_098_993, w_098_994, w_098_995, w_098_996, w_098_998, w_098_1000, w_098_1001, w_098_1003, w_098_1004, w_098_1005, w_098_1006, w_098_1008, w_098_1009, w_098_1010, w_098_1011, w_098_1013, w_098_1015, w_098_1016, w_098_1017, w_098_1019, w_098_1020, w_098_1021, w_098_1023, w_098_1024, w_098_1025, w_098_1026, w_098_1031, w_098_1032, w_098_1033, w_098_1035, w_098_1036, w_098_1037, w_098_1039, w_098_1040, w_098_1041, w_098_1042, w_098_1043, w_098_1044, w_098_1048, w_098_1049, w_098_1050, w_098_1051, w_098_1052, w_098_1055, w_098_1056, w_098_1058, w_098_1059, w_098_1060, w_098_1062, w_098_1063, w_098_1064, w_098_1065, w_098_1066, w_098_1067, w_098_1068, w_098_1070, w_098_1071, w_098_1072, w_098_1073, w_098_1074, w_098_1075, w_098_1076, w_098_1079, w_098_1083, w_098_1084, w_098_1087, w_098_1088, w_098_1089, w_098_1090, w_098_1091, w_098_1095, w_098_1096, w_098_1097, w_098_1100, w_098_1103, w_098_1106, w_098_1108, w_098_1109, w_098_1111, w_098_1112, w_098_1113, w_098_1114, w_098_1117, w_098_1119, w_098_1121, w_098_1123, w_098_1124, w_098_1126, w_098_1127, w_098_1128, w_098_1130, w_098_1131, w_098_1132, w_098_1133, w_098_1136, w_098_1137, w_098_1138, w_098_1139, w_098_1141, w_098_1142, w_098_1143, w_098_1147, w_098_1148, w_098_1149, w_098_1150, w_098_1154, w_098_1155, w_098_1156, w_098_1157, w_098_1158, w_098_1159, w_098_1163, w_098_1164, w_098_1165, w_098_1166, w_098_1168, w_098_1171, w_098_1172, w_098_1174, w_098_1176, w_098_1177, w_098_1179, w_098_1183, w_098_1185, w_098_1187, w_098_1189, w_098_1190, w_098_1191, w_098_1193, w_098_1194, w_098_1195, w_098_1196, w_098_1198, w_098_1199, w_098_1202, w_098_1204, w_098_1205, w_098_1207, w_098_1208, w_098_1213, w_098_1214, w_098_1217, w_098_1218, w_098_1222, w_098_1223, w_098_1224, w_098_1225, w_098_1226, w_098_1229, w_098_1230, w_098_1231, w_098_1232, w_098_1234, w_098_1236, w_098_1237, w_098_1238, w_098_1239, w_098_1240, w_098_1242, w_098_1243, w_098_1244, w_098_1245, w_098_1248, w_098_1249, w_098_1251, w_098_1252, w_098_1253, w_098_1254, w_098_1255, w_098_1256, w_098_1257, w_098_1258, w_098_1261, w_098_1262, w_098_1263, w_098_1264, w_098_1265, w_098_1266, w_098_1267, w_098_1268, w_098_1270, w_098_1271, w_098_1272, w_098_1273, w_098_1274, w_098_1275, w_098_1277, w_098_1278, w_098_1280, w_098_1281, w_098_1282, w_098_1284, w_098_1288, w_098_1289, w_098_1290, w_098_1291, w_098_1292, w_098_1293, w_098_1296, w_098_1300, w_098_1301, w_098_1303, w_098_1304, w_098_1305, w_098_1306, w_098_1307, w_098_1308, w_098_1309, w_098_1310, w_098_1311, w_098_1312, w_098_1314, w_098_1315, w_098_1317, w_098_1318, w_098_1320, w_098_1321, w_098_1323, w_098_1324, w_098_1325, w_098_1326, w_098_1327, w_098_1328, w_098_1331, w_098_1332, w_098_1333, w_098_1335, w_098_1336, w_098_1338, w_098_1341, w_098_1342, w_098_1344, w_098_1345, w_098_1346, w_098_1347, w_098_1348, w_098_1349, w_098_1350, w_098_1351, w_098_1352, w_098_1354, w_098_1357, w_098_1358, w_098_1359, w_098_1360, w_098_1365, w_098_1366, w_098_1367, w_098_1369, w_098_1370, w_098_1371, w_098_1372, w_098_1373, w_098_1375, w_098_1376, w_098_1377, w_098_1378, w_098_1379, w_098_1381, w_098_1382, w_098_1383, w_098_1384, w_098_1385, w_098_1386, w_098_1389, w_098_1391, w_098_1392, w_098_1393, w_098_1396, w_098_1399, w_098_1400, w_098_1401, w_098_1402, w_098_1403, w_098_1404, w_098_1405, w_098_1406, w_098_1409, w_098_1411, w_098_1412, w_098_1413, w_098_1416, w_098_1422, w_098_1424, w_098_1425, w_098_1426, w_098_1431, w_098_1432, w_098_1434, w_098_1435, w_098_1436, w_098_1438, w_098_1441, w_098_1442, w_098_1445, w_098_1447, w_098_1449, w_098_1450, w_098_1451, w_098_1452, w_098_1453, w_098_1454, w_098_1459, w_098_1460, w_098_1461, w_098_1462, w_098_1463, w_098_1464, w_098_1466, w_098_1469, w_098_1471, w_098_1474, w_098_1476, w_098_1477, w_098_1480, w_098_1481, w_098_1483, w_098_1486, w_098_1487, w_098_1488, w_098_1491, w_098_1492, w_098_1497, w_098_1498, w_098_1501, w_098_1503, w_098_1504, w_098_1505, w_098_1508, w_098_1509, w_098_1510, w_098_1512, w_098_1513, w_098_1515, w_098_1517, w_098_1518, w_098_1519, w_098_1521, w_098_1524, w_098_1526, w_098_1527, w_098_1528, w_098_1529, w_098_1530, w_098_1531, w_098_1532, w_098_1533, w_098_1534, w_098_1535, w_098_1538, w_098_1539, w_098_1541, w_098_1542, w_098_1544, w_098_1546, w_098_1547, w_098_1549, w_098_1551, w_098_1552, w_098_1553, w_098_1555, w_098_1556, w_098_1557, w_098_1558, w_098_1559, w_098_1562, w_098_1563, w_098_1565, w_098_1567, w_098_1569, w_098_1571, w_098_1574, w_098_1575, w_098_1576, w_098_1577, w_098_1578, w_098_1580, w_098_1581, w_098_1582, w_098_1583, w_098_1584, w_098_1585, w_098_1588, w_098_1590, w_098_1594, w_098_1595, w_098_1597, w_098_1599, w_098_1600, w_098_1603, w_098_1605, w_098_1607, w_098_1608, w_098_1609, w_098_1612, w_098_1614, w_098_1617, w_098_1619, w_098_1621, w_098_1623, w_098_1626, w_098_1627, w_098_1629, w_098_1630, w_098_1632, w_098_1633, w_098_1635, w_098_1636;
  wire w_099_001, w_099_003, w_099_004, w_099_006, w_099_007, w_099_011, w_099_012, w_099_013, w_099_014, w_099_019, w_099_023, w_099_024, w_099_025, w_099_026, w_099_028, w_099_030, w_099_031, w_099_036, w_099_037, w_099_039, w_099_042, w_099_043, w_099_044, w_099_045, w_099_046, w_099_050, w_099_051, w_099_054, w_099_055, w_099_059, w_099_064, w_099_066, w_099_068, w_099_071, w_099_073, w_099_081, w_099_082, w_099_083, w_099_087, w_099_088, w_099_089, w_099_090, w_099_093, w_099_097, w_099_100, w_099_101, w_099_105, w_099_107, w_099_108, w_099_109, w_099_110, w_099_111, w_099_112, w_099_117, w_099_118, w_099_119, w_099_123, w_099_124, w_099_125, w_099_130, w_099_133, w_099_134, w_099_135, w_099_138, w_099_142, w_099_147, w_099_151, w_099_154, w_099_155, w_099_156, w_099_159, w_099_163, w_099_164, w_099_166, w_099_168, w_099_170, w_099_172, w_099_174, w_099_176, w_099_178, w_099_182, w_099_183, w_099_187, w_099_190, w_099_191, w_099_194, w_099_197, w_099_200, w_099_204, w_099_205, w_099_207, w_099_208, w_099_209, w_099_211, w_099_212, w_099_213, w_099_214, w_099_217, w_099_219, w_099_225, w_099_227, w_099_230, w_099_231, w_099_233, w_099_234, w_099_235, w_099_238, w_099_239, w_099_240, w_099_244, w_099_246, w_099_247, w_099_249, w_099_250, w_099_254, w_099_255, w_099_256, w_099_257, w_099_263, w_099_269, w_099_270, w_099_271, w_099_272, w_099_275, w_099_279, w_099_280, w_099_284, w_099_285, w_099_290, w_099_292, w_099_294, w_099_296, w_099_297, w_099_299, w_099_301, w_099_303, w_099_304, w_099_305, w_099_308, w_099_311, w_099_313, w_099_314, w_099_315, w_099_316, w_099_317, w_099_323, w_099_329, w_099_330, w_099_331, w_099_333, w_099_335, w_099_340, w_099_342, w_099_343, w_099_346, w_099_347, w_099_348, w_099_349, w_099_352, w_099_354, w_099_355, w_099_358, w_099_360, w_099_362, w_099_365, w_099_371, w_099_372, w_099_374, w_099_377, w_099_380, w_099_381, w_099_382, w_099_383, w_099_385, w_099_386, w_099_387, w_099_388, w_099_389, w_099_390, w_099_391, w_099_394, w_099_396, w_099_403, w_099_405, w_099_406, w_099_408, w_099_409, w_099_410, w_099_412, w_099_413, w_099_414, w_099_415, w_099_419, w_099_421, w_099_422, w_099_424, w_099_425, w_099_426, w_099_427, w_099_431, w_099_432, w_099_433, w_099_434, w_099_436, w_099_437, w_099_438, w_099_439, w_099_441, w_099_443, w_099_445, w_099_446, w_099_447, w_099_450, w_099_451, w_099_453, w_099_455, w_099_456, w_099_461, w_099_463, w_099_465, w_099_468, w_099_469, w_099_472, w_099_474, w_099_479, w_099_483, w_099_486, w_099_487, w_099_490, w_099_494, w_099_498, w_099_499, w_099_501, w_099_503, w_099_504, w_099_505, w_099_507, w_099_513, w_099_516, w_099_519, w_099_524, w_099_526, w_099_528, w_099_529, w_099_530, w_099_531, w_099_534, w_099_540, w_099_544, w_099_546, w_099_547, w_099_548, w_099_550, w_099_551, w_099_553, w_099_555, w_099_557, w_099_558, w_099_563, w_099_566, w_099_569, w_099_571, w_099_575, w_099_576, w_099_577, w_099_578, w_099_580, w_099_581, w_099_582, w_099_583, w_099_586, w_099_588, w_099_590, w_099_592, w_099_594, w_099_597, w_099_599, w_099_600, w_099_601, w_099_602, w_099_606, w_099_608, w_099_612, w_099_613, w_099_614, w_099_616, w_099_617, w_099_623, w_099_624, w_099_627, w_099_629, w_099_630, w_099_631, w_099_632, w_099_633, w_099_634, w_099_638, w_099_640, w_099_644, w_099_645, w_099_647, w_099_651, w_099_652, w_099_654, w_099_656, w_099_661, w_099_662, w_099_667, w_099_669, w_099_670, w_099_672, w_099_674, w_099_676, w_099_678, w_099_679, w_099_680, w_099_682, w_099_684, w_099_685, w_099_687, w_099_691, w_099_694, w_099_695, w_099_696, w_099_697, w_099_698, w_099_699, w_099_700, w_099_701, w_099_705, w_099_706, w_099_708, w_099_709, w_099_710, w_099_711, w_099_712, w_099_713, w_099_716, w_099_719, w_099_721, w_099_723, w_099_729, w_099_730, w_099_732, w_099_738, w_099_741, w_099_744, w_099_749, w_099_750, w_099_752, w_099_753, w_099_756, w_099_757, w_099_762, w_099_765, w_099_767, w_099_770, w_099_773, w_099_779, w_099_780, w_099_786, w_099_787, w_099_796, w_099_797, w_099_799, w_099_801, w_099_803, w_099_808, w_099_810, w_099_811, w_099_818, w_099_824, w_099_826, w_099_827, w_099_828, w_099_831, w_099_832, w_099_834, w_099_839, w_099_840, w_099_847, w_099_854, w_099_856, w_099_858, w_099_859, w_099_864, w_099_865, w_099_866, w_099_876, w_099_880, w_099_882, w_099_883, w_099_884, w_099_888, w_099_890, w_099_892, w_099_894, w_099_895, w_099_901, w_099_905, w_099_907, w_099_909, w_099_914, w_099_918, w_099_921, w_099_922, w_099_924, w_099_925, w_099_927, w_099_928, w_099_930, w_099_933, w_099_934, w_099_935, w_099_936, w_099_948, w_099_949, w_099_952, w_099_954, w_099_957, w_099_960, w_099_961, w_099_962, w_099_963, w_099_967, w_099_974, w_099_975, w_099_982, w_099_987, w_099_990, w_099_991, w_099_992, w_099_993, w_099_994, w_099_997, w_099_1005, w_099_1012, w_099_1015, w_099_1021, w_099_1022, w_099_1024, w_099_1027, w_099_1031, w_099_1034, w_099_1036, w_099_1038, w_099_1041, w_099_1042, w_099_1044, w_099_1046, w_099_1049, w_099_1050, w_099_1053, w_099_1055, w_099_1058, w_099_1059, w_099_1065, w_099_1068, w_099_1070, w_099_1073, w_099_1075, w_099_1076, w_099_1086, w_099_1093, w_099_1099, w_099_1100, w_099_1102, w_099_1103, w_099_1106, w_099_1109, w_099_1114, w_099_1117, w_099_1123, w_099_1125, w_099_1127, w_099_1128, w_099_1133, w_099_1134, w_099_1136, w_099_1137, w_099_1140, w_099_1141, w_099_1143, w_099_1144, w_099_1146, w_099_1147, w_099_1148, w_099_1149, w_099_1152, w_099_1153, w_099_1155, w_099_1156, w_099_1157, w_099_1158, w_099_1166, w_099_1167, w_099_1170, w_099_1173, w_099_1186, w_099_1188, w_099_1191, w_099_1193, w_099_1194, w_099_1207, w_099_1208, w_099_1211, w_099_1215, w_099_1218, w_099_1222, w_099_1223, w_099_1224, w_099_1225, w_099_1226, w_099_1229, w_099_1235, w_099_1236, w_099_1242, w_099_1243, w_099_1248, w_099_1251, w_099_1254, w_099_1255, w_099_1256, w_099_1258, w_099_1262, w_099_1263, w_099_1266, w_099_1267, w_099_1273, w_099_1280, w_099_1282, w_099_1284, w_099_1285, w_099_1286, w_099_1287, w_099_1291, w_099_1297, w_099_1298, w_099_1299, w_099_1301, w_099_1304, w_099_1313, w_099_1314, w_099_1315, w_099_1317, w_099_1323, w_099_1328, w_099_1330, w_099_1331, w_099_1334, w_099_1335, w_099_1336, w_099_1341, w_099_1344, w_099_1347, w_099_1348, w_099_1351, w_099_1352, w_099_1353, w_099_1362, w_099_1365, w_099_1367, w_099_1371, w_099_1372, w_099_1376, w_099_1377, w_099_1379, w_099_1382, w_099_1386, w_099_1388, w_099_1390, w_099_1396, w_099_1397, w_099_1398, w_099_1400, w_099_1403, w_099_1404, w_099_1415, w_099_1419, w_099_1427, w_099_1428, w_099_1431, w_099_1432, w_099_1433, w_099_1436, w_099_1437, w_099_1438, w_099_1440, w_099_1441, w_099_1448, w_099_1449, w_099_1450, w_099_1457, w_099_1459, w_099_1460, w_099_1461, w_099_1464, w_099_1466, w_099_1467, w_099_1475, w_099_1476, w_099_1483, w_099_1484, w_099_1485, w_099_1486, w_099_1487, w_099_1488, w_099_1490, w_099_1506, w_099_1509, w_099_1510, w_099_1514, w_099_1515, w_099_1518, w_099_1526, w_099_1530, w_099_1532, w_099_1533, w_099_1535, w_099_1537, w_099_1540, w_099_1541, w_099_1542, w_099_1546, w_099_1549, w_099_1550, w_099_1556, w_099_1558, w_099_1562, w_099_1567, w_099_1573, w_099_1574, w_099_1575, w_099_1579, w_099_1585, w_099_1587, w_099_1588, w_099_1589, w_099_1592, w_099_1596, w_099_1597, w_099_1608, w_099_1612, w_099_1624, w_099_1625, w_099_1627, w_099_1629, w_099_1631, w_099_1635, w_099_1647, w_099_1648, w_099_1657, w_099_1659, w_099_1662, w_099_1663, w_099_1665, w_099_1669, w_099_1674, w_099_1678, w_099_1680, w_099_1681, w_099_1689, w_099_1692, w_099_1704, w_099_1705, w_099_1706, w_099_1716, w_099_1719, w_099_1720, w_099_1725, w_099_1728, w_099_1733, w_099_1735, w_099_1737, w_099_1740, w_099_1741, w_099_1750, w_099_1751, w_099_1752, w_099_1753, w_099_1756, w_099_1758, w_099_1761, w_099_1763, w_099_1765, w_099_1766, w_099_1767, w_099_1768, w_099_1769, w_099_1770, w_099_1771, w_099_1776, w_099_1783, w_099_1784, w_099_1795, w_099_1797, w_099_1799, w_099_1803, w_099_1810, w_099_1811, w_099_1814, w_099_1818, w_099_1819, w_099_1828, w_099_1829, w_099_1832, w_099_1834, w_099_1837, w_099_1840, w_099_1841, w_099_1846, w_099_1857, w_099_1858, w_099_1869, w_099_1877, w_099_1882, w_099_1885, w_099_1891, w_099_1902, w_099_1905, w_099_1910, w_099_1916, w_099_1920, w_099_1922, w_099_1924, w_099_1929, w_099_1932, w_099_1937, w_099_1939, w_099_1941, w_099_1942, w_099_1948, w_099_1951, w_099_1954, w_099_1958, w_099_1963, w_099_1969, w_099_1973, w_099_1974, w_099_1977, w_099_1979, w_099_1981, w_099_1983, w_099_1986, w_099_1989, w_099_1990, w_099_1991, w_099_1996, w_099_2005, w_099_2009, w_099_2011, w_099_2012, w_099_2015, w_099_2018, w_099_2022, w_099_2028, w_099_2032, w_099_2033, w_099_2034, w_099_2036, w_099_2039, w_099_2048, w_099_2050, w_099_2051, w_099_2063, w_099_2064, w_099_2068, w_099_2072, w_099_2076, w_099_2093, w_099_2094, w_099_2098, w_099_2101, w_099_2110, w_099_2119, w_099_2123, w_099_2129, w_099_2139, w_099_2140, w_099_2142, w_099_2144, w_099_2148, w_099_2156, w_099_2165, w_099_2170, w_099_2173, w_099_2180, w_099_2181, w_099_2183, w_099_2189, w_099_2194, w_099_2196, w_099_2197, w_099_2201, w_099_2203, w_099_2205, w_099_2212, w_099_2217, w_099_2222, w_099_2227, w_099_2229, w_099_2248, w_099_2249, w_099_2250, w_099_2259, w_099_2261, w_099_2263, w_099_2267, w_099_2268, w_099_2269, w_099_2270, w_099_2274, w_099_2282, w_099_2292, w_099_2297, w_099_2299, w_099_2300, w_099_2303, w_099_2308, w_099_2309, w_099_2310, w_099_2311, w_099_2313, w_099_2321, w_099_2322, w_099_2325, w_099_2329, w_099_2335, w_099_2337, w_099_2342, w_099_2343, w_099_2346, w_099_2353, w_099_2354, w_099_2359, w_099_2362, w_099_2364, w_099_2367, w_099_2370, w_099_2376, w_099_2384, w_099_2387, w_099_2388, w_099_2392, w_099_2396, w_099_2402, w_099_2407, w_099_2412, w_099_2413, w_099_2414, w_099_2417, w_099_2418, w_099_2421, w_099_2422, w_099_2427, w_099_2432, w_099_2434, w_099_2442, w_099_2447, w_099_2450, w_099_2452, w_099_2456, w_099_2457, w_099_2458, w_099_2459, w_099_2468, w_099_2469, w_099_2476, w_099_2478, w_099_2480, w_099_2482, w_099_2483, w_099_2484, w_099_2485, w_099_2490, w_099_2492, w_099_2496, w_099_2497, w_099_2498, w_099_2505, w_099_2508, w_099_2509, w_099_2510, w_099_2512, w_099_2516, w_099_2519, w_099_2522, w_099_2523, w_099_2526, w_099_2531, w_099_2533, w_099_2545, w_099_2547, w_099_2552, w_099_2553, w_099_2555, w_099_2556, w_099_2557, w_099_2566, w_099_2569, w_099_2571, w_099_2573, w_099_2581, w_099_2582, w_099_2583, w_099_2587, w_099_2589, w_099_2590, w_099_2591, w_099_2595, w_099_2596, w_099_2597, w_099_2598, w_099_2599, w_099_2600, w_099_2601, w_099_2602, w_099_2612, w_099_2613, w_099_2614, w_099_2622, w_099_2626, w_099_2631, w_099_2633, w_099_2636, w_099_2638, w_099_2640, w_099_2644, w_099_2645, w_099_2648, w_099_2649, w_099_2657, w_099_2663, w_099_2670, w_099_2674, w_099_2679, w_099_2682, w_099_2683, w_099_2684, w_099_2685, w_099_2688, w_099_2693, w_099_2699, w_099_2702, w_099_2705, w_099_2709, w_099_2718, w_099_2720, w_099_2723, w_099_2728, w_099_2733, w_099_2734, w_099_2736, w_099_2737, w_099_2739, w_099_2742, w_099_2745, w_099_2750, w_099_2752, w_099_2758, w_099_2759, w_099_2764, w_099_2770, w_099_2774, w_099_2775, w_099_2780, w_099_2788, w_099_2789, w_099_2792, w_099_2794, w_099_2805, w_099_2809, w_099_2811, w_099_2821, w_099_2822, w_099_2827, w_099_2828, w_099_2840, w_099_2842, w_099_2843, w_099_2844, w_099_2845, w_099_2846, w_099_2847, w_099_2849, w_099_2850, w_099_2858, w_099_2859, w_099_2861, w_099_2862, w_099_2863, w_099_2864, w_099_2865, w_099_2866, w_099_2868, w_099_2872, w_099_2876, w_099_2879, w_099_2880, w_099_2881, w_099_2883, w_099_2885, w_099_2889, w_099_2904, w_099_2907, w_099_2908, w_099_2917, w_099_2925, w_099_2926, w_099_2927, w_099_2928, w_099_2932, w_099_2936, w_099_2938, w_099_2940, w_099_2944, w_099_2955, w_099_2960, w_099_2961, w_099_2964, w_099_2968, w_099_2970, w_099_2974, w_099_2975, w_099_2978, w_099_2982, w_099_2986, w_099_2988, w_099_2990, w_099_2991, w_099_2992, w_099_2994, w_099_2997, w_099_3002, w_099_3007, w_099_3008, w_099_3015, w_099_3016, w_099_3017, w_099_3022, w_099_3026, w_099_3027, w_099_3031, w_099_3039, w_099_3041, w_099_3043, w_099_3044, w_099_3048, w_099_3054, w_099_3058, w_099_3060, w_099_3061, w_099_3066, w_099_3070, w_099_3074, w_099_3075, w_099_3078, w_099_3084, w_099_3086, w_099_3088, w_099_3089, w_099_3097, w_099_3100, w_099_3101, w_099_3106, w_099_3111, w_099_3112, w_099_3116, w_099_3122, w_099_3123, w_099_3124, w_099_3126, w_099_3131, w_099_3132, w_099_3149, w_099_3155, w_099_3159, w_099_3160, w_099_3163, w_099_3171, w_099_3177, w_099_3179, w_099_3181, w_099_3185, w_099_3186, w_099_3188, w_099_3193, w_099_3194, w_099_3198, w_099_3199, w_099_3208, w_099_3214, w_099_3224, w_099_3225, w_099_3236, w_099_3239, w_099_3242, w_099_3246, w_099_3257, w_099_3262, w_099_3265, w_099_3269, w_099_3271, w_099_3272, w_099_3275, w_099_3276, w_099_3278, w_099_3282, w_099_3285, w_099_3288, w_099_3289, w_099_3292, w_099_3298, w_099_3301, w_099_3304, w_099_3308, w_099_3309, w_099_3313, w_099_3322, w_099_3325, w_099_3326, w_099_3329, w_099_3334, w_099_3339, w_099_3341, w_099_3345, w_099_3346, w_099_3351, w_099_3356, w_099_3357, w_099_3360, w_099_3362, w_099_3366, w_099_3368, w_099_3373, w_099_3374, w_099_3377, w_099_3389, w_099_3390, w_099_3392, w_099_3393, w_099_3395, w_099_3396, w_099_3399, w_099_3404, w_099_3410, w_099_3411, w_099_3413, w_099_3414, w_099_3420, w_099_3421, w_099_3422, w_099_3427, w_099_3428, w_099_3429, w_099_3432, w_099_3433, w_099_3435, w_099_3436, w_099_3440, w_099_3441, w_099_3442, w_099_3443, w_099_3444, w_099_3446, w_099_3449, w_099_3452, w_099_3454, w_099_3465, w_099_3467, w_099_3474, w_099_3478, w_099_3479, w_099_3482, w_099_3485, w_099_3489, w_099_3490, w_099_3491, w_099_3495, w_099_3500, w_099_3502, w_099_3504, w_099_3505, w_099_3509, w_099_3510, w_099_3511, w_099_3512, w_099_3515, w_099_3518, w_099_3520, w_099_3529, w_099_3533, w_099_3544, w_099_3546, w_099_3548, w_099_3549, w_099_3552, w_099_3554, w_099_3555, w_099_3556, w_099_3567, w_099_3575, w_099_3576, w_099_3579, w_099_3585, w_099_3587, w_099_3589, w_099_3590, w_099_3594, w_099_3599, w_099_3605, w_099_3606, w_099_3611, w_099_3613, w_099_3623, w_099_3624, w_099_3625, w_099_3627, w_099_3632, w_099_3635, w_099_3637, w_099_3641, w_099_3653, w_099_3654, w_099_3657, w_099_3658, w_099_3659, w_099_3660, w_099_3661, w_099_3662, w_099_3663, w_099_3666, w_099_3669, w_099_3675, w_099_3685, w_099_3688, w_099_3695, w_099_3701, w_099_3702, w_099_3705, w_099_3708, w_099_3709, w_099_3711, w_099_3712, w_099_3714, w_099_3716, w_099_3722, w_099_3732, w_099_3734, w_099_3750, w_099_3751, w_099_3765, w_099_3769, w_099_3779, w_099_3787, w_099_3788, w_099_3789, w_099_3790, w_099_3793, w_099_3802, w_099_3804, w_099_3811, w_099_3812, w_099_3821, w_099_3827, w_099_3828, w_099_3829, w_099_3838, w_099_3845, w_099_3848, w_099_3861, w_099_3862, w_099_3864, w_099_3867, w_099_3868, w_099_3871, w_099_3873, w_099_3874, w_099_3883, w_099_3885, w_099_3889, w_099_3893, w_099_3896, w_099_3899, w_099_3900, w_099_3904, w_099_3913, w_099_3915, w_099_3919, w_099_3923, w_099_3928, w_099_3929, w_099_3933, w_099_3935, w_099_3939, w_099_3941, w_099_3945, w_099_3949, w_099_3954, w_099_3956, w_099_3957, w_099_3960, w_099_3964, w_099_3970, w_099_3974, w_099_3975, w_099_3979, w_099_3980, w_099_3982, w_099_3986, w_099_3987, w_099_3995, w_099_3999, w_099_4001, w_099_4004, w_099_4007, w_099_4009, w_099_4010, w_099_4012, w_099_4015, w_099_4017, w_099_4018, w_099_4020, w_099_4025, w_099_4027, w_099_4029, w_099_4032, w_099_4042, w_099_4044, w_099_4051, w_099_4053, w_099_4054, w_099_4056, w_099_4057, w_099_4062, w_099_4065, w_099_4066, w_099_4073, w_099_4077, w_099_4080, w_099_4082, w_099_4083, w_099_4091, w_099_4094, w_099_4096, w_099_4097, w_099_4104, w_099_4107, w_099_4109, w_099_4115, w_099_4118, w_099_4119, w_099_4122, w_099_4126, w_099_4134, w_099_4144, w_099_4147, w_099_4148, w_099_4150, w_099_4153, w_099_4154, w_099_4160, w_099_4163, w_099_4166, w_099_4167, w_099_4171, w_099_4176, w_099_4179, w_099_4186, w_099_4187, w_099_4194, w_099_4200, w_099_4202, w_099_4206, w_099_4212, w_099_4215, w_099_4217, w_099_4235, w_099_4242, w_099_4248, w_099_4249, w_099_4251, w_099_4253, w_099_4255, w_099_4256, w_099_4257, w_099_4260, w_099_4263, w_099_4265, w_099_4266, w_099_4274;
  wire w_100_000, w_100_001, w_100_002, w_100_007, w_100_008, w_100_010, w_100_011, w_100_013, w_100_016, w_100_017, w_100_025, w_100_026, w_100_027, w_100_031, w_100_032, w_100_034, w_100_035, w_100_036, w_100_037, w_100_039, w_100_040, w_100_041, w_100_044, w_100_047, w_100_052, w_100_056, w_100_057, w_100_061, w_100_063, w_100_065, w_100_066, w_100_068, w_100_069, w_100_071, w_100_072, w_100_077, w_100_080, w_100_081, w_100_082, w_100_084, w_100_086, w_100_089, w_100_090, w_100_092, w_100_094, w_100_097, w_100_098, w_100_099, w_100_102, w_100_103, w_100_105, w_100_107, w_100_108, w_100_109, w_100_110, w_100_112, w_100_113, w_100_115, w_100_117, w_100_118, w_100_120, w_100_121, w_100_123, w_100_124, w_100_125, w_100_134, w_100_136, w_100_137, w_100_139, w_100_140, w_100_145, w_100_146, w_100_147, w_100_148, w_100_149, w_100_150, w_100_154, w_100_156, w_100_157, w_100_159, w_100_162, w_100_165, w_100_169, w_100_170, w_100_171, w_100_172, w_100_174, w_100_175, w_100_176, w_100_177, w_100_178, w_100_183, w_100_184, w_100_186, w_100_190, w_100_192, w_100_193, w_100_195, w_100_196, w_100_197, w_100_200, w_100_201, w_100_202, w_100_203, w_100_204, w_100_206, w_100_208, w_100_211, w_100_219, w_100_221, w_100_222, w_100_225, w_100_227, w_100_231, w_100_232, w_100_233, w_100_238, w_100_245, w_100_247, w_100_251, w_100_258, w_100_259, w_100_261, w_100_262, w_100_263, w_100_265, w_100_266, w_100_267, w_100_269, w_100_271, w_100_278, w_100_282, w_100_284, w_100_285, w_100_286, w_100_287, w_100_289, w_100_291, w_100_296, w_100_297, w_100_303, w_100_305, w_100_306, w_100_307, w_100_309, w_100_310, w_100_311, w_100_313, w_100_314, w_100_315, w_100_318, w_100_320, w_100_323, w_100_324, w_100_325, w_100_326, w_100_327, w_100_328, w_100_333, w_100_334, w_100_335, w_100_341, w_100_343, w_100_347, w_100_349, w_100_350, w_100_352, w_100_353, w_100_355, w_100_356, w_100_358, w_100_359, w_100_360, w_100_361, w_100_363, w_100_364, w_100_365, w_100_366, w_100_367, w_100_368, w_100_369, w_100_371, w_100_373, w_100_374, w_100_378, w_100_380, w_100_383, w_100_387, w_100_389, w_100_391, w_100_392, w_100_394, w_100_397, w_100_403, w_100_406, w_100_408, w_100_409, w_100_411, w_100_413, w_100_414, w_100_415, w_100_416, w_100_419, w_100_423, w_100_424, w_100_426, w_100_430, w_100_435, w_100_437, w_100_439, w_100_440, w_100_443, w_100_444, w_100_448, w_100_449, w_100_450, w_100_452, w_100_456, w_100_457, w_100_458, w_100_459, w_100_461, w_100_462, w_100_463, w_100_464, w_100_468, w_100_471, w_100_472, w_100_474, w_100_475, w_100_476, w_100_478, w_100_482, w_100_484, w_100_488, w_100_489, w_100_492, w_100_500, w_100_501, w_100_502, w_100_503, w_100_505, w_100_508, w_100_513, w_100_516, w_100_517, w_100_518, w_100_519, w_100_521, w_100_524, w_100_530, w_100_531, w_100_533, w_100_536, w_100_538, w_100_540, w_100_544, w_100_546, w_100_547, w_100_553, w_100_560, w_100_564, w_100_565, w_100_568, w_100_569, w_100_574, w_100_576, w_100_577, w_100_582, w_100_583, w_100_589, w_100_590, w_100_596, w_100_597, w_100_599, w_100_602, w_100_603, w_100_607, w_100_609, w_100_610, w_100_611, w_100_613, w_100_614, w_100_616, w_100_617, w_100_618, w_100_620, w_100_622, w_100_623, w_100_628, w_100_629, w_100_631, w_100_632, w_100_637, w_100_638, w_100_640, w_100_643, w_100_647, w_100_648, w_100_650, w_100_654, w_100_655, w_100_656, w_100_658, w_100_660, w_100_661, w_100_662, w_100_663, w_100_665, w_100_667, w_100_672, w_100_674, w_100_676, w_100_679, w_100_681, w_100_682, w_100_683, w_100_685, w_100_690, w_100_692, w_100_694, w_100_702, w_100_703, w_100_705, w_100_706, w_100_708, w_100_710, w_100_711, w_100_712, w_100_713, w_100_718, w_100_720, w_100_722, w_100_723, w_100_726, w_100_730, w_100_734, w_100_740, w_100_744, w_100_746, w_100_747, w_100_748, w_100_749, w_100_752, w_100_754, w_100_756, w_100_758, w_100_761, w_100_762, w_100_764, w_100_766, w_100_767, w_100_768, w_100_769, w_100_776, w_100_780, w_100_781, w_100_783, w_100_784, w_100_785, w_100_786, w_100_787, w_100_789, w_100_791, w_100_793, w_100_795, w_100_796, w_100_797, w_100_798, w_100_799, w_100_800, w_100_802, w_100_803, w_100_805, w_100_806, w_100_808, w_100_810, w_100_811, w_100_814, w_100_815, w_100_816, w_100_819, w_100_824, w_100_827, w_100_828, w_100_830, w_100_832, w_100_833, w_100_834, w_100_836, w_100_838, w_100_840, w_100_841, w_100_842, w_100_843, w_100_844, w_100_847, w_100_848, w_100_849, w_100_851, w_100_852, w_100_854, w_100_855, w_100_857, w_100_858, w_100_859, w_100_861, w_100_862, w_100_863, w_100_865, w_100_867, w_100_868, w_100_870, w_100_871, w_100_872, w_100_874, w_100_875, w_100_876, w_100_877, w_100_878, w_100_879, w_100_883, w_100_886, w_100_889, w_100_891, w_100_893, w_100_896, w_100_897, w_100_900, w_100_901, w_100_902, w_100_903, w_100_904, w_100_906, w_100_907, w_100_910, w_100_912, w_100_913, w_100_915, w_100_916, w_100_920, w_100_923, w_100_927, w_100_928, w_100_930, w_100_931, w_100_933, w_100_937, w_100_941, w_100_942, w_100_945, w_100_949, w_100_952, w_100_955, w_100_956, w_100_957, w_100_962, w_100_963, w_100_965, w_100_967, w_100_968, w_100_969, w_100_970, w_100_971, w_100_973, w_100_976, w_100_977, w_100_978, w_100_980, w_100_981, w_100_982, w_100_983, w_100_984, w_100_987, w_100_989, w_100_990, w_100_991, w_100_992, w_100_993, w_100_995, w_100_996, w_100_997, w_100_999, w_100_1000, w_100_1001, w_100_1002, w_100_1005, w_100_1006, w_100_1008, w_100_1010, w_100_1012, w_100_1014, w_100_1016, w_100_1017, w_100_1020, w_100_1022, w_100_1023, w_100_1024, w_100_1028, w_100_1029, w_100_1030, w_100_1034, w_100_1035, w_100_1037, w_100_1038, w_100_1039, w_100_1040, w_100_1043, w_100_1044, w_100_1045, w_100_1046, w_100_1047, w_100_1048, w_100_1053, w_100_1056, w_100_1058, w_100_1059, w_100_1060, w_100_1062, w_100_1064, w_100_1065, w_100_1067, w_100_1068, w_100_1071, w_100_1072, w_100_1073, w_100_1075, w_100_1076, w_100_1077, w_100_1079, w_100_1082, w_100_1083, w_100_1088, w_100_1090, w_100_1091, w_100_1092, w_100_1093, w_100_1095, w_100_1096, w_100_1097, w_100_1099, w_100_1103, w_100_1105, w_100_1106, w_100_1108, w_100_1110, w_100_1112, w_100_1118, w_100_1121, w_100_1126, w_100_1128, w_100_1131, w_100_1132, w_100_1134, w_100_1135, w_100_1138, w_100_1141, w_100_1143, w_100_1144, w_100_1148, w_100_1150, w_100_1152, w_100_1153, w_100_1155, w_100_1156, w_100_1159, w_100_1163, w_100_1164, w_100_1166, w_100_1170, w_100_1171, w_100_1173, w_100_1174, w_100_1176, w_100_1177, w_100_1178, w_100_1181, w_100_1182, w_100_1192, w_100_1194, w_100_1200, w_100_1208, w_100_1210, w_100_1212, w_100_1215, w_100_1220, w_100_1224, w_100_1227, w_100_1228, w_100_1231, w_100_1236, w_100_1249, w_100_1251, w_100_1254, w_100_1255, w_100_1256, w_100_1259, w_100_1263, w_100_1265, w_100_1269, w_100_1271, w_100_1272, w_100_1279, w_100_1285, w_100_1293, w_100_1295, w_100_1296, w_100_1297, w_100_1298, w_100_1299, w_100_1301, w_100_1308, w_100_1309, w_100_1310, w_100_1313, w_100_1316, w_100_1319, w_100_1323, w_100_1326, w_100_1327, w_100_1328, w_100_1337, w_100_1338, w_100_1340, w_100_1342, w_100_1344, w_100_1346, w_100_1349, w_100_1351, w_100_1352, w_100_1354, w_100_1355, w_100_1358, w_100_1360, w_100_1362, w_100_1371, w_100_1374, w_100_1376, w_100_1379, w_100_1383, w_100_1388, w_100_1390, w_100_1395, w_100_1396, w_100_1398, w_100_1399, w_100_1402, w_100_1403, w_100_1404, w_100_1412, w_100_1417, w_100_1421, w_100_1431, w_100_1439, w_100_1441, w_100_1448, w_100_1453, w_100_1458, w_100_1461, w_100_1463, w_100_1470, w_100_1477, w_100_1483, w_100_1488, w_100_1489, w_100_1490, w_100_1495, w_100_1496, w_100_1497, w_100_1510, w_100_1511, w_100_1512, w_100_1517, w_100_1519, w_100_1520, w_100_1521, w_100_1522, w_100_1528, w_100_1538, w_100_1539, w_100_1541, w_100_1545, w_100_1549, w_100_1555, w_100_1557, w_100_1561, w_100_1562, w_100_1567, w_100_1579, w_100_1581, w_100_1585, w_100_1588, w_100_1590, w_100_1594, w_100_1611, w_100_1614, w_100_1615, w_100_1617, w_100_1618, w_100_1621, w_100_1626, w_100_1631, w_100_1633, w_100_1635, w_100_1638, w_100_1642, w_100_1643, w_100_1645, w_100_1647, w_100_1648, w_100_1651, w_100_1665, w_100_1670, w_100_1676, w_100_1679, w_100_1685, w_100_1691, w_100_1692, w_100_1693, w_100_1694, w_100_1697, w_100_1702, w_100_1709, w_100_1712, w_100_1713, w_100_1716, w_100_1725, w_100_1729, w_100_1736, w_100_1739, w_100_1740, w_100_1742, w_100_1744, w_100_1745, w_100_1747, w_100_1751, w_100_1755, w_100_1756, w_100_1758, w_100_1759, w_100_1760, w_100_1761, w_100_1763, w_100_1764, w_100_1765, w_100_1769, w_100_1773, w_100_1776, w_100_1782, w_100_1785, w_100_1794, w_100_1796, w_100_1797, w_100_1803, w_100_1804, w_100_1805, w_100_1806, w_100_1810, w_100_1817, w_100_1819, w_100_1824, w_100_1828, w_100_1829, w_100_1830, w_100_1831, w_100_1835, w_100_1838, w_100_1840, w_100_1842, w_100_1843, w_100_1844, w_100_1846, w_100_1850, w_100_1853, w_100_1855, w_100_1856, w_100_1860, w_100_1863, w_100_1864, w_100_1866, w_100_1871, w_100_1883, w_100_1884, w_100_1897, w_100_1899, w_100_1906, w_100_1908, w_100_1910, w_100_1917, w_100_1918, w_100_1920, w_100_1930, w_100_1934, w_100_1936, w_100_1937, w_100_1944, w_100_1946, w_100_1953, w_100_1956, w_100_1961, w_100_1963, w_100_1964, w_100_1965, w_100_1968, w_100_1970, w_100_1978, w_100_1986, w_100_1988, w_100_1991, w_100_1995, w_100_1996, w_100_2002, w_100_2008, w_100_2012, w_100_2016, w_100_2019, w_100_2024, w_100_2025, w_100_2034, w_100_2036, w_100_2040, w_100_2041, w_100_2042, w_100_2043, w_100_2044, w_100_2046, w_100_2056, w_100_2057, w_100_2065, w_100_2068, w_100_2069, w_100_2071, w_100_2074, w_100_2078, w_100_2080, w_100_2083, w_100_2090, w_100_2093, w_100_2102, w_100_2104, w_100_2106, w_100_2109, w_100_2110, w_100_2117, w_100_2120, w_100_2121, w_100_2123, w_100_2126, w_100_2130, w_100_2134, w_100_2136, w_100_2137, w_100_2138, w_100_2140, w_100_2145, w_100_2147, w_100_2149, w_100_2156, w_100_2159, w_100_2161, w_100_2162, w_100_2164, w_100_2166, w_100_2168, w_100_2172, w_100_2175, w_100_2176, w_100_2185, w_100_2186, w_100_2193, w_100_2197, w_100_2198, w_100_2200, w_100_2202, w_100_2210, w_100_2213, w_100_2215, w_100_2217, w_100_2219, w_100_2225, w_100_2227, w_100_2233, w_100_2239, w_100_2244, w_100_2248, w_100_2251, w_100_2252, w_100_2256, w_100_2258, w_100_2259, w_100_2265, w_100_2273, w_100_2275, w_100_2277, w_100_2289, w_100_2290, w_100_2292, w_100_2299, w_100_2300, w_100_2301, w_100_2302, w_100_2306, w_100_2309, w_100_2320, w_100_2321, w_100_2324, w_100_2325, w_100_2326, w_100_2333, w_100_2341, w_100_2351, w_100_2364, w_100_2367, w_100_2369, w_100_2385, w_100_2387, w_100_2388, w_100_2392, w_100_2394, w_100_2396, w_100_2398, w_100_2405, w_100_2411, w_100_2413, w_100_2420, w_100_2430, w_100_2432, w_100_2433, w_100_2434, w_100_2444, w_100_2453, w_100_2454, w_100_2455, w_100_2457, w_100_2463, w_100_2469, w_100_2475, w_100_2477, w_100_2479, w_100_2488, w_100_2492, w_100_2497, w_100_2502, w_100_2505, w_100_2508, w_100_2510, w_100_2511, w_100_2513, w_100_2514, w_100_2515, w_100_2518, w_100_2520, w_100_2521, w_100_2531, w_100_2532, w_100_2535, w_100_2536, w_100_2537, w_100_2539, w_100_2543, w_100_2553, w_100_2556, w_100_2558, w_100_2561, w_100_2562, w_100_2565, w_100_2566, w_100_2570, w_100_2574, w_100_2581, w_100_2583, w_100_2588, w_100_2597, w_100_2598, w_100_2599, w_100_2600, w_100_2601, w_100_2602, w_100_2603, w_100_2611, w_100_2613, w_100_2615, w_100_2618, w_100_2622, w_100_2624, w_100_2625, w_100_2629, w_100_2631, w_100_2632, w_100_2633, w_100_2635, w_100_2642, w_100_2644, w_100_2647, w_100_2648, w_100_2649, w_100_2652, w_100_2654, w_100_2667, w_100_2668, w_100_2683, w_100_2685, w_100_2697, w_100_2710, w_100_2717, w_100_2721, w_100_2722, w_100_2723, w_100_2725, w_100_2727, w_100_2728, w_100_2730, w_100_2735, w_100_2737, w_100_2738, w_100_2739, w_100_2741, w_100_2742, w_100_2743, w_100_2747, w_100_2753, w_100_2766, w_100_2767, w_100_2771, w_100_2779, w_100_2784, w_100_2787, w_100_2792, w_100_2797, w_100_2802, w_100_2803, w_100_2812, w_100_2815, w_100_2816, w_100_2818, w_100_2821, w_100_2827, w_100_2830, w_100_2832, w_100_2834, w_100_2840, w_100_2843, w_100_2849, w_100_2856, w_100_2857, w_100_2858, w_100_2860, w_100_2861, w_100_2863, w_100_2864, w_100_2865, w_100_2872, w_100_2873, w_100_2889, w_100_2904, w_100_2906, w_100_2907, w_100_2913, w_100_2914, w_100_2923, w_100_2924, w_100_2925, w_100_2927, w_100_2928, w_100_2929, w_100_2938, w_100_2939, w_100_2940, w_100_2945, w_100_2946, w_100_2949, w_100_2960, w_100_2963, w_100_2971, w_100_2975, w_100_2978, w_100_2980, w_100_2984, w_100_2986, w_100_2989, w_100_2992, w_100_3002, w_100_3003, w_100_3005, w_100_3006, w_100_3016, w_100_3022, w_100_3023, w_100_3034, w_100_3038, w_100_3041, w_100_3045, w_100_3046, w_100_3047, w_100_3049, w_100_3051, w_100_3054, w_100_3057, w_100_3062, w_100_3065, w_100_3067, w_100_3068, w_100_3070, w_100_3072, w_100_3079, w_100_3085, w_100_3086, w_100_3091, w_100_3094, w_100_3101, w_100_3102, w_100_3105, w_100_3108, w_100_3111, w_100_3114, w_100_3117, w_100_3123, w_100_3128, w_100_3133, w_100_3138, w_100_3147, w_100_3148, w_100_3150, w_100_3151, w_100_3156, w_100_3160, w_100_3162, w_100_3163, w_100_3165, w_100_3166, w_100_3169, w_100_3174, w_100_3188, w_100_3193, w_100_3201, w_100_3203, w_100_3208, w_100_3211, w_100_3215, w_100_3216, w_100_3217, w_100_3219, w_100_3221, w_100_3222, w_100_3231, w_100_3232, w_100_3240, w_100_3241, w_100_3242, w_100_3243, w_100_3246, w_100_3250, w_100_3251, w_100_3253, w_100_3255, w_100_3258, w_100_3259, w_100_3260, w_100_3261, w_100_3274, w_100_3278, w_100_3281, w_100_3297, w_100_3301, w_100_3307, w_100_3310, w_100_3312, w_100_3318, w_100_3319, w_100_3320, w_100_3335, w_100_3340, w_100_3344, w_100_3352, w_100_3355, w_100_3357, w_100_3359, w_100_3364, w_100_3365, w_100_3366, w_100_3370, w_100_3372, w_100_3380, w_100_3381, w_100_3382, w_100_3384, w_100_3391, w_100_3393, w_100_3395, w_100_3403, w_100_3406, w_100_3407, w_100_3409, w_100_3412, w_100_3419, w_100_3420, w_100_3428, w_100_3430, w_100_3432, w_100_3433, w_100_3437, w_100_3444, w_100_3446, w_100_3449, w_100_3450, w_100_3464, w_100_3467, w_100_3473, w_100_3477, w_100_3478, w_100_3482, w_100_3484, w_100_3486, w_100_3488, w_100_3491, w_100_3494, w_100_3497, w_100_3498, w_100_3511, w_100_3516, w_100_3517, w_100_3519, w_100_3521, w_100_3528, w_100_3535, w_100_3536, w_100_3537, w_100_3538, w_100_3539, w_100_3545, w_100_3547, w_100_3550, w_100_3555, w_100_3556, w_100_3561, w_100_3562, w_100_3565, w_100_3567, w_100_3568, w_100_3570, w_100_3580, w_100_3582, w_100_3585, w_100_3588, w_100_3591, w_100_3595, w_100_3598, w_100_3600, w_100_3612, w_100_3613, w_100_3624, w_100_3629, w_100_3636, w_100_3637, w_100_3639, w_100_3647, w_100_3649, w_100_3651, w_100_3654, w_100_3657, w_100_3661, w_100_3665, w_100_3666, w_100_3671, w_100_3675, w_100_3677, w_100_3685, w_100_3689, w_100_3700, w_100_3706, w_100_3708, w_100_3713, w_100_3714, w_100_3718, w_100_3722, w_100_3730, w_100_3740, w_100_3746, w_100_3749, w_100_3758, w_100_3759, w_100_3762, w_100_3764, w_100_3772, w_100_3780, w_100_3783, w_100_3788, w_100_3789, w_100_3798, w_100_3805, w_100_3806, w_100_3810, w_100_3812, w_100_3815, w_100_3816, w_100_3817, w_100_3820, w_100_3821, w_100_3822, w_100_3823, w_100_3824, w_100_3825, w_100_3826, w_100_3827, w_100_3828, w_100_3829, w_100_3830, w_100_3832;
  wire w_101_000, w_101_001, w_101_002, w_101_003, w_101_007, w_101_009, w_101_011, w_101_012, w_101_014, w_101_016, w_101_017, w_101_018, w_101_019, w_101_020, w_101_021, w_101_027, w_101_028, w_101_029, w_101_030, w_101_031, w_101_032, w_101_033, w_101_038, w_101_041, w_101_044, w_101_048, w_101_049, w_101_050, w_101_054, w_101_055, w_101_056, w_101_057, w_101_059, w_101_061, w_101_062, w_101_065, w_101_067, w_101_068, w_101_071, w_101_074, w_101_078, w_101_080, w_101_084, w_101_086, w_101_087, w_101_089, w_101_092, w_101_093, w_101_096, w_101_098, w_101_100, w_101_101, w_101_105, w_101_106, w_101_107, w_101_112, w_101_113, w_101_115, w_101_116, w_101_121, w_101_122, w_101_124, w_101_125, w_101_130, w_101_132, w_101_134, w_101_138, w_101_142, w_101_143, w_101_144, w_101_145, w_101_150, w_101_151, w_101_153, w_101_159, w_101_163, w_101_165, w_101_166, w_101_168, w_101_171, w_101_176, w_101_183, w_101_188, w_101_190, w_101_191, w_101_192, w_101_193, w_101_196, w_101_198, w_101_199, w_101_204, w_101_205, w_101_206, w_101_207, w_101_210, w_101_211, w_101_212, w_101_213, w_101_215, w_101_216, w_101_217, w_101_219, w_101_221, w_101_223, w_101_226, w_101_227, w_101_229, w_101_231, w_101_232, w_101_233, w_101_234, w_101_235, w_101_236, w_101_240, w_101_243, w_101_244, w_101_250, w_101_251, w_101_252, w_101_254, w_101_255, w_101_256, w_101_258, w_101_259, w_101_260, w_101_262, w_101_264, w_101_267, w_101_268, w_101_270, w_101_273, w_101_274, w_101_275, w_101_278, w_101_279, w_101_281, w_101_283, w_101_284, w_101_285, w_101_287, w_101_289, w_101_290, w_101_291, w_101_292, w_101_293, w_101_295, w_101_297, w_101_299, w_101_300, w_101_301, w_101_302, w_101_303, w_101_304, w_101_306, w_101_308, w_101_310, w_101_312, w_101_313, w_101_314, w_101_316, w_101_319, w_101_322, w_101_323, w_101_325, w_101_326, w_101_327, w_101_328, w_101_329, w_101_331, w_101_332, w_101_334, w_101_336, w_101_337, w_101_339, w_101_341, w_101_343, w_101_344, w_101_345, w_101_347, w_101_349, w_101_351, w_101_352, w_101_353, w_101_354, w_101_355, w_101_363, w_101_364, w_101_365, w_101_367, w_101_374, w_101_380, w_101_381, w_101_383, w_101_384, w_101_385, w_101_389, w_101_392, w_101_393, w_101_394, w_101_397, w_101_398, w_101_399, w_101_403, w_101_406, w_101_408, w_101_410, w_101_412, w_101_413, w_101_414, w_101_421, w_101_422, w_101_424, w_101_425, w_101_428, w_101_430, w_101_432, w_101_434, w_101_435, w_101_438, w_101_439, w_101_440, w_101_443, w_101_444, w_101_447, w_101_448, w_101_450, w_101_452, w_101_454, w_101_455, w_101_456, w_101_458, w_101_461, w_101_462, w_101_466, w_101_467, w_101_469, w_101_473, w_101_474, w_101_478, w_101_479, w_101_483, w_101_484, w_101_486, w_101_487, w_101_488, w_101_489, w_101_491, w_101_492, w_101_493, w_101_494, w_101_503, w_101_504, w_101_505, w_101_506, w_101_508, w_101_509, w_101_510, w_101_513, w_101_517, w_101_518, w_101_520, w_101_521, w_101_522, w_101_523, w_101_525, w_101_527, w_101_529, w_101_530, w_101_534, w_101_537, w_101_538, w_101_539, w_101_540, w_101_544, w_101_547, w_101_548, w_101_550, w_101_552, w_101_555, w_101_557, w_101_558, w_101_559, w_101_561, w_101_566, w_101_568, w_101_570, w_101_571, w_101_572, w_101_575, w_101_578, w_101_581, w_101_582, w_101_583, w_101_584, w_101_586, w_101_587, w_101_589, w_101_592, w_101_594, w_101_595, w_101_597, w_101_602, w_101_603, w_101_606, w_101_607, w_101_612, w_101_613, w_101_616, w_101_617, w_101_618, w_101_620, w_101_624, w_101_625, w_101_627, w_101_628, w_101_631, w_101_632, w_101_633, w_101_636, w_101_637, w_101_638, w_101_642, w_101_643, w_101_645, w_101_649, w_101_650, w_101_651, w_101_652, w_101_655, w_101_656, w_101_658, w_101_661, w_101_666, w_101_668, w_101_671, w_101_672, w_101_673, w_101_674, w_101_675, w_101_676, w_101_680, w_101_685, w_101_687, w_101_690, w_101_698, w_101_699, w_101_702, w_101_705, w_101_707, w_101_710, w_101_715, w_101_716, w_101_720, w_101_721, w_101_722, w_101_723, w_101_725, w_101_727, w_101_731, w_101_734, w_101_738, w_101_739, w_101_744, w_101_746, w_101_752, w_101_753, w_101_757, w_101_758, w_101_760, w_101_761, w_101_762, w_101_767, w_101_769, w_101_770, w_101_772, w_101_774, w_101_776, w_101_778, w_101_782, w_101_784, w_101_786, w_101_787, w_101_788, w_101_791, w_101_792, w_101_794, w_101_795, w_101_801, w_101_806, w_101_807, w_101_811, w_101_812, w_101_814, w_101_816, w_101_818, w_101_819, w_101_820, w_101_823, w_101_824, w_101_825, w_101_827, w_101_828, w_101_831, w_101_833, w_101_834, w_101_839, w_101_841, w_101_844, w_101_847, w_101_848, w_101_851, w_101_852, w_101_855, w_101_856, w_101_859, w_101_860, w_101_867, w_101_871, w_101_873, w_101_874, w_101_876, w_101_883, w_101_886, w_101_888, w_101_890, w_101_892, w_101_893, w_101_895, w_101_898, w_101_899, w_101_902, w_101_903, w_101_906, w_101_910, w_101_914, w_101_915, w_101_917, w_101_919, w_101_920, w_101_924, w_101_925, w_101_926, w_101_930, w_101_931, w_101_934, w_101_935, w_101_937, w_101_938, w_101_939, w_101_940, w_101_951, w_101_952, w_101_953, w_101_954, w_101_956, w_101_957, w_101_958, w_101_959, w_101_962, w_101_963, w_101_969, w_101_970, w_101_972, w_101_974, w_101_980, w_101_981, w_101_985, w_101_992, w_101_995, w_101_1000, w_101_1002, w_101_1003, w_101_1004, w_101_1007, w_101_1008, w_101_1010, w_101_1011, w_101_1013, w_101_1016, w_101_1017, w_101_1020, w_101_1023, w_101_1026, w_101_1028, w_101_1030, w_101_1032, w_101_1033, w_101_1034, w_101_1037, w_101_1040, w_101_1042, w_101_1043, w_101_1045, w_101_1051, w_101_1052, w_101_1054, w_101_1060, w_101_1062, w_101_1064, w_101_1069, w_101_1070, w_101_1073, w_101_1077, w_101_1078, w_101_1085, w_101_1086, w_101_1088, w_101_1089, w_101_1091, w_101_1092, w_101_1099, w_101_1105, w_101_1107, w_101_1111, w_101_1113, w_101_1117, w_101_1118, w_101_1119, w_101_1120, w_101_1121, w_101_1124, w_101_1125, w_101_1127, w_101_1129, w_101_1130, w_101_1132, w_101_1134, w_101_1137, w_101_1146, w_101_1147, w_101_1148, w_101_1151, w_101_1158, w_101_1163, w_101_1164, w_101_1166, w_101_1167, w_101_1168, w_101_1169, w_101_1173, w_101_1174, w_101_1175, w_101_1176, w_101_1177, w_101_1179, w_101_1181, w_101_1184, w_101_1185, w_101_1196, w_101_1197, w_101_1199, w_101_1201, w_101_1205, w_101_1206, w_101_1207, w_101_1211, w_101_1214, w_101_1219, w_101_1221, w_101_1224, w_101_1226, w_101_1229, w_101_1230, w_101_1231, w_101_1232, w_101_1234, w_101_1240, w_101_1241, w_101_1242, w_101_1244, w_101_1245, w_101_1248, w_101_1250, w_101_1252, w_101_1253, w_101_1254, w_101_1256, w_101_1258, w_101_1259, w_101_1264, w_101_1266, w_101_1268, w_101_1274, w_101_1275, w_101_1279, w_101_1283, w_101_1288, w_101_1290, w_101_1291, w_101_1293, w_101_1296, w_101_1298, w_101_1301, w_101_1302, w_101_1305, w_101_1308, w_101_1312, w_101_1313, w_101_1314, w_101_1316, w_101_1319, w_101_1322, w_101_1324, w_101_1325, w_101_1326, w_101_1327, w_101_1328, w_101_1330, w_101_1331, w_101_1332, w_101_1334, w_101_1336, w_101_1341, w_101_1342, w_101_1343, w_101_1345, w_101_1349, w_101_1350, w_101_1354, w_101_1356, w_101_1358, w_101_1365, w_101_1368, w_101_1369, w_101_1372, w_101_1373, w_101_1375, w_101_1376, w_101_1377, w_101_1379, w_101_1380, w_101_1385, w_101_1387, w_101_1389, w_101_1391, w_101_1393, w_101_1394, w_101_1397, w_101_1411, w_101_1415, w_101_1416, w_101_1417, w_101_1420, w_101_1424, w_101_1428, w_101_1433, w_101_1443, w_101_1447, w_101_1451, w_101_1453, w_101_1458, w_101_1470, w_101_1471, w_101_1474, w_101_1478, w_101_1480, w_101_1482, w_101_1496, w_101_1497, w_101_1500, w_101_1502, w_101_1504, w_101_1505, w_101_1518, w_101_1520, w_101_1521, w_101_1524, w_101_1530, w_101_1534, w_101_1535, w_101_1544, w_101_1550, w_101_1551, w_101_1554, w_101_1555, w_101_1556, w_101_1558, w_101_1559, w_101_1561, w_101_1562, w_101_1564, w_101_1576, w_101_1578, w_101_1580, w_101_1581, w_101_1583, w_101_1588, w_101_1591, w_101_1593, w_101_1595, w_101_1599, w_101_1605, w_101_1613, w_101_1623, w_101_1624, w_101_1625, w_101_1631, w_101_1632, w_101_1633, w_101_1641, w_101_1642, w_101_1645, w_101_1652, w_101_1653, w_101_1658, w_101_1661, w_101_1668, w_101_1669, w_101_1671, w_101_1674, w_101_1678, w_101_1679, w_101_1681, w_101_1697, w_101_1698, w_101_1703, w_101_1707, w_101_1708, w_101_1718, w_101_1720, w_101_1721, w_101_1723, w_101_1724, w_101_1729, w_101_1735, w_101_1739, w_101_1752, w_101_1753, w_101_1756, w_101_1765, w_101_1768, w_101_1769, w_101_1770, w_101_1774, w_101_1776, w_101_1778, w_101_1780, w_101_1781, w_101_1783, w_101_1784, w_101_1789, w_101_1793, w_101_1794, w_101_1805, w_101_1817, w_101_1825, w_101_1828, w_101_1829, w_101_1831, w_101_1836, w_101_1838, w_101_1847, w_101_1849, w_101_1853, w_101_1856, w_101_1857, w_101_1860, w_101_1861, w_101_1865, w_101_1879, w_101_1883, w_101_1884, w_101_1885, w_101_1886, w_101_1889, w_101_1890, w_101_1901, w_101_1909, w_101_1910, w_101_1914, w_101_1915, w_101_1922, w_101_1930, w_101_1939, w_101_1949, w_101_1956, w_101_1963, w_101_1965, w_101_1968, w_101_1970, w_101_1971, w_101_1972, w_101_1980, w_101_1984, w_101_1986, w_101_1987, w_101_1988, w_101_1992, w_101_1994, w_101_1996, w_101_2000, w_101_2001, w_101_2003, w_101_2006, w_101_2010, w_101_2013, w_101_2019, w_101_2020, w_101_2024, w_101_2035, w_101_2039, w_101_2040, w_101_2049, w_101_2051, w_101_2062, w_101_2063, w_101_2066, w_101_2068, w_101_2069, w_101_2071, w_101_2075, w_101_2080, w_101_2081, w_101_2083, w_101_2086, w_101_2087, w_101_2090, w_101_2092, w_101_2098, w_101_2099, w_101_2100, w_101_2104, w_101_2106, w_101_2108, w_101_2109, w_101_2112, w_101_2114, w_101_2126, w_101_2128, w_101_2129, w_101_2130, w_101_2131, w_101_2146, w_101_2151, w_101_2152, w_101_2159, w_101_2161, w_101_2167, w_101_2179, w_101_2188, w_101_2192, w_101_2193, w_101_2195, w_101_2199, w_101_2204, w_101_2211, w_101_2213, w_101_2226, w_101_2236, w_101_2238, w_101_2242, w_101_2244, w_101_2245, w_101_2246, w_101_2247, w_101_2251, w_101_2252, w_101_2254, w_101_2255, w_101_2256, w_101_2260, w_101_2261, w_101_2263, w_101_2266, w_101_2269, w_101_2271, w_101_2275, w_101_2276, w_101_2282, w_101_2283, w_101_2293, w_101_2295, w_101_2301, w_101_2304, w_101_2306, w_101_2309, w_101_2315, w_101_2316, w_101_2322, w_101_2326, w_101_2335, w_101_2346, w_101_2349, w_101_2351, w_101_2357, w_101_2359, w_101_2360, w_101_2362, w_101_2364, w_101_2365, w_101_2368, w_101_2375, w_101_2378, w_101_2387, w_101_2393, w_101_2395, w_101_2396, w_101_2397, w_101_2401, w_101_2404, w_101_2415, w_101_2417, w_101_2419, w_101_2421, w_101_2422, w_101_2424, w_101_2426, w_101_2430, w_101_2432, w_101_2434, w_101_2436, w_101_2439, w_101_2449, w_101_2452, w_101_2453, w_101_2454, w_101_2463, w_101_2469, w_101_2473, w_101_2485, w_101_2487, w_101_2489, w_101_2491, w_101_2495, w_101_2497, w_101_2500, w_101_2502, w_101_2506, w_101_2511, w_101_2513, w_101_2519, w_101_2522, w_101_2524, w_101_2525, w_101_2534, w_101_2536, w_101_2537, w_101_2541, w_101_2558, w_101_2560, w_101_2562, w_101_2570, w_101_2571, w_101_2577, w_101_2588, w_101_2592, w_101_2598, w_101_2601, w_101_2610, w_101_2615, w_101_2616, w_101_2621, w_101_2623, w_101_2636, w_101_2643, w_101_2645, w_101_2648, w_101_2650, w_101_2653, w_101_2656, w_101_2659, w_101_2660, w_101_2668, w_101_2676, w_101_2677, w_101_2678, w_101_2683, w_101_2684, w_101_2686, w_101_2689, w_101_2692, w_101_2695, w_101_2698, w_101_2706, w_101_2708, w_101_2721, w_101_2722, w_101_2726, w_101_2729, w_101_2730, w_101_2731, w_101_2737, w_101_2739, w_101_2747, w_101_2757, w_101_2758, w_101_2760, w_101_2763, w_101_2765, w_101_2767, w_101_2775, w_101_2783, w_101_2788, w_101_2791, w_101_2795, w_101_2796, w_101_2797, w_101_2798, w_101_2800, w_101_2804, w_101_2806, w_101_2809, w_101_2812, w_101_2818, w_101_2821, w_101_2826, w_101_2827, w_101_2829, w_101_2830, w_101_2832, w_101_2841, w_101_2844, w_101_2845, w_101_2846, w_101_2849, w_101_2859, w_101_2860, w_101_2865, w_101_2868, w_101_2882, w_101_2890, w_101_2894, w_101_2897, w_101_2903, w_101_2904, w_101_2906, w_101_2907, w_101_2908, w_101_2914, w_101_2923, w_101_2924, w_101_2926, w_101_2933, w_101_2935, w_101_2937, w_101_2938, w_101_2939, w_101_2940, w_101_2948, w_101_2953, w_101_2960, w_101_2963, w_101_2964, w_101_2968, w_101_2973, w_101_2975, w_101_2982, w_101_2985, w_101_2986, w_101_2988, w_101_2993, w_101_2996, w_101_3002, w_101_3006, w_101_3008, w_101_3016, w_101_3018, w_101_3021, w_101_3024, w_101_3030, w_101_3035, w_101_3036, w_101_3037, w_101_3040, w_101_3042, w_101_3048, w_101_3049, w_101_3053, w_101_3055, w_101_3056, w_101_3057, w_101_3059, w_101_3065, w_101_3066, w_101_3067, w_101_3072, w_101_3073, w_101_3076, w_101_3079, w_101_3082, w_101_3089, w_101_3095, w_101_3098, w_101_3101, w_101_3102, w_101_3108, w_101_3111, w_101_3124, w_101_3126, w_101_3127, w_101_3134, w_101_3135, w_101_3141, w_101_3156, w_101_3160, w_101_3168, w_101_3176, w_101_3179, w_101_3187, w_101_3188, w_101_3189, w_101_3193, w_101_3201, w_101_3203, w_101_3209, w_101_3214, w_101_3216, w_101_3225, w_101_3228, w_101_3231, w_101_3239, w_101_3245, w_101_3246, w_101_3249, w_101_3251, w_101_3252, w_101_3257, w_101_3260, w_101_3261, w_101_3264, w_101_3265, w_101_3287, w_101_3291, w_101_3294, w_101_3298, w_101_3299, w_101_3301, w_101_3308, w_101_3311, w_101_3313, w_101_3321, w_101_3324, w_101_3326, w_101_3329, w_101_3334, w_101_3335, w_101_3340, w_101_3343, w_101_3345, w_101_3347, w_101_3348, w_101_3349, w_101_3353, w_101_3355, w_101_3356, w_101_3357, w_101_3358, w_101_3359, w_101_3364, w_101_3365, w_101_3368, w_101_3369, w_101_3370, w_101_3376, w_101_3379, w_101_3381, w_101_3382, w_101_3383, w_101_3392, w_101_3393, w_101_3396, w_101_3397, w_101_3404, w_101_3406, w_101_3409, w_101_3411, w_101_3415, w_101_3417, w_101_3421, w_101_3426, w_101_3443, w_101_3445, w_101_3446, w_101_3460, w_101_3463, w_101_3465, w_101_3466, w_101_3468, w_101_3476, w_101_3481, w_101_3483, w_101_3486, w_101_3487, w_101_3490, w_101_3492, w_101_3501, w_101_3505, w_101_3507, w_101_3509, w_101_3513, w_101_3518, w_101_3519, w_101_3522, w_101_3523, w_101_3536, w_101_3538, w_101_3542, w_101_3549, w_101_3552, w_101_3553, w_101_3556, w_101_3561, w_101_3563, w_101_3570, w_101_3571, w_101_3574, w_101_3577, w_101_3578, w_101_3582, w_101_3590, w_101_3592, w_101_3594, w_101_3595;
  wire w_102_003, w_102_004, w_102_005, w_102_009, w_102_011, w_102_013, w_102_014, w_102_017, w_102_020, w_102_021, w_102_024, w_102_025, w_102_028, w_102_029, w_102_030, w_102_032, w_102_033, w_102_036, w_102_040, w_102_044, w_102_047, w_102_048, w_102_053, w_102_054, w_102_055, w_102_056, w_102_060, w_102_063, w_102_064, w_102_066, w_102_068, w_102_071, w_102_074, w_102_075, w_102_076, w_102_078, w_102_081, w_102_083, w_102_086, w_102_087, w_102_088, w_102_089, w_102_091, w_102_092, w_102_093, w_102_096, w_102_097, w_102_098, w_102_099, w_102_100, w_102_101, w_102_103, w_102_104, w_102_106, w_102_109, w_102_111, w_102_112, w_102_114, w_102_115, w_102_116, w_102_119, w_102_120, w_102_123, w_102_124, w_102_127, w_102_128, w_102_131, w_102_133, w_102_136, w_102_139, w_102_144, w_102_146, w_102_148, w_102_149, w_102_154, w_102_158, w_102_161, w_102_162, w_102_164, w_102_166, w_102_168, w_102_170, w_102_173, w_102_175, w_102_176, w_102_179, w_102_186, w_102_189, w_102_194, w_102_195, w_102_199, w_102_203, w_102_208, w_102_213, w_102_216, w_102_217, w_102_219, w_102_220, w_102_222, w_102_224, w_102_225, w_102_226, w_102_229, w_102_230, w_102_232, w_102_235, w_102_242, w_102_244, w_102_245, w_102_246, w_102_247, w_102_250, w_102_251, w_102_252, w_102_254, w_102_255, w_102_256, w_102_258, w_102_259, w_102_263, w_102_267, w_102_270, w_102_274, w_102_275, w_102_277, w_102_280, w_102_283, w_102_284, w_102_290, w_102_292, w_102_293, w_102_298, w_102_299, w_102_300, w_102_301, w_102_303, w_102_305, w_102_306, w_102_308, w_102_309, w_102_313, w_102_316, w_102_317, w_102_321, w_102_324, w_102_325, w_102_326, w_102_330, w_102_332, w_102_337, w_102_338, w_102_339, w_102_341, w_102_344, w_102_346, w_102_348, w_102_349, w_102_350, w_102_352, w_102_356, w_102_359, w_102_363, w_102_364, w_102_365, w_102_374, w_102_378, w_102_379, w_102_380, w_102_382, w_102_383, w_102_384, w_102_388, w_102_390, w_102_391, w_102_393, w_102_395, w_102_396, w_102_398, w_102_399, w_102_403, w_102_405, w_102_408, w_102_409, w_102_411, w_102_413, w_102_414, w_102_416, w_102_418, w_102_419, w_102_420, w_102_421, w_102_422, w_102_427, w_102_431, w_102_432, w_102_433, w_102_435, w_102_436, w_102_438, w_102_439, w_102_440, w_102_441, w_102_442, w_102_443, w_102_446, w_102_447, w_102_451, w_102_452, w_102_453, w_102_457, w_102_458, w_102_460, w_102_461, w_102_462, w_102_466, w_102_467, w_102_471, w_102_472, w_102_473, w_102_474, w_102_475, w_102_476, w_102_478, w_102_480, w_102_488, w_102_489, w_102_491, w_102_492, w_102_494, w_102_496, w_102_497, w_102_500, w_102_502, w_102_503, w_102_504, w_102_505, w_102_506, w_102_507, w_102_508, w_102_514, w_102_515, w_102_518, w_102_520, w_102_521, w_102_524, w_102_528, w_102_530, w_102_533, w_102_539, w_102_541, w_102_545, w_102_547, w_102_548, w_102_550, w_102_551, w_102_555, w_102_556, w_102_557, w_102_558, w_102_562, w_102_565, w_102_566, w_102_577, w_102_581, w_102_595, w_102_599, w_102_600, w_102_601, w_102_608, w_102_611, w_102_615, w_102_622, w_102_623, w_102_628, w_102_630, w_102_631, w_102_634, w_102_635, w_102_637, w_102_642, w_102_647, w_102_651, w_102_658, w_102_659, w_102_660, w_102_661, w_102_662, w_102_663, w_102_666, w_102_674, w_102_675, w_102_680, w_102_684, w_102_686, w_102_687, w_102_689, w_102_691, w_102_693, w_102_695, w_102_697, w_102_698, w_102_703, w_102_704, w_102_708, w_102_709, w_102_710, w_102_721, w_102_724, w_102_728, w_102_729, w_102_732, w_102_734, w_102_735, w_102_739, w_102_741, w_102_743, w_102_744, w_102_746, w_102_750, w_102_752, w_102_753, w_102_755, w_102_764, w_102_773, w_102_774, w_102_775, w_102_778, w_102_783, w_102_786, w_102_788, w_102_796, w_102_802, w_102_803, w_102_805, w_102_809, w_102_810, w_102_813, w_102_824, w_102_828, w_102_830, w_102_833, w_102_848, w_102_849, w_102_853, w_102_854, w_102_855, w_102_868, w_102_870, w_102_871, w_102_880, w_102_881, w_102_885, w_102_888, w_102_889, w_102_892, w_102_895, w_102_909, w_102_917, w_102_918, w_102_921, w_102_924, w_102_925, w_102_929, w_102_930, w_102_949, w_102_954, w_102_957, w_102_961, w_102_964, w_102_965, w_102_968, w_102_978, w_102_979, w_102_990, w_102_993, w_102_994, w_102_1012, w_102_1013, w_102_1022, w_102_1027, w_102_1028, w_102_1029, w_102_1031, w_102_1032, w_102_1033, w_102_1039, w_102_1043, w_102_1044, w_102_1046, w_102_1048, w_102_1050, w_102_1053, w_102_1073, w_102_1074, w_102_1076, w_102_1078, w_102_1081, w_102_1085, w_102_1090, w_102_1091, w_102_1093, w_102_1098, w_102_1099, w_102_1101, w_102_1106, w_102_1114, w_102_1119, w_102_1120, w_102_1123, w_102_1127, w_102_1135, w_102_1139, w_102_1140, w_102_1145, w_102_1148, w_102_1149, w_102_1150, w_102_1152, w_102_1154, w_102_1155, w_102_1157, w_102_1158, w_102_1166, w_102_1174, w_102_1177, w_102_1182, w_102_1184, w_102_1187, w_102_1188, w_102_1192, w_102_1204, w_102_1206, w_102_1207, w_102_1209, w_102_1216, w_102_1219, w_102_1221, w_102_1223, w_102_1227, w_102_1239, w_102_1241, w_102_1242, w_102_1247, w_102_1256, w_102_1260, w_102_1261, w_102_1262, w_102_1271, w_102_1274, w_102_1277, w_102_1279, w_102_1280, w_102_1283, w_102_1284, w_102_1285, w_102_1287, w_102_1288, w_102_1292, w_102_1298, w_102_1306, w_102_1308, w_102_1311, w_102_1313, w_102_1315, w_102_1320, w_102_1324, w_102_1326, w_102_1332, w_102_1335, w_102_1340, w_102_1342, w_102_1344, w_102_1348, w_102_1349, w_102_1353, w_102_1355, w_102_1358, w_102_1359, w_102_1365, w_102_1371, w_102_1373, w_102_1374, w_102_1377, w_102_1378, w_102_1391, w_102_1394, w_102_1397, w_102_1399, w_102_1400, w_102_1410, w_102_1415, w_102_1417, w_102_1418, w_102_1424, w_102_1425, w_102_1426, w_102_1427, w_102_1428, w_102_1434, w_102_1436, w_102_1443, w_102_1451, w_102_1453, w_102_1457, w_102_1459, w_102_1467, w_102_1468, w_102_1469, w_102_1470, w_102_1477, w_102_1478, w_102_1481, w_102_1483, w_102_1488, w_102_1490, w_102_1493, w_102_1497, w_102_1498, w_102_1499, w_102_1505, w_102_1507, w_102_1522, w_102_1524, w_102_1525, w_102_1530, w_102_1536, w_102_1539, w_102_1544, w_102_1549, w_102_1560, w_102_1568, w_102_1569, w_102_1570, w_102_1577, w_102_1584, w_102_1586, w_102_1590, w_102_1591, w_102_1592, w_102_1599, w_102_1602, w_102_1605, w_102_1607, w_102_1608, w_102_1610, w_102_1618, w_102_1621, w_102_1622, w_102_1623, w_102_1625, w_102_1626, w_102_1629, w_102_1631, w_102_1635, w_102_1643, w_102_1644, w_102_1650, w_102_1668, w_102_1669, w_102_1671, w_102_1672, w_102_1677, w_102_1680, w_102_1684, w_102_1694, w_102_1696, w_102_1697, w_102_1702, w_102_1706, w_102_1707, w_102_1709, w_102_1717, w_102_1720, w_102_1721, w_102_1725, w_102_1730, w_102_1733, w_102_1734, w_102_1735, w_102_1744, w_102_1747, w_102_1748, w_102_1756, w_102_1760, w_102_1764, w_102_1767, w_102_1774, w_102_1780, w_102_1781, w_102_1783, w_102_1786, w_102_1790, w_102_1792, w_102_1793, w_102_1796, w_102_1797, w_102_1799, w_102_1803, w_102_1806, w_102_1809, w_102_1812, w_102_1823, w_102_1824, w_102_1834, w_102_1840, w_102_1846, w_102_1853, w_102_1856, w_102_1857, w_102_1861, w_102_1864, w_102_1869, w_102_1871, w_102_1872, w_102_1873, w_102_1880, w_102_1884, w_102_1885, w_102_1888, w_102_1890, w_102_1893, w_102_1894, w_102_1897, w_102_1898, w_102_1911, w_102_1914, w_102_1928, w_102_1929, w_102_1931, w_102_1934, w_102_1939, w_102_1941, w_102_1949, w_102_1952, w_102_1953, w_102_1955, w_102_1963, w_102_1967, w_102_1969, w_102_1970, w_102_1974, w_102_1978, w_102_1985, w_102_1988, w_102_1994, w_102_1995, w_102_1999, w_102_2002, w_102_2005, w_102_2006, w_102_2012, w_102_2013, w_102_2024, w_102_2026, w_102_2029, w_102_2033, w_102_2037, w_102_2042, w_102_2045, w_102_2053, w_102_2055, w_102_2056, w_102_2059, w_102_2063, w_102_2071, w_102_2074, w_102_2078, w_102_2080, w_102_2081, w_102_2082, w_102_2087, w_102_2088, w_102_2091, w_102_2095, w_102_2100, w_102_2103, w_102_2107, w_102_2114, w_102_2118, w_102_2134, w_102_2137, w_102_2139, w_102_2141, w_102_2144, w_102_2157, w_102_2159, w_102_2166, w_102_2167, w_102_2171, w_102_2183, w_102_2187, w_102_2190, w_102_2192, w_102_2201, w_102_2202, w_102_2205, w_102_2206, w_102_2207, w_102_2211, w_102_2213, w_102_2216, w_102_2220, w_102_2226, w_102_2230, w_102_2233, w_102_2241, w_102_2246, w_102_2252, w_102_2256, w_102_2257, w_102_2258, w_102_2259, w_102_2261, w_102_2267, w_102_2268, w_102_2274, w_102_2275, w_102_2276, w_102_2278, w_102_2279, w_102_2281, w_102_2282, w_102_2283, w_102_2285, w_102_2286, w_102_2292, w_102_2297, w_102_2298, w_102_2299, w_102_2300, w_102_2302, w_102_2306, w_102_2308, w_102_2311, w_102_2314, w_102_2316, w_102_2319, w_102_2320, w_102_2324, w_102_2325, w_102_2334, w_102_2335, w_102_2340, w_102_2343, w_102_2345, w_102_2347, w_102_2353, w_102_2357, w_102_2361, w_102_2362, w_102_2366, w_102_2367, w_102_2370, w_102_2374, w_102_2376, w_102_2381, w_102_2383, w_102_2388, w_102_2390, w_102_2391, w_102_2399, w_102_2406, w_102_2411, w_102_2413, w_102_2414, w_102_2415, w_102_2417, w_102_2420, w_102_2433, w_102_2435, w_102_2437, w_102_2444, w_102_2448, w_102_2453, w_102_2454, w_102_2460, w_102_2462, w_102_2463, w_102_2466, w_102_2471, w_102_2473, w_102_2485, w_102_2486, w_102_2489, w_102_2492, w_102_2493, w_102_2499, w_102_2503, w_102_2507, w_102_2513, w_102_2514, w_102_2519, w_102_2520, w_102_2521, w_102_2522, w_102_2527, w_102_2528, w_102_2530, w_102_2540, w_102_2548, w_102_2549, w_102_2553, w_102_2564, w_102_2577, w_102_2580, w_102_2581, w_102_2582, w_102_2586, w_102_2594, w_102_2595, w_102_2600, w_102_2603, w_102_2605, w_102_2613, w_102_2615, w_102_2616, w_102_2618, w_102_2620, w_102_2631, w_102_2635, w_102_2637, w_102_2647, w_102_2657, w_102_2658, w_102_2659, w_102_2674, w_102_2675, w_102_2676, w_102_2680, w_102_2689, w_102_2690, w_102_2695, w_102_2699, w_102_2702, w_102_2703, w_102_2707, w_102_2708, w_102_2710, w_102_2719, w_102_2731, w_102_2735, w_102_2738, w_102_2747, w_102_2749, w_102_2753, w_102_2756, w_102_2757, w_102_2758, w_102_2759, w_102_2762, w_102_2772, w_102_2779, w_102_2781, w_102_2783, w_102_2794, w_102_2799, w_102_2801, w_102_2810, w_102_2811, w_102_2812, w_102_2816, w_102_2821, w_102_2822, w_102_2823, w_102_2830, w_102_2834, w_102_2839, w_102_2840, w_102_2841, w_102_2847, w_102_2849, w_102_2860, w_102_2864, w_102_2865, w_102_2872, w_102_2876, w_102_2879, w_102_2882, w_102_2884, w_102_2887, w_102_2890, w_102_2897, w_102_2900, w_102_2901, w_102_2903, w_102_2905, w_102_2906, w_102_2912, w_102_2915, w_102_2917, w_102_2918, w_102_2921, w_102_2924, w_102_2928, w_102_2934, w_102_2944, w_102_2957, w_102_2962, w_102_2965, w_102_2966, w_102_2971, w_102_2975, w_102_2976, w_102_2990, w_102_2992, w_102_2993, w_102_2995, w_102_2999, w_102_3008, w_102_3011, w_102_3014, w_102_3019, w_102_3020, w_102_3023, w_102_3029, w_102_3030, w_102_3032, w_102_3035, w_102_3037, w_102_3041, w_102_3046, w_102_3047, w_102_3048, w_102_3051, w_102_3056, w_102_3061, w_102_3062, w_102_3068, w_102_3071, w_102_3072, w_102_3079, w_102_3080, w_102_3084, w_102_3086, w_102_3087, w_102_3089, w_102_3098, w_102_3107, w_102_3108, w_102_3109, w_102_3123, w_102_3124, w_102_3125, w_102_3133, w_102_3134, w_102_3137, w_102_3138, w_102_3146, w_102_3147, w_102_3153, w_102_3154, w_102_3157, w_102_3161, w_102_3163, w_102_3168, w_102_3171, w_102_3175, w_102_3177, w_102_3178, w_102_3179, w_102_3181, w_102_3182, w_102_3183, w_102_3188, w_102_3189, w_102_3197, w_102_3201, w_102_3203, w_102_3205, w_102_3209, w_102_3210, w_102_3213, w_102_3214, w_102_3215, w_102_3218, w_102_3220, w_102_3224, w_102_3229, w_102_3241, w_102_3242, w_102_3244, w_102_3246, w_102_3256, w_102_3260, w_102_3262, w_102_3263, w_102_3274, w_102_3278, w_102_3281, w_102_3286, w_102_3293, w_102_3296, w_102_3297, w_102_3302, w_102_3307, w_102_3313, w_102_3318, w_102_3321, w_102_3325, w_102_3327, w_102_3328, w_102_3330, w_102_3335, w_102_3336, w_102_3337, w_102_3341, w_102_3342, w_102_3347, w_102_3349, w_102_3355, w_102_3359, w_102_3361, w_102_3366, w_102_3371, w_102_3374, w_102_3377, w_102_3378, w_102_3379, w_102_3385, w_102_3388, w_102_3397, w_102_3406, w_102_3413, w_102_3417, w_102_3419, w_102_3424, w_102_3426, w_102_3431, w_102_3434, w_102_3436, w_102_3437, w_102_3439, w_102_3440, w_102_3443, w_102_3446, w_102_3448, w_102_3451, w_102_3455, w_102_3457, w_102_3458, w_102_3461, w_102_3465, w_102_3466, w_102_3471, w_102_3477, w_102_3482, w_102_3486, w_102_3487, w_102_3488, w_102_3496, w_102_3503, w_102_3510, w_102_3517, w_102_3522, w_102_3523, w_102_3524, w_102_3527, w_102_3530, w_102_3531, w_102_3532, w_102_3535, w_102_3541, w_102_3542, w_102_3546, w_102_3548, w_102_3551, w_102_3556, w_102_3557, w_102_3559, w_102_3561, w_102_3564, w_102_3565, w_102_3569, w_102_3571, w_102_3579, w_102_3580, w_102_3582, w_102_3585, w_102_3586, w_102_3588, w_102_3590, w_102_3592, w_102_3599, w_102_3600, w_102_3603, w_102_3607, w_102_3609, w_102_3614, w_102_3620, w_102_3630, w_102_3632, w_102_3636, w_102_3640, w_102_3641, w_102_3642, w_102_3647, w_102_3648, w_102_3649, w_102_3650, w_102_3657, w_102_3659, w_102_3664, w_102_3670, w_102_3678, w_102_3680, w_102_3683, w_102_3686, w_102_3699, w_102_3704, w_102_3709, w_102_3711, w_102_3712, w_102_3715, w_102_3719, w_102_3721, w_102_3726, w_102_3731, w_102_3735, w_102_3753, w_102_3754, w_102_3755, w_102_3756, w_102_3759, w_102_3770, w_102_3772, w_102_3775, w_102_3778, w_102_3785, w_102_3787, w_102_3789, w_102_3791, w_102_3794, w_102_3798, w_102_3809, w_102_3814, w_102_3818, w_102_3819, w_102_3821, w_102_3830, w_102_3834, w_102_3836, w_102_3841, w_102_3850, w_102_3858, w_102_3859, w_102_3860, w_102_3862, w_102_3870, w_102_3875, w_102_3876, w_102_3878, w_102_3882, w_102_3883, w_102_3885, w_102_3889, w_102_3895, w_102_3899, w_102_3900, w_102_3902, w_102_3903, w_102_3904, w_102_3910, w_102_3914, w_102_3915, w_102_3916, w_102_3917, w_102_3918, w_102_3926, w_102_3930, w_102_3932, w_102_3936, w_102_3937, w_102_3944, w_102_3946, w_102_3949, w_102_3952, w_102_3955, w_102_3958, w_102_3964, w_102_3968, w_102_3969, w_102_3971, w_102_3972, w_102_3974, w_102_3982, w_102_3983, w_102_3988, w_102_3994, w_102_3996, w_102_3999, w_102_4001, w_102_4004, w_102_4008, w_102_4009, w_102_4017, w_102_4018, w_102_4022, w_102_4026, w_102_4032, w_102_4038, w_102_4041, w_102_4046, w_102_4047, w_102_4055, w_102_4056, w_102_4061, w_102_4070, w_102_4071, w_102_4072, w_102_4074, w_102_4076, w_102_4077, w_102_4080, w_102_4085, w_102_4089, w_102_4095, w_102_4108, w_102_4111, w_102_4113, w_102_4118, w_102_4122, w_102_4126, w_102_4131, w_102_4133, w_102_4135, w_102_4138, w_102_4147, w_102_4148, w_102_4149, w_102_4156, w_102_4158, w_102_4162, w_102_4164, w_102_4170, w_102_4174, w_102_4175, w_102_4181, w_102_4182, w_102_4184, w_102_4190, w_102_4195, w_102_4197, w_102_4199, w_102_4200, w_102_4204, w_102_4206, w_102_4208, w_102_4212, w_102_4229, w_102_4237, w_102_4238, w_102_4243, w_102_4248, w_102_4249, w_102_4251, w_102_4253, w_102_4257, w_102_4259, w_102_4263, w_102_4265, w_102_4268, w_102_4269, w_102_4276, w_102_4280, w_102_4281, w_102_4283, w_102_4285, w_102_4286, w_102_4287, w_102_4293, w_102_4295, w_102_4297, w_102_4299, w_102_4300, w_102_4311, w_102_4312, w_102_4314, w_102_4333, w_102_4336, w_102_4338, w_102_4339, w_102_4343, w_102_4344, w_102_4348, w_102_4350, w_102_4362, w_102_4365, w_102_4368, w_102_4373, w_102_4377, w_102_4380, w_102_4383, w_102_4387, w_102_4392, w_102_4393, w_102_4395, w_102_4402, w_102_4407, w_102_4409, w_102_4412, w_102_4417, w_102_4418, w_102_4421, w_102_4432;
  wire w_103_000, w_103_003, w_103_005, w_103_006, w_103_007, w_103_008, w_103_009, w_103_013, w_103_014, w_103_015, w_103_016, w_103_017, w_103_019, w_103_021, w_103_022, w_103_024, w_103_025, w_103_028, w_103_029, w_103_031, w_103_035, w_103_036, w_103_037, w_103_040, w_103_042, w_103_048, w_103_055, w_103_062, w_103_065, w_103_070, w_103_071, w_103_074, w_103_076, w_103_078, w_103_080, w_103_081, w_103_083, w_103_085, w_103_086, w_103_090, w_103_091, w_103_095, w_103_097, w_103_099, w_103_100, w_103_104, w_103_107, w_103_108, w_103_111, w_103_120, w_103_122, w_103_124, w_103_125, w_103_126, w_103_128, w_103_131, w_103_133, w_103_134, w_103_135, w_103_136, w_103_137, w_103_139, w_103_142, w_103_143, w_103_144, w_103_145, w_103_146, w_103_147, w_103_148, w_103_151, w_103_153, w_103_155, w_103_160, w_103_161, w_103_162, w_103_164, w_103_165, w_103_167, w_103_168, w_103_169, w_103_171, w_103_174, w_103_176, w_103_183, w_103_184, w_103_186, w_103_187, w_103_188, w_103_193, w_103_194, w_103_196, w_103_198, w_103_200, w_103_202, w_103_203, w_103_204, w_103_205, w_103_206, w_103_209, w_103_214, w_103_215, w_103_225, w_103_233, w_103_235, w_103_237, w_103_239, w_103_249, w_103_250, w_103_256, w_103_275, w_103_277, w_103_286, w_103_292, w_103_303, w_103_304, w_103_309, w_103_315, w_103_320, w_103_321, w_103_326, w_103_328, w_103_336, w_103_339, w_103_340, w_103_346, w_103_350, w_103_352, w_103_355, w_103_356, w_103_357, w_103_358, w_103_365, w_103_370, w_103_371, w_103_373, w_103_374, w_103_377, w_103_382, w_103_383, w_103_385, w_103_393, w_103_405, w_103_422, w_103_424, w_103_425, w_103_430, w_103_433, w_103_436, w_103_438, w_103_442, w_103_445, w_103_447, w_103_451, w_103_452, w_103_455, w_103_465, w_103_466, w_103_476, w_103_479, w_103_481, w_103_487, w_103_502, w_103_507, w_103_509, w_103_513, w_103_515, w_103_519, w_103_520, w_103_521, w_103_526, w_103_528, w_103_529, w_103_534, w_103_537, w_103_539, w_103_540, w_103_543, w_103_544, w_103_548, w_103_555, w_103_558, w_103_559, w_103_561, w_103_563, w_103_566, w_103_567, w_103_569, w_103_570, w_103_575, w_103_578, w_103_600, w_103_608, w_103_611, w_103_617, w_103_620, w_103_621, w_103_627, w_103_628, w_103_630, w_103_631, w_103_633, w_103_637, w_103_640, w_103_648, w_103_656, w_103_657, w_103_659, w_103_662, w_103_672, w_103_673, w_103_675, w_103_678, w_103_682, w_103_689, w_103_694, w_103_697, w_103_705, w_103_709, w_103_712, w_103_714, w_103_715, w_103_716, w_103_717, w_103_719, w_103_726, w_103_727, w_103_730, w_103_733, w_103_740, w_103_741, w_103_745, w_103_755, w_103_756, w_103_757, w_103_758, w_103_759, w_103_760, w_103_761, w_103_762, w_103_770, w_103_774, w_103_776, w_103_780, w_103_790, w_103_791, w_103_793, w_103_797, w_103_801, w_103_804, w_103_806, w_103_809, w_103_813, w_103_815, w_103_819, w_103_820, w_103_826, w_103_827, w_103_828, w_103_835, w_103_837, w_103_839, w_103_841, w_103_843, w_103_850, w_103_852, w_103_854, w_103_857, w_103_864, w_103_869, w_103_870, w_103_889, w_103_890, w_103_891, w_103_893, w_103_895, w_103_898, w_103_901, w_103_902, w_103_916, w_103_927, w_103_931, w_103_934, w_103_936, w_103_937, w_103_939, w_103_940, w_103_942, w_103_954, w_103_955, w_103_957, w_103_958, w_103_959, w_103_964, w_103_968, w_103_974, w_103_979, w_103_990, w_103_996, w_103_1006, w_103_1008, w_103_1015, w_103_1016, w_103_1017, w_103_1020, w_103_1024, w_103_1027, w_103_1032, w_103_1033, w_103_1034, w_103_1048, w_103_1055, w_103_1060, w_103_1064, w_103_1066, w_103_1068, w_103_1076, w_103_1088, w_103_1092, w_103_1103, w_103_1106, w_103_1114, w_103_1125, w_103_1131, w_103_1133, w_103_1139, w_103_1140, w_103_1142, w_103_1148, w_103_1149, w_103_1152, w_103_1159, w_103_1164, w_103_1170, w_103_1174, w_103_1179, w_103_1181, w_103_1188, w_103_1195, w_103_1201, w_103_1202, w_103_1216, w_103_1219, w_103_1221, w_103_1230, w_103_1236, w_103_1242, w_103_1249, w_103_1250, w_103_1253, w_103_1260, w_103_1261, w_103_1265, w_103_1269, w_103_1270, w_103_1273, w_103_1276, w_103_1282, w_103_1285, w_103_1295, w_103_1298, w_103_1299, w_103_1302, w_103_1303, w_103_1306, w_103_1309, w_103_1315, w_103_1316, w_103_1319, w_103_1320, w_103_1321, w_103_1323, w_103_1324, w_103_1325, w_103_1327, w_103_1329, w_103_1336, w_103_1337, w_103_1339, w_103_1348, w_103_1349, w_103_1354, w_103_1359, w_103_1367, w_103_1372, w_103_1374, w_103_1376, w_103_1379, w_103_1391, w_103_1395, w_103_1396, w_103_1397, w_103_1404, w_103_1405, w_103_1415, w_103_1417, w_103_1423, w_103_1425, w_103_1430, w_103_1438, w_103_1447, w_103_1452, w_103_1460, w_103_1469, w_103_1473, w_103_1475, w_103_1476, w_103_1479, w_103_1483, w_103_1484, w_103_1491, w_103_1496, w_103_1497, w_103_1506, w_103_1507, w_103_1509, w_103_1512, w_103_1513, w_103_1520, w_103_1522, w_103_1527, w_103_1531, w_103_1533, w_103_1535, w_103_1537, w_103_1543, w_103_1545, w_103_1551, w_103_1554, w_103_1555, w_103_1568, w_103_1571, w_103_1576, w_103_1578, w_103_1582, w_103_1584, w_103_1591, w_103_1592, w_103_1593, w_103_1599, w_103_1600, w_103_1601, w_103_1606, w_103_1612, w_103_1613, w_103_1615, w_103_1619, w_103_1625, w_103_1626, w_103_1629, w_103_1631, w_103_1632, w_103_1634, w_103_1643, w_103_1645, w_103_1647, w_103_1651, w_103_1653, w_103_1657, w_103_1660, w_103_1661, w_103_1663, w_103_1670, w_103_1673, w_103_1676, w_103_1692, w_103_1693, w_103_1694, w_103_1708, w_103_1713, w_103_1716, w_103_1718, w_103_1725, w_103_1729, w_103_1733, w_103_1737, w_103_1739, w_103_1741, w_103_1744, w_103_1745, w_103_1746, w_103_1748, w_103_1753, w_103_1754, w_103_1762, w_103_1764, w_103_1770, w_103_1771, w_103_1784, w_103_1786, w_103_1787, w_103_1791, w_103_1792, w_103_1795, w_103_1803, w_103_1805, w_103_1811, w_103_1813, w_103_1817, w_103_1819, w_103_1820, w_103_1821, w_103_1825, w_103_1830, w_103_1836, w_103_1839, w_103_1844, w_103_1845, w_103_1846, w_103_1848, w_103_1853, w_103_1856, w_103_1858, w_103_1864, w_103_1865, w_103_1868, w_103_1870, w_103_1873, w_103_1879, w_103_1881, w_103_1885, w_103_1889, w_103_1903, w_103_1904, w_103_1917, w_103_1922, w_103_1923, w_103_1926, w_103_1927, w_103_1934, w_103_1936, w_103_1940, w_103_1941, w_103_1949, w_103_1950, w_103_1951, w_103_1955, w_103_1963, w_103_1964, w_103_1968, w_103_1971, w_103_1972, w_103_1980, w_103_1990, w_103_1991, w_103_1993, w_103_1996, w_103_1999, w_103_2004, w_103_2012, w_103_2013, w_103_2014, w_103_2020, w_103_2023, w_103_2026, w_103_2027, w_103_2030, w_103_2031, w_103_2033, w_103_2035, w_103_2045, w_103_2054, w_103_2059, w_103_2061, w_103_2062, w_103_2063, w_103_2071, w_103_2073, w_103_2074, w_103_2075, w_103_2077, w_103_2084, w_103_2088, w_103_2093, w_103_2096, w_103_2097, w_103_2100, w_103_2106, w_103_2113, w_103_2114, w_103_2118, w_103_2123, w_103_2126, w_103_2127, w_103_2130, w_103_2134, w_103_2139, w_103_2145, w_103_2146, w_103_2151, w_103_2154, w_103_2156, w_103_2159, w_103_2162, w_103_2165, w_103_2168, w_103_2177, w_103_2179, w_103_2182, w_103_2183, w_103_2188, w_103_2191, w_103_2197, w_103_2199, w_103_2212, w_103_2215, w_103_2216, w_103_2221, w_103_2225, w_103_2233, w_103_2235, w_103_2238, w_103_2246, w_103_2255, w_103_2257, w_103_2259, w_103_2263, w_103_2267, w_103_2270, w_103_2279, w_103_2282, w_103_2286, w_103_2288, w_103_2290, w_103_2297, w_103_2304, w_103_2308, w_103_2313, w_103_2314, w_103_2317, w_103_2321, w_103_2322, w_103_2332, w_103_2337, w_103_2345, w_103_2348, w_103_2351, w_103_2355, w_103_2364, w_103_2366, w_103_2371, w_103_2372, w_103_2373, w_103_2374, w_103_2375, w_103_2376, w_103_2378, w_103_2380, w_103_2387, w_103_2390, w_103_2391, w_103_2393, w_103_2397, w_103_2400, w_103_2402, w_103_2407, w_103_2419, w_103_2423, w_103_2427, w_103_2428, w_103_2429, w_103_2432, w_103_2438, w_103_2444, w_103_2452, w_103_2453, w_103_2459, w_103_2465, w_103_2478, w_103_2481, w_103_2483, w_103_2487, w_103_2488, w_103_2489, w_103_2490, w_103_2501, w_103_2503, w_103_2505, w_103_2514, w_103_2515, w_103_2516, w_103_2519, w_103_2521, w_103_2522, w_103_2523, w_103_2526, w_103_2530, w_103_2531, w_103_2532, w_103_2539, w_103_2541, w_103_2542, w_103_2545, w_103_2547, w_103_2552, w_103_2558, w_103_2565, w_103_2567, w_103_2569, w_103_2589, w_103_2604, w_103_2609, w_103_2618, w_103_2620, w_103_2622, w_103_2624, w_103_2627, w_103_2631, w_103_2634, w_103_2635, w_103_2637, w_103_2638, w_103_2639, w_103_2640, w_103_2642, w_103_2647, w_103_2650, w_103_2653, w_103_2654, w_103_2662, w_103_2665, w_103_2666, w_103_2667, w_103_2669, w_103_2687, w_103_2689, w_103_2698, w_103_2705, w_103_2707, w_103_2722, w_103_2738, w_103_2739, w_103_2740, w_103_2742, w_103_2743, w_103_2745, w_103_2746, w_103_2752, w_103_2754, w_103_2759, w_103_2762, w_103_2765, w_103_2770, w_103_2771, w_103_2779, w_103_2783, w_103_2787, w_103_2788, w_103_2789, w_103_2791, w_103_2800, w_103_2803, w_103_2804, w_103_2805, w_103_2806, w_103_2814, w_103_2819, w_103_2826, w_103_2827, w_103_2828, w_103_2837, w_103_2840, w_103_2842, w_103_2843, w_103_2844, w_103_2854, w_103_2859, w_103_2861, w_103_2865, w_103_2866, w_103_2868, w_103_2871, w_103_2874, w_103_2875, w_103_2880, w_103_2884, w_103_2885, w_103_2888, w_103_2895, w_103_2897, w_103_2899, w_103_2901, w_103_2903, w_103_2904, w_103_2905, w_103_2907, w_103_2911, w_103_2916, w_103_2917, w_103_2926, w_103_2927, w_103_2929, w_103_2931, w_103_2937, w_103_2938, w_103_2948, w_103_2958, w_103_2962, w_103_2970, w_103_2977, w_103_2978, w_103_2986, w_103_2994, w_103_2995, w_103_2996, w_103_2997, w_103_3004, w_103_3011, w_103_3016, w_103_3018, w_103_3029, w_103_3035, w_103_3037, w_103_3041, w_103_3043, w_103_3050, w_103_3053, w_103_3054, w_103_3055, w_103_3058, w_103_3064, w_103_3066, w_103_3068, w_103_3069, w_103_3070, w_103_3073, w_103_3075, w_103_3076, w_103_3077, w_103_3078, w_103_3083, w_103_3090, w_103_3095, w_103_3098, w_103_3119, w_103_3129, w_103_3130, w_103_3132, w_103_3134, w_103_3137, w_103_3144, w_103_3150, w_103_3151, w_103_3154, w_103_3159, w_103_3166, w_103_3172, w_103_3174, w_103_3175, w_103_3179, w_103_3183, w_103_3186, w_103_3196, w_103_3198, w_103_3199, w_103_3200, w_103_3206, w_103_3207, w_103_3208, w_103_3209, w_103_3213, w_103_3219, w_103_3223, w_103_3224, w_103_3229, w_103_3230, w_103_3233, w_103_3251, w_103_3252, w_103_3253, w_103_3255, w_103_3260, w_103_3262, w_103_3268, w_103_3279, w_103_3282, w_103_3285, w_103_3286, w_103_3292, w_103_3300, w_103_3302, w_103_3307, w_103_3308, w_103_3312, w_103_3324, w_103_3326, w_103_3329, w_103_3331, w_103_3338, w_103_3341, w_103_3344, w_103_3349, w_103_3354, w_103_3359, w_103_3362, w_103_3363, w_103_3384, w_103_3386, w_103_3388, w_103_3395, w_103_3399, w_103_3405, w_103_3406, w_103_3407, w_103_3411, w_103_3412, w_103_3417, w_103_3419, w_103_3423, w_103_3434, w_103_3436, w_103_3439, w_103_3440, w_103_3442, w_103_3444, w_103_3447, w_103_3457, w_103_3467, w_103_3469, w_103_3470, w_103_3472, w_103_3479, w_103_3483, w_103_3486, w_103_3489, w_103_3491, w_103_3494, w_103_3497, w_103_3498, w_103_3500, w_103_3508, w_103_3509, w_103_3511, w_103_3512, w_103_3519, w_103_3525, w_103_3536, w_103_3544, w_103_3545, w_103_3548, w_103_3553, w_103_3555, w_103_3560, w_103_3563, w_103_3571, w_103_3573, w_103_3574, w_103_3575, w_103_3576, w_103_3581, w_103_3587, w_103_3592, w_103_3597, w_103_3598, w_103_3599, w_103_3601, w_103_3608, w_103_3609, w_103_3610, w_103_3612, w_103_3614, w_103_3616, w_103_3622, w_103_3624, w_103_3625, w_103_3627, w_103_3632, w_103_3635, w_103_3639, w_103_3640, w_103_3641, w_103_3644, w_103_3651, w_103_3657, w_103_3658, w_103_3660, w_103_3665, w_103_3666, w_103_3670, w_103_3673, w_103_3682, w_103_3687, w_103_3693, w_103_3695, w_103_3697, w_103_3698, w_103_3699, w_103_3700, w_103_3701, w_103_3702, w_103_3708, w_103_3710, w_103_3715, w_103_3723, w_103_3729, w_103_3731, w_103_3736, w_103_3738, w_103_3739, w_103_3740, w_103_3745, w_103_3746, w_103_3752, w_103_3753, w_103_3755, w_103_3765, w_103_3766, w_103_3768, w_103_3770, w_103_3771, w_103_3774, w_103_3775, w_103_3778, w_103_3781, w_103_3782, w_103_3785, w_103_3787, w_103_3790, w_103_3796, w_103_3799, w_103_3802, w_103_3804, w_103_3819, w_103_3821, w_103_3826, w_103_3828, w_103_3830, w_103_3834, w_103_3839, w_103_3849, w_103_3853, w_103_3857, w_103_3858, w_103_3860, w_103_3862, w_103_3864, w_103_3865, w_103_3877, w_103_3878, w_103_3888, w_103_3897, w_103_3898, w_103_3904, w_103_3909, w_103_3910, w_103_3917, w_103_3919, w_103_3922, w_103_3925, w_103_3942, w_103_3944, w_103_3953, w_103_3957, w_103_3960, w_103_3963, w_103_3971, w_103_3975, w_103_3979, w_103_3980, w_103_3986, w_103_3989, w_103_3991, w_103_4000, w_103_4001, w_103_4003, w_103_4005, w_103_4010, w_103_4014, w_103_4017, w_103_4019, w_103_4020, w_103_4021, w_103_4027, w_103_4028, w_103_4033, w_103_4037, w_103_4039, w_103_4040, w_103_4042, w_103_4049, w_103_4059, w_103_4063, w_103_4066, w_103_4070, w_103_4072, w_103_4073, w_103_4076, w_103_4077, w_103_4078, w_103_4080, w_103_4092, w_103_4099, w_103_4105, w_103_4110, w_103_4114, w_103_4116, w_103_4121, w_103_4123, w_103_4125, w_103_4127, w_103_4132, w_103_4135, w_103_4139, w_103_4141, w_103_4142, w_103_4144, w_103_4146, w_103_4148, w_103_4149, w_103_4150, w_103_4152, w_103_4155, w_103_4163, w_103_4172, w_103_4174, w_103_4182, w_103_4184, w_103_4191, w_103_4195, w_103_4196, w_103_4197, w_103_4198, w_103_4202, w_103_4205, w_103_4206, w_103_4210, w_103_4213, w_103_4215, w_103_4222, w_103_4223, w_103_4224, w_103_4227, w_103_4239, w_103_4241, w_103_4243, w_103_4251, w_103_4256, w_103_4262, w_103_4263, w_103_4267, w_103_4272, w_103_4273, w_103_4274, w_103_4277, w_103_4278, w_103_4286, w_103_4292, w_103_4296, w_103_4297, w_103_4304, w_103_4305, w_103_4310, w_103_4315, w_103_4319, w_103_4326, w_103_4327, w_103_4328, w_103_4332, w_103_4338, w_103_4340, w_103_4347, w_103_4349, w_103_4357, w_103_4364, w_103_4370, w_103_4376, w_103_4380, w_103_4389, w_103_4390, w_103_4391, w_103_4395, w_103_4399, w_103_4401, w_103_4408, w_103_4417, w_103_4426, w_103_4427, w_103_4429, w_103_4430, w_103_4441, w_103_4442, w_103_4445, w_103_4446, w_103_4456, w_103_4458, w_103_4463, w_103_4464, w_103_4480, w_103_4485, w_103_4488, w_103_4493, w_103_4494, w_103_4498, w_103_4503, w_103_4504, w_103_4512, w_103_4513, w_103_4514, w_103_4515, w_103_4520, w_103_4522, w_103_4532, w_103_4540, w_103_4543, w_103_4544, w_103_4552, w_103_4554, w_103_4562, w_103_4568, w_103_4572, w_103_4575, w_103_4584, w_103_4591, w_103_4592, w_103_4593, w_103_4597, w_103_4603, w_103_4605, w_103_4606, w_103_4607, w_103_4612, w_103_4616, w_103_4623, w_103_4631, w_103_4635, w_103_4640, w_103_4644, w_103_4646, w_103_4647, w_103_4659, w_103_4662, w_103_4664, w_103_4669, w_103_4671, w_103_4674, w_103_4679, w_103_4681, w_103_4688, w_103_4689, w_103_4693, w_103_4702, w_103_4713, w_103_4714, w_103_4719, w_103_4720, w_103_4721, w_103_4725, w_103_4726, w_103_4727, w_103_4728, w_103_4731, w_103_4734, w_103_4740, w_103_4748, w_103_4753, w_103_4758, w_103_4763, w_103_4764, w_103_4765, w_103_4767, w_103_4769, w_103_4770, w_103_4773, w_103_4774, w_103_4775, w_103_4782, w_103_4783, w_103_4784, w_103_4789, w_103_4793, w_103_4795, w_103_4798, w_103_4802, w_103_4803, w_103_4805, w_103_4806, w_103_4808;
  wire w_104_000, w_104_002, w_104_003, w_104_005, w_104_008, w_104_009, w_104_011, w_104_017, w_104_019, w_104_023, w_104_030, w_104_031, w_104_032, w_104_033, w_104_034, w_104_035, w_104_038, w_104_039, w_104_040, w_104_044, w_104_047, w_104_049, w_104_050, w_104_052, w_104_055, w_104_056, w_104_058, w_104_060, w_104_061, w_104_062, w_104_063, w_104_065, w_104_068, w_104_069, w_104_075, w_104_076, w_104_081, w_104_082, w_104_083, w_104_085, w_104_086, w_104_090, w_104_091, w_104_092, w_104_093, w_104_094, w_104_095, w_104_096, w_104_098, w_104_102, w_104_103, w_104_104, w_104_107, w_104_110, w_104_112, w_104_113, w_104_114, w_104_116, w_104_117, w_104_118, w_104_121, w_104_122, w_104_123, w_104_126, w_104_127, w_104_131, w_104_137, w_104_138, w_104_139, w_104_142, w_104_146, w_104_149, w_104_154, w_104_155, w_104_160, w_104_162, w_104_163, w_104_165, w_104_166, w_104_167, w_104_170, w_104_171, w_104_174, w_104_175, w_104_177, w_104_182, w_104_184, w_104_185, w_104_187, w_104_188, w_104_189, w_104_192, w_104_193, w_104_194, w_104_197, w_104_200, w_104_202, w_104_203, w_104_205, w_104_212, w_104_213, w_104_216, w_104_217, w_104_219, w_104_220, w_104_221, w_104_223, w_104_226, w_104_228, w_104_230, w_104_235, w_104_236, w_104_239, w_104_240, w_104_246, w_104_247, w_104_249, w_104_250, w_104_251, w_104_255, w_104_256, w_104_259, w_104_262, w_104_263, w_104_265, w_104_267, w_104_268, w_104_269, w_104_271, w_104_273, w_104_275, w_104_276, w_104_277, w_104_283, w_104_284, w_104_285, w_104_287, w_104_288, w_104_290, w_104_291, w_104_299, w_104_300, w_104_302, w_104_303, w_104_305, w_104_307, w_104_310, w_104_311, w_104_312, w_104_313, w_104_314, w_104_320, w_104_321, w_104_323, w_104_329, w_104_333, w_104_334, w_104_335, w_104_338, w_104_340, w_104_343, w_104_344, w_104_345, w_104_346, w_104_347, w_104_349, w_104_353, w_104_357, w_104_359, w_104_360, w_104_361, w_104_362, w_104_363, w_104_364, w_104_365, w_104_366, w_104_367, w_104_369, w_104_371, w_104_378, w_104_379, w_104_385, w_104_386, w_104_387, w_104_390, w_104_392, w_104_394, w_104_395, w_104_398, w_104_399, w_104_400, w_104_401, w_104_403, w_104_406, w_104_409, w_104_410, w_104_411, w_104_412, w_104_417, w_104_418, w_104_420, w_104_422, w_104_423, w_104_424, w_104_426, w_104_428, w_104_431, w_104_432, w_104_436, w_104_438, w_104_442, w_104_443, w_104_446, w_104_447, w_104_451, w_104_454, w_104_456, w_104_457, w_104_459, w_104_461, w_104_463, w_104_465, w_104_466, w_104_468, w_104_469, w_104_470, w_104_475, w_104_480, w_104_486, w_104_497, w_104_502, w_104_510, w_104_515, w_104_519, w_104_522, w_104_527, w_104_529, w_104_539, w_104_540, w_104_552, w_104_553, w_104_566, w_104_572, w_104_574, w_104_577, w_104_579, w_104_580, w_104_581, w_104_582, w_104_586, w_104_587, w_104_591, w_104_594, w_104_598, w_104_600, w_104_610, w_104_611, w_104_613, w_104_616, w_104_623, w_104_624, w_104_626, w_104_628, w_104_634, w_104_639, w_104_640, w_104_641, w_104_657, w_104_659, w_104_661, w_104_665, w_104_671, w_104_674, w_104_676, w_104_687, w_104_688, w_104_690, w_104_692, w_104_693, w_104_694, w_104_697, w_104_698, w_104_701, w_104_705, w_104_706, w_104_708, w_104_709, w_104_716, w_104_731, w_104_738, w_104_739, w_104_740, w_104_745, w_104_749, w_104_758, w_104_763, w_104_765, w_104_774, w_104_775, w_104_778, w_104_783, w_104_785, w_104_787, w_104_788, w_104_789, w_104_791, w_104_798, w_104_803, w_104_807, w_104_812, w_104_814, w_104_817, w_104_824, w_104_826, w_104_829, w_104_834, w_104_837, w_104_841, w_104_842, w_104_848, w_104_855, w_104_859, w_104_861, w_104_867, w_104_872, w_104_876, w_104_880, w_104_886, w_104_888, w_104_894, w_104_896, w_104_911, w_104_916, w_104_917, w_104_918, w_104_927, w_104_928, w_104_937, w_104_945, w_104_947, w_104_952, w_104_954, w_104_962, w_104_966, w_104_967, w_104_973, w_104_979, w_104_980, w_104_987, w_104_998, w_104_1004, w_104_1006, w_104_1009, w_104_1016, w_104_1018, w_104_1021, w_104_1022, w_104_1023, w_104_1027, w_104_1034, w_104_1037, w_104_1043, w_104_1051, w_104_1053, w_104_1055, w_104_1062, w_104_1064, w_104_1066, w_104_1070, w_104_1073, w_104_1077, w_104_1081, w_104_1084, w_104_1089, w_104_1091, w_104_1093, w_104_1101, w_104_1102, w_104_1103, w_104_1104, w_104_1107, w_104_1119, w_104_1120, w_104_1123, w_104_1132, w_104_1134, w_104_1135, w_104_1137, w_104_1140, w_104_1141, w_104_1143, w_104_1145, w_104_1147, w_104_1150, w_104_1152, w_104_1160, w_104_1161, w_104_1164, w_104_1166, w_104_1169, w_104_1172, w_104_1179, w_104_1185, w_104_1187, w_104_1189, w_104_1190, w_104_1194, w_104_1197, w_104_1198, w_104_1199, w_104_1201, w_104_1209, w_104_1213, w_104_1219, w_104_1221, w_104_1224, w_104_1225, w_104_1227, w_104_1229, w_104_1233, w_104_1236, w_104_1237, w_104_1238, w_104_1239, w_104_1242, w_104_1250, w_104_1251, w_104_1254, w_104_1257, w_104_1265, w_104_1267, w_104_1270, w_104_1285, w_104_1291, w_104_1292, w_104_1302, w_104_1303, w_104_1306, w_104_1307, w_104_1308, w_104_1316, w_104_1319, w_104_1321, w_104_1323, w_104_1324, w_104_1329, w_104_1340, w_104_1343, w_104_1348, w_104_1350, w_104_1352, w_104_1356, w_104_1357, w_104_1361, w_104_1367, w_104_1369, w_104_1374, w_104_1380, w_104_1382, w_104_1383, w_104_1391, w_104_1399, w_104_1405, w_104_1419, w_104_1422, w_104_1432, w_104_1434, w_104_1436, w_104_1437, w_104_1439, w_104_1440, w_104_1442, w_104_1445, w_104_1449, w_104_1450, w_104_1456, w_104_1463, w_104_1464, w_104_1466, w_104_1467, w_104_1472, w_104_1476, w_104_1480, w_104_1484, w_104_1487, w_104_1493, w_104_1497, w_104_1498, w_104_1499, w_104_1504, w_104_1510, w_104_1512, w_104_1513, w_104_1517, w_104_1520, w_104_1523, w_104_1524, w_104_1526, w_104_1529, w_104_1535, w_104_1539, w_104_1547, w_104_1551, w_104_1552, w_104_1553, w_104_1558, w_104_1564, w_104_1566, w_104_1577, w_104_1578, w_104_1588, w_104_1596, w_104_1602, w_104_1606, w_104_1608, w_104_1609, w_104_1612, w_104_1614, w_104_1634, w_104_1638, w_104_1642, w_104_1647, w_104_1656, w_104_1659, w_104_1662, w_104_1666, w_104_1668, w_104_1673, w_104_1675, w_104_1685, w_104_1690, w_104_1691, w_104_1693, w_104_1697, w_104_1698, w_104_1707, w_104_1712, w_104_1718, w_104_1722, w_104_1724, w_104_1725, w_104_1726, w_104_1731, w_104_1732, w_104_1735, w_104_1736, w_104_1738, w_104_1743, w_104_1750, w_104_1754, w_104_1757, w_104_1759, w_104_1768, w_104_1771, w_104_1776, w_104_1777, w_104_1778, w_104_1780, w_104_1785, w_104_1786, w_104_1790, w_104_1803, w_104_1808, w_104_1809, w_104_1814, w_104_1818, w_104_1820, w_104_1830, w_104_1833, w_104_1835, w_104_1836, w_104_1845, w_104_1846, w_104_1857, w_104_1862, w_104_1864, w_104_1888, w_104_1899, w_104_1903, w_104_1906, w_104_1914, w_104_1915, w_104_1920, w_104_1923, w_104_1929, w_104_1932, w_104_1933, w_104_1937, w_104_1940, w_104_1943, w_104_1946, w_104_1947, w_104_1951, w_104_1953, w_104_1962, w_104_1963, w_104_1966, w_104_1968, w_104_1969, w_104_1970, w_104_1971, w_104_1973, w_104_1981, w_104_1987, w_104_1992, w_104_1995, w_104_1997, w_104_1999, w_104_2000, w_104_2001, w_104_2002, w_104_2003, w_104_2005, w_104_2011, w_104_2012, w_104_2015, w_104_2022, w_104_2023, w_104_2025, w_104_2032, w_104_2034, w_104_2042, w_104_2050, w_104_2053, w_104_2057, w_104_2061, w_104_2062, w_104_2064, w_104_2067, w_104_2072, w_104_2075, w_104_2077, w_104_2081, w_104_2082, w_104_2089, w_104_2095, w_104_2098, w_104_2101, w_104_2105, w_104_2107, w_104_2108, w_104_2109, w_104_2112, w_104_2115, w_104_2123, w_104_2132, w_104_2134, w_104_2137, w_104_2140, w_104_2144, w_104_2146, w_104_2149, w_104_2150, w_104_2161, w_104_2163, w_104_2164, w_104_2166, w_104_2168, w_104_2182, w_104_2195, w_104_2204, w_104_2210, w_104_2215, w_104_2222, w_104_2223, w_104_2226, w_104_2229, w_104_2237, w_104_2239, w_104_2243, w_104_2249, w_104_2252, w_104_2254, w_104_2262, w_104_2263, w_104_2265, w_104_2268, w_104_2270, w_104_2274, w_104_2284, w_104_2290, w_104_2291, w_104_2294, w_104_2302, w_104_2304, w_104_2307, w_104_2308, w_104_2309, w_104_2314, w_104_2318, w_104_2320, w_104_2321, w_104_2323, w_104_2324, w_104_2328, w_104_2330, w_104_2331, w_104_2334, w_104_2337, w_104_2339, w_104_2350, w_104_2355, w_104_2356, w_104_2365, w_104_2369, w_104_2373, w_104_2374, w_104_2378, w_104_2383, w_104_2387, w_104_2391, w_104_2396, w_104_2398, w_104_2400, w_104_2402, w_104_2403, w_104_2411, w_104_2418, w_104_2419, w_104_2428, w_104_2430, w_104_2442, w_104_2443, w_104_2444, w_104_2445, w_104_2446, w_104_2452, w_104_2457, w_104_2465, w_104_2466, w_104_2474, w_104_2476, w_104_2477, w_104_2481, w_104_2489, w_104_2506, w_104_2509, w_104_2513, w_104_2514, w_104_2518, w_104_2521, w_104_2522, w_104_2524, w_104_2526, w_104_2528, w_104_2533, w_104_2537, w_104_2539, w_104_2541, w_104_2542, w_104_2547, w_104_2548, w_104_2549, w_104_2553, w_104_2556, w_104_2559, w_104_2563, w_104_2566, w_104_2568, w_104_2569, w_104_2572, w_104_2574, w_104_2575, w_104_2576, w_104_2578, w_104_2584, w_104_2590, w_104_2595, w_104_2596, w_104_2597, w_104_2598, w_104_2605, w_104_2614, w_104_2615, w_104_2616, w_104_2620, w_104_2621, w_104_2622, w_104_2628, w_104_2631, w_104_2634, w_104_2636, w_104_2638, w_104_2640, w_104_2641, w_104_2647, w_104_2648, w_104_2649, w_104_2651, w_104_2653, w_104_2658, w_104_2664, w_104_2666, w_104_2679, w_104_2681, w_104_2684, w_104_2685, w_104_2687, w_104_2689, w_104_2696, w_104_2702, w_104_2706, w_104_2707, w_104_2711, w_104_2716, w_104_2718, w_104_2725, w_104_2727, w_104_2729, w_104_2732, w_104_2734, w_104_2735, w_104_2736, w_104_2737, w_104_2738, w_104_2743, w_104_2745, w_104_2746, w_104_2750, w_104_2755, w_104_2757, w_104_2761, w_104_2776, w_104_2786, w_104_2789, w_104_2793, w_104_2796, w_104_2806, w_104_2807, w_104_2814, w_104_2815, w_104_2817, w_104_2818, w_104_2820, w_104_2821, w_104_2822, w_104_2824, w_104_2826, w_104_2841, w_104_2848, w_104_2849, w_104_2853, w_104_2861, w_104_2871, w_104_2872, w_104_2874, w_104_2880, w_104_2881, w_104_2883, w_104_2885, w_104_2887, w_104_2891, w_104_2893, w_104_2894, w_104_2903, w_104_2908, w_104_2910, w_104_2915, w_104_2921, w_104_2923, w_104_2924, w_104_2927, w_104_2933, w_104_2937, w_104_2941, w_104_2942, w_104_2944, w_104_2946, w_104_2952, w_104_2953, w_104_2954, w_104_2955, w_104_2956, w_104_2964, w_104_2973, w_104_2980, w_104_2983, w_104_2987, w_104_2990, w_104_2992, w_104_2993, w_104_2994, w_104_2995, w_104_2999, w_104_3024, w_104_3029, w_104_3032, w_104_3034, w_104_3038, w_104_3046, w_104_3049, w_104_3055, w_104_3063, w_104_3064, w_104_3076, w_104_3078, w_104_3080, w_104_3082, w_104_3083, w_104_3092, w_104_3104, w_104_3107, w_104_3111, w_104_3115, w_104_3119, w_104_3122, w_104_3139, w_104_3141, w_104_3144, w_104_3150, w_104_3154, w_104_3155, w_104_3159, w_104_3162, w_104_3163, w_104_3166, w_104_3170, w_104_3173, w_104_3175, w_104_3179, w_104_3181, w_104_3186, w_104_3187, w_104_3192, w_104_3193, w_104_3194, w_104_3203, w_104_3209, w_104_3213, w_104_3219, w_104_3220, w_104_3223, w_104_3226, w_104_3242, w_104_3246, w_104_3247, w_104_3255, w_104_3257, w_104_3258, w_104_3259, w_104_3266, w_104_3268, w_104_3274, w_104_3276, w_104_3284, w_104_3288, w_104_3290, w_104_3291, w_104_3296, w_104_3298, w_104_3299, w_104_3302, w_104_3307, w_104_3311, w_104_3312, w_104_3324, w_104_3332, w_104_3339, w_104_3342, w_104_3344, w_104_3346, w_104_3354, w_104_3358, w_104_3359, w_104_3360, w_104_3367, w_104_3376, w_104_3377, w_104_3379, w_104_3383, w_104_3385, w_104_3387, w_104_3391, w_104_3392, w_104_3393, w_104_3399, w_104_3402, w_104_3405, w_104_3412, w_104_3415, w_104_3420, w_104_3428, w_104_3431, w_104_3432, w_104_3435, w_104_3436, w_104_3437, w_104_3438, w_104_3441, w_104_3445, w_104_3450, w_104_3451, w_104_3453, w_104_3454, w_104_3457, w_104_3458, w_104_3466, w_104_3469, w_104_3470, w_104_3474, w_104_3476, w_104_3480, w_104_3485, w_104_3486, w_104_3496, w_104_3503, w_104_3504, w_104_3506, w_104_3510, w_104_3511, w_104_3523, w_104_3524, w_104_3526, w_104_3528, w_104_3532, w_104_3533, w_104_3537, w_104_3539, w_104_3542, w_104_3544, w_104_3545, w_104_3546, w_104_3555, w_104_3556, w_104_3559, w_104_3564, w_104_3567, w_104_3571, w_104_3574, w_104_3577, w_104_3580, w_104_3585, w_104_3588, w_104_3594, w_104_3595, w_104_3604, w_104_3605, w_104_3607, w_104_3608, w_104_3609, w_104_3615, w_104_3617, w_104_3618, w_104_3621, w_104_3626, w_104_3639, w_104_3640, w_104_3641, w_104_3644, w_104_3646, w_104_3656, w_104_3657, w_104_3662, w_104_3666, w_104_3668, w_104_3674, w_104_3681, w_104_3685, w_104_3687, w_104_3698, w_104_3700, w_104_3702, w_104_3709, w_104_3710, w_104_3713, w_104_3720, w_104_3724, w_104_3729, w_104_3737, w_104_3740, w_104_3746, w_104_3748, w_104_3754, w_104_3765, w_104_3767, w_104_3773, w_104_3780, w_104_3788, w_104_3789, w_104_3793, w_104_3795, w_104_3796, w_104_3797, w_104_3804, w_104_3806, w_104_3812, w_104_3813, w_104_3818, w_104_3820, w_104_3825, w_104_3826, w_104_3827, w_104_3830, w_104_3833, w_104_3837, w_104_3840, w_104_3841, w_104_3855, w_104_3859, w_104_3863, w_104_3864, w_104_3865, w_104_3867, w_104_3871, w_104_3872, w_104_3873, w_104_3883, w_104_3887, w_104_3889, w_104_3890, w_104_3891, w_104_3894, w_104_3895, w_104_3897, w_104_3899, w_104_3905, w_104_3909, w_104_3915, w_104_3919, w_104_3922, w_104_3923, w_104_3924, w_104_3925, w_104_3929, w_104_3930, w_104_3934, w_104_3936, w_104_3940, w_104_3946, w_104_3947, w_104_3949, w_104_3953, w_104_3957, w_104_3958, w_104_3962, w_104_3963, w_104_3964, w_104_3965, w_104_3972, w_104_3973, w_104_3974, w_104_3977, w_104_3981, w_104_3987, w_104_3992, w_104_3995, w_104_3996, w_104_3998, w_104_4001, w_104_4003, w_104_4011, w_104_4024, w_104_4028, w_104_4031, w_104_4033, w_104_4035, w_104_4042, w_104_4047, w_104_4049, w_104_4053, w_104_4058, w_104_4059, w_104_4063, w_104_4067, w_104_4070, w_104_4076, w_104_4079, w_104_4081, w_104_4082, w_104_4084, w_104_4089, w_104_4095, w_104_4101, w_104_4103, w_104_4112, w_104_4117, w_104_4121, w_104_4123, w_104_4128, w_104_4129, w_104_4130, w_104_4132, w_104_4134, w_104_4137, w_104_4138, w_104_4146, w_104_4147, w_104_4153, w_104_4154, w_104_4155, w_104_4156, w_104_4160, w_104_4162, w_104_4165, w_104_4167, w_104_4168, w_104_4174, w_104_4177, w_104_4179, w_104_4182, w_104_4194, w_104_4195, w_104_4198, w_104_4206, w_104_4207, w_104_4209, w_104_4211, w_104_4215, w_104_4224, w_104_4232, w_104_4233, w_104_4237, w_104_4240, w_104_4243, w_104_4246, w_104_4247, w_104_4250, w_104_4252, w_104_4253, w_104_4254, w_104_4255, w_104_4258, w_104_4260, w_104_4263, w_104_4273, w_104_4275, w_104_4277, w_104_4282, w_104_4284, w_104_4297, w_104_4301, w_104_4302, w_104_4305, w_104_4333, w_104_4334, w_104_4336, w_104_4340, w_104_4341, w_104_4349, w_104_4357, w_104_4361, w_104_4362, w_104_4365, w_104_4373, w_104_4374, w_104_4375, w_104_4379, w_104_4391, w_104_4396, w_104_4398, w_104_4401, w_104_4404, w_104_4406, w_104_4411, w_104_4412, w_104_4416, w_104_4418, w_104_4431, w_104_4432, w_104_4434, w_104_4442, w_104_4443, w_104_4445, w_104_4447, w_104_4455, w_104_4463, w_104_4469, w_104_4475, w_104_4476, w_104_4480, w_104_4483, w_104_4489, w_104_4493, w_104_4495, w_104_4508, w_104_4513, w_104_4514, w_104_4516, w_104_4519, w_104_4525, w_104_4526, w_104_4527, w_104_4528, w_104_4531, w_104_4535, w_104_4537, w_104_4539, w_104_4540, w_104_4541, w_104_4542, w_104_4543, w_104_4544;
  wire w_105_000, w_105_001, w_105_002, w_105_003, w_105_004, w_105_006, w_105_008, w_105_009, w_105_010, w_105_011, w_105_012, w_105_013, w_105_014, w_105_015, w_105_016, w_105_017, w_105_018, w_105_019, w_105_020, w_105_021, w_105_022, w_105_023, w_105_024, w_105_025, w_105_026, w_105_027, w_105_028, w_105_029, w_105_030, w_105_031, w_105_032, w_105_033, w_105_035, w_105_036, w_105_037, w_105_038, w_105_039, w_105_040, w_105_041, w_105_043, w_105_044, w_105_045, w_105_046, w_105_047, w_105_048, w_105_049, w_105_050, w_105_051, w_105_052, w_105_053, w_105_054, w_105_055, w_105_056, w_105_057, w_105_058, w_105_059, w_105_060, w_105_061, w_105_062, w_105_063, w_105_064, w_105_065, w_105_066, w_105_067, w_105_068, w_105_069, w_105_070, w_105_071, w_105_073, w_105_074, w_105_075, w_105_076, w_105_077, w_105_079, w_105_080, w_105_081, w_105_082, w_105_083, w_105_084, w_105_086, w_105_087, w_105_088, w_105_089, w_105_090, w_105_091, w_105_092, w_105_093, w_105_094, w_105_095, w_105_096, w_105_097, w_105_098, w_105_100, w_105_101, w_105_102, w_105_103, w_105_104, w_105_105, w_105_106, w_105_107, w_105_108, w_105_109, w_105_110, w_105_111, w_105_112, w_105_113, w_105_114, w_105_115, w_105_116, w_105_117, w_105_118, w_105_119, w_105_121, w_105_122, w_105_123, w_105_124, w_105_125, w_105_126, w_105_127, w_105_128, w_105_129, w_105_130, w_105_131, w_105_132, w_105_133, w_105_134, w_105_135, w_105_136, w_105_137, w_105_138, w_105_139, w_105_140, w_105_141, w_105_142, w_105_143, w_105_144, w_105_145, w_105_146, w_105_147, w_105_148, w_105_149, w_105_150, w_105_151, w_105_152, w_105_153, w_105_154, w_105_155, w_105_156, w_105_157, w_105_158, w_105_159, w_105_160, w_105_161, w_105_162, w_105_163, w_105_164, w_105_165, w_105_167, w_105_168, w_105_169, w_105_170, w_105_171, w_105_172, w_105_173, w_105_174, w_105_175, w_105_176, w_105_177, w_105_178, w_105_179, w_105_180, w_105_181, w_105_182, w_105_183, w_105_184, w_105_185, w_105_186, w_105_187, w_105_188, w_105_189, w_105_190, w_105_191, w_105_192, w_105_193, w_105_194, w_105_195, w_105_196, w_105_197, w_105_198, w_105_199, w_105_200, w_105_201, w_105_202, w_105_203, w_105_204, w_105_205, w_105_206, w_105_207, w_105_208, w_105_209, w_105_210, w_105_211, w_105_212, w_105_214, w_105_215, w_105_216, w_105_217, w_105_218, w_105_219, w_105_220, w_105_221, w_105_222, w_105_223, w_105_224, w_105_225, w_105_226, w_105_229, w_105_230, w_105_231, w_105_232, w_105_233, w_105_234, w_105_235, w_105_236, w_105_237, w_105_238, w_105_239, w_105_241, w_105_242, w_105_243, w_105_244, w_105_245, w_105_246, w_105_247, w_105_248, w_105_249, w_105_250, w_105_251, w_105_252, w_105_253, w_105_254, w_105_255, w_105_256, w_105_257, w_105_258, w_105_259, w_105_260, w_105_261, w_105_262, w_105_263, w_105_264, w_105_265, w_105_267, w_105_268, w_105_269, w_105_270, w_105_271, w_105_272, w_105_273, w_105_274, w_105_276, w_105_277, w_105_278, w_105_279, w_105_280, w_105_281, w_105_282, w_105_283, w_105_284, w_105_285, w_105_286, w_105_287, w_105_288, w_105_289, w_105_290, w_105_291, w_105_292, w_105_293, w_105_294, w_105_295, w_105_296, w_105_297, w_105_298, w_105_299, w_105_300, w_105_301, w_105_302, w_105_303, w_105_304, w_105_305, w_105_306, w_105_307, w_105_308, w_105_309, w_105_310, w_105_311, w_105_312, w_105_313, w_105_314, w_105_315, w_105_316, w_105_317, w_105_318, w_105_319, w_105_320, w_105_321, w_105_322, w_105_323, w_105_324, w_105_325, w_105_326, w_105_327, w_105_328, w_105_329, w_105_330, w_105_331, w_105_332, w_105_333, w_105_334, w_105_335, w_105_336, w_105_337, w_105_338, w_105_339, w_105_340, w_105_341, w_105_342, w_105_343, w_105_344, w_105_345, w_105_346, w_105_347, w_105_348, w_105_349, w_105_350, w_105_351, w_105_352, w_105_353, w_105_354, w_105_355, w_105_356, w_105_357, w_105_358, w_105_359, w_105_360, w_105_361, w_105_362, w_105_363, w_105_364, w_105_365, w_105_366, w_105_367, w_105_368, w_105_369, w_105_370, w_105_371, w_105_372, w_105_373, w_105_374, w_105_375, w_105_376, w_105_377, w_105_378, w_105_379, w_105_380, w_105_381, w_105_382, w_105_383, w_105_384, w_105_385, w_105_386, w_105_387, w_105_388, w_105_389, w_105_392, w_105_393, w_105_394, w_105_395, w_105_396, w_105_397, w_105_398, w_105_399, w_105_400, w_105_401, w_105_402, w_105_403, w_105_404, w_105_405, w_105_406, w_105_407, w_105_408, w_105_409, w_105_410, w_105_411, w_105_412, w_105_413, w_105_414, w_105_415, w_105_416, w_105_417, w_105_418, w_105_419, w_105_420, w_105_421, w_105_422, w_105_423, w_105_424, w_105_426, w_105_427, w_105_428, w_105_430, w_105_431, w_105_432, w_105_433, w_105_434, w_105_435, w_105_436, w_105_437, w_105_438, w_105_439, w_105_441, w_105_442, w_105_443, w_105_444, w_105_445, w_105_446, w_105_447, w_105_448, w_105_449, w_105_450, w_105_451, w_105_452, w_105_453, w_105_454, w_105_455, w_105_456, w_105_457, w_105_458, w_105_459, w_105_460, w_105_461, w_105_462, w_105_463, w_105_464, w_105_465, w_105_466, w_105_467, w_105_468, w_105_469, w_105_470, w_105_471, w_105_472, w_105_473, w_105_474, w_105_475, w_105_476, w_105_477, w_105_478, w_105_479, w_105_480, w_105_481, w_105_482, w_105_483, w_105_484, w_105_485, w_105_486, w_105_487, w_105_488, w_105_489, w_105_490, w_105_491, w_105_492, w_105_493, w_105_494, w_105_496, w_105_497, w_105_498, w_105_499, w_105_500, w_105_501, w_105_502, w_105_503, w_105_504, w_105_505, w_105_506, w_105_507, w_105_508, w_105_509, w_105_510, w_105_511, w_105_512, w_105_513, w_105_514, w_105_515, w_105_516, w_105_517, w_105_518, w_105_519, w_105_520, w_105_521, w_105_522, w_105_523, w_105_524, w_105_525, w_105_526, w_105_527, w_105_529, w_105_530, w_105_531, w_105_532, w_105_533, w_105_534, w_105_535, w_105_536, w_105_537, w_105_538, w_105_539, w_105_540, w_105_541, w_105_542, w_105_543, w_105_544, w_105_545, w_105_546, w_105_547;
  wire w_106_000, w_106_004, w_106_005, w_106_006, w_106_007, w_106_008, w_106_012, w_106_014, w_106_015, w_106_016, w_106_019, w_106_020, w_106_023, w_106_027, w_106_028, w_106_031, w_106_032, w_106_034, w_106_037, w_106_039, w_106_042, w_106_043, w_106_044, w_106_045, w_106_046, w_106_047, w_106_048, w_106_049, w_106_052, w_106_053, w_106_054, w_106_056, w_106_057, w_106_058, w_106_061, w_106_062, w_106_063, w_106_064, w_106_065, w_106_067, w_106_068, w_106_069, w_106_073, w_106_075, w_106_076, w_106_079, w_106_082, w_106_083, w_106_084, w_106_085, w_106_086, w_106_087, w_106_089, w_106_091, w_106_093, w_106_094, w_106_095, w_106_097, w_106_098, w_106_099, w_106_100, w_106_104, w_106_105, w_106_106, w_106_107, w_106_109, w_106_110, w_106_115, w_106_121, w_106_122, w_106_126, w_106_128, w_106_139, w_106_142, w_106_143, w_106_145, w_106_149, w_106_150, w_106_154, w_106_155, w_106_156, w_106_158, w_106_160, w_106_162, w_106_163, w_106_165, w_106_166, w_106_168, w_106_173, w_106_174, w_106_176, w_106_178, w_106_180, w_106_183, w_106_185, w_106_186, w_106_195, w_106_198, w_106_199, w_106_207, w_106_209, w_106_213, w_106_215, w_106_220, w_106_222, w_106_232, w_106_234, w_106_235, w_106_236, w_106_237, w_106_238, w_106_239, w_106_244, w_106_245, w_106_246, w_106_249, w_106_250, w_106_251, w_106_253, w_106_254, w_106_260, w_106_261, w_106_264, w_106_265, w_106_267, w_106_268, w_106_270, w_106_271, w_106_275, w_106_278, w_106_280, w_106_283, w_106_284, w_106_285, w_106_287, w_106_288, w_106_289, w_106_290, w_106_293, w_106_294, w_106_299, w_106_301, w_106_302, w_106_304, w_106_309, w_106_311, w_106_316, w_106_319, w_106_321, w_106_323, w_106_326, w_106_327, w_106_332, w_106_334, w_106_337, w_106_338, w_106_339, w_106_341, w_106_344, w_106_350, w_106_351, w_106_352, w_106_354, w_106_355, w_106_367, w_106_368, w_106_371, w_106_373, w_106_378, w_106_379, w_106_380, w_106_382, w_106_384, w_106_385, w_106_387, w_106_388, w_106_389, w_106_393, w_106_399, w_106_402, w_106_405, w_106_409, w_106_410, w_106_411, w_106_412, w_106_414, w_106_416, w_106_418, w_106_425, w_106_426, w_106_430, w_106_431, w_106_432, w_106_433, w_106_440, w_106_443, w_106_446, w_106_447, w_106_448, w_106_449, w_106_452, w_106_453, w_106_455, w_106_458, w_106_460, w_106_465, w_106_466, w_106_467, w_106_473, w_106_475, w_106_479, w_106_480, w_106_481, w_106_483, w_106_485, w_106_486, w_106_490, w_106_493, w_106_497, w_106_502, w_106_503, w_106_504, w_106_506, w_106_507, w_106_508, w_106_509, w_106_512, w_106_513, w_106_516, w_106_518, w_106_519, w_106_520, w_106_521, w_106_525, w_106_526, w_106_530, w_106_531, w_106_534, w_106_535, w_106_539, w_106_541, w_106_543, w_106_544, w_106_546, w_106_547, w_106_550, w_106_551, w_106_553, w_106_556, w_106_560, w_106_564, w_106_566, w_106_567, w_106_569, w_106_570, w_106_574, w_106_577, w_106_579, w_106_581, w_106_584, w_106_586, w_106_588, w_106_589, w_106_590, w_106_591, w_106_592, w_106_594, w_106_595, w_106_600, w_106_601, w_106_602, w_106_608, w_106_609, w_106_611, w_106_613, w_106_614, w_106_615, w_106_616, w_106_618, w_106_622, w_106_625, w_106_629, w_106_630, w_106_631, w_106_633, w_106_634, w_106_635, w_106_637, w_106_638, w_106_639, w_106_645, w_106_646, w_106_648, w_106_649, w_106_654, w_106_657, w_106_660, w_106_663, w_106_665, w_106_666, w_106_667, w_106_669, w_106_673, w_106_674, w_106_677, w_106_681, w_106_682, w_106_683, w_106_684, w_106_687, w_106_688, w_106_689, w_106_693, w_106_695, w_106_697, w_106_698, w_106_699, w_106_700, w_106_701, w_106_704, w_106_705, w_106_706, w_106_708, w_106_710, w_106_711, w_106_720, w_106_723, w_106_725, w_106_727, w_106_735, w_106_736, w_106_737, w_106_738, w_106_740, w_106_742, w_106_743, w_106_747, w_106_750, w_106_751, w_106_754, w_106_756, w_106_758, w_106_759, w_106_761, w_106_762, w_106_763, w_106_764, w_106_767, w_106_768, w_106_770, w_106_771, w_106_773, w_106_777, w_106_779, w_106_781, w_106_783, w_106_785, w_106_787, w_106_788, w_106_790, w_106_791, w_106_792, w_106_795, w_106_796, w_106_798, w_106_800, w_106_803, w_106_806, w_106_811, w_106_813, w_106_815, w_106_816, w_106_817, w_106_818, w_106_819, w_106_822, w_106_823, w_106_824, w_106_825, w_106_826, w_106_827, w_106_833, w_106_837, w_106_838, w_106_841, w_106_842, w_106_847, w_106_849, w_106_851, w_106_853, w_106_854, w_106_857, w_106_858, w_106_861, w_106_866, w_106_868, w_106_869, w_106_870, w_106_871, w_106_875, w_106_879, w_106_881, w_106_883, w_106_886, w_106_887, w_106_888, w_106_889, w_106_892, w_106_893, w_106_895, w_106_897, w_106_901, w_106_903, w_106_907, w_106_909, w_106_913, w_106_914, w_106_917, w_106_918, w_106_919, w_106_920, w_106_921, w_106_923, w_106_926, w_106_928, w_106_933, w_106_934, w_106_940, w_106_943, w_106_946, w_106_947, w_106_951, w_106_956, w_106_957, w_106_958, w_106_959, w_106_964, w_106_965, w_106_966, w_106_968, w_106_969, w_106_973, w_106_975, w_106_979, w_106_981, w_106_982, w_106_985, w_106_986, w_106_988, w_106_992, w_106_994, w_106_995, w_106_996, w_106_997, w_106_998, w_106_1000, w_106_1003, w_106_1005, w_106_1007, w_106_1010, w_106_1012, w_106_1018, w_106_1019, w_106_1020, w_106_1022, w_106_1023, w_106_1026, w_106_1028, w_106_1030, w_106_1036, w_106_1037, w_106_1041, w_106_1047, w_106_1050, w_106_1053, w_106_1055, w_106_1057, w_106_1061, w_106_1062, w_106_1065, w_106_1068, w_106_1071, w_106_1074, w_106_1076, w_106_1080, w_106_1083, w_106_1084, w_106_1086, w_106_1087, w_106_1088, w_106_1090, w_106_1091, w_106_1094, w_106_1096, w_106_1097, w_106_1098, w_106_1101, w_106_1102, w_106_1105, w_106_1107, w_106_1108, w_106_1111, w_106_1112, w_106_1115, w_106_1116, w_106_1118, w_106_1119, w_106_1124, w_106_1125, w_106_1129, w_106_1130, w_106_1132, w_106_1134, w_106_1135, w_106_1136, w_106_1138, w_106_1141, w_106_1142, w_106_1145, w_106_1146, w_106_1148, w_106_1150, w_106_1151, w_106_1152, w_106_1154, w_106_1155, w_106_1157, w_106_1162, w_106_1165, w_106_1166, w_106_1169, w_106_1172, w_106_1175, w_106_1176, w_106_1177, w_106_1180, w_106_1183, w_106_1192, w_106_1194, w_106_1196, w_106_1198, w_106_1199, w_106_1204, w_106_1205, w_106_1207, w_106_1208, w_106_1209, w_106_1211, w_106_1213, w_106_1214, w_106_1215, w_106_1216, w_106_1217, w_106_1218, w_106_1222, w_106_1223, w_106_1224, w_106_1226, w_106_1227, w_106_1232, w_106_1233, w_106_1234, w_106_1235, w_106_1237, w_106_1238, w_106_1239, w_106_1240, w_106_1244, w_106_1245, w_106_1246, w_106_1247, w_106_1249, w_106_1250, w_106_1251, w_106_1252, w_106_1253, w_106_1254, w_106_1257, w_106_1258, w_106_1261, w_106_1263, w_106_1264, w_106_1266, w_106_1269, w_106_1272, w_106_1274, w_106_1277, w_106_1281, w_106_1282, w_106_1284, w_106_1285, w_106_1286, w_106_1288, w_106_1289, w_106_1291, w_106_1292, w_106_1294, w_106_1296, w_106_1297, w_106_1298, w_106_1306, w_106_1307, w_106_1308, w_106_1309, w_106_1314, w_106_1316, w_106_1326, w_106_1328, w_106_1331, w_106_1332, w_106_1335, w_106_1336, w_106_1338, w_106_1340, w_106_1341, w_106_1345, w_106_1352, w_106_1354, w_106_1356, w_106_1357, w_106_1361, w_106_1362, w_106_1364, w_106_1368, w_106_1370, w_106_1371, w_106_1373, w_106_1376, w_106_1377, w_106_1382, w_106_1384, w_106_1388, w_106_1389, w_106_1390, w_106_1391, w_106_1399, w_106_1402, w_106_1403, w_106_1406, w_106_1408, w_106_1410, w_106_1413, w_106_1414, w_106_1419, w_106_1422, w_106_1425, w_106_1426, w_106_1427, w_106_1428, w_106_1432, w_106_1434, w_106_1439, w_106_1444, w_106_1445, w_106_1447, w_106_1448, w_106_1451, w_106_1454, w_106_1455, w_106_1461, w_106_1463, w_106_1465, w_106_1466, w_106_1467, w_106_1470, w_106_1472, w_106_1473, w_106_1476, w_106_1480, w_106_1481, w_106_1483, w_106_1485, w_106_1487, w_106_1488, w_106_1489, w_106_1490, w_106_1491, w_106_1494, w_106_1495, w_106_1497, w_106_1498, w_106_1501, w_106_1503, w_106_1505, w_106_1507, w_106_1508, w_106_1509, w_106_1513, w_106_1521, w_106_1524, w_106_1525, w_106_1527, w_106_1529, w_106_1532, w_106_1533, w_106_1534, w_106_1535, w_106_1537, w_106_1539, w_106_1540, w_106_1542, w_106_1543, w_106_1546, w_106_1547, w_106_1552, w_106_1553, w_106_1555, w_106_1556, w_106_1560, w_106_1563, w_106_1564, w_106_1565, w_106_1566, w_106_1568, w_106_1569, w_106_1570, w_106_1574, w_106_1575, w_106_1576, w_106_1579, w_106_1581, w_106_1586, w_106_1587, w_106_1590, w_106_1591, w_106_1594, w_106_1595, w_106_1597, w_106_1599, w_106_1600, w_106_1602, w_106_1604, w_106_1608, w_106_1609, w_106_1610, w_106_1613, w_106_1615, w_106_1616, w_106_1617, w_106_1618, w_106_1619, w_106_1623, w_106_1627, w_106_1629, w_106_1632, w_106_1636, w_106_1637, w_106_1638, w_106_1639, w_106_1641, w_106_1642, w_106_1645, w_106_1646, w_106_1647, w_106_1648, w_106_1650, w_106_1651, w_106_1653, w_106_1655, w_106_1658, w_106_1662, w_106_1668, w_106_1669, w_106_1671, w_106_1672, w_106_1673, w_106_1674, w_106_1677, w_106_1680, w_106_1681, w_106_1687, w_106_1688, w_106_1691, w_106_1692, w_106_1693, w_106_1694, w_106_1695, w_106_1696, w_106_1697, w_106_1698, w_106_1704, w_106_1705, w_106_1709, w_106_1710, w_106_1711, w_106_1719, w_106_1720, w_106_1721, w_106_1722, w_106_1723, w_106_1726, w_106_1727, w_106_1729, w_106_1730, w_106_1733, w_106_1737, w_106_1740, w_106_1742, w_106_1744, w_106_1746, w_106_1747, w_106_1750, w_106_1754, w_106_1758, w_106_1761, w_106_1764, w_106_1765, w_106_1767, w_106_1768, w_106_1769, w_106_1770, w_106_1771, w_106_1773, w_106_1775, w_106_1776, w_106_1782, w_106_1784, w_106_1785, w_106_1788, w_106_1792, w_106_1795, w_106_1797, w_106_1798, w_106_1806, w_106_1807, w_106_1808, w_106_1811, w_106_1812, w_106_1813, w_106_1815, w_106_1816, w_106_1817, w_106_1818, w_106_1819, w_106_1820, w_106_1821, w_106_1824, w_106_1825, w_106_1826, w_106_1828, w_106_1833, w_106_1834, w_106_1836, w_106_1838, w_106_1845, w_106_1847, w_106_1850, w_106_1853, w_106_1855, w_106_1858, w_106_1859, w_106_1861, w_106_1862, w_106_1864, w_106_1865, w_106_1867, w_106_1868, w_106_1872, w_106_1876, w_106_1877, w_106_1880, w_106_1884, w_106_1885, w_106_1888, w_106_1889, w_106_1893, w_106_1895, w_106_1902, w_106_1903, w_106_1905, w_106_1906, w_106_1908, w_106_1911, w_106_1924, w_106_1926, w_106_1928, w_106_1929, w_106_1932, w_106_1933, w_106_1936, w_106_1938, w_106_1939, w_106_1947, w_106_1951, w_106_1956, w_106_1971, w_106_1972, w_106_1973, w_106_1980, w_106_1982, w_106_1983, w_106_1989, w_106_1996, w_106_1999, w_106_2002, w_106_2004, w_106_2012, w_106_2016, w_106_2023, w_106_2024, w_106_2032, w_106_2036, w_106_2052, w_106_2063, w_106_2069, w_106_2077, w_106_2079, w_106_2088, w_106_2094, w_106_2099, w_106_2100, w_106_2101, w_106_2108, w_106_2111, w_106_2113, w_106_2115, w_106_2116, w_106_2121, w_106_2124, w_106_2125, w_106_2129, w_106_2130, w_106_2131, w_106_2133, w_106_2142, w_106_2150, w_106_2158, w_106_2160, w_106_2177, w_106_2178, w_106_2180, w_106_2185, w_106_2187, w_106_2188, w_106_2193, w_106_2203, w_106_2205, w_106_2210, w_106_2218, w_106_2221, w_106_2225, w_106_2226, w_106_2234, w_106_2237, w_106_2240, w_106_2246, w_106_2247, w_106_2250, w_106_2252, w_106_2256, w_106_2258, w_106_2260, w_106_2261, w_106_2265, w_106_2271, w_106_2273, w_106_2275, w_106_2289, w_106_2292, w_106_2296, w_106_2297, w_106_2302, w_106_2303, w_106_2304, w_106_2309, w_106_2310, w_106_2311, w_106_2312, w_106_2317, w_106_2320, w_106_2321, w_106_2326, w_106_2327, w_106_2329, w_106_2334, w_106_2335, w_106_2336, w_106_2344, w_106_2349, w_106_2353, w_106_2361, w_106_2363, w_106_2364, w_106_2371, w_106_2375, w_106_2376, w_106_2379, w_106_2383, w_106_2384, w_106_2386, w_106_2391, w_106_2392, w_106_2403, w_106_2405, w_106_2408, w_106_2419, w_106_2430, w_106_2433, w_106_2436, w_106_2439, w_106_2459, w_106_2463, w_106_2465, w_106_2466, w_106_2469, w_106_2470, w_106_2472, w_106_2473, w_106_2474, w_106_2479, w_106_2480, w_106_2481, w_106_2484, w_106_2489, w_106_2495, w_106_2500, w_106_2502, w_106_2504, w_106_2505, w_106_2518, w_106_2522, w_106_2523, w_106_2524, w_106_2529, w_106_2536, w_106_2537, w_106_2538, w_106_2539, w_106_2540, w_106_2543, w_106_2544, w_106_2545, w_106_2548, w_106_2554, w_106_2557, w_106_2562, w_106_2570, w_106_2573, w_106_2578, w_106_2586, w_106_2588, w_106_2592, w_106_2601, w_106_2613, w_106_2619, w_106_2620, w_106_2626, w_106_2630, w_106_2657, w_106_2663, w_106_2665, w_106_2667, w_106_2668, w_106_2669, w_106_2678, w_106_2685, w_106_2687, w_106_2689, w_106_2690, w_106_2703, w_106_2707, w_106_2708, w_106_2710, w_106_2713, w_106_2719, w_106_2725, w_106_2726, w_106_2727, w_106_2728, w_106_2730, w_106_2733, w_106_2735, w_106_2740, w_106_2745, w_106_2750, w_106_2763, w_106_2765, w_106_2768, w_106_2769, w_106_2770, w_106_2773, w_106_2775, w_106_2779, w_106_2783, w_106_2790, w_106_2792, w_106_2801, w_106_2807, w_106_2811, w_106_2816, w_106_2827, w_106_2831, w_106_2836, w_106_2837, w_106_2839, w_106_2842, w_106_2847, w_106_2849, w_106_2850, w_106_2853, w_106_2860, w_106_2863, w_106_2867, w_106_2868, w_106_2871, w_106_2877, w_106_2879, w_106_2884, w_106_2885, w_106_2891, w_106_2893, w_106_2897, w_106_2898, w_106_2900, w_106_2902, w_106_2908, w_106_2916, w_106_2939, w_106_2944, w_106_2949, w_106_2951, w_106_2953, w_106_2958, w_106_2964, w_106_2965, w_106_2967, w_106_2969, w_106_2973, w_106_2982, w_106_2984, w_106_2989, w_106_2996, w_106_2999, w_106_3001, w_106_3018, w_106_3019, w_106_3022, w_106_3031, w_106_3038, w_106_3041, w_106_3042, w_106_3045, w_106_3048, w_106_3052, w_106_3059, w_106_3062, w_106_3063, w_106_3064, w_106_3065, w_106_3066, w_106_3067, w_106_3068, w_106_3069, w_106_3070, w_106_3071, w_106_3073;
  wire w_107_001, w_107_004, w_107_007, w_107_009, w_107_011, w_107_014, w_107_015, w_107_016, w_107_024, w_107_025, w_107_026, w_107_029, w_107_032, w_107_035, w_107_038, w_107_040, w_107_041, w_107_044, w_107_046, w_107_047, w_107_050, w_107_051, w_107_054, w_107_057, w_107_058, w_107_060, w_107_062, w_107_064, w_107_071, w_107_073, w_107_074, w_107_076, w_107_078, w_107_079, w_107_081, w_107_083, w_107_084, w_107_085, w_107_086, w_107_087, w_107_094, w_107_095, w_107_098, w_107_099, w_107_103, w_107_104, w_107_105, w_107_106, w_107_107, w_107_108, w_107_110, w_107_111, w_107_112, w_107_115, w_107_116, w_107_118, w_107_119, w_107_121, w_107_122, w_107_125, w_107_127, w_107_129, w_107_131, w_107_132, w_107_134, w_107_137, w_107_141, w_107_142, w_107_144, w_107_146, w_107_148, w_107_149, w_107_152, w_107_153, w_107_154, w_107_155, w_107_158, w_107_160, w_107_164, w_107_165, w_107_166, w_107_170, w_107_173, w_107_174, w_107_178, w_107_179, w_107_181, w_107_182, w_107_191, w_107_196, w_107_197, w_107_198, w_107_199, w_107_200, w_107_203, w_107_210, w_107_212, w_107_214, w_107_216, w_107_218, w_107_220, w_107_221, w_107_223, w_107_224, w_107_230, w_107_231, w_107_234, w_107_241, w_107_243, w_107_244, w_107_245, w_107_246, w_107_248, w_107_255, w_107_256, w_107_257, w_107_258, w_107_260, w_107_261, w_107_264, w_107_265, w_107_268, w_107_270, w_107_271, w_107_273, w_107_277, w_107_282, w_107_283, w_107_284, w_107_287, w_107_290, w_107_291, w_107_294, w_107_295, w_107_297, w_107_298, w_107_300, w_107_302, w_107_305, w_107_307, w_107_308, w_107_309, w_107_310, w_107_311, w_107_313, w_107_315, w_107_318, w_107_319, w_107_320, w_107_322, w_107_325, w_107_326, w_107_327, w_107_328, w_107_330, w_107_331, w_107_332, w_107_333, w_107_336, w_107_337, w_107_338, w_107_339, w_107_340, w_107_342, w_107_343, w_107_347, w_107_349, w_107_352, w_107_353, w_107_356, w_107_357, w_107_358, w_107_362, w_107_364, w_107_366, w_107_368, w_107_369, w_107_372, w_107_373, w_107_374, w_107_376, w_107_377, w_107_383, w_107_384, w_107_385, w_107_386, w_107_388, w_107_393, w_107_395, w_107_396, w_107_399, w_107_402, w_107_406, w_107_409, w_107_414, w_107_419, w_107_421, w_107_423, w_107_427, w_107_428, w_107_430, w_107_431, w_107_437, w_107_438, w_107_444, w_107_446, w_107_447, w_107_448, w_107_450, w_107_453, w_107_456, w_107_457, w_107_461, w_107_462, w_107_465, w_107_467, w_107_472, w_107_475, w_107_477, w_107_478, w_107_479, w_107_482, w_107_486, w_107_487, w_107_489, w_107_490, w_107_493, w_107_497, w_107_498, w_107_501, w_107_504, w_107_505, w_107_506, w_107_508, w_107_510, w_107_515, w_107_516, w_107_518, w_107_520, w_107_521, w_107_522, w_107_523, w_107_526, w_107_527, w_107_529, w_107_531, w_107_532, w_107_535, w_107_536, w_107_537, w_107_538, w_107_541, w_107_545, w_107_547, w_107_548, w_107_550, w_107_551, w_107_553, w_107_557, w_107_560, w_107_564, w_107_568, w_107_569, w_107_570, w_107_576, w_107_577, w_107_578, w_107_579, w_107_580, w_107_584, w_107_585, w_107_587, w_107_588, w_107_590, w_107_591, w_107_594, w_107_595, w_107_597, w_107_603, w_107_607, w_107_609, w_107_611, w_107_613, w_107_614, w_107_615, w_107_616, w_107_619, w_107_620, w_107_624, w_107_625, w_107_629, w_107_630, w_107_631, w_107_632, w_107_633, w_107_634, w_107_636, w_107_642, w_107_644, w_107_645, w_107_646, w_107_647, w_107_648, w_107_652, w_107_658, w_107_660, w_107_661, w_107_665, w_107_667, w_107_668, w_107_669, w_107_670, w_107_672, w_107_673, w_107_676, w_107_677, w_107_678, w_107_679, w_107_680, w_107_681, w_107_684, w_107_685, w_107_688, w_107_691, w_107_693, w_107_695, w_107_696, w_107_697, w_107_698, w_107_699, w_107_700, w_107_701, w_107_703, w_107_704, w_107_705, w_107_707, w_107_708, w_107_710, w_107_711, w_107_713, w_107_714, w_107_716, w_107_717, w_107_720, w_107_721, w_107_723, w_107_726, w_107_727, w_107_728, w_107_729, w_107_733, w_107_734, w_107_738, w_107_743, w_107_748, w_107_751, w_107_752, w_107_754, w_107_756, w_107_757, w_107_759, w_107_760, w_107_761, w_107_763, w_107_768, w_107_772, w_107_775, w_107_776, w_107_777, w_107_787, w_107_788, w_107_789, w_107_791, w_107_792, w_107_793, w_107_796, w_107_797, w_107_800, w_107_806, w_107_807, w_107_808, w_107_812, w_107_814, w_107_815, w_107_816, w_107_818, w_107_819, w_107_822, w_107_829, w_107_831, w_107_832, w_107_833, w_107_834, w_107_839, w_107_840, w_107_841, w_107_845, w_107_847, w_107_852, w_107_853, w_107_855, w_107_860, w_107_864, w_107_877, w_107_880, w_107_882, w_107_898, w_107_901, w_107_909, w_107_913, w_107_920, w_107_930, w_107_934, w_107_940, w_107_941, w_107_946, w_107_952, w_107_956, w_107_958, w_107_969, w_107_971, w_107_973, w_107_975, w_107_978, w_107_980, w_107_981, w_107_984, w_107_990, w_107_991, w_107_993, w_107_994, w_107_998, w_107_1016, w_107_1024, w_107_1025, w_107_1037, w_107_1047, w_107_1048, w_107_1059, w_107_1061, w_107_1065, w_107_1069, w_107_1072, w_107_1075, w_107_1080, w_107_1082, w_107_1084, w_107_1087, w_107_1093, w_107_1096, w_107_1097, w_107_1098, w_107_1101, w_107_1103, w_107_1114, w_107_1138, w_107_1146, w_107_1148, w_107_1154, w_107_1156, w_107_1160, w_107_1170, w_107_1173, w_107_1183, w_107_1185, w_107_1190, w_107_1194, w_107_1202, w_107_1211, w_107_1212, w_107_1218, w_107_1219, w_107_1220, w_107_1221, w_107_1225, w_107_1228, w_107_1229, w_107_1230, w_107_1232, w_107_1233, w_107_1248, w_107_1251, w_107_1253, w_107_1254, w_107_1259, w_107_1262, w_107_1263, w_107_1268, w_107_1269, w_107_1270, w_107_1273, w_107_1274, w_107_1276, w_107_1277, w_107_1280, w_107_1287, w_107_1290, w_107_1301, w_107_1303, w_107_1304, w_107_1308, w_107_1311, w_107_1314, w_107_1323, w_107_1324, w_107_1325, w_107_1329, w_107_1330, w_107_1337, w_107_1338, w_107_1343, w_107_1347, w_107_1354, w_107_1361, w_107_1362, w_107_1363, w_107_1367, w_107_1369, w_107_1373, w_107_1377, w_107_1378, w_107_1389, w_107_1393, w_107_1398, w_107_1399, w_107_1401, w_107_1406, w_107_1417, w_107_1418, w_107_1431, w_107_1432, w_107_1433, w_107_1440, w_107_1445, w_107_1448, w_107_1452, w_107_1455, w_107_1460, w_107_1463, w_107_1466, w_107_1468, w_107_1469, w_107_1475, w_107_1478, w_107_1482, w_107_1489, w_107_1490, w_107_1494, w_107_1495, w_107_1497, w_107_1499, w_107_1501, w_107_1508, w_107_1509, w_107_1511, w_107_1517, w_107_1522, w_107_1527, w_107_1531, w_107_1534, w_107_1537, w_107_1540, w_107_1549, w_107_1555, w_107_1561, w_107_1562, w_107_1564, w_107_1566, w_107_1570, w_107_1571, w_107_1577, w_107_1578, w_107_1580, w_107_1581, w_107_1584, w_107_1589, w_107_1598, w_107_1599, w_107_1602, w_107_1604, w_107_1607, w_107_1611, w_107_1613, w_107_1614, w_107_1616, w_107_1619, w_107_1623, w_107_1624, w_107_1625, w_107_1628, w_107_1631, w_107_1633, w_107_1641, w_107_1642, w_107_1647, w_107_1654, w_107_1661, w_107_1667, w_107_1670, w_107_1681, w_107_1682, w_107_1685, w_107_1689, w_107_1691, w_107_1692, w_107_1694, w_107_1695, w_107_1700, w_107_1702, w_107_1708, w_107_1712, w_107_1713, w_107_1715, w_107_1716, w_107_1718, w_107_1725, w_107_1733, w_107_1735, w_107_1740, w_107_1745, w_107_1746, w_107_1751, w_107_1756, w_107_1757, w_107_1761, w_107_1762, w_107_1763, w_107_1771, w_107_1778, w_107_1779, w_107_1782, w_107_1796, w_107_1800, w_107_1802, w_107_1807, w_107_1811, w_107_1818, w_107_1819, w_107_1820, w_107_1821, w_107_1824, w_107_1827, w_107_1837, w_107_1838, w_107_1848, w_107_1849, w_107_1851, w_107_1852, w_107_1854, w_107_1858, w_107_1865, w_107_1868, w_107_1869, w_107_1872, w_107_1877, w_107_1878, w_107_1880, w_107_1881, w_107_1884, w_107_1890, w_107_1891, w_107_1897, w_107_1902, w_107_1904, w_107_1906, w_107_1910, w_107_1912, w_107_1913, w_107_1915, w_107_1917, w_107_1921, w_107_1924, w_107_1925, w_107_1926, w_107_1927, w_107_1931, w_107_1933, w_107_1934, w_107_1938, w_107_1943, w_107_1945, w_107_1948, w_107_1950, w_107_1955, w_107_1957, w_107_1964, w_107_1969, w_107_1970, w_107_1971, w_107_1973, w_107_1974, w_107_1981, w_107_1993, w_107_1994, w_107_1998, w_107_2005, w_107_2007, w_107_2008, w_107_2015, w_107_2017, w_107_2020, w_107_2021, w_107_2024, w_107_2029, w_107_2033, w_107_2042, w_107_2047, w_107_2048, w_107_2049, w_107_2050, w_107_2051, w_107_2054, w_107_2057, w_107_2058, w_107_2061, w_107_2072, w_107_2075, w_107_2077, w_107_2085, w_107_2086, w_107_2087, w_107_2089, w_107_2090, w_107_2093, w_107_2096, w_107_2098, w_107_2101, w_107_2106, w_107_2113, w_107_2119, w_107_2121, w_107_2122, w_107_2123, w_107_2126, w_107_2128, w_107_2131, w_107_2133, w_107_2136, w_107_2138, w_107_2139, w_107_2145, w_107_2146, w_107_2148, w_107_2152, w_107_2164, w_107_2166, w_107_2168, w_107_2170, w_107_2171, w_107_2173, w_107_2178, w_107_2179, w_107_2185, w_107_2192, w_107_2193, w_107_2196, w_107_2213, w_107_2219, w_107_2220, w_107_2222, w_107_2223, w_107_2225, w_107_2231, w_107_2235, w_107_2240, w_107_2241, w_107_2257, w_107_2259, w_107_2261, w_107_2266, w_107_2268, w_107_2269, w_107_2270, w_107_2272, w_107_2279, w_107_2281, w_107_2289, w_107_2290, w_107_2295, w_107_2298, w_107_2301, w_107_2302, w_107_2303, w_107_2304, w_107_2305, w_107_2306, w_107_2307, w_107_2309, w_107_2315, w_107_2318, w_107_2319, w_107_2320, w_107_2327, w_107_2332, w_107_2334, w_107_2340, w_107_2342, w_107_2349, w_107_2351, w_107_2355, w_107_2362, w_107_2364, w_107_2371, w_107_2374, w_107_2376, w_107_2380, w_107_2387, w_107_2392, w_107_2402, w_107_2403, w_107_2406, w_107_2411, w_107_2412, w_107_2413, w_107_2434, w_107_2440, w_107_2444, w_107_2447, w_107_2449, w_107_2457, w_107_2459, w_107_2464, w_107_2467, w_107_2471, w_107_2483, w_107_2484, w_107_2488, w_107_2489, w_107_2491, w_107_2496, w_107_2500, w_107_2506, w_107_2508, w_107_2509, w_107_2517, w_107_2528, w_107_2535, w_107_2541, w_107_2546, w_107_2547, w_107_2551, w_107_2559, w_107_2564, w_107_2565, w_107_2566, w_107_2569, w_107_2575, w_107_2576, w_107_2577, w_107_2578, w_107_2580, w_107_2586, w_107_2587, w_107_2588, w_107_2592, w_107_2597, w_107_2613, w_107_2616, w_107_2617, w_107_2622, w_107_2625, w_107_2634, w_107_2638, w_107_2641, w_107_2643, w_107_2649, w_107_2653, w_107_2654, w_107_2659, w_107_2662, w_107_2669, w_107_2671, w_107_2686, w_107_2696, w_107_2699, w_107_2700, w_107_2705, w_107_2717, w_107_2732, w_107_2733, w_107_2735, w_107_2739, w_107_2741, w_107_2744, w_107_2747, w_107_2748, w_107_2755, w_107_2769, w_107_2771, w_107_2774, w_107_2775, w_107_2776, w_107_2777, w_107_2778, w_107_2779, w_107_2783, w_107_2788, w_107_2795, w_107_2797, w_107_2798, w_107_2800, w_107_2804, w_107_2807, w_107_2814, w_107_2816, w_107_2817, w_107_2818, w_107_2824, w_107_2827, w_107_2828, w_107_2833, w_107_2836, w_107_2837, w_107_2840, w_107_2846, w_107_2847, w_107_2850, w_107_2852, w_107_2857, w_107_2858, w_107_2861, w_107_2863, w_107_2870, w_107_2872, w_107_2879, w_107_2883, w_107_2884, w_107_2893, w_107_2900, w_107_2908, w_107_2912, w_107_2913, w_107_2917, w_107_2921, w_107_2929, w_107_2935, w_107_2936, w_107_2957, w_107_2960, w_107_2964, w_107_2965, w_107_2966, w_107_2978, w_107_2980, w_107_2982, w_107_2983, w_107_2998, w_107_3001, w_107_3004, w_107_3005, w_107_3010, w_107_3018, w_107_3023, w_107_3025, w_107_3030, w_107_3033, w_107_3041, w_107_3042, w_107_3043, w_107_3044, w_107_3046, w_107_3048, w_107_3060, w_107_3064, w_107_3066, w_107_3068, w_107_3071, w_107_3074, w_107_3076, w_107_3083, w_107_3084, w_107_3089, w_107_3092, w_107_3095, w_107_3099, w_107_3108, w_107_3111, w_107_3113, w_107_3115, w_107_3116, w_107_3118, w_107_3119, w_107_3124, w_107_3125, w_107_3128, w_107_3134, w_107_3138, w_107_3140, w_107_3142, w_107_3145, w_107_3149, w_107_3150, w_107_3153, w_107_3154, w_107_3163, w_107_3164, w_107_3171, w_107_3172, w_107_3188, w_107_3195, w_107_3198, w_107_3208, w_107_3210, w_107_3211, w_107_3218, w_107_3222, w_107_3228, w_107_3247, w_107_3250, w_107_3251, w_107_3253, w_107_3254, w_107_3256, w_107_3259, w_107_3264, w_107_3267, w_107_3275, w_107_3278, w_107_3283, w_107_3284, w_107_3288, w_107_3290, w_107_3297, w_107_3303, w_107_3310, w_107_3311, w_107_3318, w_107_3320, w_107_3321, w_107_3335, w_107_3338, w_107_3341, w_107_3347, w_107_3349, w_107_3352, w_107_3356, w_107_3360, w_107_3362, w_107_3365, w_107_3366, w_107_3369, w_107_3370, w_107_3382, w_107_3386, w_107_3391, w_107_3402, w_107_3403, w_107_3404, w_107_3406, w_107_3412, w_107_3413, w_107_3416, w_107_3417, w_107_3422, w_107_3427, w_107_3431, w_107_3432, w_107_3436, w_107_3439, w_107_3446, w_107_3447, w_107_3448, w_107_3449, w_107_3452, w_107_3453, w_107_3456, w_107_3459, w_107_3462, w_107_3464, w_107_3465, w_107_3478, w_107_3486, w_107_3487, w_107_3491, w_107_3497, w_107_3501, w_107_3508, w_107_3514, w_107_3520, w_107_3523, w_107_3527, w_107_3528, w_107_3529, w_107_3532, w_107_3534, w_107_3539, w_107_3540, w_107_3549, w_107_3552, w_107_3560, w_107_3562, w_107_3565, w_107_3567, w_107_3568, w_107_3571, w_107_3576, w_107_3578, w_107_3587, w_107_3591, w_107_3592, w_107_3600, w_107_3611, w_107_3612, w_107_3614, w_107_3615, w_107_3631, w_107_3641, w_107_3645, w_107_3648, w_107_3654, w_107_3665, w_107_3667, w_107_3675, w_107_3678, w_107_3686, w_107_3699, w_107_3702, w_107_3705, w_107_3708, w_107_3711, w_107_3714, w_107_3719, w_107_3721, w_107_3728, w_107_3730, w_107_3733, w_107_3734, w_107_3741, w_107_3745, w_107_3747, w_107_3752, w_107_3753, w_107_3754, w_107_3765, w_107_3767, w_107_3771, w_107_3774, w_107_3785, w_107_3786, w_107_3788, w_107_3789, w_107_3796, w_107_3816, w_107_3819, w_107_3820, w_107_3832, w_107_3833, w_107_3834, w_107_3838, w_107_3844, w_107_3845, w_107_3853, w_107_3854, w_107_3857, w_107_3861, w_107_3868, w_107_3878, w_107_3884, w_107_3886, w_107_3889, w_107_3891, w_107_3893, w_107_3898, w_107_3899, w_107_3902, w_107_3903, w_107_3904, w_107_3906, w_107_3908, w_107_3909, w_107_3912, w_107_3917, w_107_3919, w_107_3927, w_107_3938, w_107_3943, w_107_3947, w_107_3950, w_107_3954, w_107_3957, w_107_3968, w_107_3971, w_107_3974, w_107_3975, w_107_3978, w_107_3983, w_107_3987, w_107_3997, w_107_4000, w_107_4004, w_107_4005, w_107_4009, w_107_4030, w_107_4033, w_107_4034, w_107_4038, w_107_4040, w_107_4047, w_107_4054, w_107_4063, w_107_4075, w_107_4078, w_107_4079, w_107_4080, w_107_4081, w_107_4085, w_107_4089, w_107_4090, w_107_4094, w_107_4095, w_107_4096, w_107_4097, w_107_4100, w_107_4103, w_107_4112, w_107_4114, w_107_4137, w_107_4138, w_107_4139, w_107_4140, w_107_4141, w_107_4145, w_107_4146, w_107_4147, w_107_4148, w_107_4149, w_107_4151;
  wire w_108_000, w_108_001, w_108_003, w_108_004, w_108_005, w_108_006, w_108_007, w_108_008, w_108_009, w_108_012, w_108_013, w_108_014, w_108_016, w_108_017, w_108_018, w_108_019, w_108_020, w_108_023, w_108_024, w_108_026, w_108_027, w_108_028, w_108_029, w_108_030, w_108_031, w_108_032, w_108_033, w_108_035, w_108_036, w_108_038, w_108_039, w_108_040, w_108_041, w_108_042, w_108_043, w_108_044, w_108_045, w_108_046, w_108_048, w_108_049, w_108_050, w_108_051, w_108_052, w_108_053, w_108_054, w_108_055, w_108_056, w_108_057, w_108_058, w_108_059, w_108_060, w_108_062, w_108_063, w_108_065, w_108_066, w_108_067, w_108_068, w_108_069, w_108_070, w_108_072, w_108_073, w_108_074, w_108_075, w_108_076, w_108_077, w_108_078, w_108_079, w_108_080, w_108_081, w_108_082, w_108_084, w_108_085, w_108_086, w_108_087, w_108_088, w_108_089, w_108_090, w_108_091, w_108_092, w_108_093, w_108_094, w_108_095, w_108_097, w_108_099, w_108_100, w_108_101, w_108_102, w_108_103, w_108_104, w_108_107, w_108_108, w_108_109, w_108_110, w_108_111, w_108_112, w_108_114, w_108_115, w_108_116, w_108_117, w_108_118, w_108_119, w_108_120, w_108_121, w_108_123, w_108_125, w_108_126, w_108_127, w_108_128, w_108_129, w_108_130, w_108_131, w_108_132, w_108_133, w_108_134, w_108_135, w_108_136, w_108_137, w_108_138, w_108_139, w_108_140, w_108_141, w_108_142, w_108_143, w_108_144, w_108_145, w_108_146, w_108_147, w_108_148, w_108_150, w_108_151, w_108_152, w_108_153, w_108_154, w_108_155, w_108_156, w_108_158, w_108_159, w_108_160, w_108_161, w_108_162, w_108_163, w_108_164, w_108_165, w_108_166, w_108_167, w_108_168, w_108_169, w_108_170, w_108_171, w_108_172, w_108_173, w_108_174, w_108_175, w_108_176, w_108_177, w_108_178, w_108_180, w_108_181, w_108_182, w_108_183, w_108_184, w_108_185, w_108_186, w_108_187, w_108_188, w_108_190, w_108_191, w_108_192, w_108_194, w_108_195, w_108_196, w_108_197, w_108_198, w_108_200, w_108_201, w_108_202, w_108_203, w_108_204, w_108_205, w_108_206, w_108_207, w_108_208, w_108_210, w_108_211, w_108_212, w_108_213, w_108_214, w_108_215, w_108_216, w_108_217, w_108_218, w_108_219, w_108_220, w_108_221, w_108_222, w_108_223, w_108_224, w_108_225, w_108_226, w_108_227, w_108_228, w_108_229, w_108_230, w_108_232, w_108_234, w_108_235, w_108_236, w_108_238, w_108_239, w_108_240, w_108_242, w_108_243, w_108_244, w_108_245, w_108_246, w_108_248, w_108_249, w_108_251, w_108_252, w_108_253, w_108_254, w_108_255, w_108_256, w_108_257, w_108_258, w_108_259, w_108_260, w_108_261, w_108_262, w_108_263, w_108_264, w_108_265, w_108_266, w_108_267, w_108_268, w_108_269, w_108_271, w_108_272, w_108_273, w_108_274, w_108_276, w_108_277, w_108_278, w_108_280, w_108_281, w_108_283, w_108_284, w_108_286, w_108_287, w_108_288, w_108_289, w_108_290, w_108_293, w_108_294, w_108_295, w_108_296, w_108_297, w_108_299, w_108_300, w_108_301, w_108_302, w_108_303, w_108_304, w_108_305, w_108_306, w_108_308, w_108_309, w_108_310, w_108_311, w_108_313, w_108_314, w_108_316, w_108_319, w_108_320, w_108_321, w_108_322, w_108_323, w_108_325, w_108_326, w_108_327, w_108_329, w_108_331, w_108_332, w_108_333, w_108_334, w_108_335, w_108_336, w_108_339, w_108_340, w_108_341, w_108_345, w_108_346, w_108_347, w_108_349, w_108_350, w_108_351, w_108_352, w_108_353, w_108_355, w_108_356, w_108_357, w_108_359, w_108_360, w_108_361, w_108_362, w_108_364, w_108_368, w_108_369, w_108_370, w_108_371, w_108_372, w_108_373, w_108_374, w_108_375, w_108_376, w_108_377, w_108_378, w_108_379, w_108_382, w_108_383, w_108_384, w_108_385, w_108_386, w_108_387, w_108_388, w_108_390, w_108_392, w_108_393, w_108_394, w_108_396, w_108_398, w_108_399, w_108_400, w_108_401, w_108_402, w_108_403, w_108_404, w_108_405, w_108_406, w_108_407, w_108_408, w_108_410, w_108_411, w_108_412, w_108_413, w_108_414, w_108_415, w_108_418, w_108_419, w_108_420, w_108_421, w_108_422, w_108_423, w_108_424, w_108_427, w_108_428, w_108_429, w_108_430, w_108_432, w_108_434, w_108_435, w_108_436, w_108_440, w_108_441, w_108_442, w_108_443, w_108_444, w_108_445, w_108_447, w_108_448, w_108_451, w_108_452, w_108_453, w_108_454, w_108_455, w_108_456, w_108_457, w_108_458, w_108_459, w_108_460, w_108_462, w_108_463, w_108_464, w_108_465, w_108_466, w_108_467, w_108_468, w_108_469, w_108_470, w_108_472, w_108_473, w_108_474, w_108_475, w_108_476, w_108_477, w_108_478, w_108_479, w_108_480, w_108_481, w_108_482, w_108_483, w_108_484, w_108_485, w_108_486, w_108_487, w_108_488, w_108_489, w_108_490, w_108_491, w_108_492, w_108_493, w_108_494, w_108_495, w_108_496, w_108_497, w_108_498, w_108_499, w_108_501, w_108_503, w_108_504, w_108_505, w_108_506, w_108_507, w_108_510, w_108_511, w_108_512, w_108_513, w_108_514, w_108_515, w_108_516, w_108_517, w_108_519, w_108_520, w_108_521, w_108_522, w_108_523, w_108_524, w_108_525, w_108_526, w_108_527, w_108_528, w_108_529, w_108_530, w_108_531, w_108_536, w_108_537, w_108_538, w_108_539, w_108_540, w_108_541, w_108_542, w_108_543, w_108_544, w_108_545, w_108_546, w_108_548, w_108_549, w_108_550, w_108_551, w_108_552, w_108_553, w_108_554, w_108_555, w_108_556, w_108_557, w_108_558, w_108_559, w_108_560, w_108_561, w_108_562, w_108_563, w_108_564, w_108_565, w_108_566, w_108_567, w_108_568, w_108_569, w_108_570, w_108_571, w_108_572, w_108_573, w_108_574, w_108_575, w_108_576, w_108_577, w_108_578, w_108_580, w_108_581, w_108_582, w_108_583, w_108_584, w_108_585, w_108_586, w_108_587, w_108_590, w_108_591, w_108_592, w_108_593, w_108_594, w_108_595, w_108_596, w_108_597, w_108_599, w_108_600, w_108_602, w_108_604, w_108_606, w_108_607, w_108_608, w_108_609, w_108_610, w_108_611, w_108_612, w_108_614, w_108_615, w_108_616, w_108_617, w_108_618, w_108_619, w_108_620, w_108_621, w_108_622, w_108_623, w_108_624, w_108_625, w_108_626, w_108_627, w_108_628, w_108_629, w_108_630, w_108_631, w_108_632, w_108_633, w_108_634, w_108_636, w_108_637, w_108_638, w_108_640, w_108_641, w_108_642, w_108_643, w_108_644, w_108_645, w_108_646, w_108_647, w_108_648, w_108_649, w_108_650, w_108_651, w_108_653, w_108_655, w_108_656, w_108_657, w_108_659, w_108_660, w_108_661, w_108_663, w_108_664, w_108_665, w_108_666, w_108_668, w_108_669, w_108_670, w_108_671, w_108_672, w_108_673, w_108_674, w_108_677, w_108_678, w_108_679, w_108_680, w_108_681, w_108_682, w_108_683, w_108_684, w_108_685, w_108_686, w_108_687, w_108_688, w_108_689, w_108_690, w_108_691, w_108_693, w_108_694, w_108_695, w_108_696, w_108_697, w_108_698, w_108_699, w_108_700, w_108_701, w_108_702, w_108_703, w_108_704, w_108_706, w_108_707, w_108_708, w_108_709, w_108_710, w_108_711, w_108_713, w_108_714, w_108_715, w_108_716, w_108_717, w_108_719, w_108_720, w_108_721, w_108_723, w_108_724, w_108_725, w_108_726, w_108_727, w_108_728, w_108_730, w_108_731, w_108_732, w_108_733, w_108_734, w_108_735, w_108_736, w_108_737, w_108_738, w_108_739, w_108_741, w_108_742, w_108_744, w_108_746, w_108_747, w_108_749, w_108_750, w_108_751, w_108_752, w_108_753, w_108_754, w_108_755, w_108_756, w_108_757, w_108_758, w_108_759, w_108_760, w_108_761, w_108_762, w_108_763, w_108_764, w_108_765, w_108_766, w_108_767, w_108_768, w_108_769, w_108_770, w_108_771, w_108_773, w_108_774, w_108_775, w_108_776, w_108_778, w_108_779, w_108_780, w_108_781, w_108_782, w_108_783, w_108_784, w_108_785, w_108_786, w_108_787, w_108_788, w_108_789, w_108_790, w_108_791, w_108_792, w_108_793, w_108_794, w_108_796, w_108_798, w_108_799, w_108_800, w_108_801, w_108_803, w_108_804, w_108_805, w_108_806, w_108_808, w_108_810, w_108_811, w_108_813, w_108_814, w_108_815, w_108_816, w_108_817, w_108_819, w_108_821, w_108_824, w_108_825, w_108_826, w_108_828, w_108_829, w_108_830, w_108_831, w_108_832, w_108_833, w_108_834, w_108_837, w_108_838, w_108_839, w_108_841, w_108_843, w_108_844, w_108_846, w_108_847, w_108_849, w_108_850, w_108_853, w_108_857, w_108_858, w_108_859, w_108_860, w_108_862, w_108_863, w_108_865, w_108_866, w_108_867, w_108_868;
  wire w_109_000, w_109_001, w_109_002, w_109_004, w_109_005, w_109_006, w_109_008, w_109_009, w_109_011, w_109_015, w_109_017, w_109_018, w_109_020, w_109_021, w_109_024, w_109_026, w_109_028, w_109_029, w_109_030, w_109_031, w_109_032, w_109_034, w_109_035, w_109_036, w_109_037, w_109_038, w_109_039, w_109_042, w_109_043, w_109_044, w_109_045, w_109_046, w_109_047, w_109_048, w_109_049, w_109_050, w_109_051, w_109_052, w_109_053, w_109_054, w_109_055, w_109_056, w_109_057, w_109_059, w_109_060, w_109_061, w_109_062, w_109_063, w_109_065, w_109_066, w_109_067, w_109_068, w_109_069, w_109_070, w_109_071, w_109_073, w_109_074, w_109_075, w_109_076, w_109_078, w_109_079, w_109_080, w_109_081, w_109_082, w_109_083, w_109_084, w_109_085, w_109_086, w_109_090, w_109_091, w_109_092, w_109_093, w_109_098, w_109_099, w_109_100, w_109_102, w_109_103, w_109_107, w_109_108, w_109_109, w_109_110, w_109_111, w_109_112, w_109_113, w_109_114, w_109_115, w_109_116, w_109_119, w_109_120, w_109_121, w_109_122, w_109_124, w_109_125, w_109_127, w_109_128, w_109_134, w_109_135, w_109_136, w_109_138, w_109_139, w_109_142, w_109_144, w_109_145, w_109_146, w_109_147, w_109_148, w_109_149, w_109_151, w_109_152, w_109_154, w_109_156, w_109_157, w_109_158, w_109_159, w_109_160, w_109_161, w_109_162, w_109_163, w_109_166, w_109_167, w_109_169, w_109_170, w_109_171, w_109_172, w_109_173, w_109_174, w_109_175, w_109_176, w_109_177, w_109_178, w_109_179, w_109_181, w_109_182, w_109_184, w_109_185, w_109_188, w_109_189, w_109_190, w_109_191, w_109_195, w_109_196, w_109_199, w_109_200, w_109_201, w_109_203, w_109_204, w_109_207, w_109_208, w_109_211, w_109_213, w_109_215, w_109_217, w_109_218, w_109_220, w_109_221, w_109_224, w_109_226, w_109_227, w_109_230, w_109_232, w_109_233, w_109_236, w_109_237, w_109_239, w_109_240, w_109_245, w_109_247, w_109_248, w_109_251, w_109_253, w_109_254, w_109_259, w_109_261, w_109_262, w_109_264, w_109_266, w_109_267, w_109_268, w_109_272, w_109_274, w_109_276, w_109_277, w_109_278, w_109_280, w_109_281, w_109_282, w_109_283, w_109_286, w_109_288, w_109_289, w_109_290, w_109_292, w_109_293, w_109_294, w_109_295, w_109_296, w_109_300, w_109_303, w_109_304, w_109_308, w_109_311, w_109_312, w_109_313, w_109_316, w_109_317, w_109_320, w_109_324, w_109_326, w_109_327, w_109_328, w_109_334, w_109_335, w_109_336, w_109_338, w_109_339, w_109_340, w_109_342, w_109_343, w_109_347, w_109_348, w_109_349, w_109_350, w_109_351, w_109_352, w_109_353, w_109_356, w_109_357, w_109_358, w_109_359, w_109_360, w_109_362, w_109_365, w_109_366, w_109_367, w_109_368, w_109_369, w_109_371, w_109_373, w_109_374, w_109_375, w_109_376, w_109_378, w_109_382, w_109_383, w_109_385, w_109_386, w_109_387, w_109_389, w_109_395, w_109_396, w_109_397, w_109_398, w_109_402, w_109_403, w_109_405, w_109_406, w_109_409, w_109_414, w_109_415, w_109_417, w_109_418, w_109_421, w_109_424, w_109_427, w_109_429, w_109_431, w_109_432, w_109_434, w_109_435, w_109_438, w_109_440, w_109_442, w_109_443, w_109_447, w_109_451, w_109_452, w_109_453, w_109_454, w_109_455, w_109_458, w_109_462, w_109_463, w_109_464, w_109_465, w_109_467, w_109_468, w_109_471, w_109_472, w_109_473, w_109_476, w_109_478, w_109_479, w_109_480, w_109_481, w_109_482, w_109_483, w_109_484, w_109_485, w_109_487, w_109_488, w_109_490, w_109_491, w_109_492, w_109_493, w_109_494, w_109_495, w_109_496, w_109_497, w_109_499, w_109_500, w_109_502, w_109_507, w_109_508, w_109_510, w_109_513, w_109_515, w_109_517, w_109_519, w_109_522, w_109_523, w_109_526, w_109_527, w_109_532, w_109_535, w_109_536, w_109_538, w_109_539, w_109_541, w_109_542, w_109_544, w_109_545, w_109_546, w_109_547, w_109_553, w_109_559, w_109_560, w_109_562, w_109_564, w_109_566, w_109_567, w_109_569, w_109_570, w_109_572, w_109_573, w_109_574, w_109_576, w_109_578, w_109_579, w_109_580, w_109_581, w_109_583, w_109_584, w_109_585, w_109_586, w_109_587, w_109_588, w_109_592, w_109_596, w_109_597, w_109_598, w_109_600, w_109_601, w_109_602, w_109_603, w_109_605, w_109_607, w_109_610, w_109_613, w_109_616, w_109_617, w_109_618, w_109_619, w_109_620, w_109_621, w_109_623, w_109_624, w_109_625, w_109_627, w_109_632, w_109_633, w_109_634, w_109_635, w_109_636, w_109_637, w_109_638, w_109_639, w_109_641, w_109_643, w_109_644, w_109_646, w_109_647, w_109_648, w_109_651, w_109_652, w_109_653, w_109_657, w_109_659, w_109_660, w_109_661, w_109_664, w_109_667, w_109_668, w_109_671, w_109_672, w_109_673, w_109_674, w_109_676, w_109_677, w_109_680, w_109_683, w_109_685, w_109_687, w_109_688, w_109_689, w_109_690, w_109_694, w_109_697, w_109_699, w_109_702, w_109_705, w_109_706, w_109_707, w_109_710, w_109_713, w_109_714, w_109_716, w_109_718, w_109_721, w_109_724, w_109_725, w_109_726, w_109_729, w_109_730, w_109_731, w_109_732, w_109_733, w_109_735, w_109_737, w_109_739, w_109_740, w_109_741, w_109_742, w_109_743, w_109_746, w_109_751, w_109_753, w_109_754, w_109_755, w_109_756, w_109_759, w_109_760, w_109_761, w_109_762, w_109_763, w_109_764, w_109_765, w_109_766, w_109_769, w_109_774, w_109_775, w_109_776, w_109_777, w_109_778, w_109_780, w_109_782, w_109_783, w_109_785, w_109_787, w_109_788, w_109_789, w_109_792, w_109_793, w_109_795, w_109_796, w_109_798, w_109_799, w_109_800, w_109_801, w_109_802, w_109_803, w_109_804, w_109_807, w_109_808, w_109_809, w_109_810, w_109_813, w_109_814, w_109_816, w_109_817, w_109_818, w_109_819, w_109_820, w_109_821, w_109_822, w_109_825, w_109_830, w_109_831, w_109_832, w_109_834, w_109_836, w_109_839, w_109_840, w_109_842, w_109_843, w_109_844, w_109_845, w_109_849, w_109_850, w_109_852, w_109_853, w_109_854, w_109_855, w_109_858, w_109_860, w_109_862, w_109_863, w_109_866, w_109_867, w_109_871, w_109_872, w_109_873, w_109_876, w_109_877, w_109_878, w_109_879, w_109_880, w_109_881, w_109_883, w_109_884, w_109_886, w_109_889, w_109_891, w_109_893, w_109_896, w_109_897, w_109_898, w_109_899, w_109_900, w_109_901, w_109_902, w_109_905, w_109_906, w_109_907, w_109_908, w_109_909, w_109_910, w_109_913, w_109_914, w_109_915, w_109_916, w_109_917, w_109_918, w_109_919, w_109_921, w_109_925, w_109_927, w_109_929, w_109_930, w_109_931, w_109_933, w_109_934, w_109_936, w_109_937, w_109_938, w_109_941, w_109_942, w_109_944, w_109_946, w_109_947, w_109_948, w_109_950, w_109_953, w_109_954, w_109_955, w_109_958, w_109_961, w_109_962, w_109_963, w_109_964, w_109_969, w_109_973, w_109_974, w_109_975, w_109_976, w_109_977, w_109_980, w_109_983, w_109_984, w_109_986, w_109_987, w_109_989, w_109_991, w_109_992, w_109_993, w_109_994, w_109_996, w_109_997, w_109_998, w_109_1000, w_109_1002, w_109_1003, w_109_1006, w_109_1007, w_109_1008, w_109_1010, w_109_1011, w_109_1012, w_109_1014, w_109_1019, w_109_1023, w_109_1024, w_109_1025, w_109_1026, w_109_1027, w_109_1028, w_109_1029, w_109_1030, w_109_1032, w_109_1033, w_109_1034, w_109_1036, w_109_1037, w_109_1038, w_109_1040, w_109_1041, w_109_1042, w_109_1045, w_109_1046, w_109_1047, w_109_1048, w_109_1051, w_109_1052, w_109_1053, w_109_1055, w_109_1056, w_109_1057, w_109_1058, w_109_1059, w_109_1060, w_109_1061, w_109_1066, w_109_1068, w_109_1070, w_109_1071, w_109_1072, w_109_1073, w_109_1074, w_109_1075, w_109_1076, w_109_1080, w_109_1081, w_109_1082, w_109_1083, w_109_1084, w_109_1086, w_109_1088, w_109_1089, w_109_1090, w_109_1091, w_109_1092, w_109_1099, w_109_1102, w_109_1103, w_109_1104, w_109_1105, w_109_1106, w_109_1107, w_109_1110, w_109_1111, w_109_1114, w_109_1115, w_109_1116, w_109_1118, w_109_1119, w_109_1120, w_109_1121, w_109_1122, w_109_1123, w_109_1124, w_109_1125, w_109_1126, w_109_1127, w_109_1129, w_109_1130, w_109_1131, w_109_1132, w_109_1133, w_109_1135, w_109_1136, w_109_1137, w_109_1139, w_109_1140, w_109_1141, w_109_1144, w_109_1145, w_109_1146, w_109_1147, w_109_1148, w_109_1149, w_109_1150, w_109_1154, w_109_1157, w_109_1158, w_109_1160, w_109_1164, w_109_1165, w_109_1168, w_109_1169, w_109_1170, w_109_1172, w_109_1173, w_109_1175, w_109_1176, w_109_1177, w_109_1178, w_109_1179, w_109_1180, w_109_1181, w_109_1182, w_109_1185, w_109_1187, w_109_1188, w_109_1189, w_109_1190, w_109_1192, w_109_1198, w_109_1202, w_109_1203, w_109_1204, w_109_1206, w_109_1208, w_109_1209, w_109_1210, w_109_1211, w_109_1212, w_109_1214, w_109_1215, w_109_1216, w_109_1217, w_109_1218, w_109_1219, w_109_1223, w_109_1224, w_109_1225, w_109_1227, w_109_1228, w_109_1229, w_109_1230, w_109_1232, w_109_1233, w_109_1234, w_109_1235, w_109_1237, w_109_1240, w_109_1241, w_109_1243, w_109_1244, w_109_1245, w_109_1250, w_109_1251, w_109_1254, w_109_1255, w_109_1259, w_109_1262, w_109_1266, w_109_1267, w_109_1268, w_109_1271, w_109_1272, w_109_1275, w_109_1277, w_109_1278, w_109_1280, w_109_1281, w_109_1282, w_109_1284, w_109_1287, w_109_1289, w_109_1290, w_109_1291, w_109_1292, w_109_1295, w_109_1297, w_109_1299, w_109_1300, w_109_1302, w_109_1303, w_109_1304, w_109_1305, w_109_1306, w_109_1308, w_109_1311, w_109_1315, w_109_1316, w_109_1317, w_109_1318, w_109_1323, w_109_1324, w_109_1325, w_109_1326, w_109_1327, w_109_1328, w_109_1330, w_109_1332, w_109_1334, w_109_1335, w_109_1336, w_109_1338, w_109_1339, w_109_1341, w_109_1342, w_109_1343, w_109_1344, w_109_1345, w_109_1348, w_109_1350, w_109_1354, w_109_1355, w_109_1357, w_109_1358, w_109_1359, w_109_1361, w_109_1362, w_109_1363, w_109_1365, w_109_1366, w_109_1367, w_109_1368, w_109_1371, w_109_1372, w_109_1373, w_109_1374, w_109_1377, w_109_1380, w_109_1383, w_109_1385, w_109_1389, w_109_1390, w_109_1391, w_109_1392, w_109_1393, w_109_1394, w_109_1396, w_109_1400, w_109_1403, w_109_1404, w_109_1405, w_109_1406, w_109_1408, w_109_1409, w_109_1413, w_109_1418, w_109_1425, w_109_1426, w_109_1427, w_109_1429, w_109_1431, w_109_1432, w_109_1434, w_109_1437, w_109_1438, w_109_1439, w_109_1441, w_109_1442, w_109_1445, w_109_1446, w_109_1448, w_109_1449, w_109_1453, w_109_1454, w_109_1455, w_109_1457, w_109_1461, w_109_1466, w_109_1472, w_109_1473, w_109_1474, w_109_1478, w_109_1479, w_109_1480, w_109_1481, w_109_1482, w_109_1487, w_109_1489, w_109_1490, w_109_1491, w_109_1492, w_109_1493, w_109_1494, w_109_1496, w_109_1497, w_109_1498, w_109_1499, w_109_1500, w_109_1501, w_109_1505, w_109_1507, w_109_1510, w_109_1514, w_109_1516, w_109_1517, w_109_1519, w_109_1520, w_109_1521, w_109_1524, w_109_1528, w_109_1529, w_109_1532, w_109_1533, w_109_1534, w_109_1535, w_109_1536, w_109_1537, w_109_1539, w_109_1540, w_109_1542, w_109_1543, w_109_1545, w_109_1546, w_109_1547, w_109_1548, w_109_1552, w_109_1554, w_109_1555, w_109_1556, w_109_1559, w_109_1561, w_109_1562, w_109_1564, w_109_1566, w_109_1567, w_109_1568, w_109_1569, w_109_1570, w_109_1572, w_109_1575, w_109_1576, w_109_1577, w_109_1578, w_109_1579, w_109_1582, w_109_1583, w_109_1585, w_109_1590, w_109_1593, w_109_1597, w_109_1598, w_109_1602, w_109_1603, w_109_1604, w_109_1605, w_109_1606, w_109_1607, w_109_1608, w_109_1609, w_109_1610, w_109_1614, w_109_1615, w_109_1616, w_109_1617, w_109_1618, w_109_1619, w_109_1620, w_109_1621, w_109_1625, w_109_1626, w_109_1627, w_109_1629;
  wire w_110_000, w_110_001, w_110_002, w_110_003, w_110_005, w_110_006, w_110_007, w_110_008, w_110_009, w_110_010, w_110_011, w_110_012, w_110_013, w_110_014, w_110_015, w_110_016, w_110_017, w_110_018, w_110_019, w_110_020, w_110_021, w_110_022, w_110_023, w_110_024, w_110_025, w_110_026, w_110_027, w_110_028, w_110_029, w_110_030, w_110_031, w_110_032, w_110_033, w_110_035, w_110_037, w_110_038, w_110_039, w_110_040, w_110_041, w_110_043, w_110_044, w_110_045, w_110_047, w_110_048, w_110_050, w_110_051, w_110_052, w_110_053, w_110_054, w_110_055, w_110_057, w_110_058, w_110_059, w_110_060, w_110_061, w_110_062, w_110_063, w_110_064, w_110_065, w_110_068, w_110_069, w_110_070, w_110_071, w_110_072, w_110_073, w_110_074, w_110_075, w_110_076, w_110_078, w_110_079, w_110_080, w_110_081, w_110_082, w_110_083, w_110_084, w_110_085, w_110_086, w_110_087, w_110_088, w_110_089, w_110_090, w_110_091, w_110_092, w_110_093, w_110_095, w_110_096, w_110_097, w_110_098, w_110_099, w_110_100, w_110_102, w_110_104, w_110_105, w_110_107, w_110_108, w_110_109, w_110_110, w_110_111, w_110_112, w_110_113, w_110_114, w_110_115, w_110_116, w_110_117, w_110_118, w_110_119, w_110_120, w_110_121, w_110_122, w_110_123, w_110_124, w_110_125, w_110_127, w_110_128, w_110_129, w_110_130, w_110_131, w_110_133, w_110_134, w_110_135, w_110_136, w_110_138, w_110_139, w_110_140, w_110_141, w_110_144, w_110_145, w_110_147, w_110_148, w_110_149, w_110_150, w_110_151, w_110_152, w_110_153, w_110_154, w_110_155, w_110_156, w_110_157, w_110_159, w_110_162, w_110_164, w_110_165, w_110_166, w_110_167, w_110_169, w_110_170, w_110_171, w_110_172, w_110_173, w_110_174, w_110_175, w_110_176, w_110_177, w_110_178, w_110_179, w_110_180, w_110_181, w_110_182, w_110_184, w_110_185, w_110_187, w_110_188, w_110_189, w_110_190, w_110_191, w_110_192, w_110_193, w_110_194, w_110_195, w_110_196, w_110_197, w_110_199, w_110_200, w_110_201, w_110_202, w_110_203, w_110_204, w_110_205, w_110_206, w_110_207, w_110_208, w_110_209, w_110_210, w_110_211, w_110_212, w_110_213, w_110_214, w_110_215, w_110_216, w_110_217, w_110_218, w_110_219, w_110_221, w_110_222, w_110_223, w_110_224, w_110_225, w_110_226, w_110_227, w_110_229, w_110_230, w_110_231, w_110_232, w_110_233, w_110_234, w_110_235, w_110_236, w_110_237, w_110_238, w_110_239, w_110_240, w_110_241, w_110_242, w_110_243, w_110_244, w_110_245, w_110_246, w_110_247, w_110_248, w_110_249, w_110_250, w_110_251, w_110_252, w_110_253, w_110_254, w_110_255, w_110_256, w_110_257, w_110_258, w_110_259, w_110_260, w_110_261, w_110_262, w_110_263, w_110_264, w_110_265, w_110_266, w_110_267, w_110_268, w_110_269, w_110_270, w_110_271, w_110_274, w_110_276, w_110_277, w_110_278, w_110_279, w_110_280, w_110_281, w_110_282, w_110_283, w_110_285, w_110_286, w_110_287, w_110_288, w_110_289, w_110_290, w_110_291, w_110_293, w_110_294, w_110_295, w_110_298, w_110_299, w_110_300, w_110_301, w_110_302, w_110_303, w_110_304, w_110_305, w_110_306, w_110_307, w_110_308, w_110_309, w_110_311, w_110_312, w_110_313, w_110_315, w_110_316, w_110_317, w_110_318, w_110_319, w_110_321, w_110_323, w_110_324, w_110_326, w_110_328, w_110_329, w_110_331, w_110_332, w_110_334, w_110_335, w_110_336, w_110_337, w_110_338, w_110_339, w_110_340, w_110_342, w_110_343, w_110_345, w_110_346, w_110_347, w_110_348, w_110_349, w_110_351, w_110_352, w_110_353, w_110_354, w_110_355, w_110_356, w_110_358, w_110_360, w_110_361, w_110_362, w_110_363, w_110_364, w_110_365, w_110_366, w_110_367, w_110_368, w_110_369, w_110_370, w_110_371, w_110_372, w_110_373, w_110_374, w_110_375, w_110_376, w_110_377, w_110_379, w_110_380, w_110_381, w_110_383, w_110_384, w_110_385, w_110_386, w_110_388, w_110_389, w_110_390, w_110_391, w_110_392, w_110_393, w_110_395, w_110_396, w_110_397, w_110_398, w_110_399, w_110_401, w_110_402, w_110_403, w_110_404, w_110_406, w_110_407, w_110_409, w_110_410, w_110_411, w_110_412, w_110_413, w_110_414, w_110_415, w_110_416, w_110_417, w_110_418, w_110_419, w_110_420, w_110_421, w_110_422, w_110_423, w_110_425, w_110_426, w_110_427, w_110_429, w_110_430, w_110_433, w_110_434, w_110_435, w_110_436, w_110_437, w_110_438, w_110_439, w_110_440, w_110_441, w_110_444, w_110_446, w_110_447, w_110_448, w_110_450, w_110_451, w_110_453, w_110_454, w_110_455, w_110_457, w_110_458, w_110_459, w_110_460, w_110_461, w_110_463, w_110_464, w_110_465, w_110_466, w_110_467, w_110_472, w_110_473, w_110_475, w_110_476, w_110_478, w_110_479, w_110_480, w_110_481, w_110_482, w_110_484, w_110_485, w_110_486, w_110_487, w_110_488, w_110_489, w_110_491, w_110_492, w_110_493, w_110_494, w_110_496, w_110_497, w_110_498, w_110_499, w_110_500, w_110_501, w_110_502, w_110_503, w_110_504, w_110_506, w_110_507, w_110_508, w_110_509, w_110_510, w_110_511, w_110_512, w_110_513, w_110_514, w_110_515, w_110_516, w_110_517, w_110_518, w_110_519, w_110_520, w_110_521, w_110_522, w_110_523, w_110_524, w_110_525, w_110_526, w_110_528, w_110_529, w_110_530, w_110_531, w_110_532, w_110_533, w_110_534, w_110_535, w_110_537, w_110_539, w_110_540, w_110_541, w_110_542, w_110_544, w_110_545, w_110_546, w_110_547, w_110_548, w_110_549, w_110_550, w_110_551, w_110_552, w_110_554, w_110_555, w_110_556, w_110_557, w_110_558, w_110_560, w_110_561, w_110_563, w_110_564, w_110_565, w_110_567, w_110_568, w_110_569, w_110_571, w_110_572, w_110_574, w_110_575, w_110_576, w_110_578, w_110_579, w_110_580, w_110_581, w_110_582, w_110_583, w_110_584, w_110_585, w_110_587, w_110_590, w_110_591, w_110_593, w_110_594, w_110_595, w_110_596, w_110_597, w_110_600, w_110_601, w_110_603, w_110_605, w_110_608, w_110_609, w_110_610, w_110_611, w_110_612, w_110_613, w_110_614, w_110_615, w_110_616, w_110_617, w_110_619, w_110_620, w_110_621, w_110_622, w_110_623, w_110_624, w_110_626, w_110_627, w_110_628, w_110_629, w_110_630, w_110_631, w_110_632, w_110_633, w_110_634, w_110_635, w_110_636, w_110_637, w_110_638, w_110_640, w_110_641, w_110_642, w_110_643, w_110_644, w_110_646, w_110_648, w_110_649, w_110_650, w_110_652, w_110_653, w_110_655, w_110_656, w_110_657, w_110_658, w_110_659, w_110_661, w_110_662, w_110_663, w_110_664, w_110_665, w_110_666, w_110_667, w_110_669, w_110_671, w_110_673, w_110_674, w_110_675, w_110_676, w_110_677, w_110_678, w_110_679, w_110_680, w_110_682, w_110_683, w_110_684, w_110_685, w_110_690, w_110_691, w_110_693, w_110_694, w_110_695, w_110_696, w_110_698, w_110_699, w_110_700, w_110_701, w_110_702, w_110_703, w_110_705, w_110_706, w_110_707, w_110_709, w_110_710, w_110_711, w_110_712, w_110_713, w_110_714, w_110_715, w_110_716, w_110_717, w_110_718, w_110_720, w_110_723, w_110_724, w_110_725, w_110_727, w_110_729, w_110_730, w_110_731, w_110_733, w_110_734, w_110_736, w_110_737, w_110_739, w_110_740, w_110_742, w_110_743, w_110_744, w_110_745, w_110_748, w_110_749, w_110_750, w_110_751, w_110_752, w_110_753, w_110_756, w_110_757, w_110_758, w_110_759, w_110_761, w_110_762, w_110_763, w_110_764, w_110_766, w_110_767, w_110_768, w_110_769, w_110_771, w_110_772, w_110_774, w_110_775, w_110_777, w_110_778, w_110_779, w_110_780, w_110_781, w_110_783, w_110_784, w_110_785, w_110_786, w_110_787, w_110_788, w_110_789, w_110_790, w_110_791, w_110_792, w_110_796, w_110_797, w_110_798, w_110_799, w_110_800, w_110_801, w_110_802, w_110_803, w_110_804, w_110_805, w_110_807;
  wire w_111_000, w_111_002, w_111_005, w_111_007, w_111_008, w_111_011, w_111_012, w_111_013, w_111_014, w_111_017, w_111_019, w_111_020, w_111_022, w_111_024, w_111_029, w_111_030, w_111_034, w_111_035, w_111_037, w_111_038, w_111_039, w_111_042, w_111_043, w_111_044, w_111_049, w_111_051, w_111_052, w_111_055, w_111_056, w_111_057, w_111_058, w_111_059, w_111_063, w_111_065, w_111_066, w_111_067, w_111_074, w_111_075, w_111_077, w_111_078, w_111_083, w_111_084, w_111_085, w_111_087, w_111_090, w_111_091, w_111_092, w_111_094, w_111_097, w_111_099, w_111_103, w_111_105, w_111_106, w_111_108, w_111_109, w_111_113, w_111_115, w_111_116, w_111_118, w_111_119, w_111_120, w_111_122, w_111_124, w_111_131, w_111_132, w_111_135, w_111_137, w_111_138, w_111_140, w_111_145, w_111_146, w_111_147, w_111_151, w_111_154, w_111_162, w_111_170, w_111_172, w_111_174, w_111_175, w_111_177, w_111_180, w_111_181, w_111_185, w_111_189, w_111_193, w_111_194, w_111_195, w_111_196, w_111_198, w_111_201, w_111_202, w_111_203, w_111_206, w_111_208, w_111_209, w_111_211, w_111_212, w_111_214, w_111_215, w_111_217, w_111_222, w_111_223, w_111_224, w_111_227, w_111_230, w_111_233, w_111_234, w_111_235, w_111_238, w_111_239, w_111_242, w_111_243, w_111_244, w_111_245, w_111_246, w_111_249, w_111_250, w_111_251, w_111_252, w_111_254, w_111_257, w_111_259, w_111_261, w_111_262, w_111_265, w_111_269, w_111_278, w_111_286, w_111_287, w_111_288, w_111_289, w_111_291, w_111_293, w_111_294, w_111_297, w_111_299, w_111_306, w_111_307, w_111_308, w_111_312, w_111_313, w_111_314, w_111_318, w_111_320, w_111_321, w_111_322, w_111_323, w_111_324, w_111_325, w_111_328, w_111_333, w_111_335, w_111_337, w_111_338, w_111_340, w_111_341, w_111_342, w_111_344, w_111_348, w_111_349, w_111_354, w_111_355, w_111_356, w_111_357, w_111_359, w_111_360, w_111_361, w_111_364, w_111_368, w_111_369, w_111_371, w_111_375, w_111_376, w_111_378, w_111_380, w_111_381, w_111_382, w_111_383, w_111_385, w_111_386, w_111_392, w_111_393, w_111_394, w_111_398, w_111_399, w_111_400, w_111_401, w_111_405, w_111_407, w_111_409, w_111_420, w_111_421, w_111_422, w_111_425, w_111_433, w_111_435, w_111_439, w_111_441, w_111_445, w_111_447, w_111_455, w_111_458, w_111_461, w_111_462, w_111_469, w_111_471, w_111_475, w_111_483, w_111_485, w_111_488, w_111_492, w_111_497, w_111_502, w_111_503, w_111_505, w_111_508, w_111_509, w_111_511, w_111_513, w_111_514, w_111_523, w_111_525, w_111_535, w_111_536, w_111_537, w_111_538, w_111_559, w_111_561, w_111_565, w_111_577, w_111_581, w_111_583, w_111_585, w_111_594, w_111_600, w_111_601, w_111_615, w_111_616, w_111_620, w_111_630, w_111_632, w_111_634, w_111_637, w_111_639, w_111_641, w_111_648, w_111_649, w_111_662, w_111_663, w_111_672, w_111_674, w_111_676, w_111_678, w_111_691, w_111_693, w_111_694, w_111_700, w_111_707, w_111_708, w_111_716, w_111_718, w_111_720, w_111_723, w_111_725, w_111_729, w_111_732, w_111_734, w_111_735, w_111_736, w_111_738, w_111_739, w_111_746, w_111_756, w_111_763, w_111_767, w_111_779, w_111_783, w_111_786, w_111_789, w_111_796, w_111_798, w_111_799, w_111_803, w_111_810, w_111_819, w_111_820, w_111_824, w_111_830, w_111_834, w_111_839, w_111_847, w_111_850, w_111_852, w_111_853, w_111_854, w_111_855, w_111_857, w_111_861, w_111_862, w_111_872, w_111_873, w_111_877, w_111_880, w_111_881, w_111_889, w_111_890, w_111_895, w_111_897, w_111_902, w_111_910, w_111_916, w_111_918, w_111_920, w_111_924, w_111_925, w_111_926, w_111_931, w_111_940, w_111_946, w_111_951, w_111_963, w_111_967, w_111_969, w_111_970, w_111_972, w_111_976, w_111_982, w_111_988, w_111_994, w_111_999, w_111_1002, w_111_1009, w_111_1012, w_111_1018, w_111_1027, w_111_1029, w_111_1035, w_111_1042, w_111_1063, w_111_1064, w_111_1068, w_111_1071, w_111_1072, w_111_1073, w_111_1074, w_111_1078, w_111_1081, w_111_1084, w_111_1085, w_111_1087, w_111_1091, w_111_1095, w_111_1096, w_111_1108, w_111_1111, w_111_1112, w_111_1116, w_111_1120, w_111_1125, w_111_1130, w_111_1131, w_111_1134, w_111_1135, w_111_1138, w_111_1139, w_111_1141, w_111_1145, w_111_1147, w_111_1149, w_111_1150, w_111_1152, w_111_1155, w_111_1169, w_111_1171, w_111_1181, w_111_1184, w_111_1185, w_111_1187, w_111_1188, w_111_1194, w_111_1195, w_111_1198, w_111_1199, w_111_1202, w_111_1204, w_111_1206, w_111_1210, w_111_1214, w_111_1226, w_111_1229, w_111_1232, w_111_1233, w_111_1234, w_111_1237, w_111_1239, w_111_1241, w_111_1244, w_111_1251, w_111_1252, w_111_1254, w_111_1261, w_111_1264, w_111_1268, w_111_1270, w_111_1273, w_111_1286, w_111_1294, w_111_1298, w_111_1301, w_111_1302, w_111_1304, w_111_1307, w_111_1311, w_111_1314, w_111_1315, w_111_1317, w_111_1326, w_111_1328, w_111_1329, w_111_1330, w_111_1331, w_111_1332, w_111_1333, w_111_1343, w_111_1349, w_111_1355, w_111_1364, w_111_1369, w_111_1373, w_111_1376, w_111_1381, w_111_1383, w_111_1386, w_111_1398, w_111_1407, w_111_1408, w_111_1413, w_111_1414, w_111_1420, w_111_1435, w_111_1439, w_111_1445, w_111_1448, w_111_1449, w_111_1452, w_111_1455, w_111_1457, w_111_1458, w_111_1459, w_111_1462, w_111_1465, w_111_1466, w_111_1467, w_111_1469, w_111_1470, w_111_1471, w_111_1478, w_111_1495, w_111_1498, w_111_1508, w_111_1514, w_111_1518, w_111_1524, w_111_1527, w_111_1528, w_111_1530, w_111_1532, w_111_1537, w_111_1539, w_111_1542, w_111_1551, w_111_1555, w_111_1558, w_111_1559, w_111_1560, w_111_1561, w_111_1562, w_111_1568, w_111_1569, w_111_1571, w_111_1575, w_111_1590, w_111_1592, w_111_1594, w_111_1598, w_111_1603, w_111_1618, w_111_1624, w_111_1625, w_111_1637, w_111_1640, w_111_1644, w_111_1645, w_111_1649, w_111_1655, w_111_1657, w_111_1665, w_111_1670, w_111_1673, w_111_1677, w_111_1685, w_111_1693, w_111_1694, w_111_1696, w_111_1702, w_111_1707, w_111_1710, w_111_1712, w_111_1716, w_111_1721, w_111_1733, w_111_1738, w_111_1743, w_111_1744, w_111_1745, w_111_1747, w_111_1748, w_111_1758, w_111_1762, w_111_1767, w_111_1770, w_111_1773, w_111_1775, w_111_1781, w_111_1782, w_111_1786, w_111_1791, w_111_1795, w_111_1805, w_111_1810, w_111_1812, w_111_1815, w_111_1818, w_111_1832, w_111_1840, w_111_1848, w_111_1855, w_111_1856, w_111_1857, w_111_1859, w_111_1862, w_111_1864, w_111_1870, w_111_1871, w_111_1872, w_111_1874, w_111_1878, w_111_1879, w_111_1880, w_111_1893, w_111_1894, w_111_1903, w_111_1904, w_111_1906, w_111_1908, w_111_1915, w_111_1919, w_111_1928, w_111_1931, w_111_1935, w_111_1939, w_111_1942, w_111_1950, w_111_1958, w_111_1960, w_111_1961, w_111_1962, w_111_1970, w_111_1976, w_111_1978, w_111_1985, w_111_1987, w_111_1988, w_111_1989, w_111_1991, w_111_1992, w_111_1995, w_111_1996, w_111_1997, w_111_1998, w_111_2001, w_111_2006, w_111_2009, w_111_2017, w_111_2023, w_111_2027, w_111_2028, w_111_2034, w_111_2043, w_111_2046, w_111_2049, w_111_2051, w_111_2052, w_111_2053, w_111_2068, w_111_2070, w_111_2071, w_111_2072, w_111_2075, w_111_2076, w_111_2080, w_111_2082, w_111_2083, w_111_2089, w_111_2091, w_111_2101, w_111_2103, w_111_2111, w_111_2115, w_111_2124, w_111_2125, w_111_2129, w_111_2130, w_111_2136, w_111_2148, w_111_2151, w_111_2152, w_111_2155, w_111_2159, w_111_2170, w_111_2171, w_111_2177, w_111_2183, w_111_2185, w_111_2188, w_111_2191, w_111_2193, w_111_2201, w_111_2204, w_111_2205, w_111_2212, w_111_2216, w_111_2230, w_111_2231, w_111_2247, w_111_2253, w_111_2268, w_111_2271, w_111_2272, w_111_2276, w_111_2283, w_111_2284, w_111_2292, w_111_2309, w_111_2312, w_111_2313, w_111_2316, w_111_2320, w_111_2336, w_111_2338, w_111_2339, w_111_2342, w_111_2346, w_111_2347, w_111_2348, w_111_2349, w_111_2360, w_111_2362, w_111_2373, w_111_2374, w_111_2378, w_111_2394, w_111_2395, w_111_2401, w_111_2411, w_111_2424, w_111_2427, w_111_2428, w_111_2429, w_111_2440, w_111_2443, w_111_2445, w_111_2446, w_111_2448, w_111_2458, w_111_2464, w_111_2466, w_111_2468, w_111_2475, w_111_2478, w_111_2481, w_111_2485, w_111_2487, w_111_2491, w_111_2496, w_111_2498, w_111_2502, w_111_2503, w_111_2509, w_111_2510, w_111_2512, w_111_2515, w_111_2518, w_111_2531, w_111_2545, w_111_2546, w_111_2550, w_111_2561, w_111_2563, w_111_2570, w_111_2575, w_111_2580, w_111_2581, w_111_2584, w_111_2586, w_111_2597, w_111_2600, w_111_2602, w_111_2610, w_111_2612, w_111_2613, w_111_2614, w_111_2625, w_111_2626, w_111_2629, w_111_2631, w_111_2633, w_111_2645, w_111_2646, w_111_2650, w_111_2652, w_111_2654, w_111_2660, w_111_2663, w_111_2664, w_111_2677, w_111_2682, w_111_2686, w_111_2687, w_111_2693, w_111_2694, w_111_2700, w_111_2705, w_111_2706, w_111_2710, w_111_2719, w_111_2726, w_111_2727, w_111_2729, w_111_2733, w_111_2745, w_111_2748, w_111_2754, w_111_2755, w_111_2758, w_111_2759, w_111_2760, w_111_2765, w_111_2766, w_111_2768, w_111_2776, w_111_2778, w_111_2779, w_111_2781, w_111_2790, w_111_2795, w_111_2799, w_111_2803, w_111_2815, w_111_2816, w_111_2817, w_111_2819, w_111_2833, w_111_2835, w_111_2838, w_111_2848, w_111_2854, w_111_2856, w_111_2857, w_111_2863, w_111_2868, w_111_2869, w_111_2871, w_111_2872, w_111_2879, w_111_2885, w_111_2886, w_111_2890, w_111_2891, w_111_2893, w_111_2895, w_111_2896, w_111_2897, w_111_2900, w_111_2901, w_111_2903, w_111_2908, w_111_2920, w_111_2925, w_111_2929, w_111_2933, w_111_2934, w_111_2942, w_111_2953, w_111_2961, w_111_2964, w_111_2965, w_111_2966, w_111_2969, w_111_2970, w_111_2975, w_111_2978, w_111_2984, w_111_2985, w_111_2987, w_111_2989, w_111_2992, w_111_2994, w_111_3000, w_111_3001, w_111_3002, w_111_3004, w_111_3010, w_111_3012, w_111_3016, w_111_3029, w_111_3030, w_111_3031, w_111_3036, w_111_3039, w_111_3048, w_111_3050, w_111_3051, w_111_3052, w_111_3055, w_111_3056, w_111_3058, w_111_3059, w_111_3061, w_111_3063, w_111_3065, w_111_3073, w_111_3076, w_111_3078, w_111_3086, w_111_3094, w_111_3096, w_111_3101, w_111_3108, w_111_3110, w_111_3112, w_111_3117, w_111_3122, w_111_3123, w_111_3125, w_111_3130, w_111_3131, w_111_3138, w_111_3139, w_111_3140, w_111_3143, w_111_3145, w_111_3146, w_111_3152, w_111_3154, w_111_3157, w_111_3160, w_111_3165, w_111_3171, w_111_3175, w_111_3177, w_111_3178, w_111_3181, w_111_3185, w_111_3202, w_111_3203, w_111_3205, w_111_3212, w_111_3216, w_111_3221, w_111_3225, w_111_3228, w_111_3231, w_111_3240, w_111_3251, w_111_3256, w_111_3260, w_111_3261, w_111_3270, w_111_3271, w_111_3272, w_111_3273, w_111_3274, w_111_3282, w_111_3283, w_111_3285, w_111_3293, w_111_3294, w_111_3298, w_111_3304, w_111_3305, w_111_3308, w_111_3313, w_111_3315, w_111_3323, w_111_3325, w_111_3327, w_111_3328, w_111_3329, w_111_3330, w_111_3333, w_111_3336, w_111_3338, w_111_3345, w_111_3350, w_111_3368, w_111_3379, w_111_3380, w_111_3383, w_111_3395, w_111_3402, w_111_3404, w_111_3410, w_111_3413, w_111_3414, w_111_3419, w_111_3425, w_111_3431, w_111_3433, w_111_3434, w_111_3439, w_111_3441, w_111_3451, w_111_3457, w_111_3462, w_111_3465, w_111_3468, w_111_3473, w_111_3477, w_111_3482, w_111_3488, w_111_3491, w_111_3492, w_111_3493, w_111_3494, w_111_3498, w_111_3499, w_111_3500, w_111_3501, w_111_3503, w_111_3508, w_111_3510, w_111_3516, w_111_3521, w_111_3522, w_111_3523, w_111_3530, w_111_3531, w_111_3532, w_111_3554, w_111_3566, w_111_3570, w_111_3575, w_111_3585, w_111_3594, w_111_3598, w_111_3608, w_111_3609, w_111_3611, w_111_3612, w_111_3614, w_111_3616, w_111_3623, w_111_3628, w_111_3634, w_111_3635, w_111_3636, w_111_3637, w_111_3640, w_111_3646, w_111_3651, w_111_3659, w_111_3661, w_111_3662, w_111_3665, w_111_3666, w_111_3668, w_111_3670, w_111_3672, w_111_3685, w_111_3686, w_111_3687, w_111_3689, w_111_3692, w_111_3700, w_111_3705, w_111_3715, w_111_3723, w_111_3724, w_111_3727, w_111_3734, w_111_3735, w_111_3737, w_111_3739, w_111_3740, w_111_3744, w_111_3745, w_111_3750, w_111_3754, w_111_3758, w_111_3764, w_111_3765, w_111_3767, w_111_3768, w_111_3770, w_111_3772, w_111_3773, w_111_3775, w_111_3785, w_111_3786, w_111_3790, w_111_3792, w_111_3794, w_111_3799, w_111_3801, w_111_3802, w_111_3806, w_111_3808, w_111_3812, w_111_3813, w_111_3822, w_111_3836, w_111_3837, w_111_3851, w_111_3860, w_111_3862, w_111_3872, w_111_3876, w_111_3879, w_111_3887, w_111_3888, w_111_3891, w_111_3893, w_111_3896, w_111_3899, w_111_3905, w_111_3906, w_111_3912, w_111_3922, w_111_3923, w_111_3928, w_111_3937, w_111_3941, w_111_3945, w_111_3954, w_111_3955, w_111_3956, w_111_3957, w_111_3958, w_111_3967, w_111_3968, w_111_3970, w_111_3972, w_111_3975, w_111_3977, w_111_3979, w_111_3982, w_111_3983, w_111_3994, w_111_3998, w_111_4005, w_111_4007, w_111_4008, w_111_4012, w_111_4017, w_111_4032, w_111_4035, w_111_4051, w_111_4053, w_111_4057, w_111_4059, w_111_4061, w_111_4065, w_111_4066, w_111_4075, w_111_4083, w_111_4086, w_111_4087, w_111_4089, w_111_4090, w_111_4098, w_111_4099, w_111_4105, w_111_4108, w_111_4110, w_111_4112, w_111_4118, w_111_4122, w_111_4124, w_111_4125, w_111_4134, w_111_4143, w_111_4151, w_111_4154, w_111_4157, w_111_4162, w_111_4165, w_111_4166, w_111_4171, w_111_4184, w_111_4189, w_111_4193, w_111_4197, w_111_4216, w_111_4223, w_111_4225, w_111_4227, w_111_4233, w_111_4234, w_111_4236, w_111_4237, w_111_4240, w_111_4241, w_111_4243, w_111_4244, w_111_4251, w_111_4253, w_111_4254, w_111_4255, w_111_4264, w_111_4267, w_111_4273, w_111_4285, w_111_4295, w_111_4298, w_111_4301, w_111_4302, w_111_4305, w_111_4310, w_111_4315, w_111_4318, w_111_4319, w_111_4330, w_111_4331, w_111_4333, w_111_4334, w_111_4339, w_111_4344, w_111_4345, w_111_4346, w_111_4347, w_111_4349, w_111_4351, w_111_4362, w_111_4364, w_111_4371, w_111_4376, w_111_4387, w_111_4394, w_111_4398, w_111_4399, w_111_4403, w_111_4404, w_111_4410, w_111_4412, w_111_4413, w_111_4418, w_111_4420, w_111_4423, w_111_4424, w_111_4426, w_111_4434, w_111_4436, w_111_4437, w_111_4451, w_111_4455, w_111_4457, w_111_4459, w_111_4464, w_111_4465, w_111_4468, w_111_4469, w_111_4476, w_111_4479, w_111_4485, w_111_4487, w_111_4490, w_111_4501, w_111_4505, w_111_4513, w_111_4515, w_111_4521, w_111_4523, w_111_4525, w_111_4528, w_111_4534, w_111_4535, w_111_4537, w_111_4541, w_111_4545, w_111_4551, w_111_4553, w_111_4554, w_111_4559, w_111_4564, w_111_4568, w_111_4571, w_111_4573, w_111_4574, w_111_4575, w_111_4576, w_111_4577;
  wire w_112_003, w_112_004, w_112_005, w_112_011, w_112_015, w_112_017, w_112_020, w_112_021, w_112_022, w_112_024, w_112_026, w_112_032, w_112_033, w_112_040, w_112_043, w_112_046, w_112_047, w_112_049, w_112_050, w_112_052, w_112_053, w_112_054, w_112_058, w_112_066, w_112_069, w_112_070, w_112_072, w_112_074, w_112_078, w_112_084, w_112_085, w_112_087, w_112_088, w_112_089, w_112_093, w_112_097, w_112_105, w_112_106, w_112_107, w_112_109, w_112_112, w_112_114, w_112_115, w_112_117, w_112_118, w_112_122, w_112_128, w_112_133, w_112_135, w_112_137, w_112_138, w_112_139, w_112_140, w_112_142, w_112_144, w_112_147, w_112_150, w_112_152, w_112_153, w_112_155, w_112_156, w_112_158, w_112_159, w_112_160, w_112_162, w_112_167, w_112_168, w_112_171, w_112_172, w_112_173, w_112_175, w_112_180, w_112_184, w_112_186, w_112_189, w_112_191, w_112_194, w_112_196, w_112_198, w_112_202, w_112_212, w_112_213, w_112_214, w_112_215, w_112_216, w_112_218, w_112_220, w_112_223, w_112_224, w_112_226, w_112_230, w_112_235, w_112_237, w_112_238, w_112_239, w_112_240, w_112_241, w_112_242, w_112_243, w_112_244, w_112_245, w_112_249, w_112_250, w_112_251, w_112_257, w_112_260, w_112_261, w_112_263, w_112_264, w_112_266, w_112_269, w_112_270, w_112_271, w_112_273, w_112_274, w_112_277, w_112_278, w_112_279, w_112_280, w_112_281, w_112_282, w_112_284, w_112_286, w_112_288, w_112_290, w_112_293, w_112_297, w_112_299, w_112_305, w_112_306, w_112_307, w_112_308, w_112_310, w_112_316, w_112_318, w_112_319, w_112_321, w_112_326, w_112_332, w_112_336, w_112_340, w_112_342, w_112_346, w_112_348, w_112_351, w_112_352, w_112_354, w_112_357, w_112_361, w_112_365, w_112_366, w_112_369, w_112_370, w_112_373, w_112_375, w_112_380, w_112_383, w_112_385, w_112_388, w_112_389, w_112_390, w_112_393, w_112_394, w_112_397, w_112_402, w_112_406, w_112_407, w_112_409, w_112_419, w_112_420, w_112_425, w_112_426, w_112_433, w_112_435, w_112_438, w_112_439, w_112_443, w_112_444, w_112_449, w_112_450, w_112_451, w_112_452, w_112_455, w_112_457, w_112_459, w_112_460, w_112_461, w_112_462, w_112_466, w_112_468, w_112_469, w_112_471, w_112_472, w_112_473, w_112_474, w_112_479, w_112_494, w_112_495, w_112_496, w_112_499, w_112_500, w_112_503, w_112_504, w_112_505, w_112_506, w_112_507, w_112_508, w_112_509, w_112_510, w_112_513, w_112_515, w_112_516, w_112_517, w_112_519, w_112_520, w_112_522, w_112_525, w_112_527, w_112_528, w_112_529, w_112_532, w_112_535, w_112_546, w_112_547, w_112_550, w_112_552, w_112_559, w_112_563, w_112_576, w_112_578, w_112_580, w_112_581, w_112_582, w_112_583, w_112_584, w_112_585, w_112_588, w_112_590, w_112_591, w_112_595, w_112_597, w_112_598, w_112_599, w_112_601, w_112_602, w_112_605, w_112_610, w_112_611, w_112_612, w_112_614, w_112_622, w_112_624, w_112_627, w_112_629, w_112_632, w_112_634, w_112_638, w_112_643, w_112_645, w_112_646, w_112_647, w_112_648, w_112_651, w_112_655, w_112_656, w_112_659, w_112_660, w_112_665, w_112_667, w_112_671, w_112_674, w_112_675, w_112_677, w_112_683, w_112_688, w_112_691, w_112_692, w_112_693, w_112_696, w_112_697, w_112_698, w_112_702, w_112_703, w_112_706, w_112_707, w_112_708, w_112_710, w_112_711, w_112_714, w_112_716, w_112_720, w_112_721, w_112_723, w_112_725, w_112_726, w_112_739, w_112_741, w_112_742, w_112_744, w_112_746, w_112_748, w_112_751, w_112_752, w_112_754, w_112_757, w_112_759, w_112_762, w_112_763, w_112_767, w_112_771, w_112_773, w_112_774, w_112_779, w_112_781, w_112_782, w_112_785, w_112_787, w_112_789, w_112_791, w_112_792, w_112_793, w_112_794, w_112_795, w_112_796, w_112_804, w_112_805, w_112_808, w_112_810, w_112_812, w_112_814, w_112_815, w_112_817, w_112_818, w_112_820, w_112_824, w_112_825, w_112_827, w_112_832, w_112_836, w_112_840, w_112_841, w_112_843, w_112_844, w_112_846, w_112_848, w_112_850, w_112_852, w_112_853, w_112_858, w_112_861, w_112_863, w_112_865, w_112_872, w_112_875, w_112_878, w_112_881, w_112_882, w_112_883, w_112_884, w_112_887, w_112_889, w_112_890, w_112_893, w_112_894, w_112_900, w_112_902, w_112_905, w_112_907, w_112_908, w_112_911, w_112_913, w_112_914, w_112_915, w_112_920, w_112_927, w_112_928, w_112_929, w_112_931, w_112_933, w_112_935, w_112_936, w_112_937, w_112_941, w_112_942, w_112_943, w_112_944, w_112_951, w_112_952, w_112_957, w_112_961, w_112_962, w_112_965, w_112_973, w_112_977, w_112_978, w_112_979, w_112_981, w_112_983, w_112_984, w_112_985, w_112_986, w_112_990, w_112_993, w_112_995, w_112_996, w_112_998, w_112_999, w_112_1002, w_112_1004, w_112_1005, w_112_1011, w_112_1013, w_112_1014, w_112_1018, w_112_1019, w_112_1020, w_112_1023, w_112_1024, w_112_1025, w_112_1026, w_112_1029, w_112_1032, w_112_1037, w_112_1039, w_112_1041, w_112_1045, w_112_1047, w_112_1049, w_112_1051, w_112_1052, w_112_1055, w_112_1057, w_112_1058, w_112_1059, w_112_1060, w_112_1068, w_112_1071, w_112_1072, w_112_1073, w_112_1075, w_112_1077, w_112_1081, w_112_1085, w_112_1088, w_112_1091, w_112_1092, w_112_1093, w_112_1094, w_112_1098, w_112_1103, w_112_1106, w_112_1108, w_112_1120, w_112_1131, w_112_1133, w_112_1134, w_112_1143, w_112_1145, w_112_1146, w_112_1149, w_112_1153, w_112_1154, w_112_1158, w_112_1166, w_112_1173, w_112_1177, w_112_1180, w_112_1188, w_112_1191, w_112_1195, w_112_1196, w_112_1198, w_112_1203, w_112_1211, w_112_1213, w_112_1216, w_112_1218, w_112_1223, w_112_1225, w_112_1234, w_112_1235, w_112_1241, w_112_1247, w_112_1253, w_112_1256, w_112_1258, w_112_1259, w_112_1265, w_112_1273, w_112_1274, w_112_1276, w_112_1279, w_112_1285, w_112_1286, w_112_1287, w_112_1289, w_112_1291, w_112_1296, w_112_1307, w_112_1311, w_112_1315, w_112_1323, w_112_1327, w_112_1330, w_112_1331, w_112_1332, w_112_1334, w_112_1340, w_112_1341, w_112_1344, w_112_1345, w_112_1352, w_112_1361, w_112_1363, w_112_1364, w_112_1367, w_112_1372, w_112_1373, w_112_1376, w_112_1377, w_112_1381, w_112_1386, w_112_1389, w_112_1391, w_112_1394, w_112_1396, w_112_1400, w_112_1403, w_112_1412, w_112_1417, w_112_1418, w_112_1426, w_112_1428, w_112_1429, w_112_1430, w_112_1433, w_112_1435, w_112_1438, w_112_1446, w_112_1453, w_112_1457, w_112_1463, w_112_1465, w_112_1466, w_112_1470, w_112_1479, w_112_1481, w_112_1486, w_112_1488, w_112_1491, w_112_1492, w_112_1493, w_112_1502, w_112_1516, w_112_1521, w_112_1524, w_112_1527, w_112_1529, w_112_1533, w_112_1534, w_112_1535, w_112_1537, w_112_1538, w_112_1542, w_112_1544, w_112_1545, w_112_1546, w_112_1558, w_112_1559, w_112_1563, w_112_1579, w_112_1610, w_112_1612, w_112_1613, w_112_1619, w_112_1624, w_112_1625, w_112_1627, w_112_1632, w_112_1634, w_112_1635, w_112_1639, w_112_1640, w_112_1641, w_112_1644, w_112_1647, w_112_1648, w_112_1650, w_112_1653, w_112_1656, w_112_1658, w_112_1665, w_112_1666, w_112_1670, w_112_1671, w_112_1672, w_112_1673, w_112_1675, w_112_1678, w_112_1679, w_112_1682, w_112_1687, w_112_1690, w_112_1692, w_112_1693, w_112_1700, w_112_1705, w_112_1706, w_112_1707, w_112_1711, w_112_1715, w_112_1717, w_112_1718, w_112_1719, w_112_1728, w_112_1730, w_112_1731, w_112_1734, w_112_1736, w_112_1738, w_112_1739, w_112_1741, w_112_1743, w_112_1744, w_112_1752, w_112_1757, w_112_1763, w_112_1768, w_112_1774, w_112_1777, w_112_1780, w_112_1783, w_112_1786, w_112_1801, w_112_1803, w_112_1805, w_112_1807, w_112_1811, w_112_1814, w_112_1827, w_112_1829, w_112_1833, w_112_1836, w_112_1838, w_112_1840, w_112_1841, w_112_1846, w_112_1847, w_112_1848, w_112_1852, w_112_1856, w_112_1860, w_112_1865, w_112_1866, w_112_1868, w_112_1869, w_112_1870, w_112_1871, w_112_1872, w_112_1883, w_112_1888, w_112_1889, w_112_1892, w_112_1910, w_112_1915, w_112_1916, w_112_1919, w_112_1925, w_112_1933, w_112_1936, w_112_1939, w_112_1940, w_112_1944, w_112_1945, w_112_1947, w_112_1949, w_112_1951, w_112_1952, w_112_1955, w_112_1956, w_112_1966, w_112_1970, w_112_1974, w_112_1980, w_112_1990, w_112_1994, w_112_1998, w_112_2003, w_112_2006, w_112_2023, w_112_2024, w_112_2030, w_112_2031, w_112_2032, w_112_2041, w_112_2046, w_112_2047, w_112_2051, w_112_2062, w_112_2064, w_112_2065, w_112_2066, w_112_2073, w_112_2078, w_112_2086, w_112_2088, w_112_2091, w_112_2094, w_112_2105, w_112_2109, w_112_2113, w_112_2118, w_112_2119, w_112_2120, w_112_2124, w_112_2134, w_112_2137, w_112_2149, w_112_2150, w_112_2152, w_112_2153, w_112_2156, w_112_2158, w_112_2165, w_112_2168, w_112_2172, w_112_2175, w_112_2177, w_112_2180, w_112_2181, w_112_2184, w_112_2194, w_112_2195, w_112_2201, w_112_2204, w_112_2206, w_112_2207, w_112_2215, w_112_2219, w_112_2224, w_112_2225, w_112_2227, w_112_2228, w_112_2231, w_112_2233, w_112_2234, w_112_2236, w_112_2239, w_112_2250, w_112_2259, w_112_2262, w_112_2264, w_112_2266, w_112_2268, w_112_2275, w_112_2278, w_112_2279, w_112_2285, w_112_2286, w_112_2288, w_112_2289, w_112_2290, w_112_2297, w_112_2299, w_112_2302, w_112_2309, w_112_2312, w_112_2317, w_112_2324, w_112_2325, w_112_2326, w_112_2327, w_112_2333, w_112_2346, w_112_2354, w_112_2355, w_112_2356, w_112_2364, w_112_2365, w_112_2367, w_112_2371, w_112_2373, w_112_2383, w_112_2391, w_112_2402, w_112_2408, w_112_2421, w_112_2423, w_112_2427, w_112_2430, w_112_2438, w_112_2439, w_112_2440, w_112_2444, w_112_2448, w_112_2452, w_112_2459, w_112_2461, w_112_2472, w_112_2473, w_112_2477, w_112_2478, w_112_2479, w_112_2482, w_112_2486, w_112_2489, w_112_2495, w_112_2504, w_112_2505, w_112_2508, w_112_2510, w_112_2515, w_112_2521, w_112_2522, w_112_2531, w_112_2533, w_112_2534, w_112_2538, w_112_2544, w_112_2545, w_112_2547, w_112_2556, w_112_2559, w_112_2561, w_112_2567, w_112_2569, w_112_2575, w_112_2578, w_112_2580, w_112_2581, w_112_2582, w_112_2584, w_112_2585, w_112_2588, w_112_2592, w_112_2593, w_112_2595, w_112_2600, w_112_2603, w_112_2605, w_112_2607, w_112_2610, w_112_2615, w_112_2617, w_112_2618, w_112_2619, w_112_2620, w_112_2621, w_112_2623, w_112_2631, w_112_2640, w_112_2641, w_112_2642, w_112_2643, w_112_2645, w_112_2646, w_112_2647, w_112_2648, w_112_2649, w_112_2650, w_112_2660, w_112_2665, w_112_2666, w_112_2669, w_112_2671, w_112_2674, w_112_2676, w_112_2679, w_112_2684, w_112_2686, w_112_2690, w_112_2695, w_112_2697, w_112_2701, w_112_2702, w_112_2706, w_112_2713, w_112_2718, w_112_2727, w_112_2728, w_112_2730, w_112_2733, w_112_2735, w_112_2739, w_112_2746, w_112_2747, w_112_2748, w_112_2749, w_112_2751, w_112_2752, w_112_2754, w_112_2772, w_112_2774, w_112_2779, w_112_2781, w_112_2783, w_112_2784, w_112_2789, w_112_2791, w_112_2799, w_112_2801, w_112_2806, w_112_2808, w_112_2809, w_112_2827, w_112_2831, w_112_2838, w_112_2839, w_112_2842, w_112_2846, w_112_2849, w_112_2853, w_112_2855, w_112_2856, w_112_2860, w_112_2865, w_112_2869, w_112_2871, w_112_2872, w_112_2873, w_112_2874, w_112_2877, w_112_2886, w_112_2888, w_112_2890, w_112_2901, w_112_2907, w_112_2908, w_112_2914, w_112_2923, w_112_2931, w_112_2932, w_112_2933, w_112_2936, w_112_2950, w_112_2953, w_112_2958, w_112_2963, w_112_2968, w_112_2971, w_112_2976, w_112_2978, w_112_2979, w_112_2980, w_112_2985, w_112_2991, w_112_3000, w_112_3011, w_112_3017, w_112_3024, w_112_3026, w_112_3036, w_112_3037, w_112_3042, w_112_3047, w_112_3056, w_112_3057, w_112_3060, w_112_3061, w_112_3067, w_112_3069, w_112_3072, w_112_3073, w_112_3076, w_112_3078, w_112_3080, w_112_3081, w_112_3093, w_112_3098, w_112_3099, w_112_3107, w_112_3110, w_112_3111, w_112_3115, w_112_3116, w_112_3117, w_112_3118, w_112_3121, w_112_3122, w_112_3123, w_112_3128, w_112_3130, w_112_3135, w_112_3141, w_112_3146, w_112_3153, w_112_3154, w_112_3155, w_112_3157, w_112_3161, w_112_3165, w_112_3171, w_112_3178, w_112_3182, w_112_3190, w_112_3196, w_112_3200, w_112_3223, w_112_3224, w_112_3225, w_112_3227, w_112_3228, w_112_3230, w_112_3231, w_112_3233, w_112_3240, w_112_3251, w_112_3252, w_112_3257, w_112_3262, w_112_3264, w_112_3272, w_112_3273, w_112_3275, w_112_3277, w_112_3280, w_112_3282, w_112_3295, w_112_3296, w_112_3298, w_112_3302, w_112_3303, w_112_3304, w_112_3310, w_112_3311, w_112_3322, w_112_3333, w_112_3338, w_112_3344, w_112_3351, w_112_3355, w_112_3356, w_112_3363, w_112_3366, w_112_3368, w_112_3371, w_112_3372, w_112_3376, w_112_3380, w_112_3381, w_112_3389, w_112_3395, w_112_3402, w_112_3403, w_112_3404, w_112_3408, w_112_3412, w_112_3422, w_112_3423, w_112_3425, w_112_3431, w_112_3432, w_112_3441, w_112_3443, w_112_3448, w_112_3449, w_112_3452, w_112_3457, w_112_3459, w_112_3461, w_112_3466, w_112_3471, w_112_3476, w_112_3479, w_112_3484, w_112_3486, w_112_3488, w_112_3494, w_112_3495, w_112_3500, w_112_3502, w_112_3503, w_112_3513, w_112_3516, w_112_3523, w_112_3545, w_112_3548, w_112_3552, w_112_3558, w_112_3561, w_112_3565, w_112_3583, w_112_3588, w_112_3589, w_112_3592, w_112_3604, w_112_3612, w_112_3614, w_112_3618, w_112_3632, w_112_3634, w_112_3637, w_112_3641, w_112_3643, w_112_3645, w_112_3649, w_112_3650, w_112_3651, w_112_3653, w_112_3659, w_112_3663, w_112_3672, w_112_3675, w_112_3690, w_112_3692, w_112_3701, w_112_3704, w_112_3705, w_112_3712, w_112_3717, w_112_3721, w_112_3723, w_112_3725, w_112_3731, w_112_3734, w_112_3742, w_112_3743, w_112_3744, w_112_3745, w_112_3751, w_112_3754, w_112_3759, w_112_3760, w_112_3761, w_112_3764, w_112_3765, w_112_3766, w_112_3778, w_112_3783, w_112_3784, w_112_3785, w_112_3786, w_112_3793, w_112_3794, w_112_3796, w_112_3802, w_112_3804, w_112_3807, w_112_3823, w_112_3835, w_112_3836, w_112_3838, w_112_3841, w_112_3851, w_112_3853, w_112_3856, w_112_3860, w_112_3864, w_112_3873, w_112_3875, w_112_3877, w_112_3878, w_112_3882, w_112_3883, w_112_3890, w_112_3891, w_112_3893;
  wire w_113_000, w_113_003, w_113_004, w_113_008, w_113_009, w_113_011, w_113_012, w_113_013, w_113_017, w_113_021, w_113_022, w_113_026, w_113_027, w_113_030, w_113_036, w_113_041, w_113_043, w_113_045, w_113_046, w_113_048, w_113_049, w_113_052, w_113_053, w_113_059, w_113_060, w_113_061, w_113_071, w_113_072, w_113_075, w_113_076, w_113_080, w_113_083, w_113_085, w_113_086, w_113_087, w_113_088, w_113_095, w_113_096, w_113_097, w_113_099, w_113_102, w_113_103, w_113_104, w_113_105, w_113_106, w_113_109, w_113_110, w_113_113, w_113_123, w_113_124, w_113_125, w_113_129, w_113_133, w_113_134, w_113_138, w_113_139, w_113_140, w_113_141, w_113_149, w_113_150, w_113_153, w_113_154, w_113_156, w_113_158, w_113_160, w_113_162, w_113_163, w_113_164, w_113_165, w_113_166, w_113_167, w_113_169, w_113_171, w_113_174, w_113_175, w_113_176, w_113_177, w_113_181, w_113_183, w_113_184, w_113_186, w_113_188, w_113_191, w_113_194, w_113_196, w_113_197, w_113_200, w_113_204, w_113_210, w_113_213, w_113_218, w_113_219, w_113_225, w_113_229, w_113_230, w_113_233, w_113_235, w_113_242, w_113_243, w_113_244, w_113_245, w_113_247, w_113_248, w_113_249, w_113_250, w_113_251, w_113_254, w_113_255, w_113_257, w_113_259, w_113_265, w_113_267, w_113_279, w_113_280, w_113_281, w_113_283, w_113_288, w_113_289, w_113_292, w_113_294, w_113_298, w_113_301, w_113_302, w_113_306, w_113_309, w_113_311, w_113_313, w_113_314, w_113_317, w_113_319, w_113_328, w_113_330, w_113_331, w_113_332, w_113_339, w_113_341, w_113_342, w_113_345, w_113_348, w_113_349, w_113_353, w_113_354, w_113_356, w_113_357, w_113_358, w_113_363, w_113_364, w_113_365, w_113_368, w_113_369, w_113_370, w_113_375, w_113_376, w_113_378, w_113_379, w_113_381, w_113_384, w_113_387, w_113_388, w_113_390, w_113_392, w_113_394, w_113_395, w_113_396, w_113_398, w_113_399, w_113_403, w_113_408, w_113_411, w_113_413, w_113_415, w_113_422, w_113_424, w_113_425, w_113_427, w_113_429, w_113_430, w_113_432, w_113_433, w_113_434, w_113_439, w_113_443, w_113_445, w_113_448, w_113_450, w_113_451, w_113_454, w_113_456, w_113_457, w_113_459, w_113_461, w_113_463, w_113_464, w_113_465, w_113_468, w_113_469, w_113_471, w_113_472, w_113_476, w_113_486, w_113_487, w_113_489, w_113_490, w_113_492, w_113_496, w_113_498, w_113_501, w_113_507, w_113_508, w_113_509, w_113_510, w_113_511, w_113_516, w_113_517, w_113_518, w_113_519, w_113_525, w_113_532, w_113_534, w_113_535, w_113_536, w_113_537, w_113_539, w_113_543, w_113_544, w_113_548, w_113_549, w_113_554, w_113_556, w_113_558, w_113_561, w_113_564, w_113_571, w_113_572, w_113_574, w_113_577, w_113_580, w_113_585, w_113_586, w_113_590, w_113_591, w_113_594, w_113_596, w_113_597, w_113_598, w_113_602, w_113_603, w_113_604, w_113_605, w_113_609, w_113_611, w_113_612, w_113_618, w_113_619, w_113_620, w_113_623, w_113_625, w_113_628, w_113_629, w_113_632, w_113_634, w_113_635, w_113_638, w_113_643, w_113_644, w_113_645, w_113_647, w_113_648, w_113_651, w_113_653, w_113_655, w_113_656, w_113_658, w_113_659, w_113_660, w_113_661, w_113_662, w_113_663, w_113_665, w_113_668, w_113_670, w_113_671, w_113_673, w_113_674, w_113_677, w_113_678, w_113_680, w_113_684, w_113_686, w_113_687, w_113_689, w_113_692, w_113_699, w_113_700, w_113_701, w_113_702, w_113_703, w_113_704, w_113_706, w_113_707, w_113_711, w_113_712, w_113_713, w_113_717, w_113_720, w_113_722, w_113_725, w_113_728, w_113_731, w_113_734, w_113_739, w_113_740, w_113_742, w_113_743, w_113_745, w_113_748, w_113_749, w_113_751, w_113_755, w_113_761, w_113_763, w_113_768, w_113_769, w_113_771, w_113_773, w_113_775, w_113_778, w_113_781, w_113_786, w_113_787, w_113_790, w_113_791, w_113_792, w_113_793, w_113_795, w_113_797, w_113_800, w_113_809, w_113_811, w_113_812, w_113_815, w_113_817, w_113_827, w_113_831, w_113_833, w_113_834, w_113_835, w_113_838, w_113_840, w_113_841, w_113_845, w_113_846, w_113_847, w_113_849, w_113_850, w_113_852, w_113_855, w_113_857, w_113_858, w_113_859, w_113_860, w_113_861, w_113_863, w_113_864, w_113_870, w_113_871, w_113_872, w_113_876, w_113_877, w_113_882, w_113_884, w_113_886, w_113_887, w_113_891, w_113_897, w_113_899, w_113_900, w_113_904, w_113_906, w_113_908, w_113_909, w_113_910, w_113_912, w_113_914, w_113_916, w_113_918, w_113_921, w_113_924, w_113_931, w_113_935, w_113_936, w_113_937, w_113_938, w_113_940, w_113_944, w_113_945, w_113_946, w_113_949, w_113_951, w_113_953, w_113_955, w_113_956, w_113_957, w_113_958, w_113_959, w_113_961, w_113_963, w_113_964, w_113_965, w_113_966, w_113_973, w_113_974, w_113_977, w_113_982, w_113_983, w_113_985, w_113_990, w_113_992, w_113_993, w_113_994, w_113_995, w_113_998, w_113_1000, w_113_1004, w_113_1005, w_113_1006, w_113_1007, w_113_1010, w_113_1011, w_113_1012, w_113_1013, w_113_1014, w_113_1019, w_113_1026, w_113_1029, w_113_1030, w_113_1032, w_113_1036, w_113_1037, w_113_1038, w_113_1039, w_113_1041, w_113_1042, w_113_1043, w_113_1050, w_113_1053, w_113_1054, w_113_1055, w_113_1056, w_113_1057, w_113_1061, w_113_1065, w_113_1066, w_113_1071, w_113_1078, w_113_1081, w_113_1083, w_113_1086, w_113_1087, w_113_1089, w_113_1091, w_113_1093, w_113_1095, w_113_1098, w_113_1100, w_113_1101, w_113_1102, w_113_1103, w_113_1104, w_113_1105, w_113_1106, w_113_1107, w_113_1109, w_113_1114, w_113_1115, w_113_1117, w_113_1118, w_113_1119, w_113_1123, w_113_1125, w_113_1127, w_113_1131, w_113_1137, w_113_1142, w_113_1144, w_113_1145, w_113_1147, w_113_1148, w_113_1149, w_113_1158, w_113_1162, w_113_1163, w_113_1164, w_113_1165, w_113_1167, w_113_1168, w_113_1169, w_113_1170, w_113_1172, w_113_1175, w_113_1176, w_113_1178, w_113_1180, w_113_1181, w_113_1182, w_113_1186, w_113_1188, w_113_1189, w_113_1192, w_113_1194, w_113_1196, w_113_1197, w_113_1203, w_113_1209, w_113_1213, w_113_1215, w_113_1216, w_113_1221, w_113_1223, w_113_1227, w_113_1228, w_113_1230, w_113_1231, w_113_1232, w_113_1233, w_113_1236, w_113_1242, w_113_1243, w_113_1244, w_113_1245, w_113_1248, w_113_1253, w_113_1256, w_113_1258, w_113_1261, w_113_1263, w_113_1264, w_113_1265, w_113_1268, w_113_1269, w_113_1273, w_113_1275, w_113_1276, w_113_1281, w_113_1283, w_113_1285, w_113_1286, w_113_1288, w_113_1289, w_113_1290, w_113_1301, w_113_1305, w_113_1306, w_113_1307, w_113_1308, w_113_1309, w_113_1310, w_113_1311, w_113_1315, w_113_1319, w_113_1322, w_113_1324, w_113_1325, w_113_1326, w_113_1327, w_113_1331, w_113_1336, w_113_1339, w_113_1340, w_113_1344, w_113_1346, w_113_1348, w_113_1354, w_113_1356, w_113_1360, w_113_1361, w_113_1363, w_113_1364, w_113_1365, w_113_1366, w_113_1367, w_113_1368, w_113_1369, w_113_1370, w_113_1373, w_113_1375, w_113_1380, w_113_1381, w_113_1382, w_113_1383, w_113_1385, w_113_1393, w_113_1395, w_113_1397, w_113_1400, w_113_1401, w_113_1404, w_113_1405, w_113_1409, w_113_1411, w_113_1412, w_113_1413, w_113_1415, w_113_1418, w_113_1420, w_113_1422, w_113_1423, w_113_1429, w_113_1430, w_113_1431, w_113_1433, w_113_1439, w_113_1440, w_113_1444, w_113_1445, w_113_1446, w_113_1450, w_113_1453, w_113_1455, w_113_1457, w_113_1463, w_113_1465, w_113_1466, w_113_1467, w_113_1469, w_113_1471, w_113_1474, w_113_1475, w_113_1476, w_113_1480, w_113_1483, w_113_1487, w_113_1489, w_113_1490, w_113_1491, w_113_1492, w_113_1493, w_113_1495, w_113_1496, w_113_1497, w_113_1498, w_113_1499, w_113_1501, w_113_1503, w_113_1504, w_113_1505, w_113_1513, w_113_1514, w_113_1515, w_113_1517, w_113_1520, w_113_1522, w_113_1526, w_113_1528, w_113_1529, w_113_1530, w_113_1532, w_113_1533, w_113_1534, w_113_1536, w_113_1545, w_113_1547, w_113_1551, w_113_1553, w_113_1554, w_113_1555, w_113_1556, w_113_1557, w_113_1558, w_113_1561, w_113_1563, w_113_1564, w_113_1566, w_113_1570, w_113_1571, w_113_1573, w_113_1574, w_113_1575, w_113_1576, w_113_1578, w_113_1579, w_113_1580, w_113_1584, w_113_1585, w_113_1587, w_113_1590, w_113_1594, w_113_1596, w_113_1597, w_113_1601, w_113_1602, w_113_1607, w_113_1608, w_113_1613, w_113_1615, w_113_1616, w_113_1618, w_113_1619, w_113_1620, w_113_1622, w_113_1623, w_113_1624, w_113_1627, w_113_1628, w_113_1631, w_113_1633, w_113_1634, w_113_1638, w_113_1639, w_113_1641, w_113_1642, w_113_1644, w_113_1648, w_113_1650, w_113_1653, w_113_1657, w_113_1658, w_113_1659, w_113_1660, w_113_1661, w_113_1666, w_113_1669, w_113_1672, w_113_1674, w_113_1675, w_113_1676, w_113_1677, w_113_1678, w_113_1679, w_113_1680, w_113_1681, w_113_1682, w_113_1685, w_113_1687, w_113_1688, w_113_1690, w_113_1692, w_113_1693, w_113_1696, w_113_1701, w_113_1702, w_113_1703, w_113_1706, w_113_1708, w_113_1709, w_113_1710, w_113_1714, w_113_1717, w_113_1718, w_113_1720, w_113_1723, w_113_1724, w_113_1725, w_113_1727, w_113_1731, w_113_1734, w_113_1735, w_113_1737, w_113_1739, w_113_1741, w_113_1742, w_113_1744, w_113_1750, w_113_1752, w_113_1756, w_113_1764, w_113_1765, w_113_1769, w_113_1770, w_113_1773, w_113_1781, w_113_1783, w_113_1795, w_113_1796, w_113_1798, w_113_1812, w_113_1816, w_113_1817, w_113_1826, w_113_1829, w_113_1840, w_113_1842, w_113_1852, w_113_1856, w_113_1861, w_113_1863, w_113_1870, w_113_1876, w_113_1882, w_113_1891, w_113_1892, w_113_1898, w_113_1899, w_113_1905, w_113_1906, w_113_1917, w_113_1920, w_113_1921, w_113_1923, w_113_1927, w_113_1929, w_113_1932, w_113_1934, w_113_1935, w_113_1936, w_113_1943, w_113_1951, w_113_1956, w_113_1963, w_113_1964, w_113_1966, w_113_1969, w_113_1972, w_113_1979, w_113_1980, w_113_1981, w_113_1982, w_113_1983, w_113_1985, w_113_1993, w_113_1996, w_113_2006, w_113_2008, w_113_2010, w_113_2012, w_113_2013, w_113_2014, w_113_2022, w_113_2023, w_113_2024, w_113_2025, w_113_2029, w_113_2030, w_113_2033, w_113_2036, w_113_2038, w_113_2040, w_113_2053, w_113_2055, w_113_2058, w_113_2061, w_113_2062, w_113_2066, w_113_2069, w_113_2072, w_113_2078, w_113_2083, w_113_2084, w_113_2086, w_113_2094, w_113_2097, w_113_2104, w_113_2106, w_113_2108, w_113_2109, w_113_2125, w_113_2128, w_113_2137, w_113_2139, w_113_2140, w_113_2143, w_113_2147, w_113_2148, w_113_2156, w_113_2158, w_113_2163, w_113_2168, w_113_2172, w_113_2174, w_113_2176, w_113_2184, w_113_2187, w_113_2189, w_113_2190, w_113_2192, w_113_2202, w_113_2206, w_113_2209, w_113_2214, w_113_2216, w_113_2233, w_113_2240, w_113_2267, w_113_2270, w_113_2273, w_113_2277, w_113_2284, w_113_2285, w_113_2291, w_113_2292, w_113_2294, w_113_2301, w_113_2305, w_113_2308, w_113_2310, w_113_2317, w_113_2320, w_113_2327, w_113_2331, w_113_2334, w_113_2342, w_113_2343, w_113_2346, w_113_2351, w_113_2352, w_113_2357, w_113_2362, w_113_2364, w_113_2365, w_113_2367, w_113_2369, w_113_2370, w_113_2371, w_113_2376, w_113_2381, w_113_2383, w_113_2386, w_113_2388, w_113_2389, w_113_2390, w_113_2397, w_113_2399, w_113_2401, w_113_2405, w_113_2412, w_113_2413, w_113_2415, w_113_2418, w_113_2420, w_113_2423, w_113_2427, w_113_2428, w_113_2433, w_113_2438, w_113_2444, w_113_2448, w_113_2449, w_113_2451, w_113_2452, w_113_2454, w_113_2459, w_113_2467, w_113_2468, w_113_2469, w_113_2470, w_113_2471, w_113_2474, w_113_2478, w_113_2480, w_113_2483, w_113_2486, w_113_2490, w_113_2491, w_113_2501, w_113_2504, w_113_2506, w_113_2515, w_113_2516, w_113_2517, w_113_2518, w_113_2519, w_113_2520, w_113_2531, w_113_2532, w_113_2534, w_113_2551, w_113_2556, w_113_2559, w_113_2565, w_113_2569, w_113_2576, w_113_2577, w_113_2580, w_113_2582, w_113_2593, w_113_2597, w_113_2599, w_113_2602, w_113_2603, w_113_2610, w_113_2616, w_113_2626, w_113_2629, w_113_2638, w_113_2649, w_113_2652, w_113_2653, w_113_2657, w_113_2668, w_113_2671, w_113_2672, w_113_2679, w_113_2687, w_113_2690, w_113_2700, w_113_2704, w_113_2706, w_113_2712, w_113_2715, w_113_2716, w_113_2720, w_113_2732, w_113_2737, w_113_2738, w_113_2753, w_113_2759, w_113_2764, w_113_2769, w_113_2771, w_113_2772, w_113_2776, w_113_2778, w_113_2779, w_113_2782, w_113_2784, w_113_2787, w_113_2788, w_113_2789, w_113_2791, w_113_2794, w_113_2796, w_113_2800, w_113_2801, w_113_2808, w_113_2815, w_113_2822, w_113_2829, w_113_2834, w_113_2843, w_113_2851, w_113_2853, w_113_2856, w_113_2858, w_113_2865, w_113_2869, w_113_2874, w_113_2886, w_113_2892, w_113_2895, w_113_2900, w_113_2908, w_113_2909, w_113_2914, w_113_2927, w_113_2928, w_113_2930, w_113_2935, w_113_2938, w_113_2939, w_113_2945, w_113_2946, w_113_2950, w_113_2955, w_113_2960, w_113_2961, w_113_2965, w_113_2968, w_113_2970, w_113_2972, w_113_2975, w_113_2982, w_113_2988, w_113_2998, w_113_3001, w_113_3002, w_113_3004, w_113_3010, w_113_3012, w_113_3015, w_113_3020, w_113_3022, w_113_3023, w_113_3025, w_113_3030, w_113_3034, w_113_3036, w_113_3038, w_113_3041, w_113_3043, w_113_3045, w_113_3052, w_113_3058, w_113_3061, w_113_3068, w_113_3075, w_113_3076, w_113_3077, w_113_3079, w_113_3081, w_113_3082, w_113_3089, w_113_3093, w_113_3103, w_113_3104, w_113_3105, w_113_3108, w_113_3114, w_113_3115, w_113_3120, w_113_3126, w_113_3127, w_113_3129, w_113_3130, w_113_3132, w_113_3133, w_113_3140, w_113_3141, w_113_3153, w_113_3155, w_113_3157, w_113_3160, w_113_3165, w_113_3168, w_113_3170, w_113_3172, w_113_3173, w_113_3175, w_113_3179, w_113_3207, w_113_3214, w_113_3218, w_113_3221, w_113_3223, w_113_3229, w_113_3232, w_113_3233, w_113_3236, w_113_3237, w_113_3239, w_113_3245, w_113_3249, w_113_3252, w_113_3254, w_113_3257;
  wire w_114_001, w_114_002, w_114_003, w_114_007, w_114_009, w_114_010, w_114_015, w_114_019, w_114_023, w_114_024, w_114_025, w_114_026, w_114_027, w_114_029, w_114_030, w_114_031, w_114_032, w_114_036, w_114_038, w_114_039, w_114_040, w_114_041, w_114_045, w_114_046, w_114_047, w_114_048, w_114_049, w_114_050, w_114_051, w_114_052, w_114_053, w_114_054, w_114_055, w_114_057, w_114_059, w_114_060, w_114_063, w_114_066, w_114_069, w_114_070, w_114_071, w_114_072, w_114_073, w_114_074, w_114_075, w_114_076, w_114_079, w_114_080, w_114_082, w_114_084, w_114_087, w_114_090, w_114_092, w_114_093, w_114_094, w_114_098, w_114_099, w_114_101, w_114_102, w_114_104, w_114_105, w_114_107, w_114_108, w_114_109, w_114_111, w_114_113, w_114_114, w_114_115, w_114_116, w_114_117, w_114_118, w_114_119, w_114_120, w_114_123, w_114_124, w_114_126, w_114_127, w_114_128, w_114_129, w_114_132, w_114_133, w_114_136, w_114_138, w_114_139, w_114_140, w_114_143, w_114_145, w_114_150, w_114_151, w_114_152, w_114_153, w_114_155, w_114_156, w_114_157, w_114_158, w_114_161, w_114_163, w_114_164, w_114_165, w_114_166, w_114_167, w_114_169, w_114_170, w_114_171, w_114_174, w_114_175, w_114_177, w_114_178, w_114_181, w_114_183, w_114_184, w_114_185, w_114_186, w_114_187, w_114_188, w_114_190, w_114_194, w_114_196, w_114_197, w_114_198, w_114_199, w_114_201, w_114_202, w_114_204, w_114_206, w_114_207, w_114_210, w_114_211, w_114_214, w_114_215, w_114_216, w_114_217, w_114_220, w_114_225, w_114_226, w_114_227, w_114_229, w_114_234, w_114_235, w_114_238, w_114_239, w_114_244, w_114_246, w_114_247, w_114_248, w_114_249, w_114_250, w_114_251, w_114_252, w_114_253, w_114_255, w_114_256, w_114_257, w_114_259, w_114_260, w_114_263, w_114_264, w_114_267, w_114_268, w_114_269, w_114_270, w_114_271, w_114_272, w_114_273, w_114_277, w_114_280, w_114_281, w_114_282, w_114_283, w_114_285, w_114_287, w_114_288, w_114_293, w_114_295, w_114_297, w_114_299, w_114_300, w_114_304, w_114_307, w_114_309, w_114_310, w_114_313, w_114_315, w_114_316, w_114_319, w_114_321, w_114_323, w_114_325, w_114_326, w_114_327, w_114_329, w_114_332, w_114_333, w_114_335, w_114_336, w_114_337, w_114_339, w_114_340, w_114_342, w_114_344, w_114_347, w_114_348, w_114_350, w_114_355, w_114_356, w_114_362, w_114_363, w_114_365, w_114_367, w_114_368, w_114_369, w_114_371, w_114_373, w_114_374, w_114_378, w_114_382, w_114_383, w_114_385, w_114_387, w_114_388, w_114_390, w_114_393, w_114_395, w_114_396, w_114_399, w_114_400, w_114_401, w_114_403, w_114_404, w_114_405, w_114_407, w_114_408, w_114_409, w_114_413, w_114_414, w_114_419, w_114_422, w_114_424, w_114_426, w_114_429, w_114_430, w_114_433, w_114_434, w_114_435, w_114_437, w_114_440, w_114_441, w_114_443, w_114_449, w_114_450, w_114_451, w_114_452, w_114_456, w_114_461, w_114_462, w_114_467, w_114_468, w_114_469, w_114_470, w_114_471, w_114_473, w_114_475, w_114_478, w_114_481, w_114_482, w_114_484, w_114_486, w_114_487, w_114_491, w_114_500, w_114_502, w_114_503, w_114_506, w_114_508, w_114_509, w_114_510, w_114_511, w_114_512, w_114_514, w_114_516, w_114_517, w_114_518, w_114_520, w_114_522, w_114_526, w_114_528, w_114_529, w_114_530, w_114_531, w_114_533, w_114_535, w_114_537, w_114_539, w_114_540, w_114_541, w_114_542, w_114_544, w_114_545, w_114_551, w_114_552, w_114_553, w_114_554, w_114_563, w_114_564, w_114_568, w_114_570, w_114_571, w_114_572, w_114_574, w_114_575, w_114_576, w_114_577, w_114_578, w_114_579, w_114_580, w_114_585, w_114_589, w_114_591, w_114_595, w_114_597, w_114_599, w_114_600, w_114_602, w_114_603, w_114_607, w_114_608, w_114_609, w_114_610, w_114_618, w_114_622, w_114_623, w_114_626, w_114_627, w_114_628, w_114_630, w_114_631, w_114_636, w_114_640, w_114_642, w_114_644, w_114_645, w_114_646, w_114_651, w_114_656, w_114_657, w_114_659, w_114_660, w_114_661, w_114_667, w_114_668, w_114_671, w_114_677, w_114_679, w_114_682, w_114_683, w_114_685, w_114_690, w_114_691, w_114_694, w_114_697, w_114_700, w_114_702, w_114_703, w_114_706, w_114_708, w_114_710, w_114_712, w_114_713, w_114_717, w_114_722, w_114_728, w_114_729, w_114_733, w_114_735, w_114_738, w_114_740, w_114_742, w_114_743, w_114_744, w_114_750, w_114_751, w_114_756, w_114_757, w_114_759, w_114_761, w_114_762, w_114_763, w_114_768, w_114_770, w_114_774, w_114_775, w_114_776, w_114_778, w_114_779, w_114_780, w_114_784, w_114_787, w_114_788, w_114_789, w_114_790, w_114_792, w_114_794, w_114_796, w_114_797, w_114_798, w_114_799, w_114_804, w_114_806, w_114_808, w_114_811, w_114_812, w_114_814, w_114_815, w_114_817, w_114_818, w_114_820, w_114_826, w_114_833, w_114_834, w_114_836, w_114_839, w_114_840, w_114_841, w_114_842, w_114_845, w_114_846, w_114_847, w_114_853, w_114_854, w_114_857, w_114_860, w_114_864, w_114_865, w_114_866, w_114_868, w_114_869, w_114_870, w_114_871, w_114_875, w_114_877, w_114_878, w_114_880, w_114_887, w_114_888, w_114_889, w_114_890, w_114_891, w_114_892, w_114_894, w_114_895, w_114_901, w_114_906, w_114_907, w_114_914, w_114_915, w_114_917, w_114_918, w_114_920, w_114_928, w_114_929, w_114_930, w_114_931, w_114_935, w_114_941, w_114_944, w_114_950, w_114_951, w_114_952, w_114_954, w_114_955, w_114_956, w_114_958, w_114_959, w_114_965, w_114_966, w_114_969, w_114_971, w_114_974, w_114_975, w_114_976, w_114_977, w_114_979, w_114_980, w_114_981, w_114_982, w_114_984, w_114_990, w_114_996, w_114_999, w_114_1001, w_114_1002, w_114_1003, w_114_1007, w_114_1009, w_114_1010, w_114_1011, w_114_1012, w_114_1013, w_114_1015, w_114_1017, w_114_1018, w_114_1022, w_114_1024, w_114_1025, w_114_1030, w_114_1032, w_114_1033, w_114_1034, w_114_1035, w_114_1037, w_114_1039, w_114_1040, w_114_1042, w_114_1044, w_114_1045, w_114_1046, w_114_1049, w_114_1051, w_114_1054, w_114_1056, w_114_1058, w_114_1060, w_114_1061, w_114_1062, w_114_1065, w_114_1066, w_114_1067, w_114_1069, w_114_1071, w_114_1075, w_114_1078, w_114_1079, w_114_1083, w_114_1085, w_114_1086, w_114_1087, w_114_1089, w_114_1090, w_114_1092, w_114_1095, w_114_1096, w_114_1098, w_114_1100, w_114_1104, w_114_1108, w_114_1109, w_114_1110, w_114_1111, w_114_1113, w_114_1115, w_114_1116, w_114_1118, w_114_1120, w_114_1124, w_114_1127, w_114_1129, w_114_1130, w_114_1132, w_114_1133, w_114_1136, w_114_1144, w_114_1145, w_114_1147, w_114_1149, w_114_1150, w_114_1152, w_114_1156, w_114_1158, w_114_1161, w_114_1162, w_114_1164, w_114_1166, w_114_1168, w_114_1170, w_114_1176, w_114_1179, w_114_1180, w_114_1182, w_114_1188, w_114_1189, w_114_1190, w_114_1192, w_114_1194, w_114_1195, w_114_1198, w_114_1200, w_114_1201, w_114_1203, w_114_1205, w_114_1207, w_114_1209, w_114_1211, w_114_1215, w_114_1216, w_114_1217, w_114_1220, w_114_1224, w_114_1225, w_114_1226, w_114_1227, w_114_1232, w_114_1233, w_114_1234, w_114_1235, w_114_1236, w_114_1241, w_114_1245, w_114_1247, w_114_1249, w_114_1251, w_114_1252, w_114_1257, w_114_1258, w_114_1261, w_114_1262, w_114_1267, w_114_1268, w_114_1271, w_114_1276, w_114_1278, w_114_1281, w_114_1286, w_114_1287, w_114_1290, w_114_1297, w_114_1298, w_114_1299, w_114_1300, w_114_1302, w_114_1306, w_114_1307, w_114_1309, w_114_1314, w_114_1315, w_114_1316, w_114_1318, w_114_1322, w_114_1324, w_114_1325, w_114_1326, w_114_1329, w_114_1330, w_114_1333, w_114_1334, w_114_1335, w_114_1337, w_114_1342, w_114_1343, w_114_1345, w_114_1346, w_114_1347, w_114_1348, w_114_1349, w_114_1350, w_114_1351, w_114_1352, w_114_1353, w_114_1354, w_114_1355, w_114_1356, w_114_1357, w_114_1358, w_114_1359, w_114_1360, w_114_1361, w_114_1362, w_114_1363, w_114_1368, w_114_1370, w_114_1371, w_114_1372, w_114_1375, w_114_1378, w_114_1379, w_114_1383, w_114_1385, w_114_1387, w_114_1388, w_114_1393, w_114_1398, w_114_1399, w_114_1401, w_114_1404, w_114_1407, w_114_1408, w_114_1411, w_114_1414, w_114_1416, w_114_1418, w_114_1421, w_114_1427, w_114_1428, w_114_1430, w_114_1433, w_114_1438, w_114_1440, w_114_1444, w_114_1445, w_114_1447, w_114_1450, w_114_1451, w_114_1455, w_114_1460, w_114_1462, w_114_1463, w_114_1464, w_114_1466, w_114_1468, w_114_1471, w_114_1472, w_114_1480, w_114_1484, w_114_1485, w_114_1486, w_114_1491, w_114_1492, w_114_1493, w_114_1497, w_114_1499, w_114_1504, w_114_1512, w_114_1513, w_114_1522, w_114_1523, w_114_1525, w_114_1526, w_114_1527, w_114_1528, w_114_1529, w_114_1536, w_114_1537, w_114_1538, w_114_1539, w_114_1540, w_114_1544, w_114_1545, w_114_1548, w_114_1553, w_114_1555, w_114_1556, w_114_1558, w_114_1565, w_114_1567, w_114_1568, w_114_1570, w_114_1572, w_114_1574, w_114_1578, w_114_1580, w_114_1581, w_114_1582, w_114_1586, w_114_1587, w_114_1589, w_114_1590, w_114_1591, w_114_1597, w_114_1599, w_114_1604, w_114_1605, w_114_1607, w_114_1609, w_114_1612, w_114_1613, w_114_1614, w_114_1616, w_114_1623, w_114_1624, w_114_1628, w_114_1630, w_114_1631, w_114_1632, w_114_1633, w_114_1637, w_114_1638, w_114_1639, w_114_1640, w_114_1642, w_114_1646, w_114_1647, w_114_1649, w_114_1657, w_114_1659, w_114_1660, w_114_1664, w_114_1666, w_114_1670, w_114_1678, w_114_1679, w_114_1680, w_114_1681, w_114_1682, w_114_1683, w_114_1684, w_114_1685, w_114_1691, w_114_1693, w_114_1699, w_114_1700, w_114_1703, w_114_1707, w_114_1709, w_114_1711, w_114_1713, w_114_1715, w_114_1723, w_114_1725, w_114_1729, w_114_1730, w_114_1731, w_114_1736, w_114_1737, w_114_1743, w_114_1744, w_114_1745, w_114_1750, w_114_1752, w_114_1757, w_114_1761, w_114_1763, w_114_1765, w_114_1771, w_114_1776, w_114_1779, w_114_1786, w_114_1787, w_114_1789, w_114_1792, w_114_1794, w_114_1795, w_114_1800, w_114_1802, w_114_1803, w_114_1804, w_114_1808, w_114_1813, w_114_1814, w_114_1815, w_114_1817, w_114_1818, w_114_1821, w_114_1823, w_114_1825, w_114_1826, w_114_1829, w_114_1832, w_114_1833, w_114_1834, w_114_1837, w_114_1839, w_114_1840, w_114_1842, w_114_1848, w_114_1849, w_114_1850, w_114_1851, w_114_1852, w_114_1854, w_114_1855, w_114_1858, w_114_1863, w_114_1865, w_114_1866, w_114_1871, w_114_1874, w_114_1877, w_114_1884, w_114_1889, w_114_1891, w_114_1893, w_114_1895, w_114_1896, w_114_1898, w_114_1900, w_114_1902, w_114_1903, w_114_1905, w_114_1906, w_114_1908, w_114_1909, w_114_1911, w_114_1916, w_114_1920, w_114_1927, w_114_1928, w_114_1932, w_114_1939, w_114_1940, w_114_1941, w_114_1946, w_114_1950, w_114_1951, w_114_1954, w_114_1956, w_114_1957, w_114_1958, w_114_1959, w_114_1960, w_114_1961, w_114_1968, w_114_1970, w_114_1971, w_114_1972, w_114_1975, w_114_1978, w_114_1984, w_114_1985, w_114_1987, w_114_1989, w_114_1990, w_114_1992, w_114_1996, w_114_1997, w_114_2001, w_114_2004, w_114_2007, w_114_2008, w_114_2012, w_114_2017, w_114_2018, w_114_2021, w_114_2022, w_114_2023, w_114_2028, w_114_2029, w_114_2031, w_114_2039, w_114_2041, w_114_2044, w_114_2049, w_114_2051, w_114_2052, w_114_2053, w_114_2056, w_114_2057, w_114_2059, w_114_2061, w_114_2063, w_114_2066, w_114_2067, w_114_2068, w_114_2069, w_114_2071, w_114_2072, w_114_2074, w_114_2076, w_114_2080, w_114_2081, w_114_2083, w_114_2085, w_114_2088, w_114_2089, w_114_2090, w_114_2093, w_114_2094, w_114_2095, w_114_2097, w_114_2099, w_114_2101, w_114_2102, w_114_2105, w_114_2108, w_114_2110, w_114_2112, w_114_2116, w_114_2120, w_114_2122, w_114_2123, w_114_2124, w_114_2126, w_114_2127, w_114_2128, w_114_2132, w_114_2134, w_114_2135, w_114_2136, w_114_2139, w_114_2140, w_114_2143, w_114_2144, w_114_2146, w_114_2148, w_114_2149, w_114_2153, w_114_2158, w_114_2161, w_114_2162, w_114_2163, w_114_2167, w_114_2169, w_114_2173, w_114_2179, w_114_2180, w_114_2182, w_114_2185, w_114_2189, w_114_2190, w_114_2191, w_114_2195, w_114_2197, w_114_2198, w_114_2200, w_114_2201, w_114_2205, w_114_2206, w_114_2207, w_114_2209, w_114_2211, w_114_2216, w_114_2218, w_114_2220, w_114_2230, w_114_2233, w_114_2235, w_114_2236, w_114_2242, w_114_2249, w_114_2251, w_114_2252, w_114_2254, w_114_2255, w_114_2258, w_114_2261, w_114_2263, w_114_2265, w_114_2271, w_114_2276, w_114_2278, w_114_2279, w_114_2280, w_114_2283, w_114_2285, w_114_2287, w_114_2288, w_114_2292, w_114_2295, w_114_2296, w_114_2300, w_114_2302, w_114_2303, w_114_2305, w_114_2306, w_114_2307, w_114_2309, w_114_2312, w_114_2313, w_114_2314, w_114_2318, w_114_2320, w_114_2324, w_114_2329, w_114_2331, w_114_2332, w_114_2338, w_114_2340, w_114_2346, w_114_2349, w_114_2350, w_114_2351, w_114_2353, w_114_2357, w_114_2358, w_114_2359, w_114_2361, w_114_2362, w_114_2366, w_114_2367, w_114_2368, w_114_2372, w_114_2374, w_114_2375, w_114_2376, w_114_2377, w_114_2378, w_114_2379, w_114_2380, w_114_2381, w_114_2382, w_114_2383, w_114_2384, w_114_2388, w_114_2389, w_114_2390, w_114_2391, w_114_2392, w_114_2393, w_114_2394, w_114_2396;
  wire w_115_000, w_115_002, w_115_003, w_115_004, w_115_005, w_115_006, w_115_007, w_115_008, w_115_009, w_115_010, w_115_011, w_115_012, w_115_014, w_115_015, w_115_017, w_115_018, w_115_019, w_115_020, w_115_023, w_115_024, w_115_025, w_115_026, w_115_027, w_115_029, w_115_031, w_115_032, w_115_034, w_115_035, w_115_038, w_115_040, w_115_041, w_115_043, w_115_044, w_115_047, w_115_048, w_115_049, w_115_050, w_115_051, w_115_052, w_115_053, w_115_054, w_115_055, w_115_056, w_115_057, w_115_058, w_115_062, w_115_063, w_115_064, w_115_066, w_115_067, w_115_068, w_115_070, w_115_071, w_115_072, w_115_073, w_115_075, w_115_076, w_115_077, w_115_078, w_115_079, w_115_080, w_115_081, w_115_082, w_115_084, w_115_086, w_115_088, w_115_089, w_115_090, w_115_091, w_115_093, w_115_094, w_115_095, w_115_096, w_115_097, w_115_098, w_115_099, w_115_100, w_115_101, w_115_102, w_115_103, w_115_104, w_115_105, w_115_106, w_115_107, w_115_108, w_115_110, w_115_111, w_115_114, w_115_116, w_115_118, w_115_119, w_115_121, w_115_124, w_115_125, w_115_126, w_115_127, w_115_131, w_115_134, w_115_136, w_115_139, w_115_140, w_115_141, w_115_142, w_115_143, w_115_144, w_115_145, w_115_146, w_115_148, w_115_149, w_115_150, w_115_154, w_115_155, w_115_156, w_115_158, w_115_159, w_115_160, w_115_161, w_115_162, w_115_164, w_115_165, w_115_166, w_115_167, w_115_168, w_115_169, w_115_170, w_115_171, w_115_172, w_115_173, w_115_177, w_115_178, w_115_179, w_115_180, w_115_182, w_115_184, w_115_185, w_115_186, w_115_187, w_115_191, w_115_192, w_115_193, w_115_194, w_115_195, w_115_196, w_115_197, w_115_198, w_115_200, w_115_202, w_115_204, w_115_205, w_115_206, w_115_207, w_115_208, w_115_211, w_115_213, w_115_214, w_115_215, w_115_218, w_115_220, w_115_222, w_115_223, w_115_225, w_115_226, w_115_227, w_115_229, w_115_231, w_115_232, w_115_233, w_115_235, w_115_237, w_115_238, w_115_240, w_115_241, w_115_242, w_115_243, w_115_246, w_115_247, w_115_248, w_115_249, w_115_252, w_115_253, w_115_254, w_115_257, w_115_258, w_115_259, w_115_261, w_115_262, w_115_263, w_115_264, w_115_266, w_115_267, w_115_268, w_115_270, w_115_271, w_115_274, w_115_276, w_115_277, w_115_279, w_115_280, w_115_282, w_115_283, w_115_284, w_115_285, w_115_286, w_115_287, w_115_291, w_115_292, w_115_295, w_115_296, w_115_298, w_115_299, w_115_302, w_115_305, w_115_306, w_115_307, w_115_308, w_115_309, w_115_310, w_115_312, w_115_313, w_115_314, w_115_321, w_115_324, w_115_327, w_115_328, w_115_330, w_115_331, w_115_332, w_115_333, w_115_334, w_115_335, w_115_336, w_115_337, w_115_338, w_115_339, w_115_341, w_115_342, w_115_343, w_115_345, w_115_346, w_115_347, w_115_349, w_115_350, w_115_351, w_115_352, w_115_353, w_115_354, w_115_358, w_115_359, w_115_360, w_115_361, w_115_362, w_115_364, w_115_365, w_115_366, w_115_368, w_115_371, w_115_372, w_115_373, w_115_374, w_115_375, w_115_376, w_115_380, w_115_381, w_115_382, w_115_384, w_115_385, w_115_387, w_115_388, w_115_389, w_115_390, w_115_391, w_115_393, w_115_395, w_115_397, w_115_399, w_115_400, w_115_401, w_115_402, w_115_405, w_115_406, w_115_408, w_115_410, w_115_411, w_115_412, w_115_414, w_115_416, w_115_417, w_115_418, w_115_419, w_115_420, w_115_421, w_115_422, w_115_423, w_115_424, w_115_426, w_115_428, w_115_433, w_115_434, w_115_435, w_115_436, w_115_437, w_115_442, w_115_443, w_115_444, w_115_445, w_115_446, w_115_448, w_115_449, w_115_451, w_115_453, w_115_455, w_115_456, w_115_458, w_115_460, w_115_461, w_115_462, w_115_464, w_115_465, w_115_466, w_115_467, w_115_470, w_115_471, w_115_472, w_115_474, w_115_476, w_115_478, w_115_480, w_115_481, w_115_483, w_115_486, w_115_487, w_115_489, w_115_490, w_115_491, w_115_492, w_115_493, w_115_495, w_115_496, w_115_498, w_115_500, w_115_501, w_115_502, w_115_505, w_115_506, w_115_507, w_115_508, w_115_510, w_115_511, w_115_512, w_115_513, w_115_515, w_115_523, w_115_524, w_115_525, w_115_526, w_115_528, w_115_529, w_115_530, w_115_531, w_115_532, w_115_533, w_115_535, w_115_536, w_115_537, w_115_539, w_115_540, w_115_541, w_115_543, w_115_545, w_115_547, w_115_548, w_115_549, w_115_550, w_115_551, w_115_552, w_115_553, w_115_554, w_115_555, w_115_558, w_115_559, w_115_560, w_115_564, w_115_565, w_115_566, w_115_568, w_115_569, w_115_572, w_115_573, w_115_575, w_115_576, w_115_578, w_115_581, w_115_582, w_115_583, w_115_584, w_115_585, w_115_586, w_115_590, w_115_592, w_115_593, w_115_594, w_115_595, w_115_597, w_115_598, w_115_602, w_115_603, w_115_607, w_115_608, w_115_609, w_115_610, w_115_612, w_115_614, w_115_615, w_115_616, w_115_618, w_115_619, w_115_620, w_115_621, w_115_623, w_115_624, w_115_625, w_115_628, w_115_631, w_115_632, w_115_634, w_115_636, w_115_637, w_115_638, w_115_639, w_115_641, w_115_642, w_115_644, w_115_645, w_115_646, w_115_648, w_115_651, w_115_652, w_115_653, w_115_654, w_115_655, w_115_656, w_115_657, w_115_658, w_115_659, w_115_661, w_115_662, w_115_663, w_115_664, w_115_667, w_115_669, w_115_670, w_115_671, w_115_673, w_115_674, w_115_676, w_115_677, w_115_678, w_115_679, w_115_680, w_115_681, w_115_683, w_115_686, w_115_688, w_115_690, w_115_696, w_115_697, w_115_700, w_115_702, w_115_703, w_115_709, w_115_711, w_115_712, w_115_713, w_115_714, w_115_715, w_115_716, w_115_718, w_115_721, w_115_722, w_115_723, w_115_724, w_115_725, w_115_727, w_115_729, w_115_732, w_115_733, w_115_734, w_115_736, w_115_737, w_115_738, w_115_739, w_115_741, w_115_743, w_115_744, w_115_746, w_115_748, w_115_749, w_115_751, w_115_752, w_115_753, w_115_755, w_115_756, w_115_757, w_115_758, w_115_759, w_115_760, w_115_761, w_115_762, w_115_763, w_115_764, w_115_766, w_115_767, w_115_768, w_115_769, w_115_773, w_115_774, w_115_775, w_115_779, w_115_781, w_115_785, w_115_787, w_115_788, w_115_789, w_115_791, w_115_792, w_115_794, w_115_796, w_115_797, w_115_798, w_115_800, w_115_802, w_115_803, w_115_804, w_115_806, w_115_807, w_115_808, w_115_809, w_115_815, w_115_816, w_115_817, w_115_818, w_115_819, w_115_820, w_115_821, w_115_822, w_115_823, w_115_824, w_115_828, w_115_829, w_115_830, w_115_832, w_115_833, w_115_835, w_115_836, w_115_838, w_115_839, w_115_840, w_115_842, w_115_844, w_115_846, w_115_848, w_115_852, w_115_853, w_115_854, w_115_857, w_115_858, w_115_860, w_115_861, w_115_864, w_115_865, w_115_866, w_115_868, w_115_869, w_115_870, w_115_871, w_115_874, w_115_875, w_115_882, w_115_883, w_115_884, w_115_886, w_115_887, w_115_889, w_115_890, w_115_892, w_115_895, w_115_897, w_115_899, w_115_900, w_115_901, w_115_902, w_115_903, w_115_904, w_115_905, w_115_907, w_115_908, w_115_909, w_115_910, w_115_911, w_115_913, w_115_915, w_115_916, w_115_917, w_115_918, w_115_922, w_115_923, w_115_924, w_115_925, w_115_927, w_115_929, w_115_930, w_115_932, w_115_933, w_115_934, w_115_935, w_115_936, w_115_937, w_115_940, w_115_941, w_115_944, w_115_945, w_115_947, w_115_948, w_115_951, w_115_953, w_115_956, w_115_957, w_115_958, w_115_959, w_115_960, w_115_961, w_115_966, w_115_967, w_115_969, w_115_972, w_115_982, w_115_983, w_115_984, w_115_985, w_115_986, w_115_987, w_115_988, w_115_989, w_115_990, w_115_991, w_115_992, w_115_994, w_115_997, w_115_999, w_115_1000, w_115_1002, w_115_1003, w_115_1004, w_115_1005, w_115_1006, w_115_1007, w_115_1008, w_115_1011, w_115_1012, w_115_1013, w_115_1015, w_115_1017, w_115_1023, w_115_1027, w_115_1029, w_115_1033, w_115_1034, w_115_1037, w_115_1039, w_115_1040, w_115_1042, w_115_1043, w_115_1044, w_115_1045, w_115_1046, w_115_1047, w_115_1049, w_115_1050, w_115_1051, w_115_1052, w_115_1054, w_115_1056, w_115_1057, w_115_1059, w_115_1061, w_115_1064, w_115_1069, w_115_1070, w_115_1071, w_115_1072, w_115_1074, w_115_1075, w_115_1076, w_115_1077, w_115_1081, w_115_1082, w_115_1084, w_115_1085, w_115_1087, w_115_1088, w_115_1089, w_115_1091, w_115_1093, w_115_1094, w_115_1098, w_115_1102, w_115_1108, w_115_1109, w_115_1112, w_115_1114, w_115_1115, w_115_1118, w_115_1120, w_115_1121, w_115_1122, w_115_1123, w_115_1124, w_115_1125, w_115_1127, w_115_1129, w_115_1133, w_115_1134, w_115_1136, w_115_1138, w_115_1140, w_115_1141, w_115_1142, w_115_1143, w_115_1149, w_115_1151, w_115_1152, w_115_1154, w_115_1156, w_115_1158, w_115_1159, w_115_1160, w_115_1161, w_115_1163, w_115_1164, w_115_1165, w_115_1166, w_115_1167, w_115_1168, w_115_1169, w_115_1171, w_115_1172, w_115_1173, w_115_1174, w_115_1176, w_115_1182, w_115_1184, w_115_1187, w_115_1189, w_115_1191, w_115_1193, w_115_1194, w_115_1196, w_115_1199, w_115_1202, w_115_1204, w_115_1207, w_115_1211, w_115_1212, w_115_1213, w_115_1214, w_115_1217, w_115_1218, w_115_1220, w_115_1222, w_115_1223, w_115_1225, w_115_1226, w_115_1232, w_115_1235, w_115_1236, w_115_1237, w_115_1239, w_115_1241, w_115_1242, w_115_1243, w_115_1246, w_115_1247, w_115_1250, w_115_1251, w_115_1255, w_115_1256, w_115_1257, w_115_1259, w_115_1261, w_115_1262, w_115_1269, w_115_1270, w_115_1272, w_115_1274, w_115_1275, w_115_1277, w_115_1279, w_115_1282, w_115_1284, w_115_1286, w_115_1287, w_115_1294, w_115_1295, w_115_1296, w_115_1297, w_115_1298, w_115_1299, w_115_1302, w_115_1303, w_115_1304, w_115_1308, w_115_1309, w_115_1310, w_115_1311, w_115_1312, w_115_1313, w_115_1314, w_115_1315, w_115_1317, w_115_1319, w_115_1321, w_115_1322, w_115_1323, w_115_1324, w_115_1325;
  wire w_116_000, w_116_001, w_116_004, w_116_006, w_116_012, w_116_016, w_116_018, w_116_020, w_116_021, w_116_022, w_116_023, w_116_028, w_116_029, w_116_031, w_116_033, w_116_034, w_116_037, w_116_038, w_116_039, w_116_040, w_116_041, w_116_043, w_116_044, w_116_045, w_116_046, w_116_048, w_116_049, w_116_054, w_116_055, w_116_056, w_116_058, w_116_059, w_116_060, w_116_061, w_116_062, w_116_065, w_116_066, w_116_067, w_116_071, w_116_073, w_116_074, w_116_075, w_116_077, w_116_078, w_116_079, w_116_081, w_116_083, w_116_084, w_116_086, w_116_088, w_116_095, w_116_096, w_116_097, w_116_099, w_116_103, w_116_104, w_116_111, w_116_112, w_116_115, w_116_117, w_116_121, w_116_123, w_116_124, w_116_126, w_116_130, w_116_131, w_116_133, w_116_135, w_116_136, w_116_139, w_116_142, w_116_144, w_116_146, w_116_148, w_116_149, w_116_151, w_116_155, w_116_159, w_116_160, w_116_162, w_116_163, w_116_165, w_116_166, w_116_167, w_116_170, w_116_174, w_116_175, w_116_176, w_116_177, w_116_178, w_116_180, w_116_181, w_116_184, w_116_185, w_116_186, w_116_187, w_116_188, w_116_189, w_116_191, w_116_193, w_116_194, w_116_197, w_116_199, w_116_201, w_116_202, w_116_204, w_116_205, w_116_206, w_116_211, w_116_212, w_116_213, w_116_214, w_116_215, w_116_217, w_116_221, w_116_222, w_116_224, w_116_225, w_116_227, w_116_228, w_116_231, w_116_233, w_116_235, w_116_236, w_116_237, w_116_239, w_116_240, w_116_241, w_116_242, w_116_243, w_116_244, w_116_246, w_116_248, w_116_252, w_116_253, w_116_254, w_116_255, w_116_256, w_116_258, w_116_259, w_116_260, w_116_261, w_116_262, w_116_265, w_116_268, w_116_273, w_116_274, w_116_275, w_116_277, w_116_279, w_116_282, w_116_285, w_116_286, w_116_289, w_116_290, w_116_291, w_116_293, w_116_295, w_116_298, w_116_299, w_116_300, w_116_302, w_116_304, w_116_306, w_116_307, w_116_308, w_116_312, w_116_314, w_116_315, w_116_317, w_116_318, w_116_319, w_116_320, w_116_322, w_116_329, w_116_330, w_116_332, w_116_336, w_116_337, w_116_339, w_116_340, w_116_343, w_116_344, w_116_347, w_116_348, w_116_350, w_116_352, w_116_356, w_116_358, w_116_359, w_116_360, w_116_361, w_116_363, w_116_364, w_116_365, w_116_367, w_116_368, w_116_369, w_116_371, w_116_372, w_116_374, w_116_377, w_116_378, w_116_379, w_116_380, w_116_383, w_116_385, w_116_386, w_116_389, w_116_390, w_116_391, w_116_395, w_116_396, w_116_397, w_116_398, w_116_399, w_116_401, w_116_402, w_116_403, w_116_404, w_116_405, w_116_408, w_116_409, w_116_410, w_116_411, w_116_412, w_116_414, w_116_417, w_116_420, w_116_421, w_116_423, w_116_424, w_116_427, w_116_428, w_116_429, w_116_430, w_116_431, w_116_433, w_116_434, w_116_438, w_116_439, w_116_442, w_116_443, w_116_445, w_116_447, w_116_448, w_116_449, w_116_452, w_116_454, w_116_456, w_116_459, w_116_461, w_116_464, w_116_465, w_116_466, w_116_469, w_116_470, w_116_471, w_116_473, w_116_475, w_116_477, w_116_479, w_116_480, w_116_484, w_116_485, w_116_486, w_116_487, w_116_488, w_116_490, w_116_492, w_116_497, w_116_502, w_116_505, w_116_506, w_116_508, w_116_509, w_116_510, w_116_514, w_116_517, w_116_518, w_116_519, w_116_523, w_116_524, w_116_525, w_116_526, w_116_527, w_116_528, w_116_534, w_116_535, w_116_536, w_116_537, w_116_538, w_116_540, w_116_542, w_116_544, w_116_545, w_116_548, w_116_554, w_116_556, w_116_560, w_116_564, w_116_572, w_116_573, w_116_574, w_116_575, w_116_576, w_116_577, w_116_578, w_116_581, w_116_582, w_116_583, w_116_586, w_116_587, w_116_589, w_116_590, w_116_591, w_116_598, w_116_599, w_116_600, w_116_603, w_116_607, w_116_608, w_116_610, w_116_611, w_116_612, w_116_616, w_116_618, w_116_619, w_116_621, w_116_622, w_116_623, w_116_624, w_116_625, w_116_626, w_116_627, w_116_628, w_116_629, w_116_632, w_116_633, w_116_634, w_116_635, w_116_636, w_116_637, w_116_638, w_116_640, w_116_642, w_116_643, w_116_647, w_116_649, w_116_650, w_116_652, w_116_653, w_116_654, w_116_655, w_116_656, w_116_658, w_116_659, w_116_660, w_116_662, w_116_663, w_116_664, w_116_667, w_116_668, w_116_669, w_116_671, w_116_673, w_116_674, w_116_677, w_116_680, w_116_681, w_116_682, w_116_683, w_116_684, w_116_685, w_116_686, w_116_687, w_116_688, w_116_690, w_116_691, w_116_692, w_116_693, w_116_695, w_116_697, w_116_699, w_116_700, w_116_701, w_116_703, w_116_705, w_116_708, w_116_713, w_116_714, w_116_715, w_116_716, w_116_717, w_116_718, w_116_720, w_116_723, w_116_724, w_116_725, w_116_727, w_116_729, w_116_730, w_116_731, w_116_734, w_116_735, w_116_736, w_116_738, w_116_739, w_116_740, w_116_742, w_116_746, w_116_747, w_116_748, w_116_749, w_116_751, w_116_752, w_116_754, w_116_755, w_116_757, w_116_759, w_116_760, w_116_761, w_116_762, w_116_768, w_116_770, w_116_771, w_116_773, w_116_774, w_116_775, w_116_778, w_116_779, w_116_780, w_116_781, w_116_782, w_116_783, w_116_785, w_116_786, w_116_788, w_116_790, w_116_792, w_116_793, w_116_798, w_116_801, w_116_802, w_116_803, w_116_804, w_116_805, w_116_807, w_116_808, w_116_810, w_116_812, w_116_814, w_116_815, w_116_816, w_116_817, w_116_818, w_116_823, w_116_825, w_116_827, w_116_828, w_116_829, w_116_830, w_116_833, w_116_835, w_116_837, w_116_840, w_116_841, w_116_842, w_116_845, w_116_846, w_116_849, w_116_851, w_116_853, w_116_855, w_116_861, w_116_862, w_116_863, w_116_864, w_116_866, w_116_868, w_116_869, w_116_871, w_116_872, w_116_873, w_116_874, w_116_880, w_116_883, w_116_884, w_116_887, w_116_888, w_116_889, w_116_890, w_116_892, w_116_894, w_116_896, w_116_897, w_116_898, w_116_900, w_116_901, w_116_904, w_116_905, w_116_908, w_116_909, w_116_911, w_116_913, w_116_914, w_116_918, w_116_919, w_116_920, w_116_922, w_116_923, w_116_925, w_116_927, w_116_933, w_116_935, w_116_936, w_116_937, w_116_941, w_116_944, w_116_946, w_116_948, w_116_949, w_116_950, w_116_952, w_116_957, w_116_959, w_116_960, w_116_965, w_116_967, w_116_968, w_116_969, w_116_970, w_116_971, w_116_975, w_116_976, w_116_978, w_116_981, w_116_982, w_116_983, w_116_988, w_116_989, w_116_990, w_116_991, w_116_994, w_116_996, w_116_997, w_116_999, w_116_1000, w_116_1001, w_116_1004, w_116_1008, w_116_1009, w_116_1013, w_116_1014, w_116_1016, w_116_1017, w_116_1019, w_116_1020, w_116_1021, w_116_1022, w_116_1023, w_116_1025, w_116_1027, w_116_1028, w_116_1030, w_116_1031, w_116_1032, w_116_1034, w_116_1035, w_116_1037, w_116_1038, w_116_1040, w_116_1041, w_116_1042, w_116_1043, w_116_1044, w_116_1048, w_116_1051, w_116_1052, w_116_1053, w_116_1054, w_116_1055, w_116_1056, w_116_1058, w_116_1059, w_116_1060, w_116_1061, w_116_1062, w_116_1064, w_116_1066, w_116_1067, w_116_1068, w_116_1070, w_116_1071, w_116_1072, w_116_1074, w_116_1075, w_116_1076, w_116_1077, w_116_1078, w_116_1079, w_116_1080, w_116_1081, w_116_1082, w_116_1083, w_116_1086, w_116_1087, w_116_1088, w_116_1089, w_116_1091, w_116_1093, w_116_1096, w_116_1098, w_116_1100, w_116_1102, w_116_1104, w_116_1105, w_116_1106, w_116_1107, w_116_1108, w_116_1109, w_116_1112, w_116_1114, w_116_1115, w_116_1120, w_116_1123, w_116_1124, w_116_1127, w_116_1128, w_116_1129, w_116_1130, w_116_1132, w_116_1134, w_116_1137, w_116_1139, w_116_1142, w_116_1144, w_116_1146, w_116_1148, w_116_1149, w_116_1150, w_116_1152, w_116_1154, w_116_1156, w_116_1157, w_116_1160, w_116_1161, w_116_1162, w_116_1163, w_116_1165, w_116_1166, w_116_1167, w_116_1170, w_116_1171, w_116_1174, w_116_1175, w_116_1179, w_116_1182, w_116_1186, w_116_1187, w_116_1188, w_116_1190, w_116_1192, w_116_1193, w_116_1194, w_116_1195, w_116_1196, w_116_1197, w_116_1199, w_116_1200, w_116_1201, w_116_1203, w_116_1204, w_116_1207, w_116_1211, w_116_1214, w_116_1216, w_116_1217, w_116_1220, w_116_1221, w_116_1223, w_116_1224, w_116_1225, w_116_1227, w_116_1228, w_116_1229, w_116_1230, w_116_1231, w_116_1233, w_116_1236, w_116_1239, w_116_1241, w_116_1242, w_116_1244, w_116_1246, w_116_1248, w_116_1249, w_116_1250, w_116_1251, w_116_1255, w_116_1260, w_116_1264, w_116_1267, w_116_1271, w_116_1272, w_116_1273, w_116_1279, w_116_1280, w_116_1281, w_116_1282, w_116_1284, w_116_1285, w_116_1286, w_116_1287, w_116_1288, w_116_1292, w_116_1293, w_116_1295, w_116_1297, w_116_1299, w_116_1300, w_116_1301, w_116_1302, w_116_1304, w_116_1306, w_116_1309, w_116_1310, w_116_1312, w_116_1313, w_116_1317, w_116_1319, w_116_1320, w_116_1322, w_116_1323, w_116_1324, w_116_1325, w_116_1326, w_116_1329, w_116_1330, w_116_1331, w_116_1335, w_116_1336, w_116_1337, w_116_1341, w_116_1344, w_116_1345, w_116_1346, w_116_1347, w_116_1348, w_116_1349, w_116_1351, w_116_1353, w_116_1354, w_116_1356, w_116_1358, w_116_1359, w_116_1364, w_116_1368, w_116_1370, w_116_1371, w_116_1373, w_116_1374, w_116_1375, w_116_1377, w_116_1381, w_116_1383, w_116_1386, w_116_1388, w_116_1390, w_116_1391, w_116_1392, w_116_1394, w_116_1397, w_116_1398, w_116_1399, w_116_1400, w_116_1402, w_116_1404, w_116_1405, w_116_1406, w_116_1409, w_116_1410, w_116_1411, w_116_1412, w_116_1414, w_116_1415, w_116_1416, w_116_1417, w_116_1418, w_116_1419, w_116_1420, w_116_1422, w_116_1423, w_116_1424, w_116_1426, w_116_1427, w_116_1430, w_116_1432, w_116_1434, w_116_1435, w_116_1436, w_116_1437, w_116_1438, w_116_1439, w_116_1441, w_116_1442, w_116_1443, w_116_1444, w_116_1445, w_116_1446, w_116_1449, w_116_1450, w_116_1451, w_116_1452, w_116_1455, w_116_1456, w_116_1459, w_116_1461, w_116_1463, w_116_1464, w_116_1468, w_116_1470, w_116_1471, w_116_1474, w_116_1475, w_116_1476, w_116_1477, w_116_1478, w_116_1481, w_116_1482, w_116_1483, w_116_1484, w_116_1485, w_116_1487, w_116_1488, w_116_1491, w_116_1492, w_116_1493, w_116_1495, w_116_1496, w_116_1499, w_116_1500, w_116_1501, w_116_1502, w_116_1503, w_116_1504, w_116_1505, w_116_1506, w_116_1511, w_116_1512, w_116_1513, w_116_1515, w_116_1518, w_116_1519, w_116_1521, w_116_1522, w_116_1523, w_116_1524, w_116_1527, w_116_1528, w_116_1529, w_116_1530, w_116_1531, w_116_1536, w_116_1537, w_116_1539, w_116_1540, w_116_1541, w_116_1542, w_116_1543, w_116_1544, w_116_1545, w_116_1546, w_116_1547, w_116_1553, w_116_1555, w_116_1556, w_116_1557, w_116_1558, w_116_1560, w_116_1561, w_116_1563, w_116_1564, w_116_1566, w_116_1567, w_116_1568, w_116_1569, w_116_1570, w_116_1572, w_116_1573, w_116_1574, w_116_1576, w_116_1577, w_116_1579, w_116_1583, w_116_1592, w_116_1596, w_116_1600, w_116_1601, w_116_1603, w_116_1604, w_116_1605, w_116_1606, w_116_1608, w_116_1610, w_116_1611, w_116_1613, w_116_1614, w_116_1616, w_116_1618, w_116_1619, w_116_1621, w_116_1622, w_116_1635, w_116_1639, w_116_1640, w_116_1644, w_116_1646, w_116_1649, w_116_1651, w_116_1653, w_116_1655, w_116_1656, w_116_1658, w_116_1659, w_116_1660, w_116_1662, w_116_1663, w_116_1665, w_116_1671, w_116_1673, w_116_1675, w_116_1677, w_116_1678, w_116_1679, w_116_1685, w_116_1686, w_116_1687, w_116_1688, w_116_1690, w_116_1692, w_116_1696, w_116_1697, w_116_1698, w_116_1699, w_116_1700, w_116_1701, w_116_1703, w_116_1704, w_116_1705, w_116_1706;
  wire w_117_002, w_117_007, w_117_011, w_117_013, w_117_015, w_117_018, w_117_019, w_117_021, w_117_022, w_117_024, w_117_027, w_117_028, w_117_030, w_117_033, w_117_034, w_117_035, w_117_038, w_117_041, w_117_042, w_117_043, w_117_044, w_117_047, w_117_048, w_117_054, w_117_057, w_117_058, w_117_060, w_117_065, w_117_067, w_117_068, w_117_071, w_117_073, w_117_074, w_117_081, w_117_082, w_117_088, w_117_091, w_117_094, w_117_095, w_117_100, w_117_101, w_117_106, w_117_107, w_117_111, w_117_112, w_117_115, w_117_121, w_117_124, w_117_125, w_117_126, w_117_128, w_117_129, w_117_136, w_117_140, w_117_141, w_117_143, w_117_147, w_117_149, w_117_151, w_117_153, w_117_160, w_117_163, w_117_165, w_117_167, w_117_168, w_117_170, w_117_171, w_117_172, w_117_173, w_117_174, w_117_175, w_117_177, w_117_178, w_117_179, w_117_180, w_117_181, w_117_182, w_117_183, w_117_184, w_117_186, w_117_192, w_117_194, w_117_197, w_117_199, w_117_203, w_117_207, w_117_208, w_117_209, w_117_211, w_117_213, w_117_215, w_117_218, w_117_221, w_117_225, w_117_230, w_117_236, w_117_237, w_117_238, w_117_239, w_117_246, w_117_255, w_117_256, w_117_257, w_117_259, w_117_260, w_117_261, w_117_262, w_117_264, w_117_265, w_117_266, w_117_271, w_117_272, w_117_279, w_117_282, w_117_283, w_117_287, w_117_288, w_117_289, w_117_290, w_117_291, w_117_293, w_117_295, w_117_298, w_117_300, w_117_301, w_117_306, w_117_309, w_117_311, w_117_316, w_117_318, w_117_320, w_117_321, w_117_322, w_117_325, w_117_328, w_117_329, w_117_333, w_117_338, w_117_341, w_117_344, w_117_345, w_117_346, w_117_348, w_117_349, w_117_353, w_117_354, w_117_360, w_117_364, w_117_365, w_117_366, w_117_368, w_117_370, w_117_373, w_117_378, w_117_382, w_117_383, w_117_385, w_117_386, w_117_392, w_117_397, w_117_400, w_117_401, w_117_402, w_117_403, w_117_404, w_117_406, w_117_408, w_117_410, w_117_411, w_117_415, w_117_418, w_117_419, w_117_424, w_117_427, w_117_428, w_117_430, w_117_431, w_117_433, w_117_434, w_117_438, w_117_440, w_117_443, w_117_444, w_117_447, w_117_450, w_117_451, w_117_452, w_117_454, w_117_457, w_117_461, w_117_464, w_117_465, w_117_468, w_117_470, w_117_475, w_117_476, w_117_477, w_117_479, w_117_482, w_117_484, w_117_485, w_117_489, w_117_491, w_117_492, w_117_496, w_117_499, w_117_500, w_117_501, w_117_502, w_117_510, w_117_513, w_117_514, w_117_518, w_117_519, w_117_522, w_117_526, w_117_527, w_117_528, w_117_530, w_117_533, w_117_534, w_117_535, w_117_539, w_117_541, w_117_542, w_117_543, w_117_545, w_117_546, w_117_548, w_117_556, w_117_557, w_117_562, w_117_563, w_117_565, w_117_570, w_117_572, w_117_573, w_117_575, w_117_578, w_117_580, w_117_582, w_117_585, w_117_589, w_117_591, w_117_592, w_117_598, w_117_599, w_117_600, w_117_601, w_117_602, w_117_603, w_117_610, w_117_614, w_117_618, w_117_620, w_117_623, w_117_624, w_117_625, w_117_626, w_117_628, w_117_632, w_117_637, w_117_639, w_117_641, w_117_644, w_117_645, w_117_647, w_117_650, w_117_654, w_117_657, w_117_659, w_117_663, w_117_666, w_117_667, w_117_669, w_117_672, w_117_673, w_117_677, w_117_679, w_117_682, w_117_685, w_117_686, w_117_688, w_117_689, w_117_691, w_117_699, w_117_700, w_117_701, w_117_704, w_117_708, w_117_709, w_117_710, w_117_711, w_117_712, w_117_714, w_117_715, w_117_717, w_117_718, w_117_719, w_117_720, w_117_721, w_117_722, w_117_725, w_117_727, w_117_732, w_117_734, w_117_735, w_117_736, w_117_738, w_117_741, w_117_742, w_117_746, w_117_749, w_117_751, w_117_768, w_117_771, w_117_772, w_117_773, w_117_779, w_117_784, w_117_786, w_117_798, w_117_799, w_117_802, w_117_804, w_117_805, w_117_806, w_117_808, w_117_809, w_117_811, w_117_812, w_117_818, w_117_821, w_117_825, w_117_826, w_117_828, w_117_831, w_117_833, w_117_835, w_117_836, w_117_842, w_117_843, w_117_844, w_117_845, w_117_846, w_117_847, w_117_850, w_117_851, w_117_854, w_117_861, w_117_862, w_117_864, w_117_865, w_117_870, w_117_872, w_117_878, w_117_879, w_117_881, w_117_883, w_117_884, w_117_886, w_117_889, w_117_890, w_117_892, w_117_894, w_117_896, w_117_897, w_117_898, w_117_902, w_117_909, w_117_911, w_117_914, w_117_918, w_117_923, w_117_925, w_117_928, w_117_929, w_117_930, w_117_934, w_117_935, w_117_937, w_117_940, w_117_948, w_117_950, w_117_952, w_117_953, w_117_963, w_117_964, w_117_969, w_117_970, w_117_973, w_117_977, w_117_980, w_117_982, w_117_985, w_117_987, w_117_988, w_117_993, w_117_996, w_117_999, w_117_1000, w_117_1001, w_117_1004, w_117_1008, w_117_1009, w_117_1010, w_117_1011, w_117_1016, w_117_1017, w_117_1019, w_117_1025, w_117_1026, w_117_1030, w_117_1032, w_117_1034, w_117_1036, w_117_1039, w_117_1044, w_117_1048, w_117_1049, w_117_1050, w_117_1053, w_117_1057, w_117_1058, w_117_1059, w_117_1061, w_117_1062, w_117_1065, w_117_1067, w_117_1069, w_117_1070, w_117_1071, w_117_1073, w_117_1074, w_117_1076, w_117_1078, w_117_1082, w_117_1084, w_117_1086, w_117_1087, w_117_1089, w_117_1104, w_117_1106, w_117_1107, w_117_1108, w_117_1112, w_117_1115, w_117_1117, w_117_1119, w_117_1121, w_117_1122, w_117_1125, w_117_1130, w_117_1133, w_117_1135, w_117_1140, w_117_1142, w_117_1147, w_117_1148, w_117_1153, w_117_1156, w_117_1159, w_117_1160, w_117_1162, w_117_1166, w_117_1167, w_117_1171, w_117_1178, w_117_1180, w_117_1182, w_117_1183, w_117_1187, w_117_1188, w_117_1194, w_117_1199, w_117_1200, w_117_1202, w_117_1203, w_117_1204, w_117_1206, w_117_1208, w_117_1211, w_117_1212, w_117_1213, w_117_1214, w_117_1216, w_117_1221, w_117_1223, w_117_1226, w_117_1227, w_117_1230, w_117_1232, w_117_1233, w_117_1234, w_117_1236, w_117_1237, w_117_1238, w_117_1241, w_117_1242, w_117_1243, w_117_1244, w_117_1249, w_117_1256, w_117_1258, w_117_1260, w_117_1263, w_117_1265, w_117_1266, w_117_1269, w_117_1274, w_117_1275, w_117_1279, w_117_1280, w_117_1282, w_117_1283, w_117_1289, w_117_1290, w_117_1292, w_117_1293, w_117_1299, w_117_1303, w_117_1308, w_117_1309, w_117_1317, w_117_1320, w_117_1326, w_117_1327, w_117_1328, w_117_1330, w_117_1334, w_117_1335, w_117_1336, w_117_1339, w_117_1340, w_117_1341, w_117_1342, w_117_1344, w_117_1348, w_117_1350, w_117_1352, w_117_1355, w_117_1360, w_117_1361, w_117_1362, w_117_1364, w_117_1366, w_117_1368, w_117_1369, w_117_1370, w_117_1371, w_117_1373, w_117_1376, w_117_1377, w_117_1379, w_117_1385, w_117_1394, w_117_1396, w_117_1398, w_117_1400, w_117_1401, w_117_1403, w_117_1408, w_117_1409, w_117_1412, w_117_1413, w_117_1414, w_117_1415, w_117_1416, w_117_1417, w_117_1419, w_117_1421, w_117_1424, w_117_1426, w_117_1433, w_117_1434, w_117_1436, w_117_1437, w_117_1438, w_117_1439, w_117_1442, w_117_1443, w_117_1446, w_117_1447, w_117_1452, w_117_1453, w_117_1454, w_117_1455, w_117_1456, w_117_1458, w_117_1464, w_117_1467, w_117_1469, w_117_1473, w_117_1476, w_117_1477, w_117_1479, w_117_1481, w_117_1485, w_117_1489, w_117_1493, w_117_1494, w_117_1495, w_117_1496, w_117_1499, w_117_1500, w_117_1502, w_117_1503, w_117_1507, w_117_1508, w_117_1509, w_117_1513, w_117_1514, w_117_1516, w_117_1520, w_117_1521, w_117_1522, w_117_1525, w_117_1526, w_117_1527, w_117_1529, w_117_1530, w_117_1532, w_117_1533, w_117_1534, w_117_1540, w_117_1541, w_117_1542, w_117_1547, w_117_1549, w_117_1551, w_117_1555, w_117_1556, w_117_1559, w_117_1561, w_117_1567, w_117_1573, w_117_1577, w_117_1578, w_117_1581, w_117_1582, w_117_1584, w_117_1586, w_117_1591, w_117_1604, w_117_1610, w_117_1617, w_117_1618, w_117_1619, w_117_1621, w_117_1622, w_117_1627, w_117_1628, w_117_1629, w_117_1631, w_117_1634, w_117_1637, w_117_1645, w_117_1656, w_117_1659, w_117_1663, w_117_1665, w_117_1666, w_117_1668, w_117_1674, w_117_1676, w_117_1679, w_117_1683, w_117_1687, w_117_1693, w_117_1696, w_117_1699, w_117_1701, w_117_1703, w_117_1705, w_117_1711, w_117_1720, w_117_1730, w_117_1732, w_117_1733, w_117_1737, w_117_1744, w_117_1746, w_117_1751, w_117_1752, w_117_1755, w_117_1756, w_117_1763, w_117_1764, w_117_1768, w_117_1770, w_117_1771, w_117_1773, w_117_1775, w_117_1776, w_117_1779, w_117_1780, w_117_1797, w_117_1802, w_117_1817, w_117_1823, w_117_1830, w_117_1839, w_117_1841, w_117_1842, w_117_1849, w_117_1851, w_117_1855, w_117_1860, w_117_1864, w_117_1874, w_117_1877, w_117_1879, w_117_1892, w_117_1895, w_117_1896, w_117_1898, w_117_1899, w_117_1906, w_117_1914, w_117_1916, w_117_1921, w_117_1923, w_117_1926, w_117_1928, w_117_1932, w_117_1933, w_117_1934, w_117_1937, w_117_1939, w_117_1943, w_117_1954, w_117_1959, w_117_1961, w_117_1970, w_117_1976, w_117_1981, w_117_1983, w_117_1985, w_117_1986, w_117_1995, w_117_1998, w_117_1999, w_117_2001, w_117_2010, w_117_2022, w_117_2024, w_117_2029, w_117_2047, w_117_2049, w_117_2051, w_117_2055, w_117_2060, w_117_2062, w_117_2066, w_117_2069, w_117_2072, w_117_2073, w_117_2074, w_117_2082, w_117_2085, w_117_2087, w_117_2094, w_117_2102, w_117_2109, w_117_2112, w_117_2114, w_117_2115, w_117_2119, w_117_2121, w_117_2135, w_117_2143, w_117_2148, w_117_2150, w_117_2154, w_117_2157, w_117_2160, w_117_2162, w_117_2163, w_117_2165, w_117_2167, w_117_2171, w_117_2172, w_117_2175, w_117_2177, w_117_2178, w_117_2181, w_117_2182, w_117_2183, w_117_2187, w_117_2197, w_117_2204, w_117_2211, w_117_2213, w_117_2215, w_117_2219, w_117_2220, w_117_2224, w_117_2228, w_117_2240, w_117_2254, w_117_2269, w_117_2277, w_117_2284, w_117_2292, w_117_2296, w_117_2300, w_117_2304, w_117_2306, w_117_2307, w_117_2308, w_117_2310, w_117_2312, w_117_2313, w_117_2316, w_117_2321, w_117_2323, w_117_2324, w_117_2327, w_117_2335, w_117_2339, w_117_2340, w_117_2343, w_117_2347, w_117_2350, w_117_2353, w_117_2362, w_117_2372, w_117_2373, w_117_2374, w_117_2375, w_117_2379, w_117_2390, w_117_2392, w_117_2395, w_117_2403, w_117_2417, w_117_2427, w_117_2433, w_117_2441, w_117_2449, w_117_2450, w_117_2451, w_117_2456, w_117_2458, w_117_2467, w_117_2471, w_117_2472, w_117_2473, w_117_2482, w_117_2483, w_117_2488, w_117_2489, w_117_2490, w_117_2500, w_117_2505, w_117_2506, w_117_2510, w_117_2517, w_117_2520, w_117_2522, w_117_2526, w_117_2528, w_117_2531, w_117_2533, w_117_2537, w_117_2544, w_117_2546, w_117_2548, w_117_2555, w_117_2562, w_117_2565, w_117_2568, w_117_2571, w_117_2582, w_117_2586, w_117_2593, w_117_2594, w_117_2596, w_117_2597, w_117_2603, w_117_2612, w_117_2615, w_117_2622, w_117_2625, w_117_2626, w_117_2627, w_117_2629, w_117_2632, w_117_2657, w_117_2658, w_117_2662, w_117_2663, w_117_2664, w_117_2665, w_117_2666, w_117_2668, w_117_2678, w_117_2680, w_117_2692, w_117_2706, w_117_2712, w_117_2716, w_117_2720, w_117_2721, w_117_2723, w_117_2728, w_117_2734, w_117_2737, w_117_2742, w_117_2743, w_117_2747, w_117_2748, w_117_2761, w_117_2767, w_117_2769, w_117_2772, w_117_2775, w_117_2783, w_117_2792, w_117_2797, w_117_2798, w_117_2805, w_117_2806, w_117_2810, w_117_2818, w_117_2825, w_117_2829, w_117_2837, w_117_2840, w_117_2841, w_117_2843, w_117_2844, w_117_2846, w_117_2847, w_117_2850, w_117_2852, w_117_2853, w_117_2859, w_117_2866, w_117_2870, w_117_2873, w_117_2876, w_117_2879, w_117_2880, w_117_2881, w_117_2882, w_117_2888, w_117_2899, w_117_2902, w_117_2903, w_117_2904, w_117_2909, w_117_2911, w_117_2913, w_117_2916, w_117_2921, w_117_2922, w_117_2925, w_117_2926, w_117_2927, w_117_2931, w_117_2932, w_117_2937, w_117_2941, w_117_2944, w_117_2945, w_117_2951, w_117_2952, w_117_2955, w_117_2957, w_117_2959, w_117_2969, w_117_2973, w_117_2976, w_117_2977, w_117_2983, w_117_2990, w_117_2993, w_117_2996, w_117_3003, w_117_3012, w_117_3014, w_117_3015, w_117_3017, w_117_3023, w_117_3024, w_117_3029, w_117_3039, w_117_3043, w_117_3049, w_117_3051, w_117_3052, w_117_3053, w_117_3055, w_117_3058, w_117_3075, w_117_3077, w_117_3078, w_117_3082, w_117_3083, w_117_3090, w_117_3093, w_117_3102, w_117_3106, w_117_3111, w_117_3117, w_117_3118, w_117_3122, w_117_3124, w_117_3131, w_117_3137, w_117_3140, w_117_3143, w_117_3145, w_117_3160, w_117_3162, w_117_3171, w_117_3179, w_117_3183, w_117_3195, w_117_3201, w_117_3206, w_117_3207, w_117_3213, w_117_3218, w_117_3220, w_117_3221, w_117_3227, w_117_3229, w_117_3233, w_117_3238, w_117_3239, w_117_3241, w_117_3249, w_117_3251, w_117_3253, w_117_3255, w_117_3256, w_117_3257, w_117_3268, w_117_3270, w_117_3271, w_117_3278, w_117_3280, w_117_3284, w_117_3286, w_117_3288, w_117_3296, w_117_3299, w_117_3300, w_117_3307, w_117_3324, w_117_3325, w_117_3326, w_117_3328, w_117_3329, w_117_3337, w_117_3338, w_117_3346, w_117_3354, w_117_3360, w_117_3362, w_117_3384, w_117_3388, w_117_3393, w_117_3396, w_117_3407, w_117_3409, w_117_3410, w_117_3413, w_117_3416, w_117_3419, w_117_3420, w_117_3421, w_117_3425, w_117_3428, w_117_3429, w_117_3430, w_117_3431, w_117_3434, w_117_3435, w_117_3438, w_117_3443, w_117_3447, w_117_3448, w_117_3449, w_117_3451, w_117_3452, w_117_3453, w_117_3454, w_117_3455;
  wire w_118_002, w_118_003, w_118_006, w_118_010, w_118_011, w_118_013, w_118_015, w_118_016, w_118_026, w_118_028, w_118_030, w_118_031, w_118_033, w_118_045, w_118_048, w_118_052, w_118_053, w_118_054, w_118_058, w_118_061, w_118_062, w_118_063, w_118_065, w_118_067, w_118_071, w_118_072, w_118_074, w_118_080, w_118_084, w_118_088, w_118_089, w_118_091, w_118_092, w_118_095, w_118_098, w_118_100, w_118_102, w_118_104, w_118_110, w_118_111, w_118_112, w_118_119, w_118_120, w_118_123, w_118_124, w_118_126, w_118_131, w_118_133, w_118_135, w_118_138, w_118_139, w_118_140, w_118_142, w_118_143, w_118_145, w_118_147, w_118_148, w_118_150, w_118_154, w_118_158, w_118_159, w_118_160, w_118_162, w_118_164, w_118_165, w_118_166, w_118_170, w_118_174, w_118_182, w_118_184, w_118_187, w_118_188, w_118_189, w_118_191, w_118_196, w_118_197, w_118_198, w_118_199, w_118_201, w_118_208, w_118_209, w_118_212, w_118_214, w_118_216, w_118_219, w_118_220, w_118_222, w_118_223, w_118_225, w_118_227, w_118_229, w_118_231, w_118_237, w_118_238, w_118_245, w_118_246, w_118_248, w_118_250, w_118_251, w_118_253, w_118_255, w_118_258, w_118_259, w_118_262, w_118_263, w_118_266, w_118_271, w_118_273, w_118_275, w_118_276, w_118_277, w_118_281, w_118_289, w_118_291, w_118_292, w_118_293, w_118_295, w_118_298, w_118_300, w_118_301, w_118_302, w_118_304, w_118_305, w_118_307, w_118_309, w_118_313, w_118_314, w_118_317, w_118_318, w_118_326, w_118_328, w_118_329, w_118_330, w_118_331, w_118_334, w_118_336, w_118_337, w_118_340, w_118_344, w_118_349, w_118_350, w_118_353, w_118_355, w_118_356, w_118_357, w_118_366, w_118_369, w_118_370, w_118_371, w_118_373, w_118_375, w_118_378, w_118_380, w_118_382, w_118_383, w_118_384, w_118_389, w_118_390, w_118_399, w_118_402, w_118_403, w_118_404, w_118_414, w_118_415, w_118_416, w_118_418, w_118_420, w_118_421, w_118_422, w_118_424, w_118_427, w_118_428, w_118_430, w_118_431, w_118_435, w_118_438, w_118_440, w_118_442, w_118_444, w_118_445, w_118_447, w_118_449, w_118_452, w_118_456, w_118_458, w_118_463, w_118_464, w_118_466, w_118_468, w_118_469, w_118_470, w_118_472, w_118_474, w_118_476, w_118_477, w_118_480, w_118_481, w_118_485, w_118_487, w_118_488, w_118_490, w_118_492, w_118_493, w_118_496, w_118_499, w_118_503, w_118_505, w_118_507, w_118_513, w_118_515, w_118_516, w_118_517, w_118_518, w_118_519, w_118_520, w_118_526, w_118_528, w_118_529, w_118_530, w_118_532, w_118_533, w_118_534, w_118_535, w_118_538, w_118_539, w_118_540, w_118_541, w_118_543, w_118_545, w_118_547, w_118_549, w_118_560, w_118_563, w_118_566, w_118_567, w_118_573, w_118_579, w_118_583, w_118_584, w_118_585, w_118_588, w_118_590, w_118_599, w_118_606, w_118_608, w_118_610, w_118_611, w_118_616, w_118_617, w_118_620, w_118_626, w_118_627, w_118_629, w_118_631, w_118_632, w_118_635, w_118_637, w_118_639, w_118_642, w_118_644, w_118_645, w_118_648, w_118_649, w_118_651, w_118_652, w_118_657, w_118_659, w_118_660, w_118_661, w_118_662, w_118_664, w_118_665, w_118_666, w_118_670, w_118_673, w_118_675, w_118_687, w_118_693, w_118_695, w_118_698, w_118_700, w_118_703, w_118_704, w_118_713, w_118_717, w_118_720, w_118_721, w_118_722, w_118_723, w_118_725, w_118_727, w_118_729, w_118_730, w_118_733, w_118_734, w_118_735, w_118_736, w_118_737, w_118_740, w_118_743, w_118_747, w_118_748, w_118_749, w_118_751, w_118_753, w_118_754, w_118_755, w_118_756, w_118_757, w_118_758, w_118_760, w_118_763, w_118_764, w_118_766, w_118_769, w_118_771, w_118_772, w_118_777, w_118_778, w_118_780, w_118_783, w_118_786, w_118_787, w_118_792, w_118_798, w_118_799, w_118_801, w_118_802, w_118_804, w_118_805, w_118_806, w_118_808, w_118_810, w_118_812, w_118_818, w_118_821, w_118_823, w_118_825, w_118_828, w_118_830, w_118_831, w_118_833, w_118_835, w_118_838, w_118_840, w_118_841, w_118_844, w_118_852, w_118_854, w_118_859, w_118_863, w_118_870, w_118_872, w_118_873, w_118_874, w_118_877, w_118_878, w_118_885, w_118_888, w_118_890, w_118_897, w_118_899, w_118_901, w_118_905, w_118_906, w_118_907, w_118_908, w_118_909, w_118_912, w_118_913, w_118_917, w_118_919, w_118_926, w_118_927, w_118_937, w_118_939, w_118_940, w_118_946, w_118_948, w_118_950, w_118_952, w_118_953, w_118_955, w_118_956, w_118_958, w_118_960, w_118_961, w_118_965, w_118_967, w_118_968, w_118_970, w_118_971, w_118_975, w_118_977, w_118_983, w_118_988, w_118_991, w_118_993, w_118_994, w_118_995, w_118_996, w_118_997, w_118_998, w_118_999, w_118_1001, w_118_1002, w_118_1004, w_118_1007, w_118_1008, w_118_1011, w_118_1012, w_118_1014, w_118_1016, w_118_1017, w_118_1018, w_118_1021, w_118_1023, w_118_1024, w_118_1025, w_118_1030, w_118_1034, w_118_1035, w_118_1037, w_118_1039, w_118_1041, w_118_1049, w_118_1052, w_118_1054, w_118_1056, w_118_1059, w_118_1062, w_118_1065, w_118_1077, w_118_1078, w_118_1080, w_118_1084, w_118_1085, w_118_1087, w_118_1089, w_118_1090, w_118_1092, w_118_1096, w_118_1100, w_118_1101, w_118_1103, w_118_1105, w_118_1114, w_118_1119, w_118_1120, w_118_1123, w_118_1125, w_118_1131, w_118_1134, w_118_1136, w_118_1139, w_118_1140, w_118_1143, w_118_1144, w_118_1147, w_118_1148, w_118_1150, w_118_1154, w_118_1155, w_118_1156, w_118_1157, w_118_1158, w_118_1159, w_118_1160, w_118_1163, w_118_1164, w_118_1167, w_118_1170, w_118_1175, w_118_1180, w_118_1183, w_118_1185, w_118_1186, w_118_1188, w_118_1196, w_118_1199, w_118_1203, w_118_1205, w_118_1210, w_118_1221, w_118_1222, w_118_1223, w_118_1224, w_118_1225, w_118_1226, w_118_1228, w_118_1234, w_118_1235, w_118_1237, w_118_1240, w_118_1241, w_118_1244, w_118_1246, w_118_1247, w_118_1249, w_118_1255, w_118_1257, w_118_1259, w_118_1260, w_118_1264, w_118_1267, w_118_1270, w_118_1271, w_118_1273, w_118_1275, w_118_1276, w_118_1277, w_118_1279, w_118_1283, w_118_1287, w_118_1288, w_118_1292, w_118_1294, w_118_1297, w_118_1298, w_118_1300, w_118_1302, w_118_1303, w_118_1304, w_118_1309, w_118_1315, w_118_1316, w_118_1317, w_118_1318, w_118_1319, w_118_1322, w_118_1325, w_118_1326, w_118_1328, w_118_1330, w_118_1342, w_118_1349, w_118_1351, w_118_1354, w_118_1357, w_118_1358, w_118_1359, w_118_1360, w_118_1365, w_118_1368, w_118_1369, w_118_1371, w_118_1372, w_118_1383, w_118_1384, w_118_1385, w_118_1386, w_118_1387, w_118_1389, w_118_1390, w_118_1392, w_118_1398, w_118_1399, w_118_1400, w_118_1412, w_118_1413, w_118_1420, w_118_1432, w_118_1433, w_118_1434, w_118_1436, w_118_1437, w_118_1439, w_118_1444, w_118_1449, w_118_1450, w_118_1465, w_118_1466, w_118_1468, w_118_1476, w_118_1482, w_118_1484, w_118_1485, w_118_1487, w_118_1489, w_118_1492, w_118_1496, w_118_1502, w_118_1508, w_118_1516, w_118_1518, w_118_1522, w_118_1528, w_118_1529, w_118_1544, w_118_1545, w_118_1551, w_118_1555, w_118_1558, w_118_1559, w_118_1560, w_118_1561, w_118_1563, w_118_1565, w_118_1572, w_118_1575, w_118_1580, w_118_1581, w_118_1590, w_118_1591, w_118_1598, w_118_1601, w_118_1606, w_118_1609, w_118_1610, w_118_1616, w_118_1628, w_118_1632, w_118_1633, w_118_1634, w_118_1640, w_118_1647, w_118_1648, w_118_1653, w_118_1660, w_118_1661, w_118_1664, w_118_1666, w_118_1674, w_118_1675, w_118_1683, w_118_1693, w_118_1696, w_118_1699, w_118_1703, w_118_1712, w_118_1718, w_118_1720, w_118_1721, w_118_1725, w_118_1726, w_118_1730, w_118_1731, w_118_1738, w_118_1740, w_118_1742, w_118_1749, w_118_1754, w_118_1757, w_118_1758, w_118_1761, w_118_1765, w_118_1769, w_118_1772, w_118_1775, w_118_1778, w_118_1780, w_118_1784, w_118_1789, w_118_1790, w_118_1792, w_118_1793, w_118_1799, w_118_1805, w_118_1806, w_118_1813, w_118_1818, w_118_1819, w_118_1834, w_118_1837, w_118_1846, w_118_1853, w_118_1855, w_118_1859, w_118_1863, w_118_1865, w_118_1867, w_118_1883, w_118_1897, w_118_1903, w_118_1906, w_118_1910, w_118_1914, w_118_1917, w_118_1922, w_118_1926, w_118_1928, w_118_1934, w_118_1936, w_118_1937, w_118_1944, w_118_1946, w_118_1948, w_118_1949, w_118_1950, w_118_1972, w_118_1981, w_118_1986, w_118_1987, w_118_1988, w_118_1990, w_118_1992, w_118_1996, w_118_1997, w_118_2002, w_118_2006, w_118_2007, w_118_2008, w_118_2011, w_118_2014, w_118_2020, w_118_2021, w_118_2026, w_118_2028, w_118_2033, w_118_2038, w_118_2047, w_118_2052, w_118_2053, w_118_2060, w_118_2061, w_118_2064, w_118_2067, w_118_2068, w_118_2072, w_118_2077, w_118_2080, w_118_2087, w_118_2088, w_118_2091, w_118_2099, w_118_2111, w_118_2114, w_118_2115, w_118_2116, w_118_2117, w_118_2118, w_118_2121, w_118_2124, w_118_2128, w_118_2130, w_118_2138, w_118_2147, w_118_2148, w_118_2149, w_118_2151, w_118_2153, w_118_2155, w_118_2158, w_118_2160, w_118_2162, w_118_2163, w_118_2165, w_118_2181, w_118_2184, w_118_2188, w_118_2191, w_118_2193, w_118_2197, w_118_2206, w_118_2207, w_118_2222, w_118_2225, w_118_2228, w_118_2230, w_118_2234, w_118_2236, w_118_2239, w_118_2240, w_118_2247, w_118_2254, w_118_2260, w_118_2264, w_118_2266, w_118_2268, w_118_2269, w_118_2272, w_118_2274, w_118_2281, w_118_2283, w_118_2284, w_118_2292, w_118_2297, w_118_2301, w_118_2306, w_118_2310, w_118_2311, w_118_2312, w_118_2329, w_118_2332, w_118_2337, w_118_2339, w_118_2340, w_118_2341, w_118_2347, w_118_2348, w_118_2349, w_118_2355, w_118_2368, w_118_2369, w_118_2374, w_118_2375, w_118_2378, w_118_2380, w_118_2386, w_118_2387, w_118_2394, w_118_2397, w_118_2404, w_118_2409, w_118_2412, w_118_2415, w_118_2423, w_118_2424, w_118_2428, w_118_2429, w_118_2437, w_118_2439, w_118_2443, w_118_2446, w_118_2453, w_118_2454, w_118_2458, w_118_2460, w_118_2463, w_118_2475, w_118_2485, w_118_2486, w_118_2489, w_118_2490, w_118_2491, w_118_2494, w_118_2495, w_118_2496, w_118_2502, w_118_2503, w_118_2508, w_118_2510, w_118_2514, w_118_2519, w_118_2521, w_118_2525, w_118_2526, w_118_2528, w_118_2529, w_118_2531, w_118_2543, w_118_2544, w_118_2547, w_118_2549, w_118_2553, w_118_2557, w_118_2559, w_118_2563, w_118_2567, w_118_2568, w_118_2575, w_118_2577, w_118_2587, w_118_2589, w_118_2597, w_118_2599, w_118_2600, w_118_2606, w_118_2610, w_118_2617, w_118_2621, w_118_2625, w_118_2635, w_118_2638, w_118_2644, w_118_2652, w_118_2658, w_118_2662, w_118_2663, w_118_2665, w_118_2669, w_118_2670, w_118_2675, w_118_2679, w_118_2689, w_118_2695, w_118_2700, w_118_2701, w_118_2710, w_118_2716, w_118_2717, w_118_2718, w_118_2720, w_118_2721, w_118_2722, w_118_2723, w_118_2728, w_118_2729, w_118_2734, w_118_2742, w_118_2743, w_118_2746, w_118_2762, w_118_2766, w_118_2771, w_118_2785, w_118_2792, w_118_2798, w_118_2802, w_118_2814, w_118_2815, w_118_2817, w_118_2818, w_118_2820, w_118_2826, w_118_2827, w_118_2832, w_118_2843, w_118_2846, w_118_2848, w_118_2851, w_118_2853, w_118_2857, w_118_2864, w_118_2874, w_118_2877, w_118_2878, w_118_2885, w_118_2889, w_118_2897, w_118_2900, w_118_2904, w_118_2906, w_118_2914, w_118_2916, w_118_2919, w_118_2921, w_118_2922, w_118_2926, w_118_2927, w_118_2932, w_118_2935, w_118_2941, w_118_2942, w_118_2948, w_118_2958, w_118_2965, w_118_2966, w_118_2971, w_118_2975, w_118_2986, w_118_2993, w_118_2997, w_118_3001, w_118_3002, w_118_3004, w_118_3005, w_118_3015, w_118_3016, w_118_3020, w_118_3024, w_118_3025, w_118_3027, w_118_3029, w_118_3032, w_118_3051, w_118_3059, w_118_3060, w_118_3063, w_118_3064, w_118_3065, w_118_3067, w_118_3070, w_118_3075, w_118_3077, w_118_3082, w_118_3098, w_118_3099, w_118_3103, w_118_3105, w_118_3112, w_118_3115, w_118_3119, w_118_3120, w_118_3127, w_118_3131, w_118_3136, w_118_3145, w_118_3150, w_118_3152, w_118_3157, w_118_3164, w_118_3171, w_118_3173, w_118_3174, w_118_3183, w_118_3193, w_118_3195, w_118_3203, w_118_3205, w_118_3206, w_118_3213, w_118_3224, w_118_3230, w_118_3239, w_118_3240, w_118_3244, w_118_3246, w_118_3248, w_118_3249, w_118_3250, w_118_3252, w_118_3254, w_118_3257, w_118_3258, w_118_3267, w_118_3268, w_118_3269, w_118_3272, w_118_3281, w_118_3284, w_118_3285, w_118_3291, w_118_3295, w_118_3297, w_118_3307, w_118_3310, w_118_3311, w_118_3326, w_118_3327, w_118_3330, w_118_3334, w_118_3335, w_118_3336, w_118_3341, w_118_3344, w_118_3346, w_118_3347, w_118_3349, w_118_3350, w_118_3354, w_118_3359, w_118_3366, w_118_3368, w_118_3373, w_118_3374, w_118_3381, w_118_3392, w_118_3396, w_118_3403, w_118_3405, w_118_3406, w_118_3411, w_118_3417, w_118_3421, w_118_3424, w_118_3426, w_118_3437, w_118_3442, w_118_3448, w_118_3451, w_118_3453, w_118_3458, w_118_3461, w_118_3462, w_118_3463, w_118_3467, w_118_3468, w_118_3474, w_118_3477, w_118_3483, w_118_3499, w_118_3504, w_118_3510, w_118_3511, w_118_3513, w_118_3517, w_118_3526, w_118_3531, w_118_3533, w_118_3540, w_118_3541, w_118_3548, w_118_3549, w_118_3550, w_118_3556, w_118_3564, w_118_3566, w_118_3572, w_118_3579, w_118_3584, w_118_3589, w_118_3602, w_118_3605;
  wire w_119_000, w_119_005, w_119_006, w_119_010, w_119_012, w_119_014, w_119_015, w_119_016, w_119_017, w_119_019, w_119_022, w_119_037, w_119_040, w_119_048, w_119_050, w_119_051, w_119_052, w_119_054, w_119_061, w_119_064, w_119_065, w_119_067, w_119_069, w_119_072, w_119_074, w_119_076, w_119_078, w_119_080, w_119_084, w_119_089, w_119_090, w_119_092, w_119_093, w_119_095, w_119_098, w_119_101, w_119_104, w_119_106, w_119_107, w_119_108, w_119_109, w_119_111, w_119_113, w_119_114, w_119_117, w_119_122, w_119_123, w_119_127, w_119_128, w_119_132, w_119_134, w_119_137, w_119_138, w_119_139, w_119_145, w_119_153, w_119_155, w_119_160, w_119_165, w_119_167, w_119_170, w_119_171, w_119_174, w_119_179, w_119_180, w_119_181, w_119_182, w_119_184, w_119_186, w_119_189, w_119_191, w_119_193, w_119_196, w_119_201, w_119_202, w_119_203, w_119_205, w_119_207, w_119_209, w_119_210, w_119_214, w_119_215, w_119_219, w_119_220, w_119_227, w_119_231, w_119_233, w_119_235, w_119_237, w_119_240, w_119_241, w_119_243, w_119_246, w_119_248, w_119_252, w_119_253, w_119_266, w_119_268, w_119_269, w_119_271, w_119_274, w_119_276, w_119_277, w_119_278, w_119_283, w_119_284, w_119_285, w_119_289, w_119_291, w_119_292, w_119_295, w_119_296, w_119_297, w_119_300, w_119_302, w_119_305, w_119_307, w_119_310, w_119_313, w_119_314, w_119_320, w_119_321, w_119_322, w_119_325, w_119_333, w_119_336, w_119_337, w_119_339, w_119_342, w_119_347, w_119_354, w_119_355, w_119_356, w_119_361, w_119_367, w_119_368, w_119_372, w_119_373, w_119_376, w_119_377, w_119_378, w_119_379, w_119_386, w_119_388, w_119_389, w_119_393, w_119_396, w_119_397, w_119_401, w_119_402, w_119_403, w_119_404, w_119_408, w_119_412, w_119_414, w_119_419, w_119_424, w_119_425, w_119_431, w_119_438, w_119_441, w_119_442, w_119_446, w_119_447, w_119_449, w_119_450, w_119_452, w_119_453, w_119_458, w_119_462, w_119_465, w_119_466, w_119_468, w_119_469, w_119_470, w_119_471, w_119_472, w_119_473, w_119_475, w_119_476, w_119_478, w_119_480, w_119_485, w_119_486, w_119_488, w_119_491, w_119_493, w_119_499, w_119_503, w_119_506, w_119_508, w_119_509, w_119_515, w_119_516, w_119_518, w_119_519, w_119_520, w_119_521, w_119_525, w_119_531, w_119_532, w_119_533, w_119_534, w_119_535, w_119_536, w_119_537, w_119_539, w_119_540, w_119_542, w_119_544, w_119_551, w_119_552, w_119_553, w_119_554, w_119_556, w_119_558, w_119_559, w_119_560, w_119_562, w_119_563, w_119_564, w_119_569, w_119_570, w_119_571, w_119_575, w_119_576, w_119_581, w_119_582, w_119_584, w_119_587, w_119_589, w_119_593, w_119_594, w_119_595, w_119_602, w_119_606, w_119_611, w_119_612, w_119_615, w_119_618, w_119_619, w_119_620, w_119_623, w_119_628, w_119_630, w_119_633, w_119_634, w_119_635, w_119_638, w_119_643, w_119_647, w_119_649, w_119_650, w_119_651, w_119_654, w_119_655, w_119_657, w_119_658, w_119_660, w_119_661, w_119_664, w_119_667, w_119_669, w_119_671, w_119_675, w_119_677, w_119_680, w_119_683, w_119_684, w_119_685, w_119_687, w_119_691, w_119_697, w_119_700, w_119_701, w_119_703, w_119_707, w_119_710, w_119_712, w_119_715, w_119_720, w_119_722, w_119_723, w_119_724, w_119_726, w_119_727, w_119_728, w_119_730, w_119_731, w_119_732, w_119_733, w_119_734, w_119_737, w_119_744, w_119_751, w_119_754, w_119_756, w_119_760, w_119_763, w_119_764, w_119_768, w_119_769, w_119_770, w_119_784, w_119_787, w_119_788, w_119_789, w_119_792, w_119_793, w_119_794, w_119_795, w_119_796, w_119_797, w_119_800, w_119_804, w_119_808, w_119_810, w_119_811, w_119_812, w_119_814, w_119_815, w_119_816, w_119_817, w_119_818, w_119_819, w_119_821, w_119_822, w_119_827, w_119_830, w_119_835, w_119_836, w_119_837, w_119_838, w_119_843, w_119_844, w_119_846, w_119_847, w_119_851, w_119_856, w_119_857, w_119_860, w_119_862, w_119_865, w_119_868, w_119_869, w_119_873, w_119_875, w_119_876, w_119_877, w_119_879, w_119_881, w_119_885, w_119_886, w_119_888, w_119_890, w_119_891, w_119_892, w_119_899, w_119_901, w_119_905, w_119_906, w_119_908, w_119_911, w_119_913, w_119_915, w_119_916, w_119_917, w_119_919, w_119_922, w_119_923, w_119_924, w_119_930, w_119_932, w_119_933, w_119_935, w_119_936, w_119_937, w_119_938, w_119_939, w_119_941, w_119_947, w_119_950, w_119_954, w_119_958, w_119_968, w_119_972, w_119_973, w_119_974, w_119_977, w_119_978, w_119_982, w_119_983, w_119_985, w_119_989, w_119_990, w_119_993, w_119_995, w_119_996, w_119_997, w_119_999, w_119_1004, w_119_1006, w_119_1009, w_119_1010, w_119_1011, w_119_1012, w_119_1015, w_119_1020, w_119_1026, w_119_1031, w_119_1034, w_119_1038, w_119_1042, w_119_1046, w_119_1047, w_119_1048, w_119_1050, w_119_1051, w_119_1052, w_119_1057, w_119_1059, w_119_1062, w_119_1068, w_119_1069, w_119_1071, w_119_1072, w_119_1073, w_119_1075, w_119_1078, w_119_1080, w_119_1089, w_119_1092, w_119_1093, w_119_1094, w_119_1095, w_119_1097, w_119_1098, w_119_1099, w_119_1100, w_119_1101, w_119_1104, w_119_1105, w_119_1107, w_119_1109, w_119_1116, w_119_1123, w_119_1124, w_119_1125, w_119_1127, w_119_1128, w_119_1129, w_119_1132, w_119_1133, w_119_1134, w_119_1135, w_119_1136, w_119_1138, w_119_1139, w_119_1140, w_119_1142, w_119_1153, w_119_1157, w_119_1164, w_119_1165, w_119_1168, w_119_1176, w_119_1183, w_119_1184, w_119_1186, w_119_1187, w_119_1191, w_119_1197, w_119_1198, w_119_1199, w_119_1205, w_119_1207, w_119_1212, w_119_1213, w_119_1214, w_119_1215, w_119_1225, w_119_1228, w_119_1229, w_119_1230, w_119_1232, w_119_1236, w_119_1239, w_119_1242, w_119_1247, w_119_1250, w_119_1256, w_119_1257, w_119_1259, w_119_1262, w_119_1263, w_119_1264, w_119_1266, w_119_1269, w_119_1271, w_119_1274, w_119_1275, w_119_1277, w_119_1281, w_119_1282, w_119_1283, w_119_1284, w_119_1291, w_119_1292, w_119_1294, w_119_1295, w_119_1296, w_119_1298, w_119_1299, w_119_1303, w_119_1304, w_119_1305, w_119_1313, w_119_1314, w_119_1316, w_119_1317, w_119_1318, w_119_1319, w_119_1328, w_119_1329, w_119_1331, w_119_1333, w_119_1334, w_119_1338, w_119_1339, w_119_1342, w_119_1344, w_119_1349, w_119_1350, w_119_1352, w_119_1353, w_119_1354, w_119_1355, w_119_1356, w_119_1359, w_119_1362, w_119_1363, w_119_1364, w_119_1373, w_119_1375, w_119_1377, w_119_1378, w_119_1379, w_119_1381, w_119_1383, w_119_1389, w_119_1390, w_119_1391, w_119_1393, w_119_1398, w_119_1401, w_119_1402, w_119_1403, w_119_1406, w_119_1410, w_119_1411, w_119_1413, w_119_1415, w_119_1416, w_119_1418, w_119_1419, w_119_1422, w_119_1423, w_119_1424, w_119_1425, w_119_1426, w_119_1429, w_119_1431, w_119_1435, w_119_1436, w_119_1440, w_119_1441, w_119_1442, w_119_1446, w_119_1448, w_119_1449, w_119_1450, w_119_1452, w_119_1454, w_119_1460, w_119_1462, w_119_1463, w_119_1465, w_119_1470, w_119_1473, w_119_1474, w_119_1475, w_119_1477, w_119_1481, w_119_1482, w_119_1483, w_119_1491, w_119_1495, w_119_1499, w_119_1503, w_119_1505, w_119_1509, w_119_1515, w_119_1517, w_119_1518, w_119_1527, w_119_1528, w_119_1529, w_119_1533, w_119_1534, w_119_1535, w_119_1536, w_119_1542, w_119_1543, w_119_1549, w_119_1554, w_119_1568, w_119_1569, w_119_1572, w_119_1574, w_119_1577, w_119_1579, w_119_1581, w_119_1582, w_119_1584, w_119_1585, w_119_1586, w_119_1588, w_119_1590, w_119_1591, w_119_1592, w_119_1593, w_119_1596, w_119_1598, w_119_1607, w_119_1611, w_119_1618, w_119_1628, w_119_1629, w_119_1631, w_119_1632, w_119_1634, w_119_1635, w_119_1638, w_119_1640, w_119_1644, w_119_1647, w_119_1648, w_119_1649, w_119_1650, w_119_1653, w_119_1654, w_119_1655, w_119_1657, w_119_1659, w_119_1663, w_119_1666, w_119_1668, w_119_1671, w_119_1676, w_119_1678, w_119_1679, w_119_1681, w_119_1684, w_119_1685, w_119_1686, w_119_1688, w_119_1690, w_119_1695, w_119_1697, w_119_1699, w_119_1701, w_119_1704, w_119_1710, w_119_1713, w_119_1719, w_119_1720, w_119_1721, w_119_1723, w_119_1725, w_119_1726, w_119_1727, w_119_1729, w_119_1730, w_119_1731, w_119_1733, w_119_1734, w_119_1736, w_119_1738, w_119_1740, w_119_1741, w_119_1742, w_119_1744, w_119_1745, w_119_1746, w_119_1749, w_119_1750, w_119_1754, w_119_1755, w_119_1756, w_119_1768, w_119_1771, w_119_1773, w_119_1775, w_119_1776, w_119_1779, w_119_1781, w_119_1786, w_119_1787, w_119_1789, w_119_1790, w_119_1792, w_119_1793, w_119_1797, w_119_1798, w_119_1799, w_119_1801, w_119_1804, w_119_1807, w_119_1808, w_119_1809, w_119_1810, w_119_1811, w_119_1815, w_119_1818, w_119_1819, w_119_1820, w_119_1821, w_119_1823, w_119_1826, w_119_1827, w_119_1828, w_119_1832, w_119_1839, w_119_1844, w_119_1845, w_119_1850, w_119_1857, w_119_1872, w_119_1873, w_119_1879, w_119_1881, w_119_1882, w_119_1883, w_119_1893, w_119_1896, w_119_1908, w_119_1911, w_119_1912, w_119_1922, w_119_1927, w_119_1929, w_119_1930, w_119_1942, w_119_1943, w_119_1945, w_119_1949, w_119_1950, w_119_1951, w_119_1958, w_119_1960, w_119_1961, w_119_1964, w_119_1965, w_119_1979, w_119_1980, w_119_1983, w_119_1986, w_119_1987, w_119_1988, w_119_1991, w_119_1993, w_119_2006, w_119_2007, w_119_2010, w_119_2011, w_119_2015, w_119_2017, w_119_2022, w_119_2034, w_119_2043, w_119_2046, w_119_2050, w_119_2051, w_119_2059, w_119_2061, w_119_2068, w_119_2070, w_119_2072, w_119_2073, w_119_2076, w_119_2080, w_119_2085, w_119_2091, w_119_2094, w_119_2098, w_119_2105, w_119_2108, w_119_2110, w_119_2111, w_119_2114, w_119_2116, w_119_2118, w_119_2119, w_119_2137, w_119_2139, w_119_2146, w_119_2149, w_119_2163, w_119_2165, w_119_2168, w_119_2169, w_119_2171, w_119_2177, w_119_2182, w_119_2186, w_119_2189, w_119_2193, w_119_2197, w_119_2211, w_119_2214, w_119_2216, w_119_2227, w_119_2233, w_119_2236, w_119_2238, w_119_2241, w_119_2245, w_119_2247, w_119_2248, w_119_2255, w_119_2256, w_119_2258, w_119_2267, w_119_2272, w_119_2279, w_119_2282, w_119_2286, w_119_2288, w_119_2295, w_119_2303, w_119_2310, w_119_2312, w_119_2314, w_119_2320, w_119_2337, w_119_2342, w_119_2344, w_119_2346, w_119_2349, w_119_2350, w_119_2358, w_119_2360, w_119_2363, w_119_2368, w_119_2373, w_119_2375, w_119_2380, w_119_2385, w_119_2386, w_119_2398, w_119_2399, w_119_2401, w_119_2404, w_119_2408, w_119_2410, w_119_2413, w_119_2414, w_119_2425, w_119_2427, w_119_2429, w_119_2435, w_119_2437, w_119_2444, w_119_2446, w_119_2450, w_119_2454, w_119_2457, w_119_2460, w_119_2469, w_119_2472, w_119_2483, w_119_2484, w_119_2495, w_119_2497, w_119_2498, w_119_2499, w_119_2500, w_119_2507, w_119_2509, w_119_2513, w_119_2515, w_119_2522, w_119_2523, w_119_2525, w_119_2528, w_119_2529, w_119_2531, w_119_2533, w_119_2534, w_119_2536, w_119_2538, w_119_2542, w_119_2543, w_119_2546, w_119_2553, w_119_2559, w_119_2564, w_119_2577, w_119_2578, w_119_2583, w_119_2590, w_119_2593, w_119_2596, w_119_2598, w_119_2600, w_119_2604, w_119_2612, w_119_2613, w_119_2616, w_119_2617, w_119_2623, w_119_2627, w_119_2636, w_119_2639, w_119_2642, w_119_2645, w_119_2656, w_119_2664, w_119_2675, w_119_2681, w_119_2688, w_119_2692, w_119_2694, w_119_2697, w_119_2698, w_119_2700, w_119_2702, w_119_2708, w_119_2709, w_119_2710, w_119_2713, w_119_2728, w_119_2729, w_119_2731, w_119_2732, w_119_2735, w_119_2737, w_119_2742, w_119_2743, w_119_2744, w_119_2746, w_119_2748, w_119_2750, w_119_2752, w_119_2755, w_119_2760, w_119_2765, w_119_2771, w_119_2773, w_119_2776, w_119_2778, w_119_2781, w_119_2782, w_119_2785, w_119_2792, w_119_2801, w_119_2805, w_119_2806, w_119_2807, w_119_2811, w_119_2821, w_119_2822, w_119_2824, w_119_2829, w_119_2836, w_119_2839, w_119_2842, w_119_2848, w_119_2850, w_119_2855, w_119_2870, w_119_2871, w_119_2877, w_119_2886, w_119_2888, w_119_2889, w_119_2892, w_119_2897, w_119_2900, w_119_2903, w_119_2910, w_119_2911, w_119_2920, w_119_2928, w_119_2930, w_119_2931, w_119_2935, w_119_2937, w_119_2941, w_119_2942, w_119_2946, w_119_2967, w_119_2969, w_119_2970, w_119_2980, w_119_2981, w_119_2983, w_119_2984, w_119_2997, w_119_3008, w_119_3011, w_119_3021, w_119_3022, w_119_3027, w_119_3028, w_119_3043, w_119_3055, w_119_3058, w_119_3061, w_119_3068, w_119_3071, w_119_3072, w_119_3073, w_119_3074, w_119_3080, w_119_3083, w_119_3084, w_119_3089, w_119_3093, w_119_3095, w_119_3101, w_119_3107, w_119_3112, w_119_3117, w_119_3120, w_119_3139, w_119_3147, w_119_3150, w_119_3151, w_119_3156, w_119_3159, w_119_3161, w_119_3169;
  wire w_120_000, w_120_001, w_120_002, w_120_003, w_120_004, w_120_005, w_120_006, w_120_007, w_120_008, w_120_009, w_120_010, w_120_011, w_120_012, w_120_013, w_120_014, w_120_015, w_120_016, w_120_017, w_120_018, w_120_019, w_120_020, w_120_021, w_120_022, w_120_023, w_120_024, w_120_025, w_120_026, w_120_027, w_120_028, w_120_029, w_120_030, w_120_031, w_120_032, w_120_033, w_120_034, w_120_035, w_120_036, w_120_037, w_120_038, w_120_039, w_120_040, w_120_041, w_120_042, w_120_043, w_120_044, w_120_045, w_120_046, w_120_047, w_120_048, w_120_049, w_120_050, w_120_051, w_120_052, w_120_053, w_120_054, w_120_055, w_120_056, w_120_057, w_120_058, w_120_059, w_120_060, w_120_061, w_120_062, w_120_063, w_120_064, w_120_065, w_120_066, w_120_067, w_120_068, w_120_069, w_120_070, w_120_071, w_120_072, w_120_073, w_120_074, w_120_075, w_120_076, w_120_077, w_120_078, w_120_079, w_120_080, w_120_081, w_120_082, w_120_083, w_120_084, w_120_085, w_120_086, w_120_087, w_120_088, w_120_089, w_120_090, w_120_091, w_120_092, w_120_093, w_120_094, w_120_095, w_120_096, w_120_097, w_120_098, w_120_099, w_120_100, w_120_101, w_120_102, w_120_103, w_120_104, w_120_105, w_120_106, w_120_107, w_120_108, w_120_109, w_120_110, w_120_111, w_120_112, w_120_113, w_120_114, w_120_115, w_120_116, w_120_117, w_120_118, w_120_119, w_120_120;
  wire w_121_000, w_121_001, w_121_002, w_121_006, w_121_010, w_121_011, w_121_012, w_121_015, w_121_018, w_121_021, w_121_025, w_121_030, w_121_032, w_121_036, w_121_039, w_121_045, w_121_046, w_121_047, w_121_048, w_121_054, w_121_055, w_121_056, w_121_060, w_121_061, w_121_062, w_121_063, w_121_067, w_121_069, w_121_070, w_121_072, w_121_081, w_121_082, w_121_085, w_121_086, w_121_092, w_121_093, w_121_094, w_121_096, w_121_099, w_121_101, w_121_102, w_121_103, w_121_104, w_121_108, w_121_109, w_121_110, w_121_112, w_121_114, w_121_115, w_121_117, w_121_118, w_121_125, w_121_130, w_121_134, w_121_135, w_121_139, w_121_140, w_121_147, w_121_149, w_121_157, w_121_159, w_121_168, w_121_170, w_121_172, w_121_174, w_121_175, w_121_176, w_121_178, w_121_179, w_121_180, w_121_184, w_121_196, w_121_200, w_121_201, w_121_202, w_121_203, w_121_204, w_121_208, w_121_209, w_121_212, w_121_214, w_121_215, w_121_217, w_121_222, w_121_225, w_121_226, w_121_228, w_121_232, w_121_233, w_121_236, w_121_241, w_121_242, w_121_248, w_121_249, w_121_253, w_121_254, w_121_256, w_121_258, w_121_260, w_121_262, w_121_265, w_121_266, w_121_267, w_121_269, w_121_270, w_121_271, w_121_273, w_121_276, w_121_279, w_121_280, w_121_285, w_121_286, w_121_287, w_121_288, w_121_291, w_121_294, w_121_295, w_121_301, w_121_303, w_121_307, w_121_308, w_121_309, w_121_310, w_121_311, w_121_312, w_121_313, w_121_316, w_121_318, w_121_322, w_121_324, w_121_325, w_121_329, w_121_335, w_121_336, w_121_337, w_121_340, w_121_345, w_121_347, w_121_348, w_121_349, w_121_356, w_121_357, w_121_358, w_121_361, w_121_362, w_121_363, w_121_364, w_121_366, w_121_370, w_121_372, w_121_373, w_121_381, w_121_382, w_121_385, w_121_386, w_121_394, w_121_395, w_121_397, w_121_399, w_121_407, w_121_409, w_121_411, w_121_412, w_121_419, w_121_421, w_121_426, w_121_429, w_121_433, w_121_434, w_121_437, w_121_438, w_121_442, w_121_443, w_121_450, w_121_453, w_121_454, w_121_458, w_121_461, w_121_462, w_121_463, w_121_465, w_121_467, w_121_474, w_121_475, w_121_482, w_121_483, w_121_485, w_121_489, w_121_490, w_121_491, w_121_493, w_121_496, w_121_500, w_121_501, w_121_502, w_121_504, w_121_508, w_121_515, w_121_516, w_121_525, w_121_527, w_121_532, w_121_533, w_121_534, w_121_535, w_121_536, w_121_537, w_121_542, w_121_545, w_121_546, w_121_547, w_121_550, w_121_551, w_121_553, w_121_554, w_121_555, w_121_561, w_121_565, w_121_566, w_121_568, w_121_574, w_121_575, w_121_576, w_121_577, w_121_579, w_121_580, w_121_581, w_121_582, w_121_585, w_121_586, w_121_590, w_121_594, w_121_598, w_121_600, w_121_603, w_121_607, w_121_611, w_121_612, w_121_613, w_121_614, w_121_615, w_121_617, w_121_621, w_121_622, w_121_624, w_121_628, w_121_629, w_121_631, w_121_632, w_121_634, w_121_635, w_121_636, w_121_643, w_121_645, w_121_646, w_121_649, w_121_650, w_121_651, w_121_652, w_121_659, w_121_660, w_121_663, w_121_667, w_121_669, w_121_670, w_121_672, w_121_674, w_121_675, w_121_676, w_121_677, w_121_678, w_121_682, w_121_683, w_121_689, w_121_692, w_121_695, w_121_700, w_121_719, w_121_722, w_121_724, w_121_725, w_121_726, w_121_733, w_121_739, w_121_746, w_121_761, w_121_772, w_121_774, w_121_778, w_121_779, w_121_785, w_121_786, w_121_788, w_121_789, w_121_790, w_121_791, w_121_799, w_121_800, w_121_802, w_121_805, w_121_812, w_121_816, w_121_818, w_121_820, w_121_826, w_121_827, w_121_829, w_121_833, w_121_843, w_121_845, w_121_847, w_121_854, w_121_861, w_121_864, w_121_865, w_121_867, w_121_870, w_121_882, w_121_884, w_121_886, w_121_889, w_121_894, w_121_901, w_121_904, w_121_905, w_121_914, w_121_917, w_121_919, w_121_920, w_121_924, w_121_925, w_121_926, w_121_935, w_121_936, w_121_937, w_121_944, w_121_952, w_121_957, w_121_958, w_121_961, w_121_971, w_121_972, w_121_977, w_121_980, w_121_984, w_121_990, w_121_991, w_121_993, w_121_1005, w_121_1025, w_121_1026, w_121_1030, w_121_1032, w_121_1036, w_121_1041, w_121_1044, w_121_1046, w_121_1055, w_121_1061, w_121_1065, w_121_1066, w_121_1067, w_121_1069, w_121_1072, w_121_1074, w_121_1076, w_121_1078, w_121_1081, w_121_1084, w_121_1090, w_121_1109, w_121_1114, w_121_1131, w_121_1132, w_121_1137, w_121_1139, w_121_1143, w_121_1148, w_121_1158, w_121_1161, w_121_1162, w_121_1163, w_121_1164, w_121_1172, w_121_1173, w_121_1176, w_121_1178, w_121_1183, w_121_1184, w_121_1190, w_121_1201, w_121_1203, w_121_1208, w_121_1211, w_121_1214, w_121_1219, w_121_1221, w_121_1228, w_121_1230, w_121_1231, w_121_1234, w_121_1240, w_121_1247, w_121_1248, w_121_1252, w_121_1262, w_121_1274, w_121_1279, w_121_1280, w_121_1282, w_121_1301, w_121_1313, w_121_1315, w_121_1329, w_121_1333, w_121_1335, w_121_1338, w_121_1339, w_121_1342, w_121_1347, w_121_1349, w_121_1352, w_121_1355, w_121_1358, w_121_1363, w_121_1367, w_121_1376, w_121_1378, w_121_1380, w_121_1383, w_121_1387, w_121_1393, w_121_1401, w_121_1405, w_121_1413, w_121_1415, w_121_1444, w_121_1447, w_121_1449, w_121_1450, w_121_1453, w_121_1460, w_121_1463, w_121_1466, w_121_1469, w_121_1473, w_121_1479, w_121_1483, w_121_1492, w_121_1497, w_121_1501, w_121_1504, w_121_1528, w_121_1534, w_121_1540, w_121_1542, w_121_1547, w_121_1558, w_121_1569, w_121_1575, w_121_1576, w_121_1577, w_121_1595, w_121_1597, w_121_1602, w_121_1603, w_121_1605, w_121_1610, w_121_1618, w_121_1619, w_121_1621, w_121_1622, w_121_1625, w_121_1633, w_121_1634, w_121_1635, w_121_1650, w_121_1651, w_121_1653, w_121_1654, w_121_1666, w_121_1668, w_121_1671, w_121_1674, w_121_1677, w_121_1678, w_121_1680, w_121_1684, w_121_1690, w_121_1698, w_121_1702, w_121_1705, w_121_1709, w_121_1711, w_121_1722, w_121_1724, w_121_1725, w_121_1728, w_121_1729, w_121_1734, w_121_1737, w_121_1741, w_121_1744, w_121_1755, w_121_1762, w_121_1763, w_121_1766, w_121_1769, w_121_1773, w_121_1775, w_121_1784, w_121_1785, w_121_1794, w_121_1797, w_121_1805, w_121_1806, w_121_1823, w_121_1838, w_121_1840, w_121_1841, w_121_1844, w_121_1850, w_121_1855, w_121_1858, w_121_1865, w_121_1869, w_121_1872, w_121_1874, w_121_1875, w_121_1879, w_121_1881, w_121_1882, w_121_1884, w_121_1885, w_121_1893, w_121_1895, w_121_1899, w_121_1900, w_121_1901, w_121_1902, w_121_1912, w_121_1928, w_121_1931, w_121_1936, w_121_1946, w_121_1947, w_121_1955, w_121_1956, w_121_1960, w_121_1962, w_121_1964, w_121_1966, w_121_1969, w_121_1976, w_121_1980, w_121_1982, w_121_1993, w_121_2006, w_121_2007, w_121_2011, w_121_2014, w_121_2016, w_121_2019, w_121_2029, w_121_2031, w_121_2032, w_121_2036, w_121_2040, w_121_2043, w_121_2059, w_121_2060, w_121_2075, w_121_2082, w_121_2084, w_121_2086, w_121_2088, w_121_2096, w_121_2109, w_121_2111, w_121_2113, w_121_2114, w_121_2119, w_121_2124, w_121_2127, w_121_2128, w_121_2140, w_121_2144, w_121_2148, w_121_2151, w_121_2154, w_121_2162, w_121_2174, w_121_2176, w_121_2177, w_121_2179, w_121_2180, w_121_2184, w_121_2185, w_121_2190, w_121_2191, w_121_2192, w_121_2195, w_121_2196, w_121_2199, w_121_2200, w_121_2209, w_121_2211, w_121_2213, w_121_2218, w_121_2237, w_121_2239, w_121_2250, w_121_2252, w_121_2255, w_121_2258, w_121_2262, w_121_2263, w_121_2268, w_121_2269, w_121_2279, w_121_2283, w_121_2284, w_121_2290, w_121_2293, w_121_2294, w_121_2302, w_121_2321, w_121_2331, w_121_2332, w_121_2336, w_121_2341, w_121_2342, w_121_2355, w_121_2356, w_121_2359, w_121_2362, w_121_2363, w_121_2366, w_121_2368, w_121_2371, w_121_2372, w_121_2374, w_121_2378, w_121_2379, w_121_2391, w_121_2392, w_121_2394, w_121_2395, w_121_2401, w_121_2403, w_121_2404, w_121_2405, w_121_2407, w_121_2409, w_121_2411, w_121_2414, w_121_2417, w_121_2424, w_121_2427, w_121_2444, w_121_2447, w_121_2454, w_121_2467, w_121_2473, w_121_2477, w_121_2478, w_121_2482, w_121_2489, w_121_2495, w_121_2497, w_121_2505, w_121_2507, w_121_2508, w_121_2520, w_121_2548, w_121_2551, w_121_2553, w_121_2566, w_121_2569, w_121_2572, w_121_2574, w_121_2591, w_121_2597, w_121_2613, w_121_2615, w_121_2620, w_121_2622, w_121_2624, w_121_2627, w_121_2636, w_121_2641, w_121_2642, w_121_2644, w_121_2655, w_121_2661, w_121_2668, w_121_2672, w_121_2674, w_121_2681, w_121_2685, w_121_2686, w_121_2690, w_121_2702, w_121_2705, w_121_2714, w_121_2717, w_121_2718, w_121_2721, w_121_2727, w_121_2729, w_121_2730, w_121_2741, w_121_2743, w_121_2744, w_121_2746, w_121_2751, w_121_2753, w_121_2754, w_121_2757, w_121_2764, w_121_2771, w_121_2772, w_121_2777, w_121_2783, w_121_2786, w_121_2789, w_121_2798, w_121_2800, w_121_2804, w_121_2813, w_121_2818, w_121_2820, w_121_2822, w_121_2823, w_121_2825, w_121_2832, w_121_2834, w_121_2837, w_121_2845, w_121_2846, w_121_2855, w_121_2858, w_121_2861, w_121_2866, w_121_2878, w_121_2879, w_121_2889, w_121_2914, w_121_2916, w_121_2918, w_121_2922, w_121_2931, w_121_2939, w_121_2944, w_121_2948, w_121_2950, w_121_2952, w_121_2957, w_121_2967, w_121_2971, w_121_2974, w_121_2979, w_121_2988, w_121_2996, w_121_2997, w_121_2999, w_121_3000, w_121_3001, w_121_3003, w_121_3005, w_121_3007, w_121_3013, w_121_3024, w_121_3038, w_121_3041, w_121_3053, w_121_3061, w_121_3070, w_121_3074, w_121_3076, w_121_3077, w_121_3079, w_121_3082, w_121_3084, w_121_3088, w_121_3097, w_121_3103, w_121_3108, w_121_3112, w_121_3117, w_121_3123, w_121_3126, w_121_3130, w_121_3138, w_121_3143, w_121_3144, w_121_3159, w_121_3162, w_121_3168, w_121_3169, w_121_3175, w_121_3179, w_121_3181, w_121_3187, w_121_3190, w_121_3202, w_121_3208, w_121_3215, w_121_3217, w_121_3219, w_121_3220, w_121_3223, w_121_3225, w_121_3228, w_121_3236, w_121_3238, w_121_3244, w_121_3247, w_121_3254, w_121_3264, w_121_3272, w_121_3279, w_121_3281, w_121_3282, w_121_3288, w_121_3289, w_121_3290, w_121_3294, w_121_3295, w_121_3296, w_121_3300, w_121_3302, w_121_3310, w_121_3311, w_121_3313, w_121_3319, w_121_3323, w_121_3334, w_121_3335, w_121_3336, w_121_3340, w_121_3343, w_121_3349, w_121_3358, w_121_3363, w_121_3367, w_121_3369, w_121_3371, w_121_3373, w_121_3375, w_121_3376, w_121_3383, w_121_3387, w_121_3390, w_121_3393, w_121_3394, w_121_3397, w_121_3398, w_121_3405, w_121_3413, w_121_3415, w_121_3416, w_121_3420, w_121_3424, w_121_3426, w_121_3430, w_121_3433, w_121_3438, w_121_3441, w_121_3468, w_121_3478, w_121_3480, w_121_3486, w_121_3499, w_121_3500, w_121_3505, w_121_3508, w_121_3509, w_121_3514, w_121_3546, w_121_3547, w_121_3573, w_121_3576, w_121_3582, w_121_3586, w_121_3587, w_121_3589, w_121_3593, w_121_3596, w_121_3601, w_121_3609, w_121_3614, w_121_3616, w_121_3618, w_121_3621, w_121_3623, w_121_3626, w_121_3629, w_121_3630, w_121_3633, w_121_3635, w_121_3637, w_121_3651, w_121_3666, w_121_3673, w_121_3679, w_121_3683, w_121_3684, w_121_3686, w_121_3690, w_121_3695, w_121_3700, w_121_3706, w_121_3708, w_121_3711, w_121_3714, w_121_3720, w_121_3723, w_121_3729, w_121_3734, w_121_3735, w_121_3741, w_121_3742, w_121_3744, w_121_3751, w_121_3753, w_121_3754, w_121_3757, w_121_3759, w_121_3764, w_121_3765, w_121_3767, w_121_3768, w_121_3769, w_121_3770, w_121_3771, w_121_3774, w_121_3784, w_121_3794, w_121_3796, w_121_3799, w_121_3800, w_121_3804, w_121_3805, w_121_3808, w_121_3810, w_121_3813, w_121_3820, w_121_3824, w_121_3825, w_121_3828, w_121_3833, w_121_3837, w_121_3838, w_121_3844, w_121_3845, w_121_3846, w_121_3848, w_121_3850, w_121_3855, w_121_3857, w_121_3860, w_121_3864, w_121_3879, w_121_3887, w_121_3889, w_121_3895, w_121_3899, w_121_3914, w_121_3917, w_121_3921, w_121_3933, w_121_3935, w_121_3937, w_121_3940, w_121_3956, w_121_3957, w_121_3975, w_121_3986, w_121_3987, w_121_3991, w_121_3992, w_121_4004, w_121_4005, w_121_4006, w_121_4013, w_121_4015, w_121_4019, w_121_4021, w_121_4025, w_121_4034, w_121_4036, w_121_4039, w_121_4061, w_121_4088, w_121_4101, w_121_4112, w_121_4114, w_121_4117, w_121_4126, w_121_4131, w_121_4133, w_121_4134, w_121_4139, w_121_4141, w_121_4146, w_121_4154, w_121_4156, w_121_4165, w_121_4167, w_121_4180, w_121_4181, w_121_4182, w_121_4185, w_121_4187, w_121_4188, w_121_4191, w_121_4203, w_121_4206, w_121_4207, w_121_4210, w_121_4215, w_121_4221, w_121_4224, w_121_4227, w_121_4229, w_121_4230, w_121_4234, w_121_4236, w_121_4240, w_121_4241, w_121_4242, w_121_4243, w_121_4245, w_121_4259, w_121_4266, w_121_4267, w_121_4271, w_121_4273, w_121_4280, w_121_4284, w_121_4288, w_121_4294;
  wire w_122_000, w_122_001, w_122_002, w_122_003, w_122_004, w_122_005, w_122_006, w_122_007, w_122_008, w_122_009, w_122_010, w_122_011, w_122_012, w_122_013, w_122_014, w_122_015, w_122_016, w_122_017, w_122_018, w_122_019, w_122_020, w_122_021, w_122_022, w_122_023, w_122_024, w_122_025, w_122_026, w_122_027, w_122_028, w_122_029, w_122_030, w_122_031, w_122_032, w_122_033, w_122_034, w_122_035, w_122_036, w_122_037, w_122_038, w_122_039, w_122_040, w_122_041, w_122_042, w_122_043, w_122_044, w_122_045, w_122_046, w_122_047, w_122_048, w_122_049, w_122_050, w_122_051, w_122_052, w_122_053, w_122_054, w_122_055, w_122_056, w_122_057, w_122_058, w_122_059, w_122_060, w_122_061, w_122_062, w_122_063, w_122_064, w_122_065, w_122_066, w_122_067, w_122_068, w_122_069, w_122_070, w_122_071, w_122_072, w_122_073, w_122_074, w_122_075, w_122_076, w_122_077, w_122_078, w_122_079, w_122_080, w_122_081, w_122_082, w_122_083, w_122_084, w_122_085, w_122_086, w_122_087, w_122_088, w_122_089, w_122_090, w_122_091, w_122_092, w_122_093, w_122_094, w_122_095, w_122_096, w_122_097, w_122_098, w_122_099, w_122_100, w_122_101, w_122_102, w_122_103, w_122_104, w_122_105, w_122_106, w_122_107, w_122_108, w_122_109, w_122_110, w_122_111, w_122_112, w_122_113, w_122_114, w_122_115, w_122_116, w_122_117, w_122_118, w_122_119, w_122_120, w_122_121, w_122_122, w_122_123, w_122_124, w_122_125, w_122_126, w_122_127, w_122_128, w_122_129, w_122_130, w_122_131, w_122_132, w_122_133, w_122_134, w_122_135, w_122_136, w_122_137, w_122_138, w_122_139, w_122_140, w_122_141, w_122_142, w_122_143, w_122_144, w_122_145, w_122_146, w_122_147, w_122_148, w_122_149, w_122_150, w_122_151, w_122_152, w_122_153, w_122_154, w_122_155, w_122_156, w_122_157, w_122_158, w_122_159, w_122_160, w_122_161, w_122_162, w_122_163, w_122_164, w_122_165, w_122_166, w_122_167, w_122_168, w_122_169, w_122_170, w_122_171, w_122_172, w_122_173, w_122_174, w_122_175, w_122_176, w_122_177, w_122_178, w_122_179, w_122_180, w_122_181, w_122_182, w_122_183, w_122_184, w_122_185, w_122_186, w_122_187, w_122_188, w_122_189, w_122_190, w_122_191, w_122_192, w_122_193, w_122_194, w_122_195, w_122_196, w_122_197, w_122_198, w_122_199, w_122_200, w_122_201, w_122_202, w_122_203, w_122_204, w_122_205, w_122_206, w_122_207, w_122_208, w_122_209, w_122_210, w_122_211, w_122_212, w_122_213, w_122_214, w_122_215, w_122_216, w_122_217, w_122_218, w_122_219, w_122_220, w_122_221, w_122_222, w_122_223, w_122_224, w_122_225, w_122_226, w_122_227, w_122_228, w_122_229, w_122_230, w_122_231, w_122_232, w_122_233, w_122_234, w_122_235, w_122_236, w_122_237, w_122_238, w_122_239, w_122_240, w_122_241, w_122_242, w_122_243, w_122_244, w_122_245, w_122_246, w_122_247, w_122_248, w_122_249, w_122_250, w_122_251, w_122_252, w_122_253, w_122_254, w_122_255, w_122_256, w_122_257, w_122_258, w_122_259, w_122_260, w_122_261, w_122_262, w_122_263, w_122_264, w_122_265, w_122_266, w_122_267, w_122_268, w_122_269, w_122_270, w_122_271, w_122_272, w_122_273, w_122_275;
  wire w_123_000, w_123_001, w_123_003, w_123_004, w_123_006, w_123_009, w_123_010, w_123_011, w_123_013, w_123_014, w_123_015, w_123_017, w_123_021, w_123_023, w_123_026, w_123_030, w_123_031, w_123_033, w_123_035, w_123_037, w_123_038, w_123_045, w_123_046, w_123_048, w_123_050, w_123_053, w_123_055, w_123_056, w_123_058, w_123_060, w_123_061, w_123_063, w_123_065, w_123_068, w_123_069, w_123_070, w_123_072, w_123_076, w_123_080, w_123_082, w_123_083, w_123_084, w_123_088, w_123_090, w_123_091, w_123_092, w_123_093, w_123_095, w_123_096, w_123_098, w_123_099, w_123_100, w_123_101, w_123_102, w_123_103, w_123_108, w_123_111, w_123_112, w_123_113, w_123_115, w_123_117, w_123_118, w_123_126, w_123_128, w_123_129, w_123_131, w_123_133, w_123_135, w_123_136, w_123_137, w_123_139, w_123_141, w_123_143, w_123_144, w_123_145, w_123_146, w_123_148, w_123_149, w_123_151, w_123_153, w_123_154, w_123_156, w_123_157, w_123_158, w_123_159, w_123_160, w_123_161, w_123_163, w_123_165, w_123_168, w_123_169, w_123_170, w_123_171, w_123_172, w_123_174, w_123_175, w_123_177, w_123_178, w_123_179, w_123_180, w_123_181, w_123_183, w_123_186, w_123_187, w_123_189, w_123_191, w_123_192, w_123_193, w_123_194, w_123_197, w_123_200, w_123_204, w_123_207, w_123_208, w_123_209, w_123_210, w_123_211, w_123_213, w_123_219, w_123_223, w_123_225, w_123_226, w_123_227, w_123_228, w_123_229, w_123_232, w_123_236, w_123_237, w_123_239, w_123_240, w_123_241, w_123_245, w_123_248, w_123_251, w_123_252, w_123_256, w_123_258, w_123_259, w_123_261, w_123_263, w_123_268, w_123_275, w_123_276, w_123_277, w_123_278, w_123_280, w_123_281, w_123_284, w_123_285, w_123_286, w_123_287, w_123_288, w_123_290, w_123_291, w_123_294, w_123_296, w_123_299, w_123_301, w_123_307, w_123_309, w_123_311, w_123_313, w_123_316, w_123_320, w_123_322, w_123_325, w_123_326, w_123_328, w_123_335, w_123_336, w_123_338, w_123_339, w_123_340, w_123_341, w_123_342, w_123_344, w_123_345, w_123_346, w_123_348, w_123_350, w_123_355, w_123_356, w_123_357, w_123_358, w_123_359, w_123_360, w_123_361, w_123_368, w_123_369, w_123_371, w_123_372, w_123_373, w_123_374, w_123_376, w_123_378, w_123_379, w_123_380, w_123_381, w_123_384, w_123_385, w_123_387, w_123_389, w_123_391, w_123_394, w_123_396, w_123_399, w_123_401, w_123_402, w_123_405, w_123_407, w_123_408, w_123_411, w_123_413, w_123_414, w_123_415, w_123_416, w_123_420, w_123_422, w_123_423, w_123_424, w_123_427, w_123_433, w_123_434, w_123_436, w_123_442, w_123_445, w_123_446, w_123_451, w_123_453, w_123_455, w_123_456, w_123_458, w_123_460, w_123_461, w_123_463, w_123_465, w_123_466, w_123_471, w_123_473, w_123_477, w_123_478, w_123_479, w_123_483, w_123_484, w_123_485, w_123_487, w_123_489, w_123_493, w_123_494, w_123_496, w_123_497, w_123_500, w_123_502, w_123_504, w_123_505, w_123_506, w_123_507, w_123_517, w_123_519, w_123_520, w_123_522, w_123_524, w_123_525, w_123_526, w_123_528, w_123_530, w_123_532, w_123_534, w_123_536, w_123_537, w_123_538, w_123_539, w_123_540, w_123_543, w_123_544, w_123_547, w_123_550, w_123_551, w_123_554, w_123_556, w_123_557, w_123_559, w_123_560, w_123_561, w_123_562, w_123_563, w_123_564, w_123_571, w_123_572, w_123_574, w_123_576, w_123_577, w_123_578, w_123_580, w_123_582, w_123_583, w_123_585, w_123_586, w_123_588, w_123_589, w_123_592, w_123_596, w_123_597, w_123_598, w_123_600, w_123_601, w_123_602, w_123_606, w_123_607, w_123_608, w_123_609, w_123_611, w_123_615, w_123_619, w_123_620, w_123_621, w_123_622, w_123_623, w_123_624, w_123_627, w_123_629, w_123_630, w_123_631, w_123_633, w_123_635, w_123_636, w_123_638, w_123_640, w_123_642, w_123_644, w_123_645, w_123_648, w_123_653, w_123_655, w_123_658, w_123_664, w_123_665, w_123_669, w_123_670, w_123_672, w_123_674, w_123_678, w_123_681, w_123_682, w_123_684, w_123_688, w_123_691, w_123_692, w_123_693, w_123_694, w_123_697, w_123_698, w_123_699, w_123_700, w_123_701, w_123_702, w_123_705, w_123_706, w_123_708, w_123_710, w_123_711, w_123_713, w_123_714, w_123_715, w_123_719, w_123_720, w_123_721, w_123_722, w_123_724, w_123_726, w_123_727, w_123_728, w_123_729, w_123_730, w_123_735, w_123_739, w_123_740, w_123_741, w_123_742, w_123_743, w_123_745, w_123_751, w_123_754, w_123_756, w_123_757, w_123_758, w_123_759, w_123_760, w_123_762, w_123_764, w_123_766, w_123_767, w_123_768, w_123_770, w_123_771, w_123_772, w_123_779, w_123_780, w_123_781, w_123_782, w_123_783, w_123_785, w_123_787, w_123_790, w_123_791, w_123_794, w_123_795, w_123_796, w_123_803, w_123_804, w_123_805, w_123_806, w_123_807, w_123_809, w_123_811, w_123_812, w_123_815, w_123_817, w_123_818, w_123_820, w_123_823, w_123_824, w_123_826, w_123_827, w_123_829, w_123_831, w_123_832, w_123_833, w_123_834, w_123_836, w_123_837, w_123_838, w_123_840, w_123_842, w_123_844, w_123_846, w_123_847, w_123_849, w_123_852, w_123_859, w_123_861, w_123_862, w_123_864, w_123_865, w_123_866, w_123_867, w_123_870, w_123_873, w_123_874, w_123_875, w_123_878, w_123_879, w_123_880, w_123_882, w_123_883, w_123_884, w_123_885, w_123_886, w_123_887, w_123_888, w_123_889, w_123_891, w_123_892, w_123_893, w_123_896, w_123_897, w_123_898, w_123_899, w_123_900, w_123_901, w_123_904, w_123_908, w_123_909, w_123_911, w_123_913, w_123_914, w_123_917, w_123_918, w_123_919, w_123_920, w_123_921, w_123_922, w_123_924, w_123_925, w_123_926, w_123_927, w_123_928, w_123_929, w_123_930, w_123_933, w_123_935, w_123_937, w_123_939, w_123_941, w_123_944, w_123_945, w_123_946, w_123_947, w_123_949, w_123_950, w_123_951, w_123_955, w_123_956, w_123_957, w_123_961, w_123_963, w_123_964, w_123_968, w_123_972, w_123_975, w_123_976, w_123_977, w_123_978, w_123_979, w_123_980, w_123_983, w_123_984, w_123_985, w_123_989, w_123_990, w_123_994, w_123_997, w_123_998, w_123_1004, w_123_1006, w_123_1008, w_123_1009, w_123_1010, w_123_1011, w_123_1013, w_123_1014, w_123_1015, w_123_1017, w_123_1020, w_123_1021, w_123_1022, w_123_1024, w_123_1026, w_123_1029, w_123_1030, w_123_1032, w_123_1033, w_123_1034, w_123_1035, w_123_1039, w_123_1042, w_123_1046, w_123_1051, w_123_1053, w_123_1054, w_123_1057, w_123_1059, w_123_1066, w_123_1067, w_123_1068, w_123_1071, w_123_1075, w_123_1076, w_123_1078, w_123_1081, w_123_1082, w_123_1085, w_123_1088, w_123_1091, w_123_1093, w_123_1095, w_123_1100, w_123_1104, w_123_1105, w_123_1106, w_123_1109, w_123_1111, w_123_1115, w_123_1117, w_123_1119, w_123_1121, w_123_1123, w_123_1124, w_123_1126, w_123_1128, w_123_1129, w_123_1131, w_123_1137, w_123_1140, w_123_1141, w_123_1147, w_123_1152, w_123_1153, w_123_1155, w_123_1157, w_123_1159, w_123_1162, w_123_1163, w_123_1164, w_123_1167, w_123_1169, w_123_1170, w_123_1171, w_123_1178, w_123_1181, w_123_1183, w_123_1186, w_123_1189, w_123_1191, w_123_1193, w_123_1195, w_123_1197, w_123_1198, w_123_1203, w_123_1208, w_123_1209, w_123_1210, w_123_1212, w_123_1214, w_123_1219, w_123_1220, w_123_1221, w_123_1225, w_123_1228, w_123_1231, w_123_1233, w_123_1234, w_123_1235, w_123_1237, w_123_1239, w_123_1242, w_123_1245, w_123_1248, w_123_1253, w_123_1260, w_123_1264, w_123_1266, w_123_1267, w_123_1268, w_123_1272, w_123_1281, w_123_1283, w_123_1284, w_123_1285, w_123_1288, w_123_1289, w_123_1290, w_123_1291, w_123_1293, w_123_1294, w_123_1296, w_123_1297, w_123_1298, w_123_1300, w_123_1301, w_123_1302, w_123_1304, w_123_1308, w_123_1310, w_123_1311, w_123_1316, w_123_1317, w_123_1318, w_123_1325, w_123_1326, w_123_1327, w_123_1335, w_123_1336, w_123_1338, w_123_1343, w_123_1346, w_123_1348, w_123_1353, w_123_1355, w_123_1356, w_123_1359, w_123_1360, w_123_1361, w_123_1364, w_123_1366, w_123_1370, w_123_1373, w_123_1374, w_123_1378, w_123_1379, w_123_1381, w_123_1382, w_123_1383, w_123_1384, w_123_1385, w_123_1386, w_123_1388, w_123_1389, w_123_1395, w_123_1399, w_123_1402, w_123_1409, w_123_1412, w_123_1413, w_123_1415, w_123_1416, w_123_1419, w_123_1424, w_123_1426, w_123_1428, w_123_1431, w_123_1438, w_123_1439, w_123_1443, w_123_1445, w_123_1446, w_123_1447, w_123_1451, w_123_1452, w_123_1457, w_123_1459, w_123_1461, w_123_1465, w_123_1467, w_123_1468, w_123_1470, w_123_1473, w_123_1479, w_123_1482, w_123_1483, w_123_1485, w_123_1486, w_123_1489, w_123_1491, w_123_1498, w_123_1499, w_123_1500, w_123_1504, w_123_1505, w_123_1509, w_123_1514, w_123_1519, w_123_1521, w_123_1522, w_123_1523, w_123_1524, w_123_1525, w_123_1527, w_123_1528, w_123_1532, w_123_1536, w_123_1537, w_123_1538, w_123_1539, w_123_1544, w_123_1546, w_123_1551, w_123_1552, w_123_1554, w_123_1559, w_123_1567, w_123_1570, w_123_1575, w_123_1576, w_123_1578, w_123_1580, w_123_1586, w_123_1589, w_123_1593, w_123_1595, w_123_1597, w_123_1601, w_123_1603, w_123_1609, w_123_1611, w_123_1612, w_123_1617, w_123_1618, w_123_1619, w_123_1622, w_123_1623, w_123_1628, w_123_1629, w_123_1630, w_123_1634, w_123_1636, w_123_1637, w_123_1640, w_123_1652, w_123_1659, w_123_1665, w_123_1675, w_123_1677, w_123_1679, w_123_1681, w_123_1683, w_123_1688, w_123_1689, w_123_1692, w_123_1693, w_123_1697, w_123_1698, w_123_1699, w_123_1704, w_123_1706, w_123_1709, w_123_1713, w_123_1714, w_123_1716, w_123_1718, w_123_1720, w_123_1730, w_123_1732, w_123_1733, w_123_1734, w_123_1735, w_123_1738, w_123_1743, w_123_1744, w_123_1750, w_123_1751, w_123_1757, w_123_1760, w_123_1762, w_123_1764, w_123_1772, w_123_1776, w_123_1781, w_123_1784, w_123_1786, w_123_1789, w_123_1790, w_123_1791, w_123_1793, w_123_1794, w_123_1800, w_123_1801, w_123_1803, w_123_1804, w_123_1805, w_123_1806, w_123_1808, w_123_1810, w_123_1814, w_123_1820, w_123_1822, w_123_1828, w_123_1830, w_123_1835, w_123_1836, w_123_1837, w_123_1838, w_123_1840, w_123_1841, w_123_1844, w_123_1849, w_123_1850, w_123_1851, w_123_1852, w_123_1855, w_123_1864, w_123_1866, w_123_1867, w_123_1869, w_123_1872, w_123_1875, w_123_1877, w_123_1879, w_123_1880, w_123_1887, w_123_1890, w_123_1893, w_123_1895, w_123_1899, w_123_1903, w_123_1914, w_123_1915, w_123_1916, w_123_1920, w_123_1922, w_123_1928, w_123_1933, w_123_1934, w_123_1935, w_123_1937, w_123_1939, w_123_1940, w_123_1942, w_123_1943, w_123_1945, w_123_1947, w_123_1948, w_123_1950, w_123_1955, w_123_1957, w_123_1960, w_123_1962, w_123_1965, w_123_1966, w_123_1967, w_123_1971, w_123_1988, w_123_1992, w_123_1995, w_123_1999, w_123_2004;
  wire w_124_000, w_124_001, w_124_003, w_124_006, w_124_009, w_124_013, w_124_014, w_124_015, w_124_021, w_124_024, w_124_028, w_124_032, w_124_034, w_124_037, w_124_039, w_124_041, w_124_045, w_124_050, w_124_053, w_124_054, w_124_055, w_124_056, w_124_060, w_124_064, w_124_067, w_124_068, w_124_071, w_124_072, w_124_075, w_124_076, w_124_077, w_124_078, w_124_079, w_124_083, w_124_085, w_124_089, w_124_093, w_124_094, w_124_099, w_124_100, w_124_103, w_124_104, w_124_111, w_124_114, w_124_115, w_124_116, w_124_120, w_124_121, w_124_124, w_124_126, w_124_127, w_124_128, w_124_133, w_124_134, w_124_137, w_124_138, w_124_139, w_124_140, w_124_144, w_124_145, w_124_146, w_124_149, w_124_152, w_124_153, w_124_154, w_124_157, w_124_162, w_124_163, w_124_168, w_124_171, w_124_172, w_124_174, w_124_175, w_124_176, w_124_177, w_124_178, w_124_190, w_124_198, w_124_199, w_124_204, w_124_205, w_124_206, w_124_208, w_124_210, w_124_212, w_124_226, w_124_227, w_124_230, w_124_231, w_124_232, w_124_242, w_124_247, w_124_249, w_124_252, w_124_255, w_124_258, w_124_261, w_124_265, w_124_267, w_124_268, w_124_270, w_124_271, w_124_272, w_124_273, w_124_276, w_124_278, w_124_280, w_124_283, w_124_290, w_124_291, w_124_296, w_124_297, w_124_298, w_124_299, w_124_300, w_124_301, w_124_302, w_124_308, w_124_311, w_124_313, w_124_315, w_124_319, w_124_323, w_124_328, w_124_336, w_124_337, w_124_339, w_124_341, w_124_342, w_124_344, w_124_346, w_124_348, w_124_349, w_124_354, w_124_357, w_124_358, w_124_359, w_124_361, w_124_364, w_124_367, w_124_371, w_124_372, w_124_374, w_124_376, w_124_378, w_124_379, w_124_380, w_124_381, w_124_382, w_124_386, w_124_389, w_124_391, w_124_396, w_124_399, w_124_400, w_124_402, w_124_403, w_124_406, w_124_415, w_124_416, w_124_418, w_124_420, w_124_424, w_124_428, w_124_430, w_124_431, w_124_436, w_124_437, w_124_440, w_124_441, w_124_444, w_124_447, w_124_450, w_124_451, w_124_458, w_124_461, w_124_462, w_124_464, w_124_466, w_124_469, w_124_471, w_124_473, w_124_477, w_124_480, w_124_481, w_124_486, w_124_490, w_124_492, w_124_494, w_124_496, w_124_497, w_124_500, w_124_501, w_124_502, w_124_505, w_124_512, w_124_513, w_124_515, w_124_516, w_124_518, w_124_521, w_124_526, w_124_527, w_124_528, w_124_531, w_124_533, w_124_536, w_124_539, w_124_540, w_124_542, w_124_543, w_124_546, w_124_548, w_124_549, w_124_550, w_124_553, w_124_554, w_124_558, w_124_561, w_124_563, w_124_566, w_124_571, w_124_578, w_124_579, w_124_582, w_124_584, w_124_586, w_124_589, w_124_591, w_124_597, w_124_599, w_124_600, w_124_601, w_124_603, w_124_607, w_124_608, w_124_610, w_124_613, w_124_614, w_124_620, w_124_621, w_124_623, w_124_626, w_124_627, w_124_629, w_124_631, w_124_633, w_124_636, w_124_637, w_124_645, w_124_649, w_124_651, w_124_655, w_124_658, w_124_660, w_124_663, w_124_664, w_124_665, w_124_666, w_124_667, w_124_671, w_124_672, w_124_674, w_124_678, w_124_679, w_124_681, w_124_683, w_124_690, w_124_692, w_124_693, w_124_694, w_124_697, w_124_698, w_124_699, w_124_701, w_124_702, w_124_706, w_124_708, w_124_709, w_124_712, w_124_714, w_124_716, w_124_719, w_124_720, w_124_722, w_124_723, w_124_725, w_124_728, w_124_732, w_124_737, w_124_738, w_124_739, w_124_740, w_124_741, w_124_744, w_124_745, w_124_746, w_124_749, w_124_750, w_124_752, w_124_756, w_124_757, w_124_758, w_124_759, w_124_763, w_124_764, w_124_769, w_124_771, w_124_774, w_124_775, w_124_776, w_124_780, w_124_786, w_124_788, w_124_796, w_124_797, w_124_798, w_124_803, w_124_805, w_124_808, w_124_811, w_124_815, w_124_818, w_124_819, w_124_820, w_124_822, w_124_827, w_124_828, w_124_829, w_124_831, w_124_835, w_124_836, w_124_837, w_124_841, w_124_843, w_124_844, w_124_845, w_124_846, w_124_848, w_124_849, w_124_850, w_124_852, w_124_854, w_124_856, w_124_862, w_124_863, w_124_866, w_124_867, w_124_870, w_124_875, w_124_876, w_124_880, w_124_882, w_124_884, w_124_886, w_124_888, w_124_890, w_124_893, w_124_894, w_124_899, w_124_900, w_124_901, w_124_903, w_124_906, w_124_911, w_124_914, w_124_915, w_124_925, w_124_929, w_124_933, w_124_935, w_124_936, w_124_937, w_124_939, w_124_940, w_124_942, w_124_945, w_124_946, w_124_947, w_124_948, w_124_949, w_124_952, w_124_956, w_124_959, w_124_960, w_124_962, w_124_967, w_124_968, w_124_969, w_124_973, w_124_976, w_124_982, w_124_988, w_124_992, w_124_993, w_124_995, w_124_998, w_124_1000, w_124_1003, w_124_1005, w_124_1006, w_124_1007, w_124_1010, w_124_1019, w_124_1020, w_124_1021, w_124_1023, w_124_1024, w_124_1025, w_124_1029, w_124_1033, w_124_1038, w_124_1039, w_124_1044, w_124_1046, w_124_1047, w_124_1051, w_124_1052, w_124_1056, w_124_1058, w_124_1059, w_124_1060, w_124_1062, w_124_1063, w_124_1067, w_124_1069, w_124_1072, w_124_1073, w_124_1076, w_124_1078, w_124_1079, w_124_1080, w_124_1081, w_124_1082, w_124_1083, w_124_1086, w_124_1088, w_124_1090, w_124_1094, w_124_1096, w_124_1097, w_124_1100, w_124_1103, w_124_1107, w_124_1108, w_124_1109, w_124_1110, w_124_1111, w_124_1112, w_124_1113, w_124_1115, w_124_1116, w_124_1117, w_124_1118, w_124_1121, w_124_1124, w_124_1130, w_124_1133, w_124_1137, w_124_1138, w_124_1139, w_124_1140, w_124_1145, w_124_1146, w_124_1147, w_124_1148, w_124_1149, w_124_1151, w_124_1153, w_124_1154, w_124_1157, w_124_1158, w_124_1160, w_124_1162, w_124_1166, w_124_1167, w_124_1172, w_124_1174, w_124_1181, w_124_1182, w_124_1184, w_124_1185, w_124_1192, w_124_1198, w_124_1199, w_124_1200, w_124_1203, w_124_1210, w_124_1215, w_124_1218, w_124_1223, w_124_1227, w_124_1228, w_124_1229, w_124_1230, w_124_1231, w_124_1232, w_124_1236, w_124_1241, w_124_1249, w_124_1251, w_124_1252, w_124_1255, w_124_1257, w_124_1258, w_124_1259, w_124_1260, w_124_1262, w_124_1264, w_124_1265, w_124_1266, w_124_1269, w_124_1274, w_124_1275, w_124_1278, w_124_1279, w_124_1281, w_124_1282, w_124_1284, w_124_1287, w_124_1288, w_124_1292, w_124_1308, w_124_1309, w_124_1313, w_124_1314, w_124_1315, w_124_1316, w_124_1320, w_124_1323, w_124_1324, w_124_1325, w_124_1332, w_124_1333, w_124_1334, w_124_1337, w_124_1342, w_124_1343, w_124_1344, w_124_1350, w_124_1354, w_124_1356, w_124_1359, w_124_1361, w_124_1362, w_124_1363, w_124_1366, w_124_1369, w_124_1371, w_124_1372, w_124_1375, w_124_1382, w_124_1387, w_124_1388, w_124_1389, w_124_1394, w_124_1395, w_124_1396, w_124_1401, w_124_1403, w_124_1405, w_124_1410, w_124_1414, w_124_1419, w_124_1421, w_124_1422, w_124_1423, w_124_1435, w_124_1438, w_124_1441, w_124_1442, w_124_1443, w_124_1446, w_124_1447, w_124_1448, w_124_1450, w_124_1452, w_124_1453, w_124_1454, w_124_1455, w_124_1457, w_124_1465, w_124_1470, w_124_1471, w_124_1474, w_124_1476, w_124_1477, w_124_1478, w_124_1479, w_124_1482, w_124_1484, w_124_1494, w_124_1497, w_124_1499, w_124_1500, w_124_1501, w_124_1502, w_124_1503, w_124_1504, w_124_1510, w_124_1511, w_124_1512, w_124_1514, w_124_1515, w_124_1519, w_124_1520, w_124_1521, w_124_1525, w_124_1526, w_124_1528, w_124_1531, w_124_1535, w_124_1539, w_124_1542, w_124_1546, w_124_1547, w_124_1549, w_124_1552, w_124_1553, w_124_1555, w_124_1557, w_124_1559, w_124_1562, w_124_1564, w_124_1568, w_124_1569, w_124_1575, w_124_1578, w_124_1580, w_124_1581, w_124_1588, w_124_1591, w_124_1592, w_124_1593, w_124_1594, w_124_1597, w_124_1603, w_124_1607, w_124_1612, w_124_1617, w_124_1620, w_124_1621, w_124_1623, w_124_1625, w_124_1626, w_124_1629, w_124_1631, w_124_1632, w_124_1633, w_124_1637, w_124_1638, w_124_1640, w_124_1643, w_124_1645, w_124_1652, w_124_1653, w_124_1657, w_124_1658, w_124_1663, w_124_1664, w_124_1667, w_124_1668, w_124_1673, w_124_1675, w_124_1676, w_124_1679, w_124_1681, w_124_1682, w_124_1684, w_124_1685, w_124_1686, w_124_1689, w_124_1690, w_124_1695, w_124_1696, w_124_1699, w_124_1700, w_124_1703, w_124_1705, w_124_1707, w_124_1709, w_124_1710, w_124_1712, w_124_1716, w_124_1722, w_124_1723, w_124_1726, w_124_1727, w_124_1730, w_124_1731, w_124_1734, w_124_1739, w_124_1751, w_124_1754, w_124_1757, w_124_1759, w_124_1760, w_124_1763, w_124_1764, w_124_1765, w_124_1770, w_124_1771, w_124_1772, w_124_1774, w_124_1775, w_124_1776, w_124_1779, w_124_1780, w_124_1782, w_124_1784, w_124_1785, w_124_1787, w_124_1788, w_124_1790, w_124_1791, w_124_1792, w_124_1796, w_124_1802, w_124_1803, w_124_1807, w_124_1811, w_124_1812, w_124_1814, w_124_1815, w_124_1816, w_124_1818, w_124_1819, w_124_1820, w_124_1822, w_124_1823, w_124_1824, w_124_1825, w_124_1826, w_124_1827, w_124_1828, w_124_1831, w_124_1833, w_124_1835, w_124_1840, w_124_1841, w_124_1845, w_124_1847, w_124_1848, w_124_1849, w_124_1851, w_124_1853, w_124_1860, w_124_1861, w_124_1867, w_124_1879, w_124_1881, w_124_1884, w_124_1886, w_124_1887, w_124_1888, w_124_1889, w_124_1891, w_124_1892, w_124_1894, w_124_1895, w_124_1896, w_124_1901, w_124_1908, w_124_1910, w_124_1911, w_124_1912, w_124_1914, w_124_1922, w_124_1923, w_124_1927, w_124_1928, w_124_1929, w_124_1930, w_124_1932, w_124_1934, w_124_1936, w_124_1937, w_124_1940, w_124_1944, w_124_1945, w_124_1947, w_124_1954, w_124_1955, w_124_1956, w_124_1957, w_124_1959, w_124_1960, w_124_1967, w_124_1969, w_124_1970, w_124_1977, w_124_1982, w_124_1985, w_124_1986, w_124_1990, w_124_1994, w_124_1996, w_124_2011, w_124_2016, w_124_2021, w_124_2023, w_124_2025, w_124_2029, w_124_2030, w_124_2032, w_124_2033, w_124_2035, w_124_2036, w_124_2039, w_124_2042, w_124_2043, w_124_2046, w_124_2051, w_124_2052, w_124_2055, w_124_2058, w_124_2060, w_124_2061, w_124_2066, w_124_2069, w_124_2078, w_124_2080, w_124_2084, w_124_2088, w_124_2092, w_124_2093, w_124_2095, w_124_2096, w_124_2100, w_124_2101, w_124_2102, w_124_2103, w_124_2104, w_124_2105, w_124_2107, w_124_2110, w_124_2123, w_124_2129, w_124_2131, w_124_2137, w_124_2143, w_124_2144, w_124_2151, w_124_2152, w_124_2154, w_124_2157, w_124_2159, w_124_2161, w_124_2162, w_124_2163, w_124_2165, w_124_2166, w_124_2178, w_124_2188, w_124_2190, w_124_2193, w_124_2195, w_124_2196, w_124_2197, w_124_2199, w_124_2202, w_124_2205, w_124_2206, w_124_2208, w_124_2210, w_124_2216, w_124_2218, w_124_2222, w_124_2226, w_124_2228, w_124_2230, w_124_2234, w_124_2235, w_124_2236, w_124_2237, w_124_2242, w_124_2244, w_124_2245, w_124_2246, w_124_2247, w_124_2248, w_124_2249, w_124_2256, w_124_2261, w_124_2262, w_124_2263, w_124_2267, w_124_2275, w_124_2277, w_124_2278, w_124_2281, w_124_2282, w_124_2284, w_124_2285, w_124_2288, w_124_2291, w_124_2292, w_124_2293, w_124_2301, w_124_2303, w_124_2307, w_124_2312, w_124_2314, w_124_2318, w_124_2319, w_124_2320, w_124_2321, w_124_2322, w_124_2325, w_124_2328, w_124_2331, w_124_2339, w_124_2346, w_124_2353, w_124_2354, w_124_2355, w_124_2356, w_124_2357, w_124_2360, w_124_2363, w_124_2364, w_124_2365, w_124_2366, w_124_2374, w_124_2379, w_124_2382, w_124_2386, w_124_2388, w_124_2389, w_124_2391, w_124_2394, w_124_2400, w_124_2407, w_124_2408, w_124_2411, w_124_2415, w_124_2427, w_124_2428, w_124_2435, w_124_2439, w_124_2441, w_124_2444, w_124_2451, w_124_2452, w_124_2454, w_124_2457, w_124_2464, w_124_2469, w_124_2473, w_124_2480, w_124_2483, w_124_2488, w_124_2489, w_124_2491, w_124_2494, w_124_2500, w_124_2509, w_124_2517, w_124_2535, w_124_2544, w_124_2555, w_124_2560, w_124_2568, w_124_2580, w_124_2586, w_124_2588, w_124_2590, w_124_2591, w_124_2604, w_124_2605, w_124_2611, w_124_2612, w_124_2613;
  wire w_125_002, w_125_003, w_125_004, w_125_005, w_125_007, w_125_008, w_125_011, w_125_013, w_125_016, w_125_019, w_125_020, w_125_023, w_125_026, w_125_031, w_125_033, w_125_035, w_125_036, w_125_040, w_125_041, w_125_042, w_125_043, w_125_047, w_125_049, w_125_051, w_125_052, w_125_054, w_125_055, w_125_056, w_125_057, w_125_058, w_125_061, w_125_063, w_125_070, w_125_072, w_125_076, w_125_078, w_125_081, w_125_085, w_125_092, w_125_093, w_125_100, w_125_102, w_125_103, w_125_110, w_125_112, w_125_116, w_125_117, w_125_118, w_125_122, w_125_123, w_125_125, w_125_126, w_125_130, w_125_133, w_125_138, w_125_140, w_125_143, w_125_149, w_125_153, w_125_155, w_125_159, w_125_163, w_125_164, w_125_166, w_125_173, w_125_177, w_125_180, w_125_183, w_125_190, w_125_192, w_125_193, w_125_195, w_125_197, w_125_201, w_125_202, w_125_206, w_125_208, w_125_211, w_125_214, w_125_216, w_125_217, w_125_220, w_125_224, w_125_227, w_125_229, w_125_233, w_125_234, w_125_235, w_125_236, w_125_239, w_125_240, w_125_241, w_125_243, w_125_244, w_125_245, w_125_248, w_125_250, w_125_251, w_125_254, w_125_255, w_125_257, w_125_260, w_125_264, w_125_273, w_125_274, w_125_282, w_125_285, w_125_287, w_125_291, w_125_292, w_125_295, w_125_297, w_125_299, w_125_307, w_125_311, w_125_315, w_125_318, w_125_319, w_125_320, w_125_327, w_125_328, w_125_330, w_125_331, w_125_332, w_125_333, w_125_334, w_125_339, w_125_341, w_125_342, w_125_345, w_125_348, w_125_352, w_125_353, w_125_354, w_125_355, w_125_361, w_125_365, w_125_366, w_125_369, w_125_370, w_125_372, w_125_373, w_125_376, w_125_380, w_125_383, w_125_388, w_125_393, w_125_395, w_125_398, w_125_400, w_125_401, w_125_402, w_125_404, w_125_407, w_125_409, w_125_414, w_125_415, w_125_422, w_125_424, w_125_427, w_125_428, w_125_429, w_125_430, w_125_432, w_125_433, w_125_434, w_125_435, w_125_437, w_125_443, w_125_446, w_125_449, w_125_450, w_125_451, w_125_453, w_125_456, w_125_459, w_125_465, w_125_467, w_125_468, w_125_472, w_125_473, w_125_474, w_125_477, w_125_478, w_125_480, w_125_483, w_125_484, w_125_488, w_125_491, w_125_493, w_125_495, w_125_496, w_125_503, w_125_506, w_125_508, w_125_512, w_125_514, w_125_516, w_125_519, w_125_520, w_125_521, w_125_530, w_125_531, w_125_536, w_125_537, w_125_538, w_125_540, w_125_549, w_125_556, w_125_562, w_125_566, w_125_576, w_125_577, w_125_582, w_125_583, w_125_585, w_125_586, w_125_597, w_125_606, w_125_613, w_125_614, w_125_618, w_125_619, w_125_624, w_125_632, w_125_637, w_125_641, w_125_643, w_125_645, w_125_651, w_125_655, w_125_657, w_125_665, w_125_670, w_125_671, w_125_674, w_125_676, w_125_679, w_125_681, w_125_682, w_125_683, w_125_684, w_125_696, w_125_700, w_125_711, w_125_716, w_125_718, w_125_722, w_125_726, w_125_729, w_125_730, w_125_734, w_125_743, w_125_746, w_125_747, w_125_749, w_125_753, w_125_759, w_125_761, w_125_762, w_125_763, w_125_768, w_125_778, w_125_779, w_125_784, w_125_790, w_125_794, w_125_801, w_125_804, w_125_813, w_125_817, w_125_820, w_125_823, w_125_826, w_125_829, w_125_831, w_125_832, w_125_835, w_125_837, w_125_840, w_125_848, w_125_860, w_125_862, w_125_873, w_125_874, w_125_876, w_125_877, w_125_879, w_125_883, w_125_884, w_125_899, w_125_901, w_125_902, w_125_904, w_125_927, w_125_929, w_125_930, w_125_931, w_125_932, w_125_942, w_125_943, w_125_944, w_125_945, w_125_956, w_125_961, w_125_963, w_125_976, w_125_979, w_125_984, w_125_996, w_125_997, w_125_999, w_125_1019, w_125_1022, w_125_1023, w_125_1025, w_125_1026, w_125_1027, w_125_1030, w_125_1031, w_125_1054, w_125_1055, w_125_1059, w_125_1067, w_125_1070, w_125_1077, w_125_1078, w_125_1079, w_125_1081, w_125_1094, w_125_1096, w_125_1097, w_125_1105, w_125_1106, w_125_1110, w_125_1120, w_125_1126, w_125_1132, w_125_1136, w_125_1141, w_125_1142, w_125_1144, w_125_1155, w_125_1160, w_125_1163, w_125_1165, w_125_1177, w_125_1178, w_125_1182, w_125_1184, w_125_1185, w_125_1187, w_125_1197, w_125_1198, w_125_1199, w_125_1200, w_125_1212, w_125_1216, w_125_1223, w_125_1228, w_125_1235, w_125_1236, w_125_1238, w_125_1249, w_125_1250, w_125_1254, w_125_1258, w_125_1259, w_125_1272, w_125_1281, w_125_1283, w_125_1285, w_125_1289, w_125_1295, w_125_1297, w_125_1300, w_125_1303, w_125_1306, w_125_1314, w_125_1316, w_125_1320, w_125_1322, w_125_1324, w_125_1325, w_125_1334, w_125_1335, w_125_1347, w_125_1348, w_125_1350, w_125_1354, w_125_1363, w_125_1374, w_125_1376, w_125_1385, w_125_1389, w_125_1394, w_125_1399, w_125_1403, w_125_1405, w_125_1407, w_125_1411, w_125_1415, w_125_1421, w_125_1423, w_125_1424, w_125_1432, w_125_1437, w_125_1438, w_125_1440, w_125_1442, w_125_1445, w_125_1456, w_125_1458, w_125_1462, w_125_1465, w_125_1470, w_125_1477, w_125_1487, w_125_1488, w_125_1490, w_125_1491, w_125_1495, w_125_1500, w_125_1518, w_125_1519, w_125_1520, w_125_1522, w_125_1523, w_125_1526, w_125_1531, w_125_1533, w_125_1535, w_125_1538, w_125_1541, w_125_1549, w_125_1554, w_125_1564, w_125_1576, w_125_1585, w_125_1595, w_125_1599, w_125_1611, w_125_1613, w_125_1629, w_125_1630, w_125_1635, w_125_1645, w_125_1647, w_125_1653, w_125_1655, w_125_1660, w_125_1663, w_125_1667, w_125_1668, w_125_1674, w_125_1675, w_125_1677, w_125_1684, w_125_1688, w_125_1689, w_125_1692, w_125_1702, w_125_1703, w_125_1704, w_125_1707, w_125_1710, w_125_1715, w_125_1716, w_125_1728, w_125_1731, w_125_1732, w_125_1740, w_125_1760, w_125_1769, w_125_1778, w_125_1780, w_125_1798, w_125_1800, w_125_1802, w_125_1808, w_125_1811, w_125_1814, w_125_1823, w_125_1830, w_125_1840, w_125_1841, w_125_1848, w_125_1851, w_125_1863, w_125_1864, w_125_1866, w_125_1875, w_125_1877, w_125_1881, w_125_1883, w_125_1888, w_125_1891, w_125_1894, w_125_1895, w_125_1898, w_125_1901, w_125_1903, w_125_1904, w_125_1905, w_125_1908, w_125_1912, w_125_1917, w_125_1922, w_125_1930, w_125_1935, w_125_1942, w_125_1944, w_125_1945, w_125_1948, w_125_1956, w_125_1962, w_125_1964, w_125_1973, w_125_1975, w_125_1977, w_125_1984, w_125_1987, w_125_1991, w_125_1992, w_125_1993, w_125_1995, w_125_1997, w_125_2000, w_125_2014, w_125_2018, w_125_2022, w_125_2026, w_125_2027, w_125_2028, w_125_2029, w_125_2051, w_125_2052, w_125_2056, w_125_2070, w_125_2072, w_125_2089, w_125_2091, w_125_2099, w_125_2100, w_125_2108, w_125_2109, w_125_2110, w_125_2111, w_125_2121, w_125_2131, w_125_2136, w_125_2138, w_125_2139, w_125_2154, w_125_2158, w_125_2163, w_125_2171, w_125_2173, w_125_2178, w_125_2180, w_125_2191, w_125_2198, w_125_2206, w_125_2208, w_125_2226, w_125_2228, w_125_2233, w_125_2234, w_125_2242, w_125_2244, w_125_2247, w_125_2253, w_125_2254, w_125_2256, w_125_2268, w_125_2271, w_125_2278, w_125_2279, w_125_2296, w_125_2298, w_125_2302, w_125_2311, w_125_2316, w_125_2325, w_125_2334, w_125_2337, w_125_2340, w_125_2343, w_125_2345, w_125_2346, w_125_2357, w_125_2358, w_125_2361, w_125_2366, w_125_2382, w_125_2389, w_125_2400, w_125_2407, w_125_2411, w_125_2417, w_125_2421, w_125_2426, w_125_2430, w_125_2431, w_125_2434, w_125_2435, w_125_2446, w_125_2448, w_125_2450, w_125_2452, w_125_2461, w_125_2462, w_125_2463, w_125_2466, w_125_2483, w_125_2484, w_125_2485, w_125_2486, w_125_2496, w_125_2497, w_125_2500, w_125_2505, w_125_2511, w_125_2520, w_125_2521, w_125_2522, w_125_2525, w_125_2540, w_125_2541, w_125_2542, w_125_2547, w_125_2552, w_125_2559, w_125_2561, w_125_2564, w_125_2567, w_125_2585, w_125_2587, w_125_2588, w_125_2593, w_125_2594, w_125_2595, w_125_2598, w_125_2601, w_125_2603, w_125_2604, w_125_2611, w_125_2615, w_125_2617, w_125_2619, w_125_2626, w_125_2627, w_125_2641, w_125_2642, w_125_2643, w_125_2649, w_125_2653, w_125_2666, w_125_2671, w_125_2674, w_125_2676, w_125_2677, w_125_2686, w_125_2688, w_125_2692, w_125_2693, w_125_2695, w_125_2700, w_125_2705, w_125_2707, w_125_2716, w_125_2719, w_125_2724, w_125_2728, w_125_2731, w_125_2734, w_125_2738, w_125_2741, w_125_2742, w_125_2743, w_125_2744, w_125_2747, w_125_2748, w_125_2750, w_125_2760, w_125_2761, w_125_2762, w_125_2765, w_125_2769, w_125_2770, w_125_2784, w_125_2788, w_125_2793, w_125_2794, w_125_2800, w_125_2802, w_125_2803, w_125_2809, w_125_2814, w_125_2818, w_125_2824, w_125_2834, w_125_2835, w_125_2837, w_125_2839, w_125_2843, w_125_2851, w_125_2854, w_125_2864, w_125_2865, w_125_2870, w_125_2873, w_125_2879, w_125_2883, w_125_2889, w_125_2904, w_125_2906, w_125_2908, w_125_2915, w_125_2920, w_125_2923, w_125_2931, w_125_2934, w_125_2944, w_125_2949, w_125_2950, w_125_2952, w_125_2953, w_125_2955, w_125_2961, w_125_2963, w_125_2964, w_125_2970, w_125_2971, w_125_2973, w_125_2976, w_125_2984, w_125_2986, w_125_2989, w_125_2990, w_125_2996, w_125_2998, w_125_3001, w_125_3007, w_125_3010, w_125_3026, w_125_3029, w_125_3037, w_125_3039, w_125_3045, w_125_3063, w_125_3066, w_125_3071, w_125_3074, w_125_3084, w_125_3118, w_125_3121, w_125_3134, w_125_3136, w_125_3145, w_125_3147, w_125_3162, w_125_3168, w_125_3170, w_125_3172, w_125_3180, w_125_3183, w_125_3191, w_125_3193, w_125_3199, w_125_3200, w_125_3207, w_125_3211, w_125_3226, w_125_3228, w_125_3232, w_125_3237, w_125_3239, w_125_3240, w_125_3245, w_125_3253, w_125_3255, w_125_3260, w_125_3261, w_125_3272, w_125_3273, w_125_3284, w_125_3292, w_125_3293, w_125_3303, w_125_3307, w_125_3308, w_125_3310, w_125_3314, w_125_3319, w_125_3326, w_125_3331, w_125_3332, w_125_3335, w_125_3336, w_125_3348, w_125_3350, w_125_3353, w_125_3356, w_125_3361, w_125_3366, w_125_3370, w_125_3376, w_125_3377, w_125_3389, w_125_3396, w_125_3412, w_125_3416, w_125_3417, w_125_3421, w_125_3423, w_125_3424, w_125_3425, w_125_3427, w_125_3428, w_125_3438, w_125_3443, w_125_3447, w_125_3465, w_125_3467, w_125_3478, w_125_3486, w_125_3488, w_125_3489, w_125_3491, w_125_3499, w_125_3501, w_125_3510, w_125_3516, w_125_3521, w_125_3524, w_125_3526, w_125_3527, w_125_3528, w_125_3531, w_125_3534, w_125_3538, w_125_3539, w_125_3543, w_125_3548, w_125_3550, w_125_3562, w_125_3566, w_125_3570, w_125_3573, w_125_3581, w_125_3585, w_125_3589, w_125_3591, w_125_3600, w_125_3603, w_125_3607, w_125_3608, w_125_3619, w_125_3622, w_125_3625, w_125_3627, w_125_3630, w_125_3635, w_125_3639, w_125_3641, w_125_3642, w_125_3652, w_125_3655, w_125_3657, w_125_3660, w_125_3667, w_125_3671, w_125_3681, w_125_3686, w_125_3689, w_125_3693, w_125_3694, w_125_3695, w_125_3699, w_125_3701, w_125_3704, w_125_3706, w_125_3707, w_125_3708, w_125_3713, w_125_3714, w_125_3721, w_125_3724, w_125_3739, w_125_3753, w_125_3755, w_125_3756, w_125_3759, w_125_3765, w_125_3768, w_125_3769, w_125_3770, w_125_3774, w_125_3775, w_125_3776, w_125_3785, w_125_3789, w_125_3792, w_125_3800, w_125_3806, w_125_3811, w_125_3814, w_125_3817, w_125_3819, w_125_3822, w_125_3829, w_125_3839, w_125_3841, w_125_3843, w_125_3853, w_125_3858, w_125_3862, w_125_3865, w_125_3867, w_125_3872, w_125_3879, w_125_3881, w_125_3891, w_125_3893, w_125_3894, w_125_3895, w_125_3901, w_125_3902, w_125_3919, w_125_3924, w_125_3929, w_125_3933, w_125_3934, w_125_3941, w_125_3956, w_125_3962, w_125_3971, w_125_3972, w_125_3973, w_125_3974, w_125_3975, w_125_3978, w_125_3983, w_125_3986, w_125_3991, w_125_3999, w_125_4004, w_125_4006, w_125_4012, w_125_4015, w_125_4023, w_125_4033, w_125_4034, w_125_4038, w_125_4040, w_125_4041, w_125_4044, w_125_4049, w_125_4052, w_125_4062, w_125_4063, w_125_4067, w_125_4068, w_125_4070, w_125_4071, w_125_4072, w_125_4090, w_125_4099, w_125_4101, w_125_4103, w_125_4113, w_125_4116, w_125_4123, w_125_4135, w_125_4136, w_125_4138, w_125_4146, w_125_4151, w_125_4152, w_125_4153, w_125_4160, w_125_4166, w_125_4168, w_125_4175, w_125_4176, w_125_4179, w_125_4187, w_125_4190, w_125_4197, w_125_4199, w_125_4200, w_125_4205, w_125_4215, w_125_4219, w_125_4224, w_125_4228, w_125_4230, w_125_4234, w_125_4237, w_125_4239, w_125_4243, w_125_4244, w_125_4248, w_125_4249, w_125_4253, w_125_4255, w_125_4258, w_125_4269, w_125_4271, w_125_4275, w_125_4281, w_125_4284, w_125_4287, w_125_4293, w_125_4303, w_125_4311, w_125_4312, w_125_4318, w_125_4321, w_125_4326, w_125_4328, w_125_4340, w_125_4344, w_125_4349, w_125_4355, w_125_4363, w_125_4381, w_125_4384, w_125_4388, w_125_4391, w_125_4396, w_125_4402, w_125_4404, w_125_4405, w_125_4410, w_125_4413, w_125_4416, w_125_4425, w_125_4434, w_125_4443, w_125_4452, w_125_4455, w_125_4456, w_125_4462, w_125_4466, w_125_4468, w_125_4472, w_125_4479, w_125_4481, w_125_4491, w_125_4502, w_125_4503;
  wire w_126_000, w_126_001, w_126_002, w_126_003, w_126_004, w_126_005, w_126_006, w_126_007, w_126_008, w_126_009, w_126_010, w_126_011, w_126_012, w_126_013, w_126_014, w_126_015, w_126_016, w_126_017, w_126_018, w_126_019, w_126_020, w_126_021, w_126_022, w_126_023, w_126_024, w_126_025, w_126_026, w_126_027, w_126_028, w_126_029, w_126_030, w_126_031, w_126_032, w_126_033, w_126_034, w_126_035, w_126_036, w_126_037, w_126_038, w_126_039, w_126_040, w_126_041, w_126_042, w_126_043, w_126_044, w_126_045, w_126_046, w_126_047, w_126_048, w_126_049, w_126_050, w_126_051, w_126_052, w_126_053, w_126_054, w_126_055, w_126_056, w_126_057, w_126_058, w_126_059, w_126_060, w_126_061, w_126_062, w_126_063, w_126_064, w_126_065, w_126_066, w_126_067, w_126_068, w_126_069, w_126_070, w_126_071, w_126_072, w_126_073, w_126_074, w_126_075, w_126_076, w_126_077, w_126_078, w_126_079, w_126_080, w_126_081, w_126_082, w_126_083, w_126_084, w_126_085, w_126_086, w_126_087, w_126_088, w_126_089, w_126_090, w_126_091, w_126_092, w_126_093, w_126_094, w_126_095, w_126_096, w_126_097, w_126_098, w_126_099, w_126_100, w_126_101, w_126_102, w_126_103, w_126_104, w_126_105, w_126_106, w_126_107, w_126_108, w_126_109, w_126_110, w_126_111, w_126_112, w_126_113, w_126_114, w_126_115, w_126_116, w_126_117, w_126_118, w_126_119, w_126_120, w_126_121, w_126_122, w_126_123, w_126_124, w_126_125, w_126_126, w_126_127, w_126_128, w_126_129, w_126_130, w_126_131, w_126_132, w_126_133, w_126_134, w_126_135, w_126_136, w_126_137, w_126_138, w_126_139, w_126_140, w_126_141, w_126_142, w_126_143, w_126_144, w_126_145, w_126_146, w_126_147, w_126_148, w_126_149, w_126_150, w_126_151, w_126_152, w_126_153, w_126_154, w_126_155, w_126_156, w_126_157, w_126_158, w_126_159, w_126_160, w_126_161, w_126_162, w_126_163, w_126_164, w_126_165, w_126_166, w_126_167, w_126_168, w_126_169, w_126_170, w_126_171, w_126_172, w_126_173, w_126_174, w_126_175, w_126_176, w_126_177, w_126_178, w_126_179, w_126_180, w_126_181, w_126_182, w_126_183, w_126_184, w_126_185, w_126_186, w_126_187, w_126_188, w_126_189, w_126_190, w_126_191, w_126_192, w_126_193, w_126_194;
  wire w_127_000, w_127_001, w_127_002, w_127_003, w_127_004, w_127_005, w_127_006, w_127_007, w_127_008, w_127_010, w_127_011, w_127_014, w_127_015, w_127_016, w_127_017, w_127_018, w_127_019, w_127_020, w_127_022, w_127_023, w_127_024, w_127_025, w_127_026, w_127_027, w_127_028, w_127_030, w_127_031, w_127_032, w_127_033, w_127_034, w_127_035, w_127_036, w_127_037, w_127_038, w_127_039, w_127_040, w_127_041, w_127_042, w_127_044, w_127_045, w_127_046, w_127_047, w_127_048, w_127_050, w_127_051, w_127_052, w_127_053, w_127_054, w_127_055, w_127_056, w_127_057, w_127_058, w_127_059, w_127_060, w_127_061, w_127_062, w_127_063, w_127_064, w_127_065, w_127_066, w_127_067, w_127_068, w_127_069, w_127_070, w_127_071, w_127_072, w_127_073, w_127_075, w_127_076, w_127_077, w_127_078, w_127_079, w_127_080, w_127_081, w_127_082, w_127_083, w_127_084, w_127_085, w_127_087, w_127_088, w_127_089, w_127_090, w_127_091, w_127_092, w_127_093, w_127_094, w_127_095, w_127_096, w_127_097, w_127_098, w_127_099, w_127_100, w_127_101, w_127_102, w_127_103, w_127_105, w_127_106, w_127_107, w_127_108, w_127_109, w_127_110, w_127_111, w_127_112, w_127_114, w_127_115, w_127_116, w_127_117, w_127_118, w_127_119, w_127_120, w_127_121, w_127_123, w_127_124, w_127_126, w_127_127, w_127_128, w_127_129, w_127_130, w_127_131, w_127_132, w_127_133, w_127_134, w_127_135, w_127_137, w_127_138, w_127_139, w_127_140, w_127_142, w_127_144, w_127_145, w_127_146, w_127_147, w_127_148, w_127_149, w_127_150, w_127_151, w_127_152, w_127_153, w_127_155, w_127_156, w_127_157, w_127_158, w_127_159, w_127_160, w_127_161, w_127_162, w_127_163, w_127_164, w_127_166, w_127_167, w_127_168, w_127_169, w_127_170, w_127_171, w_127_172, w_127_174, w_127_175, w_127_177, w_127_180, w_127_181, w_127_182, w_127_183, w_127_184, w_127_185, w_127_186, w_127_187, w_127_188, w_127_189, w_127_190, w_127_191, w_127_192, w_127_193, w_127_194, w_127_195, w_127_197, w_127_198, w_127_199, w_127_201, w_127_202, w_127_203, w_127_204, w_127_205, w_127_206, w_127_207, w_127_208, w_127_210, w_127_211, w_127_212, w_127_213, w_127_214, w_127_215, w_127_216, w_127_217, w_127_218, w_127_219, w_127_220, w_127_222, w_127_223, w_127_224, w_127_225, w_127_227, w_127_228, w_127_229, w_127_230, w_127_231, w_127_232, w_127_233, w_127_234, w_127_236, w_127_237, w_127_238, w_127_239, w_127_241, w_127_242, w_127_243, w_127_244, w_127_245, w_127_246, w_127_247, w_127_248, w_127_249, w_127_250, w_127_251, w_127_252, w_127_253, w_127_254, w_127_256, w_127_257, w_127_258, w_127_259, w_127_260, w_127_261, w_127_263, w_127_264, w_127_265, w_127_266, w_127_267, w_127_268, w_127_269, w_127_271, w_127_272, w_127_273, w_127_274, w_127_275, w_127_276, w_127_277, w_127_278, w_127_279, w_127_280, w_127_281, w_127_282, w_127_283, w_127_284, w_127_285, w_127_286, w_127_287, w_127_289, w_127_290, w_127_291, w_127_292, w_127_293, w_127_295, w_127_296, w_127_297, w_127_298, w_127_300, w_127_301, w_127_302, w_127_303, w_127_304, w_127_305, w_127_306, w_127_307, w_127_308, w_127_309, w_127_311, w_127_312, w_127_313, w_127_314, w_127_315, w_127_316, w_127_317, w_127_318, w_127_319, w_127_320, w_127_321, w_127_322, w_127_323, w_127_324, w_127_325, w_127_326, w_127_327, w_127_328, w_127_329, w_127_330, w_127_331, w_127_333, w_127_334, w_127_335, w_127_336, w_127_337, w_127_338, w_127_339, w_127_340, w_127_341, w_127_342, w_127_343, w_127_344, w_127_345, w_127_346, w_127_347, w_127_348, w_127_349, w_127_350, w_127_351, w_127_352, w_127_353, w_127_354, w_127_355, w_127_356, w_127_357, w_127_358, w_127_359, w_127_360, w_127_361, w_127_362, w_127_363, w_127_364, w_127_365, w_127_366, w_127_368, w_127_369, w_127_370, w_127_371, w_127_373, w_127_374, w_127_375, w_127_377, w_127_378, w_127_379, w_127_380, w_127_383, w_127_384, w_127_385, w_127_386, w_127_387, w_127_388, w_127_389, w_127_390, w_127_391, w_127_392, w_127_393, w_127_394, w_127_396, w_127_397, w_127_398, w_127_399, w_127_400, w_127_401, w_127_402, w_127_403, w_127_405, w_127_406, w_127_408, w_127_409, w_127_410, w_127_411, w_127_412, w_127_413, w_127_414, w_127_415, w_127_416, w_127_417, w_127_418, w_127_419, w_127_420, w_127_421, w_127_423, w_127_424, w_127_425, w_127_427, w_127_428, w_127_429, w_127_430, w_127_431, w_127_432, w_127_433, w_127_434, w_127_435, w_127_436, w_127_438, w_127_439, w_127_440, w_127_441, w_127_442, w_127_443, w_127_444, w_127_445, w_127_446, w_127_448, w_127_449, w_127_450, w_127_451, w_127_452, w_127_453, w_127_454, w_127_455, w_127_456, w_127_457, w_127_458, w_127_460, w_127_461, w_127_464, w_127_465, w_127_466, w_127_467, w_127_468, w_127_470, w_127_471, w_127_472, w_127_473, w_127_474, w_127_475, w_127_476, w_127_477, w_127_478, w_127_479, w_127_480, w_127_481, w_127_482, w_127_483, w_127_484, w_127_485, w_127_486, w_127_487, w_127_488, w_127_489, w_127_490, w_127_491, w_127_492, w_127_494, w_127_495, w_127_496, w_127_497, w_127_498, w_127_499, w_127_500, w_127_501, w_127_502, w_127_504, w_127_505, w_127_506, w_127_507, w_127_508, w_127_509, w_127_510, w_127_511, w_127_512, w_127_513, w_127_514, w_127_515, w_127_516, w_127_517, w_127_518, w_127_519, w_127_520, w_127_521, w_127_522, w_127_523, w_127_524, w_127_525, w_127_527, w_127_528, w_127_529, w_127_530, w_127_532, w_127_534, w_127_535, w_127_536, w_127_537, w_127_538, w_127_539, w_127_540, w_127_541, w_127_542, w_127_543, w_127_544, w_127_545, w_127_546, w_127_547, w_127_548, w_127_549, w_127_552, w_127_553, w_127_556, w_127_558, w_127_559, w_127_560, w_127_561, w_127_562, w_127_563, w_127_564, w_127_565, w_127_566, w_127_567, w_127_568, w_127_570, w_127_571, w_127_573, w_127_574, w_127_575, w_127_576, w_127_577, w_127_578, w_127_579, w_127_580, w_127_581, w_127_582, w_127_583, w_127_584, w_127_585, w_127_586, w_127_587, w_127_588, w_127_589, w_127_590, w_127_591, w_127_593, w_127_595, w_127_596, w_127_597, w_127_598, w_127_600, w_127_601, w_127_603, w_127_605, w_127_606, w_127_607, w_127_608, w_127_609, w_127_610, w_127_611, w_127_612, w_127_613, w_127_614;
  wire w_128_000, w_128_002, w_128_005, w_128_006, w_128_007, w_128_008, w_128_012, w_128_013, w_128_014, w_128_015, w_128_016, w_128_018, w_128_021, w_128_024, w_128_028, w_128_031, w_128_035, w_128_037, w_128_038, w_128_039, w_128_044, w_128_045, w_128_046, w_128_047, w_128_048, w_128_050, w_128_055, w_128_058, w_128_059, w_128_060, w_128_062, w_128_063, w_128_064, w_128_072, w_128_073, w_128_074, w_128_078, w_128_085, w_128_087, w_128_089, w_128_090, w_128_093, w_128_094, w_128_095, w_128_097, w_128_098, w_128_102, w_128_105, w_128_109, w_128_110, w_128_112, w_128_114, w_128_116, w_128_121, w_128_123, w_128_126, w_128_128, w_128_130, w_128_137, w_128_139, w_128_145, w_128_146, w_128_149, w_128_151, w_128_154, w_128_156, w_128_158, w_128_162, w_128_166, w_128_169, w_128_171, w_128_172, w_128_177, w_128_179, w_128_180, w_128_182, w_128_183, w_128_184, w_128_193, w_128_197, w_128_199, w_128_200, w_128_201, w_128_204, w_128_207, w_128_208, w_128_211, w_128_215, w_128_216, w_128_219, w_128_221, w_128_223, w_128_226, w_128_227, w_128_228, w_128_233, w_128_237, w_128_239, w_128_242, w_128_243, w_128_246, w_128_249, w_128_250, w_128_251, w_128_252, w_128_253, w_128_256, w_128_257, w_128_258, w_128_260, w_128_262, w_128_263, w_128_267, w_128_268, w_128_272, w_128_274, w_128_277, w_128_280, w_128_281, w_128_286, w_128_287, w_128_289, w_128_291, w_128_292, w_128_293, w_128_295, w_128_296, w_128_298, w_128_299, w_128_300, w_128_302, w_128_311, w_128_312, w_128_313, w_128_316, w_128_319, w_128_320, w_128_321, w_128_323, w_128_324, w_128_325, w_128_328, w_128_330, w_128_332, w_128_333, w_128_342, w_128_343, w_128_344, w_128_346, w_128_350, w_128_351, w_128_352, w_128_355, w_128_357, w_128_363, w_128_366, w_128_367, w_128_368, w_128_369, w_128_370, w_128_375, w_128_377, w_128_379, w_128_384, w_128_387, w_128_389, w_128_391, w_128_393, w_128_395, w_128_397, w_128_398, w_128_404, w_128_405, w_128_407, w_128_408, w_128_409, w_128_411, w_128_418, w_128_420, w_128_424, w_128_430, w_128_431, w_128_432, w_128_433, w_128_434, w_128_435, w_128_437, w_128_439, w_128_440, w_128_442, w_128_443, w_128_445, w_128_447, w_128_453, w_128_455, w_128_456, w_128_461, w_128_465, w_128_468, w_128_469, w_128_471, w_128_483, w_128_485, w_128_489, w_128_490, w_128_495, w_128_504, w_128_505, w_128_507, w_128_511, w_128_514, w_128_516, w_128_520, w_128_521, w_128_525, w_128_526, w_128_527, w_128_535, w_128_540, w_128_541, w_128_542, w_128_543, w_128_546, w_128_555, w_128_556, w_128_558, w_128_559, w_128_562, w_128_563, w_128_566, w_128_568, w_128_569, w_128_570, w_128_572, w_128_576, w_128_577, w_128_578, w_128_579, w_128_587, w_128_589, w_128_593, w_128_599, w_128_607, w_128_609, w_128_611, w_128_612, w_128_613, w_128_619, w_128_620, w_128_622, w_128_624, w_128_625, w_128_626, w_128_629, w_128_636, w_128_639, w_128_640, w_128_644, w_128_645, w_128_649, w_128_650, w_128_651, w_128_654, w_128_655, w_128_660, w_128_662, w_128_663, w_128_664, w_128_667, w_128_673, w_128_676, w_128_677, w_128_683, w_128_684, w_128_686, w_128_692, w_128_693, w_128_694, w_128_699, w_128_705, w_128_706, w_128_707, w_128_709, w_128_711, w_128_712, w_128_713, w_128_720, w_128_721, w_128_723, w_128_724, w_128_725, w_128_727, w_128_729, w_128_731, w_128_732, w_128_733, w_128_735, w_128_737, w_128_738, w_128_740, w_128_741, w_128_742, w_128_749, w_128_752, w_128_753, w_128_754, w_128_755, w_128_758, w_128_759, w_128_760, w_128_763, w_128_768, w_128_770, w_128_771, w_128_772, w_128_775, w_128_776, w_128_780, w_128_781, w_128_782, w_128_784, w_128_788, w_128_791, w_128_792, w_128_793, w_128_794, w_128_799, w_128_800, w_128_802, w_128_806, w_128_807, w_128_813, w_128_814, w_128_820, w_128_824, w_128_825, w_128_828, w_128_830, w_128_834, w_128_837, w_128_838, w_128_840, w_128_841, w_128_844, w_128_845, w_128_849, w_128_858, w_128_861, w_128_863, w_128_869, w_128_870, w_128_872, w_128_873, w_128_874, w_128_878, w_128_880, w_128_884, w_128_886, w_128_891, w_128_892, w_128_893, w_128_895, w_128_896, w_128_900, w_128_904, w_128_906, w_128_908, w_128_909, w_128_910, w_128_911, w_128_912, w_128_918, w_128_919, w_128_922, w_128_926, w_128_927, w_128_928, w_128_930, w_128_932, w_128_934, w_128_935, w_128_938, w_128_940, w_128_949, w_128_950, w_128_951, w_128_954, w_128_957, w_128_958, w_128_960, w_128_962, w_128_964, w_128_967, w_128_968, w_128_969, w_128_974, w_128_975, w_128_979, w_128_984, w_128_985, w_128_986, w_128_988, w_128_991, w_128_995, w_128_1006, w_128_1009, w_128_1010, w_128_1012, w_128_1021, w_128_1022, w_128_1023, w_128_1026, w_128_1027, w_128_1030, w_128_1032, w_128_1035, w_128_1042, w_128_1047, w_128_1048, w_128_1050, w_128_1053, w_128_1056, w_128_1057, w_128_1061, w_128_1064, w_128_1067, w_128_1068, w_128_1069, w_128_1071, w_128_1073, w_128_1074, w_128_1078, w_128_1081, w_128_1085, w_128_1089, w_128_1090, w_128_1093, w_128_1098, w_128_1100, w_128_1106, w_128_1113, w_128_1114, w_128_1116, w_128_1120, w_128_1125, w_128_1126, w_128_1127, w_128_1132, w_128_1136, w_128_1137, w_128_1141, w_128_1151, w_128_1152, w_128_1153, w_128_1156, w_128_1157, w_128_1158, w_128_1160, w_128_1161, w_128_1162, w_128_1165, w_128_1166, w_128_1168, w_128_1173, w_128_1174, w_128_1175, w_128_1177, w_128_1178, w_128_1181, w_128_1185, w_128_1186, w_128_1188, w_128_1189, w_128_1192, w_128_1193, w_128_1195, w_128_1196, w_128_1197, w_128_1201, w_128_1202, w_128_1203, w_128_1208, w_128_1212, w_128_1213, w_128_1215, w_128_1218, w_128_1219, w_128_1220, w_128_1225, w_128_1228, w_128_1231, w_128_1232, w_128_1234, w_128_1236, w_128_1239, w_128_1240, w_128_1247, w_128_1248, w_128_1250, w_128_1252, w_128_1255, w_128_1267, w_128_1269, w_128_1271, w_128_1273, w_128_1277, w_128_1288, w_128_1289, w_128_1290, w_128_1291, w_128_1292, w_128_1293, w_128_1294, w_128_1298, w_128_1299, w_128_1304, w_128_1307, w_128_1308, w_128_1310, w_128_1314, w_128_1317, w_128_1318, w_128_1322, w_128_1326, w_128_1331, w_128_1332, w_128_1340, w_128_1345, w_128_1347, w_128_1348, w_128_1349, w_128_1351, w_128_1354, w_128_1359, w_128_1362, w_128_1364, w_128_1365, w_128_1366, w_128_1368, w_128_1369, w_128_1371, w_128_1373, w_128_1375, w_128_1376, w_128_1383, w_128_1385, w_128_1386, w_128_1389, w_128_1398, w_128_1402, w_128_1404, w_128_1409, w_128_1410, w_128_1413, w_128_1415, w_128_1417, w_128_1418, w_128_1419, w_128_1420, w_128_1421, w_128_1424, w_128_1425, w_128_1430, w_128_1431, w_128_1433, w_128_1436, w_128_1439, w_128_1441, w_128_1444, w_128_1445, w_128_1446, w_128_1447, w_128_1448, w_128_1452, w_128_1453, w_128_1461, w_128_1465, w_128_1468, w_128_1469, w_128_1470, w_128_1472, w_128_1478, w_128_1480, w_128_1488, w_128_1490, w_128_1491, w_128_1493, w_128_1496, w_128_1497, w_128_1498, w_128_1502, w_128_1503, w_128_1504, w_128_1509, w_128_1512, w_128_1513, w_128_1514, w_128_1515, w_128_1516, w_128_1517, w_128_1518, w_128_1521, w_128_1523, w_128_1525, w_128_1528, w_128_1529, w_128_1531, w_128_1532, w_128_1533, w_128_1537, w_128_1538, w_128_1539, w_128_1540, w_128_1543, w_128_1548, w_128_1549, w_128_1550, w_128_1552, w_128_1553, w_128_1556, w_128_1557, w_128_1559, w_128_1561, w_128_1565, w_128_1566, w_128_1576, w_128_1577, w_128_1589, w_128_1593, w_128_1594, w_128_1596, w_128_1600, w_128_1602, w_128_1604, w_128_1606, w_128_1607, w_128_1608, w_128_1611, w_128_1616, w_128_1621, w_128_1622, w_128_1623, w_128_1625, w_128_1626, w_128_1630, w_128_1632, w_128_1633, w_128_1634, w_128_1635, w_128_1638, w_128_1639, w_128_1641, w_128_1643, w_128_1644, w_128_1647, w_128_1652, w_128_1655, w_128_1656, w_128_1657, w_128_1658, w_128_1659, w_128_1664, w_128_1669, w_128_1671, w_128_1673, w_128_1679, w_128_1680, w_128_1681, w_128_1683, w_128_1688, w_128_1690, w_128_1693, w_128_1694, w_128_1700, w_128_1701, w_128_1706, w_128_1708, w_128_1709, w_128_1711, w_128_1714, w_128_1715, w_128_1716, w_128_1719, w_128_1720, w_128_1722, w_128_1727, w_128_1729, w_128_1731, w_128_1735, w_128_1736, w_128_1742, w_128_1744, w_128_1745, w_128_1747, w_128_1749, w_128_1754, w_128_1755, w_128_1758, w_128_1761, w_128_1764, w_128_1767, w_128_1768, w_128_1769, w_128_1770, w_128_1771, w_128_1773, w_128_1774, w_128_1778, w_128_1784, w_128_1785, w_128_1786, w_128_1787, w_128_1790, w_128_1792, w_128_1793, w_128_1796, w_128_1801, w_128_1802, w_128_1803, w_128_1804, w_128_1806, w_128_1808, w_128_1810, w_128_1813, w_128_1814, w_128_1819, w_128_1820, w_128_1821, w_128_1823, w_128_1824, w_128_1826, w_128_1831, w_128_1832, w_128_1833, w_128_1835, w_128_1837, w_128_1839, w_128_1840, w_128_1841, w_128_1842, w_128_1850, w_128_1853, w_128_1860, w_128_1861, w_128_1862, w_128_1866, w_128_1868, w_128_1870, w_128_1871, w_128_1872, w_128_1878, w_128_1884, w_128_1888, w_128_1890, w_128_1891, w_128_1892, w_128_1903, w_128_1904, w_128_1906, w_128_1907, w_128_1909, w_128_1913, w_128_1916, w_128_1918, w_128_1919, w_128_1922, w_128_1925, w_128_1926, w_128_1927, w_128_1929, w_128_1932, w_128_1939, w_128_1941, w_128_1942, w_128_1945, w_128_1946, w_128_1948, w_128_1954, w_128_1956, w_128_1957, w_128_1958, w_128_1960, w_128_1961, w_128_1966, w_128_1967, w_128_1968, w_128_1969, w_128_1970, w_128_1973, w_128_1975, w_128_1977, w_128_1981, w_128_1984, w_128_1985, w_128_1987, w_128_1993, w_128_1997, w_128_1999, w_128_2000, w_128_2003, w_128_2004, w_128_2005, w_128_2006, w_128_2007, w_128_2010, w_128_2012, w_128_2013, w_128_2016, w_128_2022, w_128_2025, w_128_2026, w_128_2028, w_128_2033, w_128_2036, w_128_2038, w_128_2046, w_128_2048, w_128_2054, w_128_2056, w_128_2057, w_128_2061, w_128_2066, w_128_2069, w_128_2074, w_128_2076, w_128_2077, w_128_2078, w_128_2080, w_128_2082, w_128_2083, w_128_2087, w_128_2088, w_128_2095, w_128_2096, w_128_2097, w_128_2099, w_128_2100, w_128_2101, w_128_2103, w_128_2104, w_128_2106, w_128_2108, w_128_2109, w_128_2110, w_128_2113, w_128_2114, w_128_2120, w_128_2122, w_128_2126, w_128_2127, w_128_2128, w_128_2131, w_128_2135, w_128_2136, w_128_2137, w_128_2139, w_128_2141, w_128_2143, w_128_2146, w_128_2148, w_128_2150, w_128_2152, w_128_2154, w_128_2155, w_128_2157, w_128_2165, w_128_2167, w_128_2168, w_128_2172, w_128_2173, w_128_2174, w_128_2175, w_128_2180, w_128_2182, w_128_2184, w_128_2185, w_128_2190, w_128_2191, w_128_2194, w_128_2196, w_128_2197, w_128_2199, w_128_2200, w_128_2201, w_128_2202, w_128_2204, w_128_2205, w_128_2208, w_128_2211, w_128_2219, w_128_2221, w_128_2222, w_128_2223, w_128_2229, w_128_2230, w_128_2231, w_128_2234, w_128_2238, w_128_2239, w_128_2245, w_128_2253, w_128_2254, w_128_2255, w_128_2263, w_128_2268, w_128_2269, w_128_2270, w_128_2271, w_128_2275, w_128_2280, w_128_2281, w_128_2285, w_128_2287, w_128_2291, w_128_2292, w_128_2294, w_128_2296, w_128_2298, w_128_2299, w_128_2301, w_128_2302, w_128_2304, w_128_2305, w_128_2312, w_128_2315, w_128_2320, w_128_2321, w_128_2323, w_128_2325, w_128_2328, w_128_2329, w_128_2330, w_128_2331, w_128_2333, w_128_2337, w_128_2338, w_128_2340, w_128_2344, w_128_2347, w_128_2348, w_128_2350, w_128_2352, w_128_2353, w_128_2355, w_128_2357, w_128_2359, w_128_2360, w_128_2363, w_128_2366, w_128_2368, w_128_2373, w_128_2375, w_128_2378, w_128_2379, w_128_2382, w_128_2386, w_128_2387, w_128_2396, w_128_2399, w_128_2402, w_128_2413, w_128_2416, w_128_2422, w_128_2423, w_128_2424, w_128_2427, w_128_2430, w_128_2431, w_128_2437, w_128_2443, w_128_2446, w_128_2448, w_128_2453, w_128_2456, w_128_2459, w_128_2461;
  wire w_129_000, w_129_001, w_129_002, w_129_006, w_129_007, w_129_008, w_129_013, w_129_015, w_129_017, w_129_018, w_129_020, w_129_021, w_129_023, w_129_024, w_129_025, w_129_028, w_129_029, w_129_032, w_129_033, w_129_036, w_129_039, w_129_042, w_129_044, w_129_046, w_129_047, w_129_049, w_129_050, w_129_052, w_129_054, w_129_056, w_129_063, w_129_064, w_129_067, w_129_068, w_129_069, w_129_072, w_129_073, w_129_075, w_129_077, w_129_078, w_129_079, w_129_083, w_129_084, w_129_085, w_129_095, w_129_099, w_129_108, w_129_109, w_129_110, w_129_111, w_129_112, w_129_114, w_129_115, w_129_119, w_129_120, w_129_125, w_129_128, w_129_131, w_129_132, w_129_133, w_129_134, w_129_137, w_129_140, w_129_142, w_129_144, w_129_145, w_129_152, w_129_153, w_129_161, w_129_162, w_129_167, w_129_175, w_129_180, w_129_181, w_129_182, w_129_187, w_129_189, w_129_190, w_129_195, w_129_197, w_129_202, w_129_203, w_129_205, w_129_211, w_129_212, w_129_215, w_129_220, w_129_221, w_129_222, w_129_226, w_129_227, w_129_233, w_129_234, w_129_235, w_129_236, w_129_237, w_129_239, w_129_240, w_129_243, w_129_246, w_129_254, w_129_269, w_129_275, w_129_276, w_129_278, w_129_281, w_129_286, w_129_287, w_129_290, w_129_292, w_129_297, w_129_302, w_129_305, w_129_310, w_129_314, w_129_315, w_129_317, w_129_324, w_129_326, w_129_328, w_129_329, w_129_331, w_129_332, w_129_333, w_129_335, w_129_336, w_129_341, w_129_342, w_129_343, w_129_345, w_129_346, w_129_350, w_129_351, w_129_353, w_129_354, w_129_360, w_129_361, w_129_364, w_129_368, w_129_370, w_129_372, w_129_376, w_129_377, w_129_379, w_129_381, w_129_384, w_129_386, w_129_388, w_129_391, w_129_392, w_129_400, w_129_402, w_129_405, w_129_407, w_129_409, w_129_411, w_129_416, w_129_419, w_129_420, w_129_425, w_129_426, w_129_427, w_129_428, w_129_429, w_129_431, w_129_434, w_129_439, w_129_440, w_129_442, w_129_444, w_129_448, w_129_450, w_129_454, w_129_455, w_129_456, w_129_459, w_129_460, w_129_461, w_129_463, w_129_464, w_129_466, w_129_467, w_129_472, w_129_476, w_129_478, w_129_481, w_129_483, w_129_486, w_129_487, w_129_488, w_129_490, w_129_491, w_129_493, w_129_494, w_129_495, w_129_496, w_129_498, w_129_504, w_129_507, w_129_509, w_129_512, w_129_514, w_129_517, w_129_520, w_129_522, w_129_523, w_129_526, w_129_528, w_129_529, w_129_536, w_129_538, w_129_539, w_129_544, w_129_545, w_129_546, w_129_548, w_129_551, w_129_553, w_129_555, w_129_560, w_129_563, w_129_566, w_129_568, w_129_575, w_129_576, w_129_577, w_129_581, w_129_590, w_129_592, w_129_594, w_129_595, w_129_600, w_129_602, w_129_607, w_129_609, w_129_610, w_129_616, w_129_617, w_129_618, w_129_620, w_129_622, w_129_624, w_129_627, w_129_630, w_129_636, w_129_637, w_129_638, w_129_642, w_129_643, w_129_644, w_129_649, w_129_652, w_129_653, w_129_654, w_129_660, w_129_661, w_129_662, w_129_667, w_129_668, w_129_675, w_129_681, w_129_683, w_129_687, w_129_688, w_129_689, w_129_691, w_129_693, w_129_695, w_129_696, w_129_697, w_129_700, w_129_702, w_129_704, w_129_706, w_129_709, w_129_710, w_129_711, w_129_713, w_129_716, w_129_720, w_129_722, w_129_725, w_129_726, w_129_727, w_129_728, w_129_730, w_129_733, w_129_735, w_129_736, w_129_740, w_129_742, w_129_744, w_129_745, w_129_746, w_129_747, w_129_749, w_129_751, w_129_756, w_129_760, w_129_761, w_129_764, w_129_766, w_129_767, w_129_768, w_129_769, w_129_770, w_129_772, w_129_779, w_129_783, w_129_796, w_129_797, w_129_798, w_129_800, w_129_804, w_129_806, w_129_812, w_129_814, w_129_821, w_129_826, w_129_827, w_129_828, w_129_831, w_129_832, w_129_838, w_129_840, w_129_842, w_129_843, w_129_846, w_129_849, w_129_850, w_129_853, w_129_856, w_129_857, w_129_859, w_129_861, w_129_862, w_129_867, w_129_869, w_129_871, w_129_873, w_129_874, w_129_876, w_129_878, w_129_880, w_129_881, w_129_882, w_129_884, w_129_892, w_129_893, w_129_895, w_129_898, w_129_909, w_129_911, w_129_914, w_129_922, w_129_926, w_129_928, w_129_931, w_129_933, w_129_938, w_129_939, w_129_941, w_129_942, w_129_950, w_129_954, w_129_959, w_129_965, w_129_967, w_129_977, w_129_979, w_129_980, w_129_981, w_129_984, w_129_986, w_129_989, w_129_992, w_129_999, w_129_1001, w_129_1003, w_129_1010, w_129_1011, w_129_1012, w_129_1016, w_129_1017, w_129_1019, w_129_1020, w_129_1021, w_129_1023, w_129_1024, w_129_1025, w_129_1026, w_129_1028, w_129_1029, w_129_1030, w_129_1033, w_129_1040, w_129_1044, w_129_1045, w_129_1049, w_129_1050, w_129_1060, w_129_1061, w_129_1062, w_129_1063, w_129_1064, w_129_1071, w_129_1074, w_129_1075, w_129_1077, w_129_1078, w_129_1082, w_129_1085, w_129_1087, w_129_1089, w_129_1090, w_129_1098, w_129_1100, w_129_1102, w_129_1104, w_129_1106, w_129_1110, w_129_1111, w_129_1119, w_129_1122, w_129_1123, w_129_1127, w_129_1131, w_129_1132, w_129_1135, w_129_1137, w_129_1140, w_129_1142, w_129_1148, w_129_1151, w_129_1153, w_129_1159, w_129_1160, w_129_1161, w_129_1164, w_129_1165, w_129_1168, w_129_1172, w_129_1174, w_129_1175, w_129_1176, w_129_1183, w_129_1187, w_129_1189, w_129_1190, w_129_1194, w_129_1196, w_129_1199, w_129_1202, w_129_1203, w_129_1204, w_129_1206, w_129_1207, w_129_1208, w_129_1209, w_129_1210, w_129_1212, w_129_1218, w_129_1222, w_129_1226, w_129_1227, w_129_1228, w_129_1229, w_129_1230, w_129_1232, w_129_1233, w_129_1238, w_129_1239, w_129_1240, w_129_1242, w_129_1244, w_129_1249, w_129_1257, w_129_1262, w_129_1268, w_129_1278, w_129_1279, w_129_1283, w_129_1293, w_129_1294, w_129_1300, w_129_1304, w_129_1305, w_129_1306, w_129_1312, w_129_1325, w_129_1336, w_129_1341, w_129_1342, w_129_1343, w_129_1344, w_129_1346, w_129_1349, w_129_1351, w_129_1352, w_129_1356, w_129_1370, w_129_1373, w_129_1377, w_129_1381, w_129_1383, w_129_1389, w_129_1391, w_129_1392, w_129_1397, w_129_1400, w_129_1418, w_129_1419, w_129_1422, w_129_1425, w_129_1441, w_129_1445, w_129_1446, w_129_1447, w_129_1449, w_129_1454, w_129_1456, w_129_1458, w_129_1468, w_129_1477, w_129_1478, w_129_1483, w_129_1484, w_129_1496, w_129_1497, w_129_1499, w_129_1500, w_129_1502, w_129_1508, w_129_1513, w_129_1517, w_129_1518, w_129_1527, w_129_1554, w_129_1560, w_129_1563, w_129_1570, w_129_1573, w_129_1575, w_129_1579, w_129_1587, w_129_1588, w_129_1589, w_129_1607, w_129_1613, w_129_1614, w_129_1619, w_129_1622, w_129_1624, w_129_1629, w_129_1641, w_129_1642, w_129_1656, w_129_1671, w_129_1673, w_129_1679, w_129_1680, w_129_1685, w_129_1697, w_129_1702, w_129_1703, w_129_1720, w_129_1721, w_129_1726, w_129_1729, w_129_1740, w_129_1741, w_129_1748, w_129_1777, w_129_1782, w_129_1784, w_129_1792, w_129_1793, w_129_1797, w_129_1803, w_129_1805, w_129_1806, w_129_1808, w_129_1811, w_129_1820, w_129_1823, w_129_1824, w_129_1825, w_129_1827, w_129_1831, w_129_1840, w_129_1844, w_129_1851, w_129_1855, w_129_1860, w_129_1873, w_129_1875, w_129_1882, w_129_1883, w_129_1898, w_129_1899, w_129_1904, w_129_1917, w_129_1920, w_129_1921, w_129_1930, w_129_1941, w_129_1945, w_129_1946, w_129_1954, w_129_1960, w_129_1966, w_129_1967, w_129_1968, w_129_1971, w_129_1976, w_129_1994, w_129_1996, w_129_2000, w_129_2001, w_129_2009, w_129_2019, w_129_2032, w_129_2036, w_129_2038, w_129_2039, w_129_2043, w_129_2046, w_129_2052, w_129_2063, w_129_2064, w_129_2065, w_129_2067, w_129_2080, w_129_2083, w_129_2087, w_129_2089, w_129_2096, w_129_2102, w_129_2105, w_129_2111, w_129_2113, w_129_2116, w_129_2117, w_129_2128, w_129_2131, w_129_2132, w_129_2140, w_129_2143, w_129_2145, w_129_2160, w_129_2162, w_129_2163, w_129_2164, w_129_2170, w_129_2188, w_129_2199, w_129_2206, w_129_2215, w_129_2219, w_129_2222, w_129_2223, w_129_2227, w_129_2233, w_129_2234, w_129_2236, w_129_2244, w_129_2250, w_129_2252, w_129_2260, w_129_2261, w_129_2262, w_129_2279, w_129_2283, w_129_2290, w_129_2294, w_129_2295, w_129_2299, w_129_2306, w_129_2307, w_129_2315, w_129_2317, w_129_2320, w_129_2325, w_129_2329, w_129_2333, w_129_2335, w_129_2337, w_129_2340, w_129_2342, w_129_2344, w_129_2346, w_129_2347, w_129_2352, w_129_2358, w_129_2359, w_129_2361, w_129_2369, w_129_2374, w_129_2381, w_129_2384, w_129_2386, w_129_2389, w_129_2398, w_129_2401, w_129_2406, w_129_2407, w_129_2411, w_129_2421, w_129_2425, w_129_2427, w_129_2428, w_129_2431, w_129_2446, w_129_2459, w_129_2461, w_129_2468, w_129_2474, w_129_2475, w_129_2481, w_129_2483, w_129_2486, w_129_2487, w_129_2492, w_129_2495, w_129_2500, w_129_2502, w_129_2507, w_129_2513, w_129_2516, w_129_2517, w_129_2522, w_129_2529, w_129_2534, w_129_2545, w_129_2546, w_129_2555, w_129_2563, w_129_2569, w_129_2575, w_129_2576, w_129_2578, w_129_2583, w_129_2587, w_129_2594, w_129_2598, w_129_2602, w_129_2606, w_129_2609, w_129_2610, w_129_2616, w_129_2628, w_129_2630, w_129_2638, w_129_2639, w_129_2644, w_129_2651, w_129_2653, w_129_2659, w_129_2660, w_129_2661, w_129_2665, w_129_2668, w_129_2677, w_129_2681, w_129_2684, w_129_2692, w_129_2695, w_129_2706, w_129_2707, w_129_2719, w_129_2720, w_129_2737, w_129_2741, w_129_2748, w_129_2751, w_129_2752, w_129_2759, w_129_2774, w_129_2777, w_129_2778, w_129_2779, w_129_2787, w_129_2788, w_129_2793, w_129_2794, w_129_2796, w_129_2806, w_129_2807, w_129_2813, w_129_2814, w_129_2815, w_129_2825, w_129_2826, w_129_2833, w_129_2836, w_129_2840, w_129_2841, w_129_2850, w_129_2856, w_129_2857, w_129_2862, w_129_2873, w_129_2876, w_129_2885, w_129_2891, w_129_2893, w_129_2896, w_129_2905, w_129_2906, w_129_2910, w_129_2922, w_129_2928, w_129_2929, w_129_2940, w_129_2943, w_129_2946, w_129_2953, w_129_2954, w_129_2961, w_129_2964, w_129_2967, w_129_2972, w_129_2973, w_129_2981, w_129_2986, w_129_2988, w_129_2990, w_129_2993, w_129_3004, w_129_3006, w_129_3008, w_129_3009, w_129_3018, w_129_3025, w_129_3031, w_129_3033, w_129_3034, w_129_3037, w_129_3040, w_129_3050, w_129_3051, w_129_3052, w_129_3054, w_129_3055, w_129_3067, w_129_3072, w_129_3074, w_129_3076, w_129_3083, w_129_3087, w_129_3090, w_129_3103, w_129_3111, w_129_3115, w_129_3118, w_129_3124, w_129_3127, w_129_3134, w_129_3143, w_129_3145, w_129_3153, w_129_3154, w_129_3156, w_129_3161, w_129_3163, w_129_3175, w_129_3176, w_129_3182, w_129_3183, w_129_3187, w_129_3201, w_129_3202, w_129_3212, w_129_3213, w_129_3214, w_129_3217, w_129_3218, w_129_3219, w_129_3225, w_129_3229, w_129_3238, w_129_3242, w_129_3244, w_129_3246, w_129_3247, w_129_3254, w_129_3258, w_129_3262, w_129_3268, w_129_3275, w_129_3278, w_129_3282, w_129_3296, w_129_3297, w_129_3302, w_129_3309, w_129_3310, w_129_3313, w_129_3314, w_129_3317, w_129_3319, w_129_3323, w_129_3324, w_129_3330, w_129_3337, w_129_3340, w_129_3349, w_129_3350, w_129_3351, w_129_3358, w_129_3361, w_129_3370, w_129_3374, w_129_3376, w_129_3380, w_129_3385, w_129_3386, w_129_3393, w_129_3394, w_129_3395, w_129_3396, w_129_3398, w_129_3403, w_129_3409, w_129_3418, w_129_3419, w_129_3420, w_129_3424, w_129_3427, w_129_3431, w_129_3432, w_129_3434, w_129_3443, w_129_3448, w_129_3450, w_129_3451, w_129_3454, w_129_3459, w_129_3460, w_129_3470, w_129_3473, w_129_3477, w_129_3478, w_129_3480, w_129_3481, w_129_3484, w_129_3485, w_129_3506, w_129_3511, w_129_3512, w_129_3520, w_129_3524, w_129_3525, w_129_3529, w_129_3530, w_129_3544, w_129_3549, w_129_3550, w_129_3556, w_129_3560, w_129_3562, w_129_3565, w_129_3566, w_129_3567, w_129_3573, w_129_3574, w_129_3579, w_129_3581, w_129_3584, w_129_3589, w_129_3616, w_129_3619, w_129_3622, w_129_3625, w_129_3627, w_129_3635, w_129_3650, w_129_3651, w_129_3657, w_129_3664, w_129_3666, w_129_3670, w_129_3678, w_129_3679, w_129_3681, w_129_3682, w_129_3690, w_129_3691, w_129_3692, w_129_3699, w_129_3702, w_129_3703, w_129_3713, w_129_3715, w_129_3723, w_129_3725, w_129_3730, w_129_3746, w_129_3748;
  wire w_130_006, w_130_007, w_130_011, w_130_014, w_130_017, w_130_020, w_130_024, w_130_025, w_130_026, w_130_027, w_130_031, w_130_034, w_130_035, w_130_036, w_130_041, w_130_042, w_130_043, w_130_052, w_130_054, w_130_059, w_130_060, w_130_062, w_130_068, w_130_071, w_130_076, w_130_077, w_130_078, w_130_083, w_130_084, w_130_088, w_130_096, w_130_101, w_130_102, w_130_105, w_130_107, w_130_109, w_130_110, w_130_112, w_130_114, w_130_116, w_130_117, w_130_119, w_130_121, w_130_122, w_130_127, w_130_129, w_130_132, w_130_134, w_130_135, w_130_138, w_130_140, w_130_141, w_130_146, w_130_148, w_130_150, w_130_151, w_130_152, w_130_158, w_130_164, w_130_165, w_130_166, w_130_170, w_130_172, w_130_175, w_130_178, w_130_179, w_130_182, w_130_184, w_130_190, w_130_194, w_130_197, w_130_198, w_130_203, w_130_206, w_130_207, w_130_208, w_130_211, w_130_214, w_130_217, w_130_224, w_130_225, w_130_226, w_130_230, w_130_238, w_130_243, w_130_245, w_130_246, w_130_248, w_130_251, w_130_254, w_130_257, w_130_262, w_130_264, w_130_266, w_130_267, w_130_270, w_130_271, w_130_273, w_130_274, w_130_276, w_130_277, w_130_279, w_130_283, w_130_284, w_130_285, w_130_290, w_130_291, w_130_292, w_130_293, w_130_296, w_130_297, w_130_299, w_130_300, w_130_303, w_130_306, w_130_308, w_130_309, w_130_315, w_130_317, w_130_318, w_130_320, w_130_321, w_130_322, w_130_323, w_130_324, w_130_325, w_130_327, w_130_330, w_130_332, w_130_337, w_130_339, w_130_341, w_130_355, w_130_356, w_130_357, w_130_358, w_130_360, w_130_365, w_130_366, w_130_367, w_130_374, w_130_376, w_130_381, w_130_384, w_130_385, w_130_391, w_130_394, w_130_398, w_130_402, w_130_403, w_130_404, w_130_405, w_130_407, w_130_414, w_130_418, w_130_419, w_130_423, w_130_424, w_130_429, w_130_430, w_130_431, w_130_437, w_130_439, w_130_440, w_130_444, w_130_446, w_130_448, w_130_450, w_130_452, w_130_453, w_130_460, w_130_461, w_130_465, w_130_467, w_130_468, w_130_469, w_130_474, w_130_480, w_130_481, w_130_484, w_130_485, w_130_487, w_130_489, w_130_490, w_130_491, w_130_492, w_130_497, w_130_499, w_130_500, w_130_501, w_130_502, w_130_503, w_130_504, w_130_505, w_130_506, w_130_509, w_130_515, w_130_516, w_130_517, w_130_518, w_130_520, w_130_529, w_130_530, w_130_534, w_130_538, w_130_546, w_130_550, w_130_551, w_130_559, w_130_566, w_130_567, w_130_569, w_130_571, w_130_572, w_130_574, w_130_576, w_130_577, w_130_579, w_130_581, w_130_582, w_130_585, w_130_587, w_130_591, w_130_592, w_130_601, w_130_602, w_130_604, w_130_605, w_130_606, w_130_608, w_130_609, w_130_610, w_130_611, w_130_612, w_130_613, w_130_614, w_130_617, w_130_618, w_130_619, w_130_623, w_130_627, w_130_629, w_130_631, w_130_637, w_130_639, w_130_642, w_130_657, w_130_666, w_130_670, w_130_672, w_130_676, w_130_679, w_130_683, w_130_684, w_130_685, w_130_686, w_130_687, w_130_689, w_130_693, w_130_695, w_130_701, w_130_707, w_130_708, w_130_709, w_130_710, w_130_711, w_130_721, w_130_723, w_130_725, w_130_726, w_130_727, w_130_730, w_130_732, w_130_734, w_130_740, w_130_746, w_130_747, w_130_748, w_130_752, w_130_756, w_130_758, w_130_763, w_130_764, w_130_765, w_130_769, w_130_770, w_130_771, w_130_780, w_130_781, w_130_782, w_130_787, w_130_788, w_130_793, w_130_796, w_130_797, w_130_799, w_130_802, w_130_803, w_130_806, w_130_808, w_130_810, w_130_812, w_130_815, w_130_816, w_130_817, w_130_819, w_130_827, w_130_828, w_130_836, w_130_838, w_130_846, w_130_849, w_130_854, w_130_857, w_130_860, w_130_865, w_130_867, w_130_870, w_130_871, w_130_873, w_130_874, w_130_876, w_130_880, w_130_882, w_130_884, w_130_885, w_130_886, w_130_887, w_130_890, w_130_894, w_130_897, w_130_898, w_130_899, w_130_901, w_130_904, w_130_905, w_130_908, w_130_911, w_130_912, w_130_913, w_130_914, w_130_917, w_130_919, w_130_920, w_130_921, w_130_923, w_130_927, w_130_928, w_130_930, w_130_934, w_130_937, w_130_942, w_130_943, w_130_944, w_130_945, w_130_954, w_130_960, w_130_962, w_130_964, w_130_965, w_130_966, w_130_969, w_130_970, w_130_976, w_130_977, w_130_979, w_130_980, w_130_981, w_130_982, w_130_984, w_130_985, w_130_986, w_130_987, w_130_988, w_130_990, w_130_992, w_130_996, w_130_997, w_130_998, w_130_1002, w_130_1004, w_130_1007, w_130_1012, w_130_1014, w_130_1016, w_130_1018, w_130_1021, w_130_1025, w_130_1027, w_130_1028, w_130_1035, w_130_1038, w_130_1049, w_130_1051, w_130_1060, w_130_1067, w_130_1068, w_130_1070, w_130_1072, w_130_1073, w_130_1079, w_130_1081, w_130_1085, w_130_1086, w_130_1091, w_130_1094, w_130_1096, w_130_1100, w_130_1103, w_130_1106, w_130_1109, w_130_1110, w_130_1123, w_130_1127, w_130_1128, w_130_1129, w_130_1131, w_130_1134, w_130_1135, w_130_1138, w_130_1139, w_130_1140, w_130_1141, w_130_1150, w_130_1151, w_130_1154, w_130_1159, w_130_1160, w_130_1164, w_130_1167, w_130_1168, w_130_1169, w_130_1176, w_130_1179, w_130_1181, w_130_1183, w_130_1184, w_130_1187, w_130_1188, w_130_1189, w_130_1191, w_130_1195, w_130_1199, w_130_1200, w_130_1202, w_130_1206, w_130_1207, w_130_1210, w_130_1211, w_130_1213, w_130_1215, w_130_1218, w_130_1220, w_130_1224, w_130_1230, w_130_1232, w_130_1238, w_130_1252, w_130_1260, w_130_1265, w_130_1266, w_130_1269, w_130_1271, w_130_1278, w_130_1280, w_130_1281, w_130_1287, w_130_1289, w_130_1294, w_130_1295, w_130_1297, w_130_1298, w_130_1301, w_130_1304, w_130_1306, w_130_1308, w_130_1313, w_130_1320, w_130_1326, w_130_1327, w_130_1330, w_130_1334, w_130_1341, w_130_1343, w_130_1346, w_130_1349, w_130_1351, w_130_1353, w_130_1354, w_130_1374, w_130_1379, w_130_1387, w_130_1389, w_130_1392, w_130_1399, w_130_1407, w_130_1421, w_130_1424, w_130_1426, w_130_1428, w_130_1429, w_130_1432, w_130_1433, w_130_1435, w_130_1442, w_130_1444, w_130_1445, w_130_1455, w_130_1458, w_130_1463, w_130_1472, w_130_1479, w_130_1480, w_130_1493, w_130_1496, w_130_1498, w_130_1502, w_130_1506, w_130_1518, w_130_1521, w_130_1524, w_130_1532, w_130_1533, w_130_1534, w_130_1540, w_130_1547, w_130_1550, w_130_1554, w_130_1561, w_130_1567, w_130_1569, w_130_1571, w_130_1576, w_130_1581, w_130_1583, w_130_1589, w_130_1590, w_130_1592, w_130_1602, w_130_1603, w_130_1607, w_130_1619, w_130_1624, w_130_1628, w_130_1631, w_130_1633, w_130_1639, w_130_1643, w_130_1645, w_130_1647, w_130_1653, w_130_1658, w_130_1661, w_130_1662, w_130_1663, w_130_1664, w_130_1665, w_130_1668, w_130_1669, w_130_1676, w_130_1682, w_130_1688, w_130_1691, w_130_1702, w_130_1703, w_130_1707, w_130_1708, w_130_1710, w_130_1713, w_130_1715, w_130_1717, w_130_1720, w_130_1721, w_130_1724, w_130_1728, w_130_1732, w_130_1734, w_130_1736, w_130_1738, w_130_1742, w_130_1747, w_130_1757, w_130_1764, w_130_1771, w_130_1773, w_130_1777, w_130_1781, w_130_1784, w_130_1795, w_130_1796, w_130_1800, w_130_1810, w_130_1816, w_130_1820, w_130_1821, w_130_1825, w_130_1827, w_130_1832, w_130_1833, w_130_1834, w_130_1839, w_130_1850, w_130_1856, w_130_1859, w_130_1866, w_130_1867, w_130_1875, w_130_1876, w_130_1883, w_130_1887, w_130_1888, w_130_1900, w_130_1904, w_130_1905, w_130_1907, w_130_1908, w_130_1914, w_130_1916, w_130_1928, w_130_1934, w_130_1941, w_130_1942, w_130_1944, w_130_1948, w_130_1950, w_130_1952, w_130_1958, w_130_1964, w_130_1968, w_130_1969, w_130_1971, w_130_1982, w_130_1992, w_130_2001, w_130_2004, w_130_2006, w_130_2009, w_130_2013, w_130_2014, w_130_2015, w_130_2025, w_130_2026, w_130_2033, w_130_2039, w_130_2040, w_130_2041, w_130_2042, w_130_2047, w_130_2051, w_130_2055, w_130_2058, w_130_2060, w_130_2063, w_130_2064, w_130_2065, w_130_2067, w_130_2070, w_130_2075, w_130_2076, w_130_2092, w_130_2094, w_130_2101, w_130_2103, w_130_2110, w_130_2116, w_130_2117, w_130_2143, w_130_2144, w_130_2148, w_130_2149, w_130_2154, w_130_2179, w_130_2181, w_130_2193, w_130_2197, w_130_2201, w_130_2216, w_130_2221, w_130_2230, w_130_2235, w_130_2238, w_130_2247, w_130_2253, w_130_2256, w_130_2257, w_130_2265, w_130_2267, w_130_2268, w_130_2276, w_130_2281, w_130_2283, w_130_2287, w_130_2288, w_130_2289, w_130_2290, w_130_2297, w_130_2298, w_130_2299, w_130_2307, w_130_2309, w_130_2310, w_130_2312, w_130_2313, w_130_2315, w_130_2317, w_130_2318, w_130_2322, w_130_2337, w_130_2338, w_130_2342, w_130_2345, w_130_2349, w_130_2361, w_130_2362, w_130_2364, w_130_2367, w_130_2370, w_130_2371, w_130_2373, w_130_2385, w_130_2387, w_130_2391, w_130_2408, w_130_2419, w_130_2420, w_130_2424, w_130_2432, w_130_2436, w_130_2437, w_130_2444, w_130_2451, w_130_2452, w_130_2454, w_130_2460, w_130_2463, w_130_2482, w_130_2484, w_130_2485, w_130_2489, w_130_2490, w_130_2495, w_130_2497, w_130_2498, w_130_2510, w_130_2511, w_130_2514, w_130_2517, w_130_2522, w_130_2523, w_130_2525, w_130_2538, w_130_2540, w_130_2541, w_130_2543, w_130_2545, w_130_2548, w_130_2557, w_130_2561, w_130_2576, w_130_2577, w_130_2578, w_130_2579, w_130_2582, w_130_2585, w_130_2587, w_130_2591, w_130_2604, w_130_2606, w_130_2613, w_130_2616, w_130_2624, w_130_2628, w_130_2646, w_130_2648, w_130_2653, w_130_2654, w_130_2660, w_130_2663, w_130_2665, w_130_2666, w_130_2669, w_130_2670, w_130_2674, w_130_2677, w_130_2679, w_130_2683, w_130_2698, w_130_2705, w_130_2711, w_130_2713, w_130_2721, w_130_2724, w_130_2731, w_130_2733, w_130_2735, w_130_2736, w_130_2750, w_130_2751, w_130_2752, w_130_2753, w_130_2759, w_130_2761, w_130_2766, w_130_2769, w_130_2775, w_130_2783, w_130_2793, w_130_2799, w_130_2801, w_130_2803, w_130_2810, w_130_2813, w_130_2817, w_130_2821, w_130_2825, w_130_2831, w_130_2833, w_130_2834, w_130_2846, w_130_2848, w_130_2850, w_130_2851, w_130_2862, w_130_2863, w_130_2871, w_130_2876, w_130_2877, w_130_2879, w_130_2887, w_130_2898, w_130_2905, w_130_2906, w_130_2914, w_130_2916, w_130_2918, w_130_2925, w_130_2932, w_130_2941, w_130_2945, w_130_2946, w_130_2947, w_130_2954, w_130_2958, w_130_2960, w_130_2967, w_130_2971, w_130_2974, w_130_2978, w_130_2982, w_130_2985, w_130_2996, w_130_3001, w_130_3002, w_130_3004, w_130_3007, w_130_3008, w_130_3012, w_130_3029, w_130_3030, w_130_3031, w_130_3032, w_130_3037, w_130_3041, w_130_3044, w_130_3051, w_130_3078, w_130_3080, w_130_3088, w_130_3101, w_130_3105, w_130_3107, w_130_3109, w_130_3117, w_130_3120, w_130_3121, w_130_3123, w_130_3128, w_130_3131, w_130_3141, w_130_3143, w_130_3156, w_130_3161, w_130_3163, w_130_3168, w_130_3171, w_130_3180, w_130_3183, w_130_3184, w_130_3187, w_130_3189, w_130_3194, w_130_3195, w_130_3203, w_130_3207, w_130_3208, w_130_3209, w_130_3210, w_130_3213, w_130_3214, w_130_3215, w_130_3221, w_130_3223, w_130_3235, w_130_3240, w_130_3248, w_130_3257, w_130_3262, w_130_3263, w_130_3267, w_130_3269, w_130_3275, w_130_3276, w_130_3282, w_130_3304, w_130_3312, w_130_3313, w_130_3323, w_130_3329, w_130_3331, w_130_3333, w_130_3339, w_130_3345, w_130_3347, w_130_3357, w_130_3358, w_130_3361, w_130_3362, w_130_3373, w_130_3374, w_130_3379, w_130_3382, w_130_3383, w_130_3385, w_130_3386, w_130_3389, w_130_3398, w_130_3399, w_130_3403, w_130_3411, w_130_3414, w_130_3418, w_130_3420, w_130_3426, w_130_3436, w_130_3438, w_130_3440, w_130_3443, w_130_3444, w_130_3446, w_130_3461, w_130_3466, w_130_3467, w_130_3468, w_130_3479, w_130_3486, w_130_3490, w_130_3508, w_130_3510, w_130_3514, w_130_3522, w_130_3532, w_130_3534, w_130_3539, w_130_3541, w_130_3545, w_130_3549, w_130_3556, w_130_3559, w_130_3570, w_130_3579, w_130_3582, w_130_3588, w_130_3590, w_130_3591, w_130_3594, w_130_3595, w_130_3624, w_130_3628, w_130_3632, w_130_3633, w_130_3638, w_130_3645, w_130_3652, w_130_3657, w_130_3658, w_130_3659, w_130_3668, w_130_3669, w_130_3675, w_130_3691, w_130_3695, w_130_3708, w_130_3710, w_130_3713, w_130_3715, w_130_3731, w_130_3732, w_130_3742, w_130_3756, w_130_3757, w_130_3762, w_130_3763, w_130_3767, w_130_3770, w_130_3771, w_130_3772, w_130_3773, w_130_3774, w_130_3775, w_130_3776, w_130_3777, w_130_3778, w_130_3779, w_130_3780, w_130_3784, w_130_3785, w_130_3786, w_130_3790, w_130_3791, w_130_3792, w_130_3793, w_130_3794, w_130_3795, w_130_3796, w_130_3797, w_130_3798, w_130_3799, w_130_3800, w_130_3801, w_130_3803;
  wire w_131_005, w_131_007, w_131_010, w_131_012, w_131_019, w_131_020, w_131_021, w_131_026, w_131_027, w_131_032, w_131_033, w_131_038, w_131_042, w_131_047, w_131_048, w_131_051, w_131_052, w_131_055, w_131_058, w_131_059, w_131_060, w_131_062, w_131_069, w_131_071, w_131_074, w_131_076, w_131_081, w_131_082, w_131_085, w_131_087, w_131_091, w_131_092, w_131_098, w_131_101, w_131_104, w_131_105, w_131_106, w_131_107, w_131_108, w_131_111, w_131_114, w_131_115, w_131_120, w_131_124, w_131_125, w_131_128, w_131_130, w_131_132, w_131_133, w_131_135, w_131_139, w_131_142, w_131_144, w_131_145, w_131_148, w_131_149, w_131_151, w_131_152, w_131_153, w_131_158, w_131_159, w_131_161, w_131_166, w_131_169, w_131_170, w_131_171, w_131_172, w_131_174, w_131_175, w_131_176, w_131_179, w_131_182, w_131_183, w_131_187, w_131_188, w_131_190, w_131_196, w_131_197, w_131_209, w_131_212, w_131_216, w_131_218, w_131_220, w_131_223, w_131_228, w_131_230, w_131_232, w_131_237, w_131_240, w_131_242, w_131_249, w_131_257, w_131_259, w_131_260, w_131_261, w_131_267, w_131_268, w_131_269, w_131_275, w_131_279, w_131_284, w_131_286, w_131_287, w_131_290, w_131_291, w_131_298, w_131_299, w_131_300, w_131_301, w_131_306, w_131_308, w_131_309, w_131_311, w_131_312, w_131_313, w_131_315, w_131_320, w_131_325, w_131_326, w_131_330, w_131_338, w_131_339, w_131_341, w_131_342, w_131_343, w_131_346, w_131_349, w_131_353, w_131_354, w_131_355, w_131_357, w_131_360, w_131_362, w_131_365, w_131_366, w_131_369, w_131_373, w_131_375, w_131_377, w_131_378, w_131_379, w_131_380, w_131_381, w_131_382, w_131_387, w_131_388, w_131_393, w_131_394, w_131_395, w_131_404, w_131_414, w_131_415, w_131_416, w_131_417, w_131_420, w_131_424, w_131_426, w_131_429, w_131_432, w_131_436, w_131_437, w_131_438, w_131_443, w_131_446, w_131_447, w_131_450, w_131_451, w_131_455, w_131_459, w_131_461, w_131_463, w_131_468, w_131_473, w_131_477, w_131_478, w_131_487, w_131_488, w_131_493, w_131_501, w_131_506, w_131_509, w_131_512, w_131_515, w_131_517, w_131_518, w_131_519, w_131_523, w_131_526, w_131_528, w_131_532, w_131_535, w_131_536, w_131_537, w_131_538, w_131_540, w_131_541, w_131_543, w_131_546, w_131_547, w_131_549, w_131_550, w_131_556, w_131_557, w_131_577, w_131_579, w_131_581, w_131_583, w_131_588, w_131_589, w_131_593, w_131_595, w_131_598, w_131_601, w_131_603, w_131_607, w_131_608, w_131_611, w_131_613, w_131_617, w_131_620, w_131_627, w_131_629, w_131_632, w_131_642, w_131_643, w_131_646, w_131_647, w_131_649, w_131_650, w_131_654, w_131_655, w_131_657, w_131_665, w_131_667, w_131_670, w_131_671, w_131_672, w_131_676, w_131_679, w_131_685, w_131_687, w_131_689, w_131_692, w_131_694, w_131_695, w_131_700, w_131_701, w_131_702, w_131_703, w_131_706, w_131_707, w_131_708, w_131_709, w_131_716, w_131_717, w_131_721, w_131_722, w_131_724, w_131_729, w_131_731, w_131_735, w_131_737, w_131_748, w_131_757, w_131_760, w_131_762, w_131_764, w_131_765, w_131_769, w_131_771, w_131_772, w_131_773, w_131_790, w_131_795, w_131_800, w_131_801, w_131_803, w_131_805, w_131_812, w_131_816, w_131_818, w_131_831, w_131_834, w_131_840, w_131_841, w_131_844, w_131_847, w_131_848, w_131_849, w_131_851, w_131_852, w_131_857, w_131_858, w_131_861, w_131_863, w_131_867, w_131_868, w_131_886, w_131_887, w_131_891, w_131_893, w_131_911, w_131_912, w_131_913, w_131_918, w_131_921, w_131_923, w_131_927, w_131_934, w_131_935, w_131_936, w_131_941, w_131_961, w_131_962, w_131_971, w_131_977, w_131_983, w_131_984, w_131_986, w_131_989, w_131_992, w_131_993, w_131_994, w_131_1005, w_131_1007, w_131_1010, w_131_1014, w_131_1017, w_131_1019, w_131_1024, w_131_1026, w_131_1036, w_131_1043, w_131_1049, w_131_1068, w_131_1080, w_131_1084, w_131_1099, w_131_1100, w_131_1104, w_131_1106, w_131_1118, w_131_1124, w_131_1126, w_131_1127, w_131_1128, w_131_1132, w_131_1143, w_131_1144, w_131_1146, w_131_1147, w_131_1148, w_131_1152, w_131_1153, w_131_1155, w_131_1169, w_131_1170, w_131_1172, w_131_1189, w_131_1190, w_131_1196, w_131_1205, w_131_1213, w_131_1231, w_131_1233, w_131_1234, w_131_1239, w_131_1244, w_131_1245, w_131_1246, w_131_1248, w_131_1250, w_131_1251, w_131_1258, w_131_1273, w_131_1274, w_131_1279, w_131_1283, w_131_1288, w_131_1293, w_131_1294, w_131_1295, w_131_1297, w_131_1298, w_131_1300, w_131_1308, w_131_1309, w_131_1310, w_131_1333, w_131_1338, w_131_1339, w_131_1347, w_131_1350, w_131_1351, w_131_1358, w_131_1359, w_131_1365, w_131_1367, w_131_1374, w_131_1375, w_131_1384, w_131_1385, w_131_1391, w_131_1393, w_131_1396, w_131_1405, w_131_1415, w_131_1416, w_131_1418, w_131_1420, w_131_1421, w_131_1423, w_131_1435, w_131_1437, w_131_1444, w_131_1448, w_131_1450, w_131_1455, w_131_1456, w_131_1458, w_131_1459, w_131_1469, w_131_1476, w_131_1480, w_131_1486, w_131_1489, w_131_1498, w_131_1501, w_131_1503, w_131_1506, w_131_1507, w_131_1511, w_131_1515, w_131_1530, w_131_1534, w_131_1535, w_131_1536, w_131_1545, w_131_1551, w_131_1554, w_131_1558, w_131_1568, w_131_1576, w_131_1578, w_131_1583, w_131_1584, w_131_1588, w_131_1590, w_131_1607, w_131_1616, w_131_1617, w_131_1623, w_131_1626, w_131_1627, w_131_1628, w_131_1629, w_131_1639, w_131_1641, w_131_1646, w_131_1647, w_131_1648, w_131_1655, w_131_1673, w_131_1680, w_131_1681, w_131_1686, w_131_1687, w_131_1694, w_131_1700, w_131_1708, w_131_1711, w_131_1714, w_131_1716, w_131_1727, w_131_1731, w_131_1739, w_131_1743, w_131_1748, w_131_1764, w_131_1768, w_131_1779, w_131_1792, w_131_1795, w_131_1796, w_131_1797, w_131_1801, w_131_1809, w_131_1810, w_131_1813, w_131_1818, w_131_1823, w_131_1825, w_131_1833, w_131_1836, w_131_1837, w_131_1849, w_131_1853, w_131_1859, w_131_1861, w_131_1880, w_131_1882, w_131_1885, w_131_1887, w_131_1900, w_131_1902, w_131_1905, w_131_1917, w_131_1922, w_131_1924, w_131_1929, w_131_1930, w_131_1932, w_131_1933, w_131_1938, w_131_1940, w_131_1942, w_131_1943, w_131_1944, w_131_1954, w_131_1956, w_131_1957, w_131_1958, w_131_1961, w_131_1965, w_131_1976, w_131_1979, w_131_1980, w_131_1983, w_131_1984, w_131_1991, w_131_1992, w_131_1994, w_131_1995, w_131_2005, w_131_2007, w_131_2018, w_131_2022, w_131_2026, w_131_2027, w_131_2039, w_131_2041, w_131_2042, w_131_2044, w_131_2048, w_131_2049, w_131_2055, w_131_2057, w_131_2062, w_131_2064, w_131_2070, w_131_2077, w_131_2083, w_131_2088, w_131_2092, w_131_2097, w_131_2110, w_131_2111, w_131_2113, w_131_2115, w_131_2116, w_131_2117, w_131_2123, w_131_2126, w_131_2134, w_131_2146, w_131_2151, w_131_2162, w_131_2173, w_131_2190, w_131_2192, w_131_2193, w_131_2200, w_131_2201, w_131_2206, w_131_2210, w_131_2214, w_131_2216, w_131_2218, w_131_2222, w_131_2223, w_131_2224, w_131_2225, w_131_2228, w_131_2239, w_131_2243, w_131_2245, w_131_2252, w_131_2260, w_131_2264, w_131_2265, w_131_2270, w_131_2275, w_131_2276, w_131_2280, w_131_2292, w_131_2293, w_131_2296, w_131_2297, w_131_2298, w_131_2300, w_131_2304, w_131_2305, w_131_2307, w_131_2308, w_131_2310, w_131_2319, w_131_2322, w_131_2326, w_131_2331, w_131_2335, w_131_2347, w_131_2349, w_131_2355, w_131_2361, w_131_2365, w_131_2371, w_131_2379, w_131_2382, w_131_2402, w_131_2415, w_131_2418, w_131_2425, w_131_2428, w_131_2429, w_131_2432, w_131_2434, w_131_2439, w_131_2441, w_131_2448, w_131_2451, w_131_2454, w_131_2456, w_131_2457, w_131_2460, w_131_2461, w_131_2463, w_131_2469, w_131_2471, w_131_2481, w_131_2488, w_131_2504, w_131_2509, w_131_2525, w_131_2541, w_131_2543, w_131_2545, w_131_2553, w_131_2556, w_131_2557, w_131_2566, w_131_2569, w_131_2576, w_131_2577, w_131_2580, w_131_2584, w_131_2594, w_131_2597, w_131_2598, w_131_2604, w_131_2607, w_131_2609, w_131_2616, w_131_2623, w_131_2628, w_131_2629, w_131_2645, w_131_2650, w_131_2654, w_131_2655, w_131_2659, w_131_2665, w_131_2670, w_131_2674, w_131_2679, w_131_2685, w_131_2689, w_131_2692, w_131_2696, w_131_2707, w_131_2711, w_131_2716, w_131_2721, w_131_2730, w_131_2731, w_131_2734, w_131_2735, w_131_2744, w_131_2746, w_131_2752, w_131_2754, w_131_2755, w_131_2770, w_131_2783, w_131_2786, w_131_2789, w_131_2790, w_131_2792, w_131_2793, w_131_2799, w_131_2800, w_131_2802, w_131_2810, w_131_2812, w_131_2818, w_131_2822, w_131_2829, w_131_2832, w_131_2833, w_131_2834, w_131_2837, w_131_2838, w_131_2839, w_131_2844, w_131_2850, w_131_2851, w_131_2853, w_131_2855, w_131_2858, w_131_2863, w_131_2864, w_131_2867, w_131_2874, w_131_2875, w_131_2880, w_131_2884, w_131_2886, w_131_2888, w_131_2889, w_131_2895, w_131_2897, w_131_2902, w_131_2903, w_131_2909, w_131_2914, w_131_2927, w_131_2941, w_131_2942, w_131_2943, w_131_2947, w_131_2949, w_131_2952, w_131_2954, w_131_2959, w_131_2960, w_131_2967, w_131_2969, w_131_2977, w_131_2986, w_131_2987, w_131_2993, w_131_2994, w_131_3002, w_131_3004, w_131_3014, w_131_3021, w_131_3024, w_131_3030, w_131_3035, w_131_3039, w_131_3041, w_131_3044, w_131_3048, w_131_3050, w_131_3056, w_131_3057, w_131_3067, w_131_3070, w_131_3078, w_131_3079, w_131_3083, w_131_3088, w_131_3096, w_131_3098, w_131_3099, w_131_3100, w_131_3105, w_131_3108, w_131_3111, w_131_3115, w_131_3117, w_131_3120, w_131_3125, w_131_3129, w_131_3156, w_131_3165, w_131_3167, w_131_3170, w_131_3185, w_131_3188, w_131_3189, w_131_3191, w_131_3192, w_131_3194, w_131_3199, w_131_3205, w_131_3213, w_131_3214, w_131_3215, w_131_3219, w_131_3220, w_131_3221, w_131_3225, w_131_3248, w_131_3257, w_131_3258, w_131_3265, w_131_3269, w_131_3271, w_131_3272, w_131_3310, w_131_3312, w_131_3317, w_131_3320, w_131_3323, w_131_3332, w_131_3333, w_131_3345, w_131_3347, w_131_3348, w_131_3358, w_131_3361, w_131_3371, w_131_3376, w_131_3377, w_131_3378, w_131_3385, w_131_3392, w_131_3395, w_131_3399, w_131_3407, w_131_3411, w_131_3413, w_131_3418, w_131_3427, w_131_3429, w_131_3431, w_131_3433, w_131_3437, w_131_3441, w_131_3448, w_131_3449, w_131_3451, w_131_3454, w_131_3460, w_131_3465, w_131_3469, w_131_3470, w_131_3474, w_131_3479, w_131_3482, w_131_3485, w_131_3488, w_131_3489, w_131_3490, w_131_3495, w_131_3502, w_131_3504, w_131_3509, w_131_3510, w_131_3513, w_131_3518, w_131_3520, w_131_3522, w_131_3534, w_131_3542, w_131_3545, w_131_3550, w_131_3555, w_131_3556, w_131_3563, w_131_3571, w_131_3572, w_131_3578, w_131_3580, w_131_3589, w_131_3593, w_131_3599, w_131_3610, w_131_3613, w_131_3621, w_131_3626, w_131_3632, w_131_3638, w_131_3642, w_131_3645, w_131_3647, w_131_3651, w_131_3654, w_131_3655, w_131_3656, w_131_3675, w_131_3679, w_131_3680, w_131_3688, w_131_3694, w_131_3695, w_131_3698, w_131_3706, w_131_3707, w_131_3711, w_131_3717, w_131_3719, w_131_3722, w_131_3728, w_131_3744, w_131_3748, w_131_3751, w_131_3755, w_131_3756, w_131_3757, w_131_3759, w_131_3764, w_131_3765, w_131_3772, w_131_3778, w_131_3780, w_131_3783, w_131_3786, w_131_3787, w_131_3790, w_131_3797, w_131_3804, w_131_3814, w_131_3815, w_131_3817, w_131_3824, w_131_3825, w_131_3827, w_131_3829, w_131_3835, w_131_3838, w_131_3858, w_131_3865, w_131_3868, w_131_3869, w_131_3883, w_131_3886, w_131_3889, w_131_3895, w_131_3898, w_131_3902, w_131_3905, w_131_3914, w_131_3915, w_131_3918, w_131_3926, w_131_3929, w_131_3935, w_131_3936, w_131_3952, w_131_3954, w_131_3957, w_131_3963, w_131_3969, w_131_3971, w_131_3977, w_131_3984, w_131_3986, w_131_3987, w_131_3996, w_131_3997, w_131_4005, w_131_4006, w_131_4008, w_131_4016, w_131_4019, w_131_4021, w_131_4026, w_131_4033, w_131_4035, w_131_4054, w_131_4056, w_131_4059, w_131_4064, w_131_4065, w_131_4068, w_131_4070, w_131_4088, w_131_4102, w_131_4104, w_131_4106, w_131_4109, w_131_4110, w_131_4112, w_131_4122, w_131_4133, w_131_4134, w_131_4139, w_131_4142, w_131_4144, w_131_4148, w_131_4152, w_131_4158, w_131_4160, w_131_4165, w_131_4167, w_131_4177, w_131_4185, w_131_4195, w_131_4207, w_131_4214, w_131_4218, w_131_4223, w_131_4226, w_131_4228, w_131_4237, w_131_4238, w_131_4239, w_131_4244, w_131_4246, w_131_4247, w_131_4250, w_131_4255, w_131_4256, w_131_4257, w_131_4258, w_131_4259, w_131_4260, w_131_4264, w_131_4265, w_131_4266, w_131_4267, w_131_4269;
  wire w_132_001, w_132_002, w_132_003, w_132_005, w_132_009, w_132_011, w_132_012, w_132_014, w_132_016, w_132_020, w_132_021, w_132_023, w_132_025, w_132_026, w_132_029, w_132_032, w_132_034, w_132_037, w_132_038, w_132_039, w_132_040, w_132_041, w_132_042, w_132_045, w_132_049, w_132_050, w_132_051, w_132_053, w_132_054, w_132_056, w_132_057, w_132_058, w_132_061, w_132_064, w_132_066, w_132_067, w_132_069, w_132_071, w_132_073, w_132_075, w_132_076, w_132_079, w_132_080, w_132_085, w_132_086, w_132_088, w_132_090, w_132_092, w_132_098, w_132_100, w_132_102, w_132_103, w_132_105, w_132_108, w_132_109, w_132_110, w_132_112, w_132_116, w_132_118, w_132_119, w_132_121, w_132_123, w_132_124, w_132_126, w_132_127, w_132_128, w_132_129, w_132_131, w_132_136, w_132_141, w_132_147, w_132_150, w_132_152, w_132_155, w_132_157, w_132_159, w_132_160, w_132_161, w_132_163, w_132_164, w_132_165, w_132_167, w_132_169, w_132_172, w_132_173, w_132_174, w_132_180, w_132_185, w_132_186, w_132_188, w_132_189, w_132_190, w_132_191, w_132_194, w_132_195, w_132_197, w_132_199, w_132_200, w_132_201, w_132_202, w_132_206, w_132_208, w_132_210, w_132_211, w_132_214, w_132_217, w_132_218, w_132_220, w_132_222, w_132_225, w_132_228, w_132_229, w_132_233, w_132_234, w_132_236, w_132_237, w_132_238, w_132_240, w_132_243, w_132_244, w_132_246, w_132_247, w_132_250, w_132_251, w_132_252, w_132_253, w_132_259, w_132_261, w_132_262, w_132_263, w_132_265, w_132_266, w_132_271, w_132_272, w_132_275, w_132_276, w_132_278, w_132_279, w_132_288, w_132_290, w_132_291, w_132_293, w_132_297, w_132_298, w_132_299, w_132_302, w_132_303, w_132_304, w_132_305, w_132_306, w_132_307, w_132_309, w_132_311, w_132_316, w_132_318, w_132_321, w_132_322, w_132_323, w_132_324, w_132_327, w_132_329, w_132_332, w_132_333, w_132_336, w_132_339, w_132_342, w_132_344, w_132_345, w_132_346, w_132_348, w_132_349, w_132_351, w_132_352, w_132_354, w_132_355, w_132_356, w_132_357, w_132_359, w_132_361, w_132_362, w_132_364, w_132_365, w_132_368, w_132_370, w_132_372, w_132_373, w_132_374, w_132_376, w_132_377, w_132_379, w_132_381, w_132_383, w_132_384, w_132_385, w_132_387, w_132_393, w_132_394, w_132_396, w_132_397, w_132_398, w_132_399, w_132_401, w_132_403, w_132_404, w_132_409, w_132_413, w_132_414, w_132_415, w_132_419, w_132_420, w_132_421, w_132_422, w_132_423, w_132_426, w_132_429, w_132_431, w_132_434, w_132_435, w_132_436, w_132_437, w_132_439, w_132_441, w_132_442, w_132_444, w_132_445, w_132_446, w_132_447, w_132_449, w_132_450, w_132_451, w_132_452, w_132_453, w_132_455, w_132_457, w_132_458, w_132_460, w_132_461, w_132_463, w_132_465, w_132_467, w_132_469, w_132_471, w_132_472, w_132_473, w_132_476, w_132_477, w_132_478, w_132_480, w_132_481, w_132_482, w_132_483, w_132_484, w_132_486, w_132_487, w_132_488, w_132_489, w_132_491, w_132_494, w_132_495, w_132_496, w_132_499, w_132_504, w_132_506, w_132_508, w_132_510, w_132_512, w_132_513, w_132_514, w_132_516, w_132_517, w_132_518, w_132_519, w_132_522, w_132_523, w_132_524, w_132_527, w_132_529, w_132_531, w_132_532, w_132_534, w_132_535, w_132_536, w_132_537, w_132_539, w_132_546, w_132_548, w_132_549, w_132_552, w_132_553, w_132_554, w_132_557, w_132_561, w_132_562, w_132_566, w_132_567, w_132_569, w_132_573, w_132_574, w_132_575, w_132_577, w_132_578, w_132_579, w_132_580, w_132_583, w_132_584, w_132_586, w_132_587, w_132_588, w_132_589, w_132_591, w_132_592, w_132_598, w_132_600, w_132_601, w_132_602, w_132_604, w_132_605, w_132_606, w_132_607, w_132_611, w_132_612, w_132_615, w_132_616, w_132_618, w_132_619, w_132_621, w_132_623, w_132_624, w_132_628, w_132_631, w_132_634, w_132_635, w_132_636, w_132_637, w_132_638, w_132_640, w_132_641, w_132_643, w_132_644, w_132_648, w_132_649, w_132_654, w_132_658, w_132_659, w_132_660, w_132_661, w_132_664, w_132_665, w_132_669, w_132_672, w_132_673, w_132_676, w_132_678, w_132_679, w_132_680, w_132_683, w_132_687, w_132_689, w_132_693, w_132_695, w_132_698, w_132_699, w_132_701, w_132_704, w_132_707, w_132_708, w_132_714, w_132_717, w_132_718, w_132_719, w_132_721, w_132_722, w_132_732, w_132_733, w_132_734, w_132_735, w_132_736, w_132_740, w_132_741, w_132_743, w_132_744, w_132_745, w_132_746, w_132_747, w_132_749, w_132_753, w_132_754, w_132_759, w_132_760, w_132_761, w_132_764, w_132_766, w_132_769, w_132_770, w_132_774, w_132_775, w_132_778, w_132_779, w_132_781, w_132_782, w_132_784, w_132_785, w_132_787, w_132_789, w_132_793, w_132_794, w_132_795, w_132_798, w_132_799, w_132_801, w_132_802, w_132_807, w_132_808, w_132_811, w_132_815, w_132_817, w_132_818, w_132_820, w_132_823, w_132_824, w_132_825, w_132_826, w_132_828, w_132_831, w_132_833, w_132_836, w_132_837, w_132_838, w_132_840, w_132_841, w_132_844, w_132_845, w_132_846, w_132_848, w_132_850, w_132_851, w_132_852, w_132_857, w_132_858, w_132_860, w_132_864, w_132_867, w_132_870, w_132_872, w_132_877, w_132_879, w_132_880, w_132_881, w_132_882, w_132_883, w_132_885, w_132_888, w_132_889, w_132_890, w_132_891, w_132_894, w_132_895, w_132_896, w_132_898, w_132_899, w_132_900, w_132_905, w_132_907, w_132_908, w_132_909, w_132_910, w_132_912, w_132_914, w_132_915, w_132_918, w_132_919, w_132_920, w_132_921, w_132_922, w_132_924, w_132_928, w_132_930, w_132_931, w_132_932, w_132_933, w_132_934, w_132_935, w_132_939, w_132_940, w_132_942, w_132_943, w_132_945, w_132_950, w_132_951, w_132_952, w_132_958, w_132_962, w_132_964, w_132_965, w_132_966, w_132_967, w_132_970, w_132_974, w_132_975, w_132_976, w_132_977, w_132_978, w_132_979, w_132_981, w_132_982, w_132_983, w_132_985, w_132_987, w_132_988, w_132_989, w_132_990, w_132_991, w_132_992, w_132_1000, w_132_1001, w_132_1003, w_132_1004, w_132_1005, w_132_1006, w_132_1008, w_132_1011, w_132_1012, w_132_1014, w_132_1016, w_132_1017, w_132_1019, w_132_1020, w_132_1021, w_132_1022, w_132_1026, w_132_1027, w_132_1028, w_132_1029, w_132_1030, w_132_1032, w_132_1038, w_132_1040, w_132_1044, w_132_1045, w_132_1048, w_132_1050, w_132_1051, w_132_1053, w_132_1054, w_132_1057, w_132_1058, w_132_1059, w_132_1064, w_132_1065, w_132_1066, w_132_1067, w_132_1068, w_132_1070, w_132_1072, w_132_1073, w_132_1075, w_132_1076, w_132_1077, w_132_1078, w_132_1079, w_132_1080, w_132_1081, w_132_1082, w_132_1083, w_132_1084, w_132_1087, w_132_1088, w_132_1089, w_132_1090, w_132_1092, w_132_1095, w_132_1096, w_132_1097, w_132_1100, w_132_1104, w_132_1105, w_132_1107, w_132_1108, w_132_1109, w_132_1112, w_132_1120, w_132_1122, w_132_1124, w_132_1127, w_132_1128, w_132_1130, w_132_1131, w_132_1132, w_132_1133, w_132_1134, w_132_1135, w_132_1137, w_132_1141, w_132_1142, w_132_1144, w_132_1148, w_132_1150, w_132_1152, w_132_1153, w_132_1154, w_132_1155, w_132_1157, w_132_1159, w_132_1164, w_132_1165, w_132_1167, w_132_1169, w_132_1172, w_132_1173, w_132_1178, w_132_1180, w_132_1181, w_132_1184, w_132_1186, w_132_1187, w_132_1192, w_132_1193, w_132_1194, w_132_1195, w_132_1196, w_132_1198, w_132_1200, w_132_1203, w_132_1204, w_132_1211, w_132_1212, w_132_1213, w_132_1216, w_132_1217, w_132_1222, w_132_1227, w_132_1231, w_132_1233, w_132_1234, w_132_1237, w_132_1241, w_132_1245, w_132_1246, w_132_1247, w_132_1248, w_132_1250, w_132_1251, w_132_1253, w_132_1254, w_132_1259, w_132_1260, w_132_1266, w_132_1268, w_132_1270, w_132_1277, w_132_1279, w_132_1280, w_132_1281, w_132_1282, w_132_1285, w_132_1289, w_132_1291, w_132_1293, w_132_1296, w_132_1299, w_132_1304, w_132_1307, w_132_1311, w_132_1312, w_132_1322, w_132_1323, w_132_1324, w_132_1328, w_132_1331, w_132_1332, w_132_1333, w_132_1334, w_132_1336, w_132_1342, w_132_1343, w_132_1346, w_132_1348, w_132_1353, w_132_1354, w_132_1355, w_132_1366, w_132_1367, w_132_1369, w_132_1370, w_132_1373, w_132_1375, w_132_1379, w_132_1385, w_132_1386, w_132_1388, w_132_1389, w_132_1396, w_132_1401, w_132_1402, w_132_1403, w_132_1404, w_132_1407, w_132_1408, w_132_1409, w_132_1416, w_132_1427, w_132_1431, w_132_1432, w_132_1438, w_132_1440, w_132_1441, w_132_1444, w_132_1445, w_132_1446, w_132_1447, w_132_1448, w_132_1450, w_132_1451, w_132_1457, w_132_1458, w_132_1459, w_132_1464, w_132_1465, w_132_1473, w_132_1475, w_132_1477, w_132_1478, w_132_1481, w_132_1486, w_132_1487, w_132_1488, w_132_1496, w_132_1501, w_132_1502, w_132_1505, w_132_1509, w_132_1511, w_132_1514, w_132_1515, w_132_1516, w_132_1518, w_132_1519, w_132_1523, w_132_1525, w_132_1527, w_132_1530, w_132_1538, w_132_1539, w_132_1543, w_132_1544, w_132_1547, w_132_1548, w_132_1549, w_132_1552, w_132_1556, w_132_1558, w_132_1561, w_132_1562, w_132_1563, w_132_1566, w_132_1569, w_132_1571, w_132_1575, w_132_1577, w_132_1578, w_132_1579, w_132_1580, w_132_1585, w_132_1586, w_132_1588, w_132_1589, w_132_1590, w_132_1591, w_132_1592, w_132_1597, w_132_1599, w_132_1601, w_132_1606, w_132_1612, w_132_1613, w_132_1617, w_132_1619, w_132_1624, w_132_1627, w_132_1633, w_132_1636, w_132_1637, w_132_1643, w_132_1648, w_132_1650, w_132_1651, w_132_1652, w_132_1654, w_132_1661, w_132_1662, w_132_1667, w_132_1668, w_132_1672, w_132_1673, w_132_1678, w_132_1680, w_132_1684, w_132_1686, w_132_1688, w_132_1692, w_132_1696, w_132_1697, w_132_1698, w_132_1700, w_132_1702, w_132_1704, w_132_1706, w_132_1707, w_132_1710, w_132_1717, w_132_1719, w_132_1720, w_132_1721, w_132_1722, w_132_1725, w_132_1728, w_132_1731, w_132_1736, w_132_1737, w_132_1741, w_132_1743, w_132_1746, w_132_1748, w_132_1750, w_132_1752, w_132_1755, w_132_1757, w_132_1759, w_132_1764, w_132_1766, w_132_1769, w_132_1770, w_132_1771, w_132_1773, w_132_1774, w_132_1775, w_132_1776, w_132_1778, w_132_1780, w_132_1782, w_132_1785, w_132_1793, w_132_1794, w_132_1795, w_132_1798, w_132_1801, w_132_1802, w_132_1804, w_132_1807, w_132_1812, w_132_1816, w_132_1818, w_132_1824, w_132_1830, w_132_1831, w_132_1832, w_132_1833, w_132_1836, w_132_1838, w_132_1840, w_132_1841, w_132_1842, w_132_1843, w_132_1845, w_132_1848, w_132_1849, w_132_1855, w_132_1858, w_132_1859, w_132_1860, w_132_1861, w_132_1864, w_132_1865, w_132_1866, w_132_1867, w_132_1868, w_132_1875, w_132_1876, w_132_1877, w_132_1878, w_132_1879, w_132_1880, w_132_1881, w_132_1882, w_132_1886, w_132_1887, w_132_1888, w_132_1889, w_132_1890, w_132_1891, w_132_1893, w_132_1895, w_132_1896, w_132_1897, w_132_1898, w_132_1899, w_132_1900, w_132_1901, w_132_1902, w_132_1903, w_132_1905;
  wire w_133_000, w_133_006, w_133_007, w_133_008, w_133_009, w_133_010, w_133_012, w_133_013, w_133_014, w_133_015, w_133_016, w_133_018, w_133_019, w_133_020, w_133_021, w_133_024, w_133_026, w_133_027, w_133_028, w_133_029, w_133_032, w_133_034, w_133_035, w_133_036, w_133_037, w_133_039, w_133_041, w_133_042, w_133_043, w_133_044, w_133_045, w_133_046, w_133_047, w_133_049, w_133_050, w_133_051, w_133_053, w_133_055, w_133_056, w_133_057, w_133_058, w_133_059, w_133_060, w_133_061, w_133_062, w_133_064, w_133_065, w_133_067, w_133_068, w_133_069, w_133_070, w_133_072, w_133_073, w_133_074, w_133_075, w_133_076, w_133_077, w_133_078, w_133_079, w_133_080, w_133_081, w_133_082, w_133_083, w_133_085, w_133_086, w_133_087, w_133_088, w_133_089, w_133_090, w_133_091, w_133_092, w_133_093, w_133_094, w_133_095, w_133_096, w_133_098, w_133_099, w_133_102, w_133_103, w_133_104, w_133_106, w_133_108, w_133_111, w_133_112, w_133_114, w_133_116, w_133_117, w_133_118, w_133_120, w_133_121, w_133_122, w_133_124, w_133_127, w_133_128, w_133_129, w_133_130, w_133_131, w_133_133, w_133_134, w_133_135, w_133_136, w_133_137, w_133_139, w_133_140, w_133_141, w_133_143, w_133_144, w_133_147, w_133_149, w_133_150, w_133_152, w_133_153, w_133_154, w_133_155, w_133_156, w_133_157, w_133_158, w_133_159, w_133_160, w_133_161, w_133_162, w_133_164, w_133_165, w_133_166, w_133_167, w_133_168, w_133_172, w_133_173, w_133_174, w_133_175, w_133_176, w_133_178, w_133_179, w_133_180, w_133_181, w_133_182, w_133_185, w_133_186, w_133_187, w_133_188, w_133_189, w_133_190, w_133_193, w_133_194, w_133_198, w_133_201, w_133_202, w_133_204, w_133_205, w_133_206, w_133_207, w_133_208, w_133_211, w_133_212, w_133_213, w_133_214, w_133_216, w_133_218, w_133_219, w_133_221, w_133_222, w_133_223, w_133_224, w_133_225, w_133_226, w_133_227, w_133_229, w_133_232, w_133_233, w_133_234, w_133_235, w_133_236, w_133_237, w_133_238, w_133_239, w_133_240, w_133_242, w_133_245, w_133_246, w_133_247, w_133_248, w_133_249, w_133_250, w_133_251, w_133_252, w_133_253, w_133_254, w_133_255, w_133_256, w_133_260, w_133_262, w_133_263, w_133_264, w_133_265, w_133_266, w_133_267, w_133_268, w_133_269, w_133_270, w_133_271, w_133_272, w_133_273, w_133_275, w_133_276, w_133_277, w_133_278, w_133_283, w_133_286, w_133_288, w_133_289, w_133_290, w_133_292, w_133_293, w_133_294, w_133_295, w_133_296, w_133_297, w_133_298, w_133_299, w_133_301, w_133_303, w_133_304, w_133_305, w_133_306, w_133_307, w_133_308, w_133_309, w_133_310, w_133_312, w_133_313, w_133_314, w_133_315, w_133_316, w_133_317, w_133_319, w_133_321, w_133_322, w_133_323, w_133_324, w_133_325, w_133_328, w_133_330, w_133_331, w_133_332, w_133_333, w_133_335, w_133_337, w_133_338, w_133_340, w_133_342, w_133_344, w_133_345, w_133_346, w_133_347, w_133_348, w_133_349, w_133_350, w_133_351, w_133_353, w_133_357, w_133_359, w_133_360, w_133_361, w_133_366, w_133_367, w_133_368, w_133_369, w_133_371, w_133_372, w_133_373, w_133_374, w_133_375, w_133_376, w_133_378, w_133_379, w_133_380, w_133_382, w_133_384, w_133_386, w_133_387, w_133_388, w_133_393, w_133_394, w_133_395, w_133_396, w_133_399, w_133_401, w_133_402, w_133_403, w_133_405, w_133_408, w_133_410, w_133_411, w_133_412, w_133_413, w_133_414, w_133_415, w_133_416, w_133_417, w_133_420, w_133_422, w_133_423, w_133_424, w_133_425, w_133_427, w_133_428, w_133_432, w_133_433, w_133_434, w_133_435, w_133_438, w_133_439, w_133_441, w_133_443, w_133_444, w_133_446, w_133_447, w_133_448, w_133_449, w_133_450, w_133_451, w_133_452, w_133_454, w_133_459, w_133_461, w_133_462, w_133_464, w_133_466, w_133_467, w_133_469, w_133_471, w_133_472, w_133_473, w_133_474, w_133_476, w_133_477, w_133_478, w_133_479, w_133_480, w_133_481, w_133_482, w_133_484, w_133_485, w_133_486, w_133_487, w_133_489, w_133_490, w_133_492, w_133_494, w_133_495, w_133_497, w_133_498, w_133_499, w_133_500, w_133_501, w_133_503, w_133_504, w_133_505, w_133_506, w_133_507, w_133_509, w_133_512, w_133_513, w_133_518, w_133_522, w_133_523, w_133_525, w_133_526, w_133_528, w_133_529, w_133_531, w_133_533, w_133_534, w_133_535, w_133_536, w_133_538, w_133_539, w_133_540, w_133_541, w_133_542, w_133_543, w_133_544, w_133_545, w_133_546, w_133_547, w_133_548, w_133_549, w_133_550, w_133_551, w_133_552, w_133_553, w_133_555, w_133_556, w_133_557, w_133_558, w_133_559, w_133_561, w_133_562, w_133_563, w_133_569, w_133_570, w_133_571, w_133_572, w_133_573, w_133_574, w_133_577, w_133_578, w_133_580, w_133_581, w_133_582, w_133_583, w_133_584, w_133_588, w_133_589, w_133_591, w_133_592, w_133_593, w_133_594, w_133_596, w_133_597, w_133_599, w_133_601, w_133_603, w_133_605, w_133_606, w_133_608, w_133_609, w_133_610, w_133_613, w_133_614, w_133_615, w_133_616, w_133_618, w_133_620, w_133_622, w_133_623, w_133_624, w_133_625, w_133_626, w_133_627, w_133_629, w_133_630, w_133_632, w_133_633, w_133_634, w_133_635, w_133_636, w_133_637, w_133_638, w_133_640, w_133_641, w_133_642, w_133_643, w_133_645, w_133_646, w_133_648, w_133_650, w_133_651, w_133_652, w_133_653, w_133_658, w_133_659, w_133_661, w_133_662, w_133_663, w_133_664, w_133_665, w_133_666, w_133_667, w_133_668, w_133_669, w_133_671, w_133_672, w_133_674, w_133_675, w_133_676, w_133_679, w_133_680, w_133_681, w_133_683, w_133_684, w_133_685, w_133_686, w_133_688, w_133_689, w_133_690, w_133_693, w_133_695, w_133_696, w_133_697, w_133_698, w_133_699, w_133_700, w_133_701, w_133_703, w_133_705, w_133_706, w_133_707, w_133_708, w_133_709, w_133_710, w_133_711, w_133_712, w_133_713, w_133_714, w_133_715, w_133_716, w_133_718, w_133_719, w_133_720, w_133_721, w_133_722, w_133_723, w_133_724, w_133_726, w_133_727, w_133_728, w_133_730, w_133_732, w_133_733, w_133_736, w_133_738, w_133_739, w_133_740, w_133_743, w_133_745, w_133_746, w_133_747, w_133_748, w_133_749, w_133_751, w_133_752, w_133_753, w_133_754, w_133_755, w_133_756, w_133_757, w_133_758, w_133_759, w_133_762, w_133_764, w_133_765, w_133_766, w_133_767, w_133_769, w_133_770, w_133_771, w_133_772, w_133_774, w_133_775, w_133_776, w_133_777, w_133_778, w_133_780, w_133_781, w_133_783, w_133_784, w_133_785, w_133_786, w_133_787, w_133_790, w_133_791, w_133_793, w_133_794, w_133_795, w_133_796, w_133_797, w_133_799, w_133_802, w_133_803, w_133_804, w_133_805, w_133_806, w_133_807, w_133_808, w_133_809, w_133_812, w_133_813, w_133_815, w_133_818, w_133_819, w_133_820, w_133_822, w_133_823, w_133_824, w_133_825, w_133_826, w_133_827, w_133_828, w_133_830, w_133_831, w_133_834, w_133_836, w_133_838, w_133_839, w_133_841, w_133_842, w_133_843, w_133_844, w_133_845, w_133_846, w_133_847, w_133_848, w_133_849, w_133_850, w_133_851, w_133_852, w_133_853, w_133_855, w_133_856, w_133_857, w_133_858, w_133_859, w_133_860, w_133_862, w_133_864, w_133_867, w_133_868, w_133_869, w_133_874, w_133_875, w_133_876, w_133_878, w_133_884, w_133_885, w_133_887, w_133_888, w_133_889, w_133_891, w_133_894, w_133_895, w_133_898, w_133_899, w_133_901, w_133_902, w_133_903, w_133_904, w_133_907, w_133_908, w_133_909, w_133_910, w_133_912, w_133_914, w_133_916, w_133_917, w_133_918, w_133_919, w_133_920, w_133_921, w_133_927, w_133_929, w_133_930, w_133_931, w_133_932, w_133_933, w_133_934, w_133_936, w_133_938, w_133_940, w_133_941, w_133_943, w_133_944, w_133_945, w_133_946, w_133_947, w_133_949, w_133_951, w_133_952, w_133_953, w_133_954, w_133_955, w_133_956, w_133_957, w_133_959, w_133_960, w_133_961, w_133_962, w_133_963, w_133_964, w_133_965, w_133_967, w_133_968, w_133_969, w_133_970, w_133_971, w_133_972, w_133_974, w_133_975, w_133_980;
  wire w_134_004, w_134_008, w_134_012, w_134_016, w_134_017, w_134_021, w_134_022, w_134_024, w_134_025, w_134_027, w_134_031, w_134_032, w_134_034, w_134_035, w_134_037, w_134_042, w_134_048, w_134_052, w_134_054, w_134_056, w_134_058, w_134_065, w_134_067, w_134_073, w_134_082, w_134_087, w_134_096, w_134_097, w_134_103, w_134_104, w_134_107, w_134_108, w_134_109, w_134_110, w_134_113, w_134_118, w_134_121, w_134_122, w_134_125, w_134_126, w_134_127, w_134_128, w_134_131, w_134_133, w_134_134, w_134_139, w_134_145, w_134_146, w_134_149, w_134_150, w_134_151, w_134_153, w_134_160, w_134_161, w_134_163, w_134_165, w_134_168, w_134_169, w_134_182, w_134_187, w_134_191, w_134_192, w_134_194, w_134_196, w_134_197, w_134_203, w_134_208, w_134_212, w_134_215, w_134_220, w_134_221, w_134_227, w_134_229, w_134_232, w_134_234, w_134_235, w_134_241, w_134_246, w_134_247, w_134_254, w_134_258, w_134_263, w_134_268, w_134_272, w_134_273, w_134_276, w_134_277, w_134_278, w_134_281, w_134_283, w_134_285, w_134_286, w_134_287, w_134_288, w_134_289, w_134_291, w_134_292, w_134_293, w_134_294, w_134_296, w_134_298, w_134_299, w_134_301, w_134_306, w_134_309, w_134_310, w_134_312, w_134_314, w_134_315, w_134_322, w_134_329, w_134_330, w_134_331, w_134_332, w_134_333, w_134_335, w_134_337, w_134_338, w_134_339, w_134_340, w_134_342, w_134_343, w_134_344, w_134_346, w_134_350, w_134_352, w_134_356, w_134_357, w_134_361, w_134_362, w_134_363, w_134_369, w_134_370, w_134_377, w_134_379, w_134_385, w_134_386, w_134_387, w_134_390, w_134_392, w_134_396, w_134_397, w_134_401, w_134_407, w_134_408, w_134_411, w_134_412, w_134_413, w_134_415, w_134_416, w_134_423, w_134_431, w_134_432, w_134_433, w_134_436, w_134_437, w_134_440, w_134_441, w_134_444, w_134_447, w_134_448, w_134_449, w_134_453, w_134_455, w_134_457, w_134_460, w_134_461, w_134_465, w_134_470, w_134_476, w_134_480, w_134_487, w_134_492, w_134_496, w_134_499, w_134_502, w_134_504, w_134_506, w_134_507, w_134_509, w_134_510, w_134_513, w_134_515, w_134_520, w_134_523, w_134_527, w_134_530, w_134_532, w_134_533, w_134_535, w_134_536, w_134_537, w_134_538, w_134_541, w_134_543, w_134_547, w_134_548, w_134_551, w_134_552, w_134_553, w_134_555, w_134_556, w_134_557, w_134_558, w_134_561, w_134_563, w_134_566, w_134_567, w_134_568, w_134_573, w_134_576, w_134_579, w_134_584, w_134_585, w_134_586, w_134_589, w_134_593, w_134_594, w_134_596, w_134_597, w_134_598, w_134_603, w_134_605, w_134_607, w_134_609, w_134_611, w_134_613, w_134_614, w_134_616, w_134_617, w_134_618, w_134_621, w_134_623, w_134_624, w_134_625, w_134_626, w_134_632, w_134_639, w_134_640, w_134_644, w_134_648, w_134_656, w_134_664, w_134_667, w_134_670, w_134_671, w_134_674, w_134_679, w_134_680, w_134_684, w_134_688, w_134_702, w_134_704, w_134_707, w_134_711, w_134_715, w_134_716, w_134_723, w_134_729, w_134_730, w_134_731, w_134_733, w_134_739, w_134_740, w_134_742, w_134_746, w_134_750, w_134_752, w_134_755, w_134_756, w_134_758, w_134_759, w_134_762, w_134_764, w_134_767, w_134_770, w_134_777, w_134_780, w_134_783, w_134_784, w_134_787, w_134_788, w_134_789, w_134_790, w_134_791, w_134_797, w_134_803, w_134_804, w_134_806, w_134_807, w_134_814, w_134_822, w_134_827, w_134_829, w_134_834, w_134_835, w_134_840, w_134_841, w_134_842, w_134_846, w_134_852, w_134_853, w_134_854, w_134_856, w_134_858, w_134_859, w_134_860, w_134_863, w_134_865, w_134_869, w_134_870, w_134_871, w_134_876, w_134_877, w_134_881, w_134_883, w_134_886, w_134_888, w_134_890, w_134_899, w_134_902, w_134_903, w_134_904, w_134_906, w_134_908, w_134_910, w_134_914, w_134_920, w_134_931, w_134_932, w_134_933, w_134_936, w_134_938, w_134_945, w_134_948, w_134_952, w_134_955, w_134_956, w_134_959, w_134_961, w_134_964, w_134_966, w_134_969, w_134_970, w_134_971, w_134_974, w_134_979, w_134_982, w_134_987, w_134_988, w_134_989, w_134_994, w_134_998, w_134_1003, w_134_1007, w_134_1008, w_134_1014, w_134_1016, w_134_1017, w_134_1020, w_134_1026, w_134_1028, w_134_1037, w_134_1047, w_134_1049, w_134_1054, w_134_1055, w_134_1057, w_134_1062, w_134_1064, w_134_1066, w_134_1068, w_134_1069, w_134_1070, w_134_1076, w_134_1078, w_134_1080, w_134_1087, w_134_1088, w_134_1090, w_134_1098, w_134_1099, w_134_1101, w_134_1105, w_134_1106, w_134_1107, w_134_1112, w_134_1115, w_134_1117, w_134_1118, w_134_1122, w_134_1124, w_134_1133, w_134_1134, w_134_1135, w_134_1138, w_134_1139, w_134_1140, w_134_1143, w_134_1144, w_134_1149, w_134_1151, w_134_1159, w_134_1160, w_134_1162, w_134_1163, w_134_1165, w_134_1169, w_134_1177, w_134_1180, w_134_1183, w_134_1184, w_134_1186, w_134_1188, w_134_1190, w_134_1194, w_134_1196, w_134_1199, w_134_1201, w_134_1202, w_134_1206, w_134_1208, w_134_1212, w_134_1214, w_134_1216, w_134_1221, w_134_1229, w_134_1230, w_134_1235, w_134_1240, w_134_1242, w_134_1243, w_134_1245, w_134_1246, w_134_1247, w_134_1248, w_134_1249, w_134_1251, w_134_1254, w_134_1257, w_134_1258, w_134_1259, w_134_1262, w_134_1264, w_134_1266, w_134_1267, w_134_1270, w_134_1273, w_134_1275, w_134_1276, w_134_1280, w_134_1286, w_134_1292, w_134_1293, w_134_1294, w_134_1295, w_134_1296, w_134_1299, w_134_1307, w_134_1308, w_134_1310, w_134_1313, w_134_1314, w_134_1316, w_134_1319, w_134_1324, w_134_1326, w_134_1334, w_134_1337, w_134_1338, w_134_1339, w_134_1340, w_134_1342, w_134_1345, w_134_1347, w_134_1348, w_134_1353, w_134_1356, w_134_1358, w_134_1360, w_134_1361, w_134_1362, w_134_1363, w_134_1366, w_134_1368, w_134_1375, w_134_1376, w_134_1378, w_134_1379, w_134_1380, w_134_1383, w_134_1384, w_134_1387, w_134_1391, w_134_1392, w_134_1396, w_134_1399, w_134_1401, w_134_1403, w_134_1405, w_134_1408, w_134_1409, w_134_1414, w_134_1415, w_134_1417, w_134_1419, w_134_1420, w_134_1423, w_134_1425, w_134_1429, w_134_1430, w_134_1434, w_134_1435, w_134_1437, w_134_1443, w_134_1444, w_134_1449, w_134_1450, w_134_1451, w_134_1453, w_134_1454, w_134_1455, w_134_1458, w_134_1459, w_134_1461, w_134_1462, w_134_1466, w_134_1467, w_134_1468, w_134_1469, w_134_1473, w_134_1476, w_134_1478, w_134_1481, w_134_1487, w_134_1488, w_134_1490, w_134_1495, w_134_1496, w_134_1497, w_134_1500, w_134_1501, w_134_1505, w_134_1506, w_134_1508, w_134_1509, w_134_1512, w_134_1519, w_134_1522, w_134_1524, w_134_1529, w_134_1535, w_134_1537, w_134_1541, w_134_1543, w_134_1551, w_134_1553, w_134_1554, w_134_1557, w_134_1561, w_134_1567, w_134_1570, w_134_1576, w_134_1579, w_134_1584, w_134_1585, w_134_1588, w_134_1591, w_134_1592, w_134_1596, w_134_1601, w_134_1602, w_134_1603, w_134_1604, w_134_1606, w_134_1608, w_134_1618, w_134_1619, w_134_1621, w_134_1622, w_134_1630, w_134_1631, w_134_1632, w_134_1634, w_134_1638, w_134_1644, w_134_1645, w_134_1647, w_134_1649, w_134_1652, w_134_1653, w_134_1655, w_134_1657, w_134_1658, w_134_1661, w_134_1666, w_134_1668, w_134_1669, w_134_1676, w_134_1679, w_134_1680, w_134_1688, w_134_1694, w_134_1697, w_134_1698, w_134_1702, w_134_1703, w_134_1704, w_134_1706, w_134_1707, w_134_1709, w_134_1712, w_134_1714, w_134_1715, w_134_1716, w_134_1717, w_134_1718, w_134_1719, w_134_1722, w_134_1725, w_134_1727, w_134_1728, w_134_1729, w_134_1730, w_134_1731, w_134_1736, w_134_1740, w_134_1742, w_134_1747, w_134_1749, w_134_1753, w_134_1755, w_134_1756, w_134_1757, w_134_1767, w_134_1769, w_134_1772, w_134_1778, w_134_1779, w_134_1782, w_134_1783, w_134_1785, w_134_1789, w_134_1790, w_134_1791, w_134_1793, w_134_1796, w_134_1797, w_134_1804, w_134_1809, w_134_1810, w_134_1815, w_134_1816, w_134_1817, w_134_1820, w_134_1822, w_134_1823, w_134_1834, w_134_1835, w_134_1836, w_134_1841, w_134_1844, w_134_1845, w_134_1846, w_134_1847, w_134_1850, w_134_1853, w_134_1854, w_134_1857, w_134_1858, w_134_1861, w_134_1863, w_134_1864, w_134_1867, w_134_1869, w_134_1870, w_134_1871, w_134_1873, w_134_1879, w_134_1880, w_134_1882, w_134_1886, w_134_1889, w_134_1893, w_134_1894, w_134_1896, w_134_1899, w_134_1904, w_134_1906, w_134_1908, w_134_1911, w_134_1914, w_134_1915, w_134_1924, w_134_1925, w_134_1926, w_134_1936, w_134_1939, w_134_1940, w_134_1941, w_134_1942, w_134_1944, w_134_1948, w_134_1949, w_134_1950, w_134_1953, w_134_1954, w_134_1959, w_134_1961, w_134_1962, w_134_1964, w_134_1969, w_134_1973, w_134_1974, w_134_1976, w_134_1981, w_134_1982, w_134_1983, w_134_1986, w_134_1990, w_134_1997, w_134_1999, w_134_2000, w_134_2010, w_134_2013, w_134_2019, w_134_2022, w_134_2026, w_134_2029, w_134_2036, w_134_2038, w_134_2041, w_134_2042, w_134_2051, w_134_2056, w_134_2057, w_134_2058, w_134_2068, w_134_2074, w_134_2078, w_134_2085, w_134_2091, w_134_2092, w_134_2093, w_134_2094, w_134_2098, w_134_2099, w_134_2101, w_134_2102, w_134_2106, w_134_2110, w_134_2111, w_134_2114, w_134_2115, w_134_2116, w_134_2118, w_134_2119, w_134_2121, w_134_2123, w_134_2125, w_134_2129, w_134_2132, w_134_2137, w_134_2138, w_134_2141, w_134_2144, w_134_2157, w_134_2162, w_134_2163, w_134_2165, w_134_2169, w_134_2179, w_134_2180, w_134_2182, w_134_2188, w_134_2194, w_134_2195, w_134_2198, w_134_2201, w_134_2205, w_134_2208, w_134_2211, w_134_2214, w_134_2216, w_134_2222, w_134_2231, w_134_2233, w_134_2244, w_134_2245, w_134_2251, w_134_2255, w_134_2257, w_134_2262, w_134_2265, w_134_2267, w_134_2272, w_134_2274, w_134_2282, w_134_2293, w_134_2297, w_134_2298, w_134_2302, w_134_2309, w_134_2317, w_134_2319, w_134_2320, w_134_2322, w_134_2324, w_134_2327, w_134_2332, w_134_2335, w_134_2337, w_134_2343, w_134_2345, w_134_2346, w_134_2357, w_134_2366, w_134_2367, w_134_2383, w_134_2392, w_134_2394, w_134_2399, w_134_2401, w_134_2409, w_134_2410, w_134_2414, w_134_2417, w_134_2421, w_134_2430, w_134_2432, w_134_2433, w_134_2435, w_134_2438, w_134_2443, w_134_2446, w_134_2454, w_134_2460, w_134_2463, w_134_2464, w_134_2469, w_134_2480, w_134_2483, w_134_2485, w_134_2487, w_134_2490, w_134_2494, w_134_2504, w_134_2505, w_134_2508, w_134_2512, w_134_2513, w_134_2514, w_134_2515, w_134_2520, w_134_2521, w_134_2539, w_134_2541, w_134_2552, w_134_2562, w_134_2564, w_134_2588, w_134_2590, w_134_2607, w_134_2608, w_134_2609, w_134_2610, w_134_2611, w_134_2619, w_134_2629, w_134_2636, w_134_2637, w_134_2640, w_134_2645, w_134_2649, w_134_2652, w_134_2656, w_134_2660, w_134_2662, w_134_2666, w_134_2667, w_134_2669, w_134_2674, w_134_2675, w_134_2682, w_134_2683, w_134_2687, w_134_2689, w_134_2691, w_134_2692, w_134_2693, w_134_2695, w_134_2696, w_134_2697, w_134_2700, w_134_2703, w_134_2707, w_134_2708, w_134_2712, w_134_2715, w_134_2717, w_134_2720, w_134_2721, w_134_2722, w_134_2723, w_134_2763, w_134_2767, w_134_2768, w_134_2769, w_134_2771, w_134_2775, w_134_2780, w_134_2781, w_134_2782, w_134_2783, w_134_2784, w_134_2785, w_134_2786;
  wire w_135_001, w_135_005, w_135_009, w_135_011, w_135_013, w_135_018, w_135_021, w_135_025, w_135_027, w_135_028, w_135_029, w_135_032, w_135_035, w_135_037, w_135_041, w_135_042, w_135_043, w_135_044, w_135_048, w_135_050, w_135_057, w_135_058, w_135_061, w_135_063, w_135_069, w_135_070, w_135_071, w_135_072, w_135_074, w_135_086, w_135_091, w_135_093, w_135_097, w_135_098, w_135_101, w_135_102, w_135_106, w_135_108, w_135_112, w_135_117, w_135_119, w_135_127, w_135_128, w_135_129, w_135_132, w_135_138, w_135_139, w_135_140, w_135_143, w_135_144, w_135_146, w_135_147, w_135_154, w_135_157, w_135_158, w_135_159, w_135_160, w_135_162, w_135_165, w_135_169, w_135_172, w_135_174, w_135_175, w_135_177, w_135_185, w_135_187, w_135_188, w_135_190, w_135_191, w_135_192, w_135_193, w_135_197, w_135_198, w_135_204, w_135_206, w_135_207, w_135_209, w_135_214, w_135_216, w_135_217, w_135_222, w_135_224, w_135_225, w_135_226, w_135_229, w_135_231, w_135_233, w_135_234, w_135_237, w_135_240, w_135_249, w_135_252, w_135_253, w_135_254, w_135_255, w_135_262, w_135_268, w_135_271, w_135_274, w_135_275, w_135_276, w_135_279, w_135_281, w_135_288, w_135_289, w_135_292, w_135_294, w_135_295, w_135_299, w_135_301, w_135_302, w_135_307, w_135_310, w_135_311, w_135_312, w_135_315, w_135_325, w_135_326, w_135_330, w_135_334, w_135_342, w_135_343, w_135_344, w_135_351, w_135_353, w_135_354, w_135_357, w_135_359, w_135_360, w_135_361, w_135_362, w_135_367, w_135_368, w_135_369, w_135_370, w_135_373, w_135_374, w_135_376, w_135_377, w_135_379, w_135_393, w_135_397, w_135_398, w_135_400, w_135_401, w_135_410, w_135_412, w_135_416, w_135_418, w_135_420, w_135_422, w_135_432, w_135_437, w_135_438, w_135_440, w_135_445, w_135_448, w_135_457, w_135_459, w_135_461, w_135_462, w_135_464, w_135_466, w_135_467, w_135_468, w_135_474, w_135_475, w_135_476, w_135_486, w_135_488, w_135_489, w_135_491, w_135_497, w_135_498, w_135_506, w_135_508, w_135_514, w_135_524, w_135_526, w_135_527, w_135_530, w_135_531, w_135_538, w_135_542, w_135_548, w_135_550, w_135_554, w_135_556, w_135_558, w_135_559, w_135_560, w_135_563, w_135_565, w_135_566, w_135_567, w_135_573, w_135_580, w_135_583, w_135_584, w_135_587, w_135_589, w_135_592, w_135_595, w_135_599, w_135_601, w_135_603, w_135_605, w_135_609, w_135_611, w_135_612, w_135_613, w_135_617, w_135_619, w_135_624, w_135_626, w_135_627, w_135_628, w_135_633, w_135_635, w_135_644, w_135_646, w_135_647, w_135_650, w_135_651, w_135_653, w_135_657, w_135_660, w_135_661, w_135_666, w_135_668, w_135_675, w_135_681, w_135_683, w_135_685, w_135_688, w_135_691, w_135_692, w_135_694, w_135_696, w_135_697, w_135_699, w_135_704, w_135_707, w_135_710, w_135_711, w_135_712, w_135_714, w_135_715, w_135_716, w_135_722, w_135_726, w_135_729, w_135_730, w_135_731, w_135_736, w_135_751, w_135_752, w_135_753, w_135_757, w_135_763, w_135_766, w_135_769, w_135_770, w_135_771, w_135_773, w_135_775, w_135_780, w_135_781, w_135_785, w_135_787, w_135_789, w_135_791, w_135_792, w_135_800, w_135_805, w_135_806, w_135_810, w_135_811, w_135_815, w_135_819, w_135_820, w_135_821, w_135_824, w_135_827, w_135_828, w_135_831, w_135_832, w_135_834, w_135_835, w_135_838, w_135_842, w_135_847, w_135_849, w_135_850, w_135_851, w_135_853, w_135_855, w_135_859, w_135_860, w_135_862, w_135_867, w_135_875, w_135_876, w_135_877, w_135_878, w_135_881, w_135_882, w_135_884, w_135_888, w_135_890, w_135_892, w_135_895, w_135_896, w_135_898, w_135_899, w_135_900, w_135_904, w_135_907, w_135_909, w_135_913, w_135_915, w_135_917, w_135_919, w_135_924, w_135_925, w_135_928, w_135_931, w_135_932, w_135_934, w_135_937, w_135_940, w_135_941, w_135_945, w_135_947, w_135_948, w_135_949, w_135_966, w_135_969, w_135_971, w_135_975, w_135_976, w_135_980, w_135_983, w_135_984, w_135_987, w_135_988, w_135_989, w_135_993, w_135_994, w_135_998, w_135_1002, w_135_1005, w_135_1010, w_135_1015, w_135_1017, w_135_1019, w_135_1020, w_135_1022, w_135_1024, w_135_1025, w_135_1027, w_135_1030, w_135_1031, w_135_1038, w_135_1039, w_135_1043, w_135_1046, w_135_1050, w_135_1057, w_135_1063, w_135_1065, w_135_1067, w_135_1069, w_135_1071, w_135_1073, w_135_1074, w_135_1084, w_135_1089, w_135_1091, w_135_1095, w_135_1097, w_135_1101, w_135_1102, w_135_1103, w_135_1104, w_135_1106, w_135_1107, w_135_1108, w_135_1109, w_135_1110, w_135_1112, w_135_1113, w_135_1116, w_135_1119, w_135_1121, w_135_1125, w_135_1130, w_135_1133, w_135_1134, w_135_1137, w_135_1138, w_135_1139, w_135_1141, w_135_1143, w_135_1144, w_135_1147, w_135_1149, w_135_1150, w_135_1151, w_135_1153, w_135_1155, w_135_1157, w_135_1158, w_135_1160, w_135_1163, w_135_1164, w_135_1168, w_135_1169, w_135_1172, w_135_1176, w_135_1181, w_135_1182, w_135_1183, w_135_1184, w_135_1185, w_135_1186, w_135_1190, w_135_1191, w_135_1196, w_135_1198, w_135_1200, w_135_1201, w_135_1202, w_135_1203, w_135_1204, w_135_1206, w_135_1207, w_135_1210, w_135_1212, w_135_1215, w_135_1216, w_135_1217, w_135_1218, w_135_1221, w_135_1222, w_135_1224, w_135_1226, w_135_1228, w_135_1232, w_135_1237, w_135_1240, w_135_1242, w_135_1243, w_135_1248, w_135_1249, w_135_1250, w_135_1256, w_135_1258, w_135_1259, w_135_1261, w_135_1262, w_135_1267, w_135_1268, w_135_1271, w_135_1274, w_135_1277, w_135_1279, w_135_1281, w_135_1283, w_135_1285, w_135_1286, w_135_1290, w_135_1293, w_135_1299, w_135_1301, w_135_1303, w_135_1307, w_135_1309, w_135_1310, w_135_1313, w_135_1315, w_135_1316, w_135_1317, w_135_1324, w_135_1325, w_135_1328, w_135_1332, w_135_1334, w_135_1337, w_135_1339, w_135_1340, w_135_1341, w_135_1342, w_135_1344, w_135_1347, w_135_1348, w_135_1349, w_135_1354, w_135_1356, w_135_1358, w_135_1359, w_135_1364, w_135_1367, w_135_1371, w_135_1376, w_135_1379, w_135_1380, w_135_1381, w_135_1383, w_135_1391, w_135_1392, w_135_1394, w_135_1395, w_135_1396, w_135_1397, w_135_1399, w_135_1400, w_135_1402, w_135_1404, w_135_1407, w_135_1410, w_135_1412, w_135_1414, w_135_1415, w_135_1425, w_135_1428, w_135_1431, w_135_1434, w_135_1437, w_135_1441, w_135_1444, w_135_1445, w_135_1447, w_135_1448, w_135_1450, w_135_1457, w_135_1459, w_135_1461, w_135_1462, w_135_1463, w_135_1467, w_135_1470, w_135_1471, w_135_1474, w_135_1475, w_135_1477, w_135_1479, w_135_1480, w_135_1485, w_135_1488, w_135_1492, w_135_1493, w_135_1494, w_135_1497, w_135_1500, w_135_1504, w_135_1506, w_135_1508, w_135_1509, w_135_1510, w_135_1512, w_135_1515, w_135_1521, w_135_1524, w_135_1527, w_135_1530, w_135_1533, w_135_1535, w_135_1539, w_135_1542, w_135_1544, w_135_1545, w_135_1547, w_135_1548, w_135_1554, w_135_1555, w_135_1559, w_135_1562, w_135_1563, w_135_1564, w_135_1566, w_135_1569, w_135_1572, w_135_1576, w_135_1577, w_135_1582, w_135_1583, w_135_1584, w_135_1588, w_135_1593, w_135_1594, w_135_1599, w_135_1602, w_135_1604, w_135_1605, w_135_1606, w_135_1610, w_135_1613, w_135_1614, w_135_1617, w_135_1624, w_135_1629, w_135_1631, w_135_1632, w_135_1634, w_135_1636, w_135_1638, w_135_1641, w_135_1645, w_135_1647, w_135_1651, w_135_1653, w_135_1655, w_135_1657, w_135_1659, w_135_1660, w_135_1661, w_135_1662, w_135_1666, w_135_1668, w_135_1671, w_135_1672, w_135_1673, w_135_1678, w_135_1686, w_135_1687, w_135_1689, w_135_1690, w_135_1695, w_135_1697, w_135_1701, w_135_1703, w_135_1704, w_135_1705, w_135_1706, w_135_1709, w_135_1711, w_135_1712, w_135_1713, w_135_1714, w_135_1716, w_135_1717, w_135_1721, w_135_1723, w_135_1724, w_135_1725, w_135_1726, w_135_1728, w_135_1731, w_135_1732, w_135_1733, w_135_1735, w_135_1737, w_135_1738, w_135_1745, w_135_1751, w_135_1752, w_135_1753, w_135_1754, w_135_1756, w_135_1757, w_135_1759, w_135_1761, w_135_1763, w_135_1764, w_135_1765, w_135_1773, w_135_1777, w_135_1778, w_135_1779, w_135_1781, w_135_1789, w_135_1793, w_135_1794, w_135_1797, w_135_1799, w_135_1801, w_135_1804, w_135_1806, w_135_1813, w_135_1815, w_135_1817, w_135_1818, w_135_1823, w_135_1824, w_135_1829, w_135_1839, w_135_1850, w_135_1856, w_135_1860, w_135_1861, w_135_1866, w_135_1870, w_135_1874, w_135_1875, w_135_1878, w_135_1883, w_135_1885, w_135_1890, w_135_1899, w_135_1901, w_135_1902, w_135_1903, w_135_1905, w_135_1908, w_135_1918, w_135_1933, w_135_1934, w_135_1940, w_135_1944, w_135_1945, w_135_1947, w_135_1948, w_135_1949, w_135_1950, w_135_1961, w_135_1965, w_135_1967, w_135_1969, w_135_1972, w_135_1983, w_135_1984, w_135_1987, w_135_1996, w_135_1998, w_135_2005, w_135_2008, w_135_2013, w_135_2030, w_135_2037, w_135_2040, w_135_2042, w_135_2055, w_135_2057, w_135_2059, w_135_2064, w_135_2072, w_135_2076, w_135_2078, w_135_2080, w_135_2086, w_135_2094, w_135_2098, w_135_2102, w_135_2105, w_135_2112, w_135_2113, w_135_2116, w_135_2119, w_135_2123, w_135_2127, w_135_2130, w_135_2137, w_135_2138, w_135_2139, w_135_2149, w_135_2155, w_135_2157, w_135_2165, w_135_2180, w_135_2184, w_135_2187, w_135_2190, w_135_2198, w_135_2205, w_135_2213, w_135_2220, w_135_2225, w_135_2229, w_135_2233, w_135_2236, w_135_2243, w_135_2247, w_135_2250, w_135_2254, w_135_2256, w_135_2267, w_135_2274, w_135_2275, w_135_2279, w_135_2287, w_135_2288, w_135_2289, w_135_2290, w_135_2297, w_135_2300, w_135_2307, w_135_2310, w_135_2321, w_135_2322, w_135_2328, w_135_2330, w_135_2340, w_135_2345, w_135_2346, w_135_2348, w_135_2352, w_135_2353, w_135_2356, w_135_2359, w_135_2361, w_135_2362, w_135_2363, w_135_2365, w_135_2376, w_135_2378, w_135_2388, w_135_2397, w_135_2400, w_135_2402, w_135_2406, w_135_2412, w_135_2416, w_135_2422, w_135_2425, w_135_2427, w_135_2436, w_135_2447, w_135_2452, w_135_2456, w_135_2465, w_135_2468, w_135_2473, w_135_2480, w_135_2482, w_135_2487, w_135_2494, w_135_2499, w_135_2502, w_135_2509, w_135_2510, w_135_2513, w_135_2519, w_135_2522, w_135_2532, w_135_2536, w_135_2538, w_135_2539, w_135_2541, w_135_2542, w_135_2545, w_135_2546, w_135_2553, w_135_2554, w_135_2559, w_135_2564, w_135_2569, w_135_2573, w_135_2578, w_135_2584, w_135_2594, w_135_2595, w_135_2596, w_135_2602, w_135_2604, w_135_2606, w_135_2627, w_135_2630, w_135_2635, w_135_2651, w_135_2658, w_135_2681, w_135_2683, w_135_2689, w_135_2695, w_135_2705, w_135_2707, w_135_2710, w_135_2711, w_135_2717, w_135_2722, w_135_2723, w_135_2732, w_135_2733, w_135_2735, w_135_2746, w_135_2748, w_135_2750, w_135_2764, w_135_2765, w_135_2768, w_135_2770, w_135_2774, w_135_2776, w_135_2782, w_135_2786, w_135_2789, w_135_2792, w_135_2794, w_135_2795, w_135_2800, w_135_2803, w_135_2806, w_135_2809, w_135_2811, w_135_2813, w_135_2815, w_135_2816, w_135_2838, w_135_2840, w_135_2843, w_135_2848, w_135_2849, w_135_2868, w_135_2869, w_135_2872, w_135_2874, w_135_2876, w_135_2899, w_135_2912, w_135_2913, w_135_2914, w_135_2923, w_135_2927, w_135_2928, w_135_2936, w_135_2939, w_135_2942, w_135_2952, w_135_2953, w_135_2956, w_135_2957, w_135_2961, w_135_2970, w_135_2971, w_135_2974, w_135_2984, w_135_2985, w_135_2996, w_135_3006, w_135_3013, w_135_3026, w_135_3030, w_135_3035, w_135_3038, w_135_3048, w_135_3052, w_135_3056, w_135_3058, w_135_3074, w_135_3082, w_135_3086, w_135_3088, w_135_3093, w_135_3102, w_135_3105, w_135_3123, w_135_3131, w_135_3142, w_135_3143, w_135_3145, w_135_3151, w_135_3156, w_135_3159, w_135_3160, w_135_3163, w_135_3164, w_135_3166, w_135_3170, w_135_3173, w_135_3176, w_135_3178, w_135_3184, w_135_3187, w_135_3191, w_135_3192, w_135_3193, w_135_3197, w_135_3198, w_135_3199, w_135_3200, w_135_3201, w_135_3202, w_135_3203, w_135_3204, w_135_3205, w_135_3206, w_135_3207, w_135_3209;
  wire w_136_001, w_136_002, w_136_003, w_136_004, w_136_005, w_136_009, w_136_010, w_136_011, w_136_012, w_136_014, w_136_017, w_136_021, w_136_022, w_136_023, w_136_024, w_136_029, w_136_030, w_136_032, w_136_033, w_136_035, w_136_037, w_136_038, w_136_039, w_136_041, w_136_044, w_136_046, w_136_047, w_136_048, w_136_049, w_136_050, w_136_052, w_136_054, w_136_058, w_136_059, w_136_060, w_136_062, w_136_063, w_136_067, w_136_069, w_136_072, w_136_073, w_136_078, w_136_079, w_136_083, w_136_086, w_136_088, w_136_090, w_136_091, w_136_093, w_136_095, w_136_098, w_136_100, w_136_101, w_136_103, w_136_104, w_136_106, w_136_108, w_136_110, w_136_111, w_136_112, w_136_113, w_136_117, w_136_119, w_136_121, w_136_123, w_136_126, w_136_127, w_136_128, w_136_130, w_136_133, w_136_134, w_136_139, w_136_140, w_136_141, w_136_142, w_136_143, w_136_149, w_136_152, w_136_153, w_136_154, w_136_156, w_136_157, w_136_158, w_136_159, w_136_161, w_136_162, w_136_163, w_136_164, w_136_165, w_136_166, w_136_167, w_136_168, w_136_169, w_136_170, w_136_172, w_136_175, w_136_177, w_136_182, w_136_183, w_136_184, w_136_185, w_136_186, w_136_187, w_136_191, w_136_193, w_136_198, w_136_202, w_136_203, w_136_209, w_136_210, w_136_213, w_136_214, w_136_218, w_136_220, w_136_221, w_136_222, w_136_224, w_136_228, w_136_231, w_136_234, w_136_237, w_136_240, w_136_242, w_136_243, w_136_244, w_136_246, w_136_247, w_136_250, w_136_252, w_136_253, w_136_254, w_136_257, w_136_258, w_136_260, w_136_262, w_136_265, w_136_266, w_136_267, w_136_268, w_136_271, w_136_272, w_136_275, w_136_276, w_136_277, w_136_278, w_136_283, w_136_287, w_136_290, w_136_292, w_136_295, w_136_297, w_136_298, w_136_299, w_136_302, w_136_303, w_136_305, w_136_307, w_136_312, w_136_317, w_136_318, w_136_319, w_136_322, w_136_330, w_136_334, w_136_335, w_136_336, w_136_337, w_136_338, w_136_340, w_136_341, w_136_342, w_136_343, w_136_344, w_136_346, w_136_348, w_136_352, w_136_356, w_136_362, w_136_366, w_136_367, w_136_369, w_136_370, w_136_372, w_136_376, w_136_384, w_136_392, w_136_393, w_136_394, w_136_397, w_136_398, w_136_399, w_136_400, w_136_401, w_136_404, w_136_405, w_136_408, w_136_414, w_136_417, w_136_419, w_136_421, w_136_427, w_136_428, w_136_432, w_136_435, w_136_437, w_136_438, w_136_447, w_136_449, w_136_460, w_136_461, w_136_466, w_136_468, w_136_473, w_136_474, w_136_476, w_136_477, w_136_478, w_136_480, w_136_481, w_136_482, w_136_488, w_136_490, w_136_496, w_136_497, w_136_498, w_136_503, w_136_507, w_136_509, w_136_512, w_136_515, w_136_516, w_136_518, w_136_519, w_136_525, w_136_531, w_136_532, w_136_537, w_136_542, w_136_546, w_136_549, w_136_552, w_136_553, w_136_555, w_136_556, w_136_560, w_136_561, w_136_565, w_136_566, w_136_570, w_136_572, w_136_581, w_136_585, w_136_587, w_136_593, w_136_595, w_136_599, w_136_602, w_136_603, w_136_606, w_136_609, w_136_610, w_136_613, w_136_615, w_136_616, w_136_618, w_136_620, w_136_622, w_136_623, w_136_624, w_136_625, w_136_627, w_136_628, w_136_632, w_136_633, w_136_637, w_136_638, w_136_639, w_136_640, w_136_643, w_136_647, w_136_650, w_136_651, w_136_652, w_136_653, w_136_658, w_136_659, w_136_662, w_136_665, w_136_666, w_136_672, w_136_675, w_136_677, w_136_680, w_136_681, w_136_682, w_136_683, w_136_684, w_136_687, w_136_688, w_136_691, w_136_696, w_136_697, w_136_699, w_136_701, w_136_702, w_136_705, w_136_706, w_136_708, w_136_709, w_136_710, w_136_713, w_136_716, w_136_717, w_136_722, w_136_723, w_136_726, w_136_727, w_136_733, w_136_734, w_136_739, w_136_745, w_136_747, w_136_750, w_136_751, w_136_752, w_136_754, w_136_762, w_136_763, w_136_764, w_136_765, w_136_769, w_136_771, w_136_779, w_136_780, w_136_781, w_136_784, w_136_785, w_136_787, w_136_795, w_136_796, w_136_802, w_136_803, w_136_813, w_136_814, w_136_816, w_136_817, w_136_819, w_136_823, w_136_829, w_136_830, w_136_841, w_136_845, w_136_853, w_136_854, w_136_855, w_136_856, w_136_859, w_136_865, w_136_866, w_136_870, w_136_873, w_136_875, w_136_877, w_136_878, w_136_881, w_136_882, w_136_886, w_136_887, w_136_895, w_136_899, w_136_901, w_136_910, w_136_912, w_136_916, w_136_918, w_136_920, w_136_928, w_136_931, w_136_932, w_136_935, w_136_938, w_136_939, w_136_945, w_136_946, w_136_949, w_136_952, w_136_959, w_136_963, w_136_966, w_136_968, w_136_972, w_136_973, w_136_975, w_136_976, w_136_980, w_136_981, w_136_983, w_136_988, w_136_990, w_136_996, w_136_997, w_136_998, w_136_1000, w_136_1001, w_136_1002, w_136_1006, w_136_1007, w_136_1010, w_136_1012, w_136_1013, w_136_1017, w_136_1018, w_136_1023, w_136_1025, w_136_1027, w_136_1029, w_136_1031, w_136_1035, w_136_1040, w_136_1048, w_136_1050, w_136_1055, w_136_1056, w_136_1057, w_136_1059, w_136_1061, w_136_1062, w_136_1063, w_136_1065, w_136_1071, w_136_1074, w_136_1077, w_136_1078, w_136_1080, w_136_1082, w_136_1087, w_136_1090, w_136_1092, w_136_1093, w_136_1094, w_136_1095, w_136_1103, w_136_1109, w_136_1110, w_136_1116, w_136_1118, w_136_1119, w_136_1121, w_136_1122, w_136_1124, w_136_1129, w_136_1130, w_136_1133, w_136_1141, w_136_1144, w_136_1145, w_136_1149, w_136_1156, w_136_1159, w_136_1161, w_136_1165, w_136_1166, w_136_1168, w_136_1170, w_136_1172, w_136_1177, w_136_1178, w_136_1183, w_136_1187, w_136_1197, w_136_1199, w_136_1201, w_136_1202, w_136_1204, w_136_1205, w_136_1206, w_136_1207, w_136_1209, w_136_1217, w_136_1218, w_136_1221, w_136_1222, w_136_1223, w_136_1234, w_136_1235, w_136_1237, w_136_1239, w_136_1241, w_136_1242, w_136_1250, w_136_1257, w_136_1260, w_136_1261, w_136_1262, w_136_1263, w_136_1265, w_136_1273, w_136_1275, w_136_1277, w_136_1281, w_136_1289, w_136_1294, w_136_1297, w_136_1304, w_136_1305, w_136_1307, w_136_1308, w_136_1309, w_136_1311, w_136_1313, w_136_1318, w_136_1319, w_136_1320, w_136_1321, w_136_1327, w_136_1329, w_136_1333, w_136_1334, w_136_1341, w_136_1344, w_136_1348, w_136_1351, w_136_1354, w_136_1359, w_136_1370, w_136_1372, w_136_1374, w_136_1376, w_136_1377, w_136_1381, w_136_1382, w_136_1385, w_136_1386, w_136_1389, w_136_1390, w_136_1392, w_136_1396, w_136_1402, w_136_1403, w_136_1404, w_136_1406, w_136_1410, w_136_1413, w_136_1417, w_136_1419, w_136_1420, w_136_1423, w_136_1427, w_136_1434, w_136_1435, w_136_1436, w_136_1441, w_136_1442, w_136_1444, w_136_1448, w_136_1449, w_136_1451, w_136_1453, w_136_1455, w_136_1457, w_136_1460, w_136_1466, w_136_1467, w_136_1468, w_136_1469, w_136_1477, w_136_1478, w_136_1480, w_136_1485, w_136_1486, w_136_1487, w_136_1488, w_136_1493, w_136_1496, w_136_1497, w_136_1498, w_136_1499, w_136_1503, w_136_1508, w_136_1510, w_136_1512, w_136_1514, w_136_1517, w_136_1525, w_136_1530, w_136_1531, w_136_1532, w_136_1533, w_136_1534, w_136_1535, w_136_1537, w_136_1538, w_136_1541, w_136_1555, w_136_1556, w_136_1557, w_136_1560, w_136_1563, w_136_1564, w_136_1565, w_136_1567, w_136_1571, w_136_1574, w_136_1580, w_136_1582, w_136_1585, w_136_1591, w_136_1592, w_136_1594, w_136_1596, w_136_1601, w_136_1604, w_136_1617, w_136_1618, w_136_1619, w_136_1620, w_136_1622, w_136_1625, w_136_1626, w_136_1628, w_136_1629, w_136_1635, w_136_1636, w_136_1637, w_136_1642, w_136_1644, w_136_1646, w_136_1649, w_136_1655, w_136_1660, w_136_1661, w_136_1662, w_136_1664, w_136_1666, w_136_1669, w_136_1671, w_136_1672, w_136_1678, w_136_1681, w_136_1686, w_136_1695, w_136_1698, w_136_1713, w_136_1716, w_136_1717, w_136_1723, w_136_1724, w_136_1727, w_136_1731, w_136_1732, w_136_1734, w_136_1736, w_136_1745, w_136_1746, w_136_1747, w_136_1748, w_136_1749, w_136_1751, w_136_1753, w_136_1756, w_136_1757, w_136_1758, w_136_1759, w_136_1762, w_136_1763, w_136_1768, w_136_1769, w_136_1771, w_136_1775, w_136_1776, w_136_1782, w_136_1785, w_136_1787, w_136_1788, w_136_1789, w_136_1791, w_136_1792, w_136_1793, w_136_1794, w_136_1799, w_136_1801, w_136_1804, w_136_1805, w_136_1807, w_136_1808, w_136_1809, w_136_1811, w_136_1813, w_136_1816, w_136_1818, w_136_1822, w_136_1824, w_136_1828, w_136_1831, w_136_1833, w_136_1834, w_136_1836, w_136_1837, w_136_1838, w_136_1839, w_136_1851, w_136_1852, w_136_1853, w_136_1855, w_136_1863, w_136_1866, w_136_1869, w_136_1882, w_136_1883, w_136_1888, w_136_1894, w_136_1895, w_136_1901, w_136_1902, w_136_1906, w_136_1910, w_136_1918, w_136_1919, w_136_1920, w_136_1924, w_136_1926, w_136_1929, w_136_1932, w_136_1935, w_136_1942, w_136_1945, w_136_1948, w_136_1949, w_136_1951, w_136_1952, w_136_1953, w_136_1954, w_136_1959, w_136_1960, w_136_1968, w_136_1969, w_136_1979, w_136_1981, w_136_1983, w_136_1984, w_136_1987, w_136_1990, w_136_1993, w_136_1995, w_136_1996, w_136_1997, w_136_1999, w_136_2003, w_136_2009, w_136_2021, w_136_2030, w_136_2035, w_136_2039, w_136_2043, w_136_2051, w_136_2054, w_136_2055, w_136_2058, w_136_2059, w_136_2060, w_136_2065, w_136_2067, w_136_2069, w_136_2075, w_136_2079, w_136_2081, w_136_2083, w_136_2084, w_136_2085, w_136_2087, w_136_2089, w_136_2091, w_136_2092, w_136_2095, w_136_2097, w_136_2100, w_136_2104, w_136_2107, w_136_2111, w_136_2114, w_136_2116, w_136_2118, w_136_2120, w_136_2122, w_136_2123, w_136_2126, w_136_2127, w_136_2132, w_136_2133, w_136_2134, w_136_2138, w_136_2139, w_136_2143, w_136_2144, w_136_2146, w_136_2148, w_136_2150, w_136_2153, w_136_2155, w_136_2159, w_136_2165, w_136_2167, w_136_2168, w_136_2172, w_136_2174, w_136_2175, w_136_2177, w_136_2180, w_136_2181, w_136_2183, w_136_2188, w_136_2190, w_136_2191, w_136_2194, w_136_2197, w_136_2199, w_136_2201, w_136_2203, w_136_2204, w_136_2205, w_136_2208, w_136_2212, w_136_2213, w_136_2217, w_136_2218, w_136_2219, w_136_2222, w_136_2223, w_136_2226, w_136_2232, w_136_2234, w_136_2240, w_136_2242, w_136_2243, w_136_2249, w_136_2251, w_136_2253, w_136_2256, w_136_2259, w_136_2263, w_136_2272, w_136_2273, w_136_2274, w_136_2279, w_136_2280, w_136_2281, w_136_2285, w_136_2287, w_136_2292, w_136_2294, w_136_2296, w_136_2299, w_136_2300, w_136_2301, w_136_2309, w_136_2310, w_136_2311, w_136_2312, w_136_2318, w_136_2319, w_136_2324, w_136_2325, w_136_2326, w_136_2327, w_136_2330, w_136_2331, w_136_2332, w_136_2333, w_136_2334, w_136_2337;
  wire w_137_002, w_137_007, w_137_008, w_137_009, w_137_019, w_137_020, w_137_021, w_137_026, w_137_029, w_137_030, w_137_031, w_137_032, w_137_033, w_137_036, w_137_039, w_137_047, w_137_049, w_137_053, w_137_054, w_137_055, w_137_056, w_137_064, w_137_066, w_137_071, w_137_073, w_137_078, w_137_087, w_137_092, w_137_097, w_137_106, w_137_107, w_137_110, w_137_114, w_137_124, w_137_125, w_137_133, w_137_134, w_137_142, w_137_145, w_137_149, w_137_151, w_137_153, w_137_160, w_137_161, w_137_163, w_137_164, w_137_165, w_137_169, w_137_170, w_137_176, w_137_178, w_137_179, w_137_181, w_137_184, w_137_185, w_137_186, w_137_187, w_137_188, w_137_189, w_137_191, w_137_199, w_137_201, w_137_206, w_137_208, w_137_212, w_137_221, w_137_222, w_137_225, w_137_227, w_137_228, w_137_229, w_137_230, w_137_233, w_137_240, w_137_241, w_137_243, w_137_250, w_137_253, w_137_257, w_137_260, w_137_262, w_137_263, w_137_265, w_137_268, w_137_270, w_137_272, w_137_273, w_137_274, w_137_280, w_137_288, w_137_302, w_137_312, w_137_313, w_137_320, w_137_322, w_137_325, w_137_327, w_137_328, w_137_329, w_137_332, w_137_336, w_137_337, w_137_339, w_137_341, w_137_343, w_137_344, w_137_347, w_137_353, w_137_354, w_137_362, w_137_367, w_137_368, w_137_375, w_137_382, w_137_384, w_137_385, w_137_392, w_137_393, w_137_401, w_137_403, w_137_406, w_137_409, w_137_410, w_137_419, w_137_434, w_137_436, w_137_450, w_137_452, w_137_458, w_137_464, w_137_476, w_137_491, w_137_496, w_137_497, w_137_501, w_137_510, w_137_514, w_137_516, w_137_520, w_137_532, w_137_533, w_137_534, w_137_538, w_137_542, w_137_544, w_137_546, w_137_557, w_137_558, w_137_562, w_137_566, w_137_572, w_137_576, w_137_579, w_137_600, w_137_605, w_137_612, w_137_623, w_137_630, w_137_637, w_137_640, w_137_644, w_137_651, w_137_659, w_137_660, w_137_666, w_137_668, w_137_669, w_137_670, w_137_672, w_137_680, w_137_684, w_137_686, w_137_697, w_137_711, w_137_726, w_137_731, w_137_735, w_137_739, w_137_746, w_137_748, w_137_752, w_137_763, w_137_767, w_137_769, w_137_771, w_137_778, w_137_782, w_137_789, w_137_793, w_137_794, w_137_795, w_137_802, w_137_804, w_137_805, w_137_807, w_137_814, w_137_816, w_137_827, w_137_833, w_137_841, w_137_844, w_137_850, w_137_851, w_137_855, w_137_857, w_137_858, w_137_859, w_137_872, w_137_880, w_137_882, w_137_883, w_137_886, w_137_887, w_137_889, w_137_890, w_137_923, w_137_930, w_137_936, w_137_943, w_137_946, w_137_953, w_137_967, w_137_968, w_137_973, w_137_974, w_137_979, w_137_987, w_137_998, w_137_1013, w_137_1015, w_137_1016, w_137_1019, w_137_1030, w_137_1036, w_137_1037, w_137_1043, w_137_1053, w_137_1064, w_137_1066, w_137_1073, w_137_1076, w_137_1080, w_137_1081, w_137_1082, w_137_1086, w_137_1093, w_137_1104, w_137_1106, w_137_1110, w_137_1114, w_137_1115, w_137_1123, w_137_1129, w_137_1132, w_137_1133, w_137_1136, w_137_1138, w_137_1162, w_137_1165, w_137_1173, w_137_1175, w_137_1184, w_137_1186, w_137_1187, w_137_1195, w_137_1198, w_137_1199, w_137_1217, w_137_1223, w_137_1227, w_137_1232, w_137_1234, w_137_1240, w_137_1242, w_137_1248, w_137_1252, w_137_1260, w_137_1271, w_137_1275, w_137_1278, w_137_1294, w_137_1313, w_137_1324, w_137_1331, w_137_1333, w_137_1336, w_137_1337, w_137_1341, w_137_1344, w_137_1356, w_137_1360, w_137_1366, w_137_1367, w_137_1369, w_137_1382, w_137_1385, w_137_1392, w_137_1396, w_137_1400, w_137_1407, w_137_1408, w_137_1414, w_137_1416, w_137_1420, w_137_1438, w_137_1440, w_137_1442, w_137_1448, w_137_1450, w_137_1453, w_137_1457, w_137_1459, w_137_1460, w_137_1464, w_137_1465, w_137_1466, w_137_1468, w_137_1476, w_137_1482, w_137_1483, w_137_1496, w_137_1501, w_137_1511, w_137_1517, w_137_1527, w_137_1549, w_137_1552, w_137_1558, w_137_1562, w_137_1564, w_137_1572, w_137_1582, w_137_1590, w_137_1593, w_137_1597, w_137_1599, w_137_1600, w_137_1605, w_137_1611, w_137_1637, w_137_1641, w_137_1649, w_137_1650, w_137_1656, w_137_1664, w_137_1678, w_137_1681, w_137_1683, w_137_1685, w_137_1689, w_137_1692, w_137_1693, w_137_1700, w_137_1702, w_137_1703, w_137_1704, w_137_1711, w_137_1713, w_137_1716, w_137_1723, w_137_1724, w_137_1727, w_137_1732, w_137_1748, w_137_1764, w_137_1768, w_137_1789, w_137_1791, w_137_1794, w_137_1797, w_137_1804, w_137_1805, w_137_1807, w_137_1815, w_137_1819, w_137_1829, w_137_1834, w_137_1842, w_137_1847, w_137_1857, w_137_1860, w_137_1861, w_137_1866, w_137_1871, w_137_1874, w_137_1878, w_137_1882, w_137_1896, w_137_1905, w_137_1917, w_137_1925, w_137_1931, w_137_1938, w_137_1945, w_137_1946, w_137_1948, w_137_1949, w_137_1950, w_137_1956, w_137_1960, w_137_1961, w_137_1969, w_137_1974, w_137_1984, w_137_1994, w_137_1997, w_137_1998, w_137_2007, w_137_2018, w_137_2031, w_137_2044, w_137_2053, w_137_2054, w_137_2057, w_137_2058, w_137_2067, w_137_2075, w_137_2096, w_137_2104, w_137_2106, w_137_2126, w_137_2134, w_137_2135, w_137_2136, w_137_2138, w_137_2141, w_137_2152, w_137_2155, w_137_2158, w_137_2161, w_137_2162, w_137_2168, w_137_2175, w_137_2186, w_137_2187, w_137_2191, w_137_2193, w_137_2199, w_137_2200, w_137_2202, w_137_2206, w_137_2225, w_137_2233, w_137_2236, w_137_2237, w_137_2239, w_137_2245, w_137_2264, w_137_2270, w_137_2271, w_137_2276, w_137_2283, w_137_2288, w_137_2290, w_137_2298, w_137_2299, w_137_2300, w_137_2305, w_137_2312, w_137_2317, w_137_2318, w_137_2320, w_137_2339, w_137_2343, w_137_2345, w_137_2346, w_137_2354, w_137_2355, w_137_2360, w_137_2362, w_137_2366, w_137_2367, w_137_2372, w_137_2374, w_137_2375, w_137_2377, w_137_2379, w_137_2381, w_137_2383, w_137_2387, w_137_2392, w_137_2397, w_137_2403, w_137_2405, w_137_2407, w_137_2412, w_137_2413, w_137_2419, w_137_2420, w_137_2428, w_137_2430, w_137_2431, w_137_2435, w_137_2436, w_137_2443, w_137_2444, w_137_2447, w_137_2460, w_137_2464, w_137_2470, w_137_2487, w_137_2488, w_137_2489, w_137_2491, w_137_2492, w_137_2504, w_137_2505, w_137_2506, w_137_2513, w_137_2516, w_137_2517, w_137_2530, w_137_2533, w_137_2534, w_137_2538, w_137_2541, w_137_2545, w_137_2549, w_137_2550, w_137_2551, w_137_2553, w_137_2571, w_137_2587, w_137_2590, w_137_2593, w_137_2598, w_137_2609, w_137_2610, w_137_2619, w_137_2628, w_137_2635, w_137_2637, w_137_2640, w_137_2647, w_137_2648, w_137_2649, w_137_2654, w_137_2658, w_137_2660, w_137_2661, w_137_2669, w_137_2672, w_137_2687, w_137_2689, w_137_2691, w_137_2692, w_137_2696, w_137_2703, w_137_2707, w_137_2714, w_137_2715, w_137_2722, w_137_2730, w_137_2761, w_137_2765, w_137_2778, w_137_2785, w_137_2786, w_137_2787, w_137_2790, w_137_2795, w_137_2804, w_137_2807, w_137_2815, w_137_2820, w_137_2829, w_137_2832, w_137_2834, w_137_2836, w_137_2837, w_137_2838, w_137_2842, w_137_2844, w_137_2849, w_137_2850, w_137_2853, w_137_2855, w_137_2856, w_137_2861, w_137_2873, w_137_2879, w_137_2883, w_137_2885, w_137_2888, w_137_2893, w_137_2895, w_137_2903, w_137_2915, w_137_2924, w_137_2929, w_137_2936, w_137_2938, w_137_2943, w_137_2952, w_137_2958, w_137_2974, w_137_2981, w_137_2990, w_137_2998, w_137_3016, w_137_3017, w_137_3025, w_137_3027, w_137_3035, w_137_3049, w_137_3050, w_137_3051, w_137_3056, w_137_3062, w_137_3071, w_137_3081, w_137_3082, w_137_3084, w_137_3085, w_137_3092, w_137_3105, w_137_3106, w_137_3107, w_137_3112, w_137_3118, w_137_3124, w_137_3125, w_137_3126, w_137_3149, w_137_3150, w_137_3152, w_137_3157, w_137_3163, w_137_3178, w_137_3182, w_137_3203, w_137_3211, w_137_3224, w_137_3230, w_137_3231, w_137_3236, w_137_3240, w_137_3244, w_137_3257, w_137_3260, w_137_3276, w_137_3290, w_137_3292, w_137_3296, w_137_3297, w_137_3299, w_137_3301, w_137_3307, w_137_3312, w_137_3324, w_137_3327, w_137_3335, w_137_3337, w_137_3341, w_137_3356, w_137_3357, w_137_3358, w_137_3362, w_137_3364, w_137_3366, w_137_3368, w_137_3384, w_137_3387, w_137_3388, w_137_3389, w_137_3390, w_137_3394, w_137_3408, w_137_3414, w_137_3423, w_137_3436, w_137_3441, w_137_3454, w_137_3469, w_137_3470, w_137_3484, w_137_3497, w_137_3503, w_137_3505, w_137_3507, w_137_3508, w_137_3509, w_137_3513, w_137_3514, w_137_3515, w_137_3518, w_137_3519, w_137_3520, w_137_3528, w_137_3532, w_137_3540, w_137_3544, w_137_3545, w_137_3549, w_137_3552, w_137_3554, w_137_3558, w_137_3564, w_137_3575, w_137_3583, w_137_3590, w_137_3591, w_137_3594, w_137_3596, w_137_3599, w_137_3602, w_137_3604, w_137_3606, w_137_3622, w_137_3623, w_137_3628, w_137_3632, w_137_3637, w_137_3639, w_137_3645, w_137_3650, w_137_3653, w_137_3656, w_137_3662, w_137_3669, w_137_3680, w_137_3688, w_137_3692, w_137_3700, w_137_3702, w_137_3707, w_137_3714, w_137_3719, w_137_3722, w_137_3725, w_137_3727, w_137_3734, w_137_3736, w_137_3741, w_137_3750, w_137_3759, w_137_3765, w_137_3771, w_137_3773, w_137_3775, w_137_3779, w_137_3782, w_137_3786, w_137_3790, w_137_3796, w_137_3799, w_137_3801, w_137_3802, w_137_3804, w_137_3805, w_137_3809, w_137_3817, w_137_3832, w_137_3834, w_137_3835, w_137_3836, w_137_3841, w_137_3850, w_137_3851, w_137_3859, w_137_3867, w_137_3869, w_137_3872, w_137_3879, w_137_3882, w_137_3901, w_137_3906, w_137_3907, w_137_3918, w_137_3924, w_137_3927, w_137_3936, w_137_3948, w_137_3966, w_137_3969, w_137_3972, w_137_3974, w_137_3975, w_137_3978, w_137_3979, w_137_3983, w_137_3989, w_137_3991, w_137_3993, w_137_3995, w_137_3997, w_137_4004, w_137_4005, w_137_4006, w_137_4008, w_137_4015, w_137_4021, w_137_4025, w_137_4027, w_137_4028, w_137_4031, w_137_4037, w_137_4038, w_137_4056, w_137_4062, w_137_4071, w_137_4073, w_137_4076, w_137_4079, w_137_4096, w_137_4106, w_137_4109, w_137_4113, w_137_4149, w_137_4151, w_137_4154, w_137_4160, w_137_4169, w_137_4174, w_137_4177, w_137_4185, w_137_4187, w_137_4188, w_137_4193, w_137_4198, w_137_4199, w_137_4200, w_137_4217, w_137_4220, w_137_4225, w_137_4226, w_137_4229, w_137_4231, w_137_4237, w_137_4240, w_137_4247, w_137_4260, w_137_4262, w_137_4268, w_137_4279, w_137_4281, w_137_4289, w_137_4291, w_137_4297, w_137_4301, w_137_4303, w_137_4313, w_137_4314, w_137_4318, w_137_4327, w_137_4338, w_137_4353, w_137_4360, w_137_4361, w_137_4365, w_137_4366, w_137_4370, w_137_4374, w_137_4379, w_137_4382, w_137_4383, w_137_4392, w_137_4393, w_137_4396, w_137_4407, w_137_4414, w_137_4417, w_137_4421, w_137_4422, w_137_4425, w_137_4428, w_137_4433, w_137_4443, w_137_4446, w_137_4447, w_137_4448, w_137_4454, w_137_4456, w_137_4458, w_137_4463, w_137_4467, w_137_4473, w_137_4485, w_137_4492, w_137_4495, w_137_4496, w_137_4497, w_137_4500, w_137_4501, w_137_4503, w_137_4506, w_137_4508, w_137_4509, w_137_4517, w_137_4520, w_137_4521, w_137_4525, w_137_4530, w_137_4533, w_137_4536, w_137_4538, w_137_4542, w_137_4544, w_137_4545, w_137_4549, w_137_4555, w_137_4558, w_137_4564, w_137_4565, w_137_4566, w_137_4567, w_137_4572, w_137_4575, w_137_4576, w_137_4585, w_137_4588, w_137_4590, w_137_4600, w_137_4601, w_137_4606, w_137_4609, w_137_4622, w_137_4627, w_137_4634, w_137_4645, w_137_4646, w_137_4648, w_137_4651, w_137_4660, w_137_4661, w_137_4675, w_137_4684, w_137_4685, w_137_4696, w_137_4698, w_137_4701, w_137_4709, w_137_4716;
  wire w_138_000, w_138_001, w_138_002, w_138_003, w_138_004, w_138_005, w_138_009, w_138_010, w_138_012, w_138_014, w_138_015, w_138_016, w_138_017, w_138_018, w_138_019, w_138_020, w_138_021, w_138_022, w_138_023, w_138_026, w_138_027, w_138_030, w_138_033, w_138_035, w_138_036, w_138_038, w_138_039, w_138_040, w_138_043, w_138_044, w_138_046, w_138_047, w_138_048, w_138_050, w_138_052, w_138_053, w_138_057, w_138_058, w_138_059, w_138_060, w_138_061, w_138_062, w_138_065, w_138_067, w_138_068, w_138_069, w_138_070, w_138_072, w_138_075, w_138_077, w_138_079, w_138_081, w_138_082, w_138_083, w_138_085, w_138_086, w_138_092, w_138_093, w_138_096, w_138_098, w_138_099, w_138_100, w_138_101, w_138_103, w_138_104, w_138_105, w_138_106, w_138_107, w_138_109, w_138_110, w_138_111, w_138_112, w_138_114, w_138_115, w_138_116, w_138_118, w_138_125, w_138_126, w_138_130, w_138_133, w_138_134, w_138_136, w_138_137, w_138_141, w_138_142, w_138_143, w_138_144, w_138_145, w_138_146, w_138_148, w_138_151, w_138_153, w_138_154, w_138_155, w_138_156, w_138_157, w_138_160, w_138_161, w_138_162, w_138_163, w_138_167, w_138_173, w_138_174, w_138_176, w_138_177, w_138_180, w_138_181, w_138_182, w_138_183, w_138_185, w_138_190, w_138_192, w_138_193, w_138_194, w_138_195, w_138_197, w_138_198, w_138_199, w_138_200, w_138_201, w_138_204, w_138_205, w_138_206, w_138_210, w_138_211, w_138_212, w_138_216, w_138_218, w_138_219, w_138_221, w_138_222, w_138_223, w_138_224, w_138_227, w_138_228, w_138_229, w_138_231, w_138_236, w_138_239, w_138_240, w_138_241, w_138_242, w_138_244, w_138_245, w_138_246, w_138_248, w_138_249, w_138_250, w_138_251, w_138_253, w_138_254, w_138_255, w_138_256, w_138_257, w_138_258, w_138_259, w_138_261, w_138_263, w_138_265, w_138_266, w_138_267, w_138_268, w_138_270, w_138_271, w_138_272, w_138_273, w_138_274, w_138_276, w_138_277, w_138_278, w_138_279, w_138_280, w_138_281, w_138_283, w_138_284, w_138_286, w_138_287, w_138_288, w_138_289, w_138_290, w_138_294, w_138_295, w_138_297, w_138_301, w_138_302, w_138_303, w_138_304, w_138_305, w_138_309, w_138_311, w_138_313, w_138_314, w_138_315, w_138_316, w_138_317, w_138_318, w_138_319, w_138_320, w_138_321, w_138_323, w_138_324, w_138_325, w_138_326, w_138_327, w_138_328, w_138_329, w_138_331, w_138_334, w_138_336, w_138_337, w_138_339, w_138_340, w_138_344, w_138_345, w_138_346, w_138_347, w_138_348, w_138_350, w_138_351, w_138_355, w_138_356, w_138_357, w_138_359, w_138_360, w_138_361, w_138_362, w_138_364, w_138_366, w_138_368, w_138_370, w_138_371, w_138_372, w_138_374, w_138_376, w_138_380, w_138_381, w_138_382, w_138_384, w_138_385, w_138_386, w_138_387, w_138_389, w_138_390, w_138_391, w_138_393, w_138_394, w_138_395, w_138_397, w_138_398, w_138_400, w_138_401, w_138_405, w_138_407, w_138_413, w_138_414, w_138_415, w_138_416, w_138_417, w_138_418, w_138_419, w_138_420, w_138_423, w_138_425, w_138_427, w_138_428, w_138_429, w_138_430, w_138_431, w_138_432, w_138_433, w_138_434, w_138_437, w_138_438, w_138_441, w_138_442, w_138_443, w_138_444, w_138_446, w_138_448, w_138_449, w_138_450, w_138_451, w_138_454, w_138_455, w_138_456, w_138_458, w_138_459, w_138_462, w_138_463, w_138_464, w_138_466, w_138_467, w_138_468, w_138_470, w_138_471, w_138_475, w_138_476, w_138_477, w_138_479, w_138_480, w_138_481, w_138_482, w_138_483, w_138_485, w_138_486, w_138_487, w_138_489, w_138_490, w_138_492, w_138_494, w_138_495, w_138_496, w_138_497, w_138_500, w_138_501, w_138_505, w_138_507, w_138_508, w_138_512, w_138_513, w_138_514, w_138_515, w_138_519, w_138_520, w_138_526, w_138_528, w_138_531, w_138_533, w_138_534, w_138_535, w_138_536, w_138_537, w_138_540, w_138_542, w_138_544, w_138_546, w_138_549, w_138_550, w_138_552, w_138_554, w_138_557, w_138_559, w_138_562, w_138_564, w_138_567, w_138_568, w_138_570, w_138_571, w_138_572, w_138_573, w_138_575, w_138_578, w_138_579, w_138_580, w_138_583, w_138_585, w_138_586, w_138_588, w_138_589, w_138_590, w_138_591, w_138_594, w_138_595, w_138_596, w_138_597, w_138_598, w_138_599, w_138_600, w_138_601, w_138_603, w_138_604, w_138_605, w_138_606, w_138_608, w_138_611, w_138_614, w_138_615, w_138_616, w_138_617, w_138_618, w_138_623, w_138_624, w_138_625, w_138_626, w_138_633, w_138_636, w_138_637, w_138_638, w_138_640, w_138_641, w_138_642, w_138_644, w_138_646, w_138_647, w_138_648, w_138_649, w_138_650, w_138_651, w_138_653, w_138_655, w_138_656, w_138_658, w_138_660, w_138_662, w_138_664, w_138_666, w_138_668, w_138_669, w_138_671, w_138_676, w_138_678, w_138_679, w_138_680, w_138_681, w_138_682, w_138_683, w_138_690, w_138_692, w_138_693, w_138_696, w_138_700, w_138_701, w_138_703, w_138_704, w_138_705, w_138_708, w_138_709, w_138_710, w_138_713, w_138_714, w_138_715, w_138_722, w_138_724, w_138_726, w_138_727, w_138_730, w_138_734, w_138_735, w_138_739, w_138_740, w_138_741, w_138_742, w_138_744, w_138_745, w_138_746, w_138_747, w_138_748, w_138_749, w_138_750, w_138_753, w_138_754, w_138_756, w_138_757, w_138_758, w_138_760, w_138_761, w_138_762, w_138_763, w_138_764, w_138_766, w_138_767, w_138_773, w_138_774, w_138_775, w_138_776, w_138_779, w_138_780, w_138_781, w_138_782, w_138_783, w_138_785, w_138_786, w_138_787, w_138_789, w_138_790, w_138_792, w_138_793, w_138_796, w_138_797, w_138_800, w_138_802, w_138_805, w_138_806, w_138_808, w_138_809, w_138_812, w_138_813, w_138_814, w_138_815, w_138_816, w_138_817, w_138_818, w_138_820, w_138_821, w_138_822, w_138_826, w_138_827, w_138_829, w_138_830, w_138_832, w_138_833, w_138_834, w_138_835, w_138_836, w_138_838, w_138_840, w_138_842, w_138_843, w_138_846, w_138_847, w_138_848, w_138_850, w_138_851, w_138_852, w_138_853, w_138_854, w_138_855, w_138_862, w_138_864, w_138_865, w_138_868, w_138_871, w_138_873, w_138_876, w_138_877, w_138_878, w_138_879, w_138_880, w_138_881, w_138_882, w_138_885, w_138_886, w_138_890, w_138_891, w_138_893, w_138_895, w_138_898, w_138_902, w_138_905, w_138_906, w_138_907, w_138_908, w_138_909, w_138_910, w_138_911, w_138_913, w_138_914, w_138_916, w_138_918, w_138_919, w_138_920, w_138_922, w_138_924, w_138_926, w_138_929, w_138_930, w_138_932, w_138_933, w_138_934, w_138_935, w_138_936, w_138_937, w_138_938, w_138_939, w_138_940, w_138_941, w_138_946, w_138_947, w_138_948, w_138_950, w_138_951, w_138_953, w_138_954, w_138_957, w_138_958, w_138_961, w_138_962, w_138_966, w_138_972, w_138_975, w_138_976, w_138_978, w_138_980, w_138_981, w_138_982, w_138_983, w_138_984, w_138_985, w_138_988, w_138_989, w_138_990, w_138_992, w_138_993, w_138_994, w_138_996, w_138_1000, w_138_1001, w_138_1002, w_138_1003, w_138_1008, w_138_1014, w_138_1019, w_138_1020, w_138_1021, w_138_1022, w_138_1023, w_138_1025, w_138_1027, w_138_1028, w_138_1029, w_138_1030, w_138_1031, w_138_1032, w_138_1035, w_138_1036, w_138_1037, w_138_1038, w_138_1040, w_138_1042, w_138_1043, w_138_1045, w_138_1049, w_138_1052, w_138_1053, w_138_1054, w_138_1059, w_138_1060, w_138_1064, w_138_1065, w_138_1067, w_138_1068, w_138_1069, w_138_1070, w_138_1071, w_138_1074, w_138_1075, w_138_1076, w_138_1079, w_138_1080, w_138_1081, w_138_1083, w_138_1086, w_138_1088, w_138_1089, w_138_1092, w_138_1093, w_138_1094, w_138_1095, w_138_1096, w_138_1097, w_138_1099, w_138_1102, w_138_1106, w_138_1107, w_138_1108, w_138_1109, w_138_1110, w_138_1114, w_138_1115, w_138_1116, w_138_1117, w_138_1119, w_138_1120, w_138_1121, w_138_1124, w_138_1125, w_138_1130, w_138_1131, w_138_1132, w_138_1133, w_138_1134, w_138_1135, w_138_1136, w_138_1137, w_138_1140, w_138_1141, w_138_1142, w_138_1143, w_138_1144, w_138_1145, w_138_1147, w_138_1149, w_138_1153, w_138_1155, w_138_1156, w_138_1159, w_138_1160, w_138_1163, w_138_1164, w_138_1165, w_138_1166, w_138_1167, w_138_1168, w_138_1169, w_138_1171, w_138_1172, w_138_1173, w_138_1174, w_138_1175, w_138_1177, w_138_1180, w_138_1181, w_138_1182, w_138_1183, w_138_1184, w_138_1185, w_138_1186, w_138_1188, w_138_1189, w_138_1190, w_138_1191, w_138_1192, w_138_1194, w_138_1195, w_138_1202, w_138_1204, w_138_1209, w_138_1211, w_138_1213, w_138_1217, w_138_1219, w_138_1220, w_138_1222, w_138_1223, w_138_1225, w_138_1226, w_138_1229, w_138_1231, w_138_1232, w_138_1233, w_138_1234, w_138_1236, w_138_1237, w_138_1241, w_138_1242, w_138_1244, w_138_1247, w_138_1248, w_138_1250, w_138_1251, w_138_1253, w_138_1257, w_138_1258, w_138_1260, w_138_1262, w_138_1265;
  wire w_139_000, w_139_001, w_139_002, w_139_003, w_139_004, w_139_005, w_139_006, w_139_007, w_139_008, w_139_009, w_139_010, w_139_011, w_139_012, w_139_013, w_139_014, w_139_015, w_139_016, w_139_017, w_139_018, w_139_019, w_139_020, w_139_021, w_139_022, w_139_023, w_139_024, w_139_025, w_139_026, w_139_027, w_139_028, w_139_029, w_139_030, w_139_031, w_139_032, w_139_033, w_139_034, w_139_035, w_139_036, w_139_037, w_139_038, w_139_039, w_139_040, w_139_041, w_139_042, w_139_043, w_139_044, w_139_045, w_139_046, w_139_047, w_139_048, w_139_049, w_139_050, w_139_051, w_139_052, w_139_053, w_139_054, w_139_055, w_139_056, w_139_057, w_139_058, w_139_059, w_139_060, w_139_061, w_139_062, w_139_063, w_139_064, w_139_065, w_139_066, w_139_067, w_139_068, w_139_069, w_139_070, w_139_071, w_139_072, w_139_073, w_139_074, w_139_075, w_139_076, w_139_077, w_139_078, w_139_079, w_139_080, w_139_081, w_139_082, w_139_084, w_139_085, w_139_086, w_139_087, w_139_088, w_139_089, w_139_090, w_139_091, w_139_092, w_139_093, w_139_094, w_139_095, w_139_096, w_139_097, w_139_098, w_139_099, w_139_100, w_139_101, w_139_102, w_139_103, w_139_104, w_139_105, w_139_106, w_139_107, w_139_108, w_139_109, w_139_110, w_139_111, w_139_112, w_139_113, w_139_114, w_139_115, w_139_116, w_139_117, w_139_118, w_139_119, w_139_120, w_139_121, w_139_122, w_139_123, w_139_124, w_139_125, w_139_126, w_139_127, w_139_128, w_139_129, w_139_130, w_139_131, w_139_133, w_139_134, w_139_135, w_139_136, w_139_137, w_139_138, w_139_141, w_139_142, w_139_143, w_139_144, w_139_145, w_139_146, w_139_147, w_139_148, w_139_149, w_139_150, w_139_151, w_139_152, w_139_153, w_139_154, w_139_155, w_139_156, w_139_157, w_139_158, w_139_159, w_139_160, w_139_161, w_139_162, w_139_163, w_139_164, w_139_165, w_139_166, w_139_168, w_139_170, w_139_171, w_139_172, w_139_173, w_139_174, w_139_175, w_139_176, w_139_177, w_139_178, w_139_179, w_139_180, w_139_181, w_139_182, w_139_183, w_139_184, w_139_185, w_139_186, w_139_187, w_139_188, w_139_189, w_139_190, w_139_191, w_139_192, w_139_193, w_139_194, w_139_195, w_139_196, w_139_197, w_139_198, w_139_199, w_139_200, w_139_201, w_139_202, w_139_203, w_139_204, w_139_205, w_139_206, w_139_207, w_139_209, w_139_210, w_139_211, w_139_212, w_139_213, w_139_214, w_139_215, w_139_216, w_139_217, w_139_218, w_139_219, w_139_220, w_139_221, w_139_222, w_139_223, w_139_224, w_139_225, w_139_226, w_139_227, w_139_228, w_139_229, w_139_230, w_139_231, w_139_232, w_139_233, w_139_235, w_139_236, w_139_238, w_139_239, w_139_240, w_139_241, w_139_242, w_139_243, w_139_244, w_139_245, w_139_246, w_139_247, w_139_248, w_139_249, w_139_250, w_139_251, w_139_252, w_139_253, w_139_254, w_139_255, w_139_257, w_139_258, w_139_259, w_139_260, w_139_261, w_139_262, w_139_263, w_139_264, w_139_265, w_139_266, w_139_267, w_139_268, w_139_269, w_139_270, w_139_271, w_139_272, w_139_273, w_139_274, w_139_275, w_139_276, w_139_277, w_139_278, w_139_279, w_139_280, w_139_281, w_139_282, w_139_283, w_139_284, w_139_285, w_139_286, w_139_287, w_139_288, w_139_289, w_139_290, w_139_292, w_139_293, w_139_294, w_139_295, w_139_296, w_139_297, w_139_298, w_139_299, w_139_300, w_139_301, w_139_302, w_139_303, w_139_304, w_139_305, w_139_306, w_139_307, w_139_308, w_139_309, w_139_310, w_139_312, w_139_313, w_139_314, w_139_315, w_139_316;
  wire w_140_000, w_140_006, w_140_007, w_140_009, w_140_012, w_140_013, w_140_014, w_140_017, w_140_018, w_140_021, w_140_024, w_140_025, w_140_026, w_140_032, w_140_033, w_140_034, w_140_039, w_140_042, w_140_044, w_140_045, w_140_057, w_140_058, w_140_062, w_140_069, w_140_074, w_140_077, w_140_081, w_140_083, w_140_084, w_140_094, w_140_096, w_140_097, w_140_099, w_140_102, w_140_103, w_140_105, w_140_106, w_140_108, w_140_110, w_140_115, w_140_116, w_140_117, w_140_119, w_140_120, w_140_124, w_140_127, w_140_129, w_140_131, w_140_132, w_140_133, w_140_139, w_140_146, w_140_147, w_140_161, w_140_164, w_140_166, w_140_167, w_140_170, w_140_172, w_140_173, w_140_174, w_140_177, w_140_179, w_140_180, w_140_184, w_140_187, w_140_188, w_140_198, w_140_201, w_140_205, w_140_206, w_140_208, w_140_215, w_140_216, w_140_217, w_140_226, w_140_227, w_140_230, w_140_231, w_140_233, w_140_234, w_140_237, w_140_239, w_140_240, w_140_247, w_140_249, w_140_250, w_140_251, w_140_254, w_140_259, w_140_260, w_140_261, w_140_263, w_140_269, w_140_274, w_140_283, w_140_284, w_140_286, w_140_290, w_140_291, w_140_296, w_140_300, w_140_302, w_140_303, w_140_304, w_140_305, w_140_307, w_140_310, w_140_311, w_140_312, w_140_313, w_140_317, w_140_318, w_140_320, w_140_321, w_140_323, w_140_324, w_140_331, w_140_332, w_140_333, w_140_334, w_140_337, w_140_339, w_140_344, w_140_348, w_140_352, w_140_359, w_140_361, w_140_365, w_140_366, w_140_369, w_140_371, w_140_373, w_140_376, w_140_379, w_140_386, w_140_387, w_140_389, w_140_392, w_140_394, w_140_395, w_140_397, w_140_398, w_140_400, w_140_405, w_140_406, w_140_408, w_140_409, w_140_412, w_140_417, w_140_423, w_140_425, w_140_426, w_140_428, w_140_430, w_140_434, w_140_436, w_140_437, w_140_438, w_140_440, w_140_441, w_140_442, w_140_443, w_140_444, w_140_447, w_140_448, w_140_450, w_140_455, w_140_463, w_140_464, w_140_470, w_140_475, w_140_477, w_140_479, w_140_487, w_140_488, w_140_495, w_140_496, w_140_497, w_140_503, w_140_504, w_140_505, w_140_506, w_140_509, w_140_515, w_140_516, w_140_517, w_140_527, w_140_530, w_140_533, w_140_541, w_140_543, w_140_544, w_140_545, w_140_546, w_140_549, w_140_551, w_140_554, w_140_562, w_140_563, w_140_574, w_140_576, w_140_577, w_140_582, w_140_586, w_140_587, w_140_590, w_140_592, w_140_595, w_140_599, w_140_604, w_140_609, w_140_610, w_140_611, w_140_612, w_140_614, w_140_615, w_140_618, w_140_620, w_140_621, w_140_622, w_140_628, w_140_630, w_140_632, w_140_633, w_140_636, w_140_638, w_140_641, w_140_642, w_140_649, w_140_650, w_140_651, w_140_652, w_140_656, w_140_661, w_140_666, w_140_667, w_140_668, w_140_670, w_140_673, w_140_675, w_140_679, w_140_680, w_140_684, w_140_685, w_140_690, w_140_694, w_140_696, w_140_697, w_140_703, w_140_705, w_140_709, w_140_712, w_140_714, w_140_725, w_140_735, w_140_736, w_140_740, w_140_742, w_140_743, w_140_744, w_140_747, w_140_750, w_140_751, w_140_757, w_140_758, w_140_759, w_140_760, w_140_766, w_140_768, w_140_769, w_140_771, w_140_775, w_140_778, w_140_780, w_140_782, w_140_783, w_140_785, w_140_797, w_140_803, w_140_805, w_140_807, w_140_809, w_140_810, w_140_813, w_140_814, w_140_815, w_140_818, w_140_823, w_140_826, w_140_831, w_140_835, w_140_839, w_140_840, w_140_842, w_140_846, w_140_849, w_140_851, w_140_852, w_140_854, w_140_858, w_140_863, w_140_864, w_140_866, w_140_867, w_140_870, w_140_875, w_140_876, w_140_878, w_140_879, w_140_883, w_140_884, w_140_886, w_140_888, w_140_890, w_140_894, w_140_900, w_140_901, w_140_908, w_140_912, w_140_914, w_140_915, w_140_918, w_140_927, w_140_931, w_140_933, w_140_935, w_140_943, w_140_944, w_140_947, w_140_948, w_140_950, w_140_954, w_140_960, w_140_961, w_140_963, w_140_964, w_140_965, w_140_967, w_140_969, w_140_980, w_140_982, w_140_997, w_140_998, w_140_1000, w_140_1002, w_140_1003, w_140_1006, w_140_1010, w_140_1011, w_140_1013, w_140_1015, w_140_1016, w_140_1022, w_140_1023, w_140_1026, w_140_1029, w_140_1030, w_140_1031, w_140_1033, w_140_1036, w_140_1043, w_140_1044, w_140_1045, w_140_1048, w_140_1051, w_140_1058, w_140_1061, w_140_1065, w_140_1066, w_140_1073, w_140_1077, w_140_1079, w_140_1085, w_140_1089, w_140_1091, w_140_1096, w_140_1097, w_140_1099, w_140_1104, w_140_1108, w_140_1110, w_140_1114, w_140_1116, w_140_1118, w_140_1121, w_140_1123, w_140_1125, w_140_1130, w_140_1135, w_140_1137, w_140_1141, w_140_1142, w_140_1144, w_140_1146, w_140_1147, w_140_1149, w_140_1151, w_140_1152, w_140_1153, w_140_1154, w_140_1164, w_140_1165, w_140_1167, w_140_1169, w_140_1172, w_140_1176, w_140_1178, w_140_1181, w_140_1182, w_140_1189, w_140_1192, w_140_1194, w_140_1195, w_140_1196, w_140_1198, w_140_1201, w_140_1202, w_140_1204, w_140_1207, w_140_1209, w_140_1210, w_140_1211, w_140_1213, w_140_1214, w_140_1215, w_140_1216, w_140_1218, w_140_1227, w_140_1231, w_140_1233, w_140_1235, w_140_1238, w_140_1239, w_140_1240, w_140_1241, w_140_1247, w_140_1248, w_140_1250, w_140_1252, w_140_1256, w_140_1260, w_140_1262, w_140_1268, w_140_1277, w_140_1283, w_140_1284, w_140_1285, w_140_1286, w_140_1290, w_140_1297, w_140_1299, w_140_1306, w_140_1307, w_140_1310, w_140_1312, w_140_1313, w_140_1314, w_140_1316, w_140_1320, w_140_1324, w_140_1326, w_140_1328, w_140_1329, w_140_1332, w_140_1336, w_140_1339, w_140_1341, w_140_1343, w_140_1344, w_140_1345, w_140_1348, w_140_1350, w_140_1351, w_140_1353, w_140_1364, w_140_1365, w_140_1367, w_140_1370, w_140_1374, w_140_1376, w_140_1377, w_140_1379, w_140_1385, w_140_1387, w_140_1394, w_140_1396, w_140_1398, w_140_1399, w_140_1402, w_140_1407, w_140_1411, w_140_1414, w_140_1415, w_140_1417, w_140_1423, w_140_1424, w_140_1425, w_140_1426, w_140_1427, w_140_1430, w_140_1432, w_140_1438, w_140_1441, w_140_1444, w_140_1447, w_140_1450, w_140_1453, w_140_1456, w_140_1460, w_140_1465, w_140_1468, w_140_1469, w_140_1472, w_140_1477, w_140_1480, w_140_1485, w_140_1489, w_140_1500, w_140_1502, w_140_1505, w_140_1506, w_140_1509, w_140_1516, w_140_1519, w_140_1522, w_140_1523, w_140_1524, w_140_1527, w_140_1528, w_140_1530, w_140_1540, w_140_1542, w_140_1547, w_140_1548, w_140_1549, w_140_1555, w_140_1562, w_140_1567, w_140_1571, w_140_1572, w_140_1577, w_140_1580, w_140_1581, w_140_1583, w_140_1589, w_140_1597, w_140_1599, w_140_1605, w_140_1610, w_140_1611, w_140_1616, w_140_1617, w_140_1622, w_140_1624, w_140_1625, w_140_1626, w_140_1631, w_140_1635, w_140_1641, w_140_1643, w_140_1644, w_140_1650, w_140_1654, w_140_1657, w_140_1660, w_140_1662, w_140_1670, w_140_1671, w_140_1678, w_140_1679, w_140_1680, w_140_1681, w_140_1692, w_140_1693, w_140_1698, w_140_1699, w_140_1705, w_140_1706, w_140_1707, w_140_1708, w_140_1709, w_140_1711, w_140_1715, w_140_1718, w_140_1719, w_140_1720, w_140_1724, w_140_1726, w_140_1727, w_140_1730, w_140_1732, w_140_1734, w_140_1735, w_140_1741, w_140_1742, w_140_1747, w_140_1750, w_140_1751, w_140_1752, w_140_1753, w_140_1755, w_140_1760, w_140_1762, w_140_1765, w_140_1766, w_140_1767, w_140_1769, w_140_1770, w_140_1774, w_140_1776, w_140_1782, w_140_1787, w_140_1788, w_140_1789, w_140_1792, w_140_1797, w_140_1798, w_140_1799, w_140_1800, w_140_1801, w_140_1805, w_140_1807, w_140_1812, w_140_1814, w_140_1815, w_140_1816, w_140_1819, w_140_1820, w_140_1827, w_140_1830, w_140_1835, w_140_1837, w_140_1838, w_140_1843, w_140_1844, w_140_1846, w_140_1852, w_140_1853, w_140_1855, w_140_1859, w_140_1863, w_140_1865, w_140_1867, w_140_1868, w_140_1869, w_140_1871, w_140_1876, w_140_1877, w_140_1878, w_140_1885, w_140_1887, w_140_1890, w_140_1893, w_140_1896, w_140_1897, w_140_1900, w_140_1906, w_140_1907, w_140_1908, w_140_1911, w_140_1912, w_140_1916, w_140_1926, w_140_1929, w_140_1931, w_140_1932, w_140_1933, w_140_1938, w_140_1939, w_140_1944, w_140_1945, w_140_1947, w_140_1950, w_140_1951, w_140_1953, w_140_1956, w_140_1966, w_140_1967, w_140_1969, w_140_1970, w_140_1975, w_140_1977, w_140_1979, w_140_1988, w_140_1989, w_140_1992, w_140_1996, w_140_2001, w_140_2005, w_140_2007, w_140_2008, w_140_2010, w_140_2012, w_140_2014, w_140_2015, w_140_2018, w_140_2024, w_140_2025, w_140_2029, w_140_2031, w_140_2032, w_140_2040, w_140_2042, w_140_2056, w_140_2060, w_140_2063, w_140_2065, w_140_2068, w_140_2070, w_140_2072, w_140_2074, w_140_2077, w_140_2083, w_140_2085, w_140_2086, w_140_2088, w_140_2089, w_140_2093, w_140_2096, w_140_2098, w_140_2106, w_140_2107, w_140_2109, w_140_2113, w_140_2114, w_140_2125, w_140_2128, w_140_2132, w_140_2133, w_140_2134, w_140_2139, w_140_2141, w_140_2142, w_140_2143, w_140_2150, w_140_2151, w_140_2156, w_140_2161, w_140_2162, w_140_2165, w_140_2167, w_140_2169, w_140_2171, w_140_2172, w_140_2174, w_140_2177, w_140_2184, w_140_2194, w_140_2198, w_140_2200, w_140_2201, w_140_2203, w_140_2204, w_140_2207, w_140_2208, w_140_2209, w_140_2213, w_140_2218, w_140_2221, w_140_2222, w_140_2224, w_140_2229, w_140_2240, w_140_2245, w_140_2246, w_140_2248, w_140_2254, w_140_2259, w_140_2261, w_140_2268, w_140_2270, w_140_2271, w_140_2281, w_140_2282, w_140_2283, w_140_2284, w_140_2289, w_140_2290, w_140_2299, w_140_2302, w_140_2303, w_140_2307, w_140_2311, w_140_2313, w_140_2315, w_140_2318, w_140_2321, w_140_2322, w_140_2330, w_140_2332, w_140_2336, w_140_2338, w_140_2348, w_140_2350, w_140_2352, w_140_2354, w_140_2359, w_140_2361, w_140_2368, w_140_2369, w_140_2372, w_140_2375, w_140_2379, w_140_2380, w_140_2383, w_140_2385, w_140_2398, w_140_2400, w_140_2401, w_140_2404, w_140_2419, w_140_2427, w_140_2429, w_140_2431, w_140_2438, w_140_2439, w_140_2442, w_140_2443, w_140_2448, w_140_2452, w_140_2453, w_140_2454, w_140_2458, w_140_2460, w_140_2463, w_140_2471, w_140_2472, w_140_2481, w_140_2493, w_140_2511, w_140_2513, w_140_2518, w_140_2520, w_140_2521, w_140_2525, w_140_2527, w_140_2540, w_140_2545, w_140_2553, w_140_2556, w_140_2557, w_140_2558, w_140_2561, w_140_2562, w_140_2572, w_140_2580, w_140_2581, w_140_2588, w_140_2590, w_140_2592, w_140_2594, w_140_2599, w_140_2604, w_140_2605, w_140_2612, w_140_2622, w_140_2628;
  wire w_141_000, w_141_001, w_141_002, w_141_006, w_141_009, w_141_010, w_141_011, w_141_017, w_141_022, w_141_024, w_141_028, w_141_031, w_141_035, w_141_036, w_141_037, w_141_038, w_141_041, w_141_043, w_141_048, w_141_050, w_141_051, w_141_052, w_141_060, w_141_063, w_141_064, w_141_065, w_141_066, w_141_067, w_141_068, w_141_069, w_141_070, w_141_073, w_141_076, w_141_077, w_141_079, w_141_081, w_141_085, w_141_088, w_141_089, w_141_093, w_141_098, w_141_101, w_141_103, w_141_105, w_141_108, w_141_110, w_141_111, w_141_113, w_141_114, w_141_116, w_141_128, w_141_129, w_141_131, w_141_132, w_141_134, w_141_136, w_141_137, w_141_139, w_141_141, w_141_145, w_141_146, w_141_147, w_141_150, w_141_152, w_141_154, w_141_155, w_141_156, w_141_157, w_141_158, w_141_160, w_141_161, w_141_162, w_141_165, w_141_169, w_141_171, w_141_172, w_141_173, w_141_175, w_141_176, w_141_177, w_141_179, w_141_180, w_141_181, w_141_182, w_141_183, w_141_184, w_141_186, w_141_187, w_141_189, w_141_190, w_141_192, w_141_193, w_141_195, w_141_203, w_141_204, w_141_206, w_141_211, w_141_213, w_141_214, w_141_215, w_141_216, w_141_219, w_141_222, w_141_224, w_141_228, w_141_235, w_141_236, w_141_240, w_141_242, w_141_247, w_141_251, w_141_253, w_141_256, w_141_257, w_141_260, w_141_262, w_141_264, w_141_267, w_141_270, w_141_273, w_141_275, w_141_280, w_141_281, w_141_282, w_141_283, w_141_284, w_141_285, w_141_286, w_141_288, w_141_289, w_141_290, w_141_291, w_141_292, w_141_297, w_141_298, w_141_299, w_141_300, w_141_303, w_141_304, w_141_305, w_141_307, w_141_308, w_141_312, w_141_313, w_141_316, w_141_317, w_141_318, w_141_319, w_141_322, w_141_328, w_141_329, w_141_335, w_141_336, w_141_337, w_141_338, w_141_339, w_141_340, w_141_345, w_141_347, w_141_351, w_141_353, w_141_356, w_141_357, w_141_358, w_141_359, w_141_360, w_141_361, w_141_364, w_141_365, w_141_368, w_141_370, w_141_371, w_141_372, w_141_377, w_141_379, w_141_380, w_141_383, w_141_384, w_141_385, w_141_386, w_141_387, w_141_388, w_141_396, w_141_401, w_141_404, w_141_405, w_141_406, w_141_408, w_141_411, w_141_413, w_141_416, w_141_420, w_141_422, w_141_423, w_141_425, w_141_429, w_141_432, w_141_434, w_141_437, w_141_438, w_141_439, w_141_441, w_141_443, w_141_444, w_141_451, w_141_452, w_141_453, w_141_455, w_141_461, w_141_466, w_141_467, w_141_472, w_141_474, w_141_475, w_141_477, w_141_479, w_141_480, w_141_481, w_141_483, w_141_484, w_141_487, w_141_490, w_141_493, w_141_494, w_141_495, w_141_498, w_141_502, w_141_503, w_141_506, w_141_507, w_141_508, w_141_509, w_141_510, w_141_511, w_141_512, w_141_515, w_141_518, w_141_519, w_141_520, w_141_523, w_141_524, w_141_526, w_141_527, w_141_528, w_141_529, w_141_533, w_141_534, w_141_535, w_141_537, w_141_538, w_141_543, w_141_545, w_141_546, w_141_549, w_141_550, w_141_551, w_141_552, w_141_553, w_141_554, w_141_555, w_141_556, w_141_558, w_141_559, w_141_560, w_141_561, w_141_563, w_141_566, w_141_567, w_141_570, w_141_571, w_141_572, w_141_574, w_141_575, w_141_576, w_141_580, w_141_582, w_141_587, w_141_588, w_141_592, w_141_597, w_141_598, w_141_599, w_141_600, w_141_601, w_141_602, w_141_603, w_141_604, w_141_605, w_141_611, w_141_612, w_141_615, w_141_617, w_141_621, w_141_622, w_141_624, w_141_626, w_141_627, w_141_628, w_141_629, w_141_630, w_141_631, w_141_633, w_141_634, w_141_637, w_141_638, w_141_639, w_141_640, w_141_644, w_141_646, w_141_648, w_141_649, w_141_650, w_141_651, w_141_652, w_141_653, w_141_654, w_141_658, w_141_660, w_141_668, w_141_671, w_141_673, w_141_676, w_141_678, w_141_680, w_141_683, w_141_687, w_141_689, w_141_690, w_141_691, w_141_693, w_141_696, w_141_700, w_141_704, w_141_706, w_141_707, w_141_708, w_141_710, w_141_711, w_141_713, w_141_716, w_141_717, w_141_719, w_141_721, w_141_723, w_141_724, w_141_727, w_141_728, w_141_731, w_141_733, w_141_734, w_141_736, w_141_737, w_141_741, w_141_744, w_141_745, w_141_748, w_141_751, w_141_754, w_141_755, w_141_756, w_141_760, w_141_761, w_141_763, w_141_764, w_141_765, w_141_772, w_141_775, w_141_776, w_141_777, w_141_780, w_141_786, w_141_787, w_141_789, w_141_792, w_141_795, w_141_797, w_141_798, w_141_799, w_141_800, w_141_803, w_141_805, w_141_810, w_141_811, w_141_816, w_141_822, w_141_824, w_141_825, w_141_826, w_141_828, w_141_831, w_141_832, w_141_833, w_141_834, w_141_835, w_141_836, w_141_841, w_141_842, w_141_845, w_141_848, w_141_849, w_141_850, w_141_851, w_141_852, w_141_854, w_141_855, w_141_857, w_141_859, w_141_862, w_141_865, w_141_868, w_141_871, w_141_872, w_141_873, w_141_877, w_141_880, w_141_882, w_141_884, w_141_887, w_141_888, w_141_898, w_141_899, w_141_900, w_141_901, w_141_902, w_141_903, w_141_909, w_141_910, w_141_911, w_141_913, w_141_917, w_141_918, w_141_919, w_141_922, w_141_923, w_141_928, w_141_929, w_141_935, w_141_939, w_141_940, w_141_944, w_141_945, w_141_949, w_141_950, w_141_951, w_141_958, w_141_959, w_141_961, w_141_962, w_141_964, w_141_965, w_141_966, w_141_969, w_141_970, w_141_971, w_141_972, w_141_975, w_141_979, w_141_984, w_141_985, w_141_987, w_141_988, w_141_991, w_141_993, w_141_996, w_141_997, w_141_1000, w_141_1001, w_141_1002, w_141_1006, w_141_1010, w_141_1013, w_141_1016, w_141_1020, w_141_1021, w_141_1025, w_141_1027, w_141_1028, w_141_1029, w_141_1032, w_141_1035, w_141_1037, w_141_1039, w_141_1040, w_141_1041, w_141_1043, w_141_1044, w_141_1048, w_141_1051, w_141_1053, w_141_1058, w_141_1066, w_141_1070, w_141_1071, w_141_1076, w_141_1077, w_141_1078, w_141_1080, w_141_1081, w_141_1082, w_141_1086, w_141_1087, w_141_1088, w_141_1089, w_141_1090, w_141_1093, w_141_1094, w_141_1096, w_141_1098, w_141_1101, w_141_1102, w_141_1103, w_141_1104, w_141_1108, w_141_1112, w_141_1113, w_141_1114, w_141_1116, w_141_1117, w_141_1118, w_141_1119, w_141_1121, w_141_1123, w_141_1124, w_141_1128, w_141_1130, w_141_1131, w_141_1132, w_141_1133, w_141_1134, w_141_1136, w_141_1137, w_141_1138, w_141_1140, w_141_1141, w_141_1142, w_141_1143, w_141_1145, w_141_1147, w_141_1148, w_141_1151, w_141_1152, w_141_1153, w_141_1154, w_141_1156, w_141_1158, w_141_1160, w_141_1162, w_141_1163, w_141_1164, w_141_1169, w_141_1173, w_141_1174, w_141_1176, w_141_1178, w_141_1180, w_141_1181, w_141_1182, w_141_1185, w_141_1187, w_141_1188, w_141_1189, w_141_1190, w_141_1194, w_141_1196, w_141_1197, w_141_1198, w_141_1200, w_141_1202, w_141_1207, w_141_1208, w_141_1209, w_141_1210, w_141_1219, w_141_1220, w_141_1224, w_141_1226, w_141_1228, w_141_1229, w_141_1230, w_141_1235, w_141_1237, w_141_1239, w_141_1240, w_141_1242, w_141_1246, w_141_1248, w_141_1249, w_141_1250, w_141_1251, w_141_1257, w_141_1261, w_141_1262, w_141_1263, w_141_1265, w_141_1273, w_141_1276, w_141_1278, w_141_1287, w_141_1288, w_141_1291, w_141_1293, w_141_1294, w_141_1300, w_141_1302, w_141_1303, w_141_1305, w_141_1306, w_141_1307, w_141_1309, w_141_1312, w_141_1316, w_141_1317, w_141_1318, w_141_1319, w_141_1320, w_141_1323, w_141_1325, w_141_1326, w_141_1328, w_141_1333, w_141_1335, w_141_1337, w_141_1339, w_141_1341, w_141_1344, w_141_1345, w_141_1346, w_141_1347, w_141_1349, w_141_1350, w_141_1351, w_141_1353, w_141_1354, w_141_1355, w_141_1357, w_141_1358, w_141_1359, w_141_1361, w_141_1363, w_141_1364, w_141_1365, w_141_1366, w_141_1368, w_141_1369, w_141_1372, w_141_1373, w_141_1374, w_141_1377, w_141_1379, w_141_1382, w_141_1385, w_141_1393, w_141_1394, w_141_1399, w_141_1403, w_141_1407, w_141_1408, w_141_1410, w_141_1412, w_141_1415, w_141_1416, w_141_1421, w_141_1424, w_141_1425, w_141_1426, w_141_1428, w_141_1432, w_141_1433, w_141_1436, w_141_1440, w_141_1445, w_141_1452, w_141_1456, w_141_1460, w_141_1461, w_141_1462, w_141_1465, w_141_1468, w_141_1470, w_141_1473, w_141_1475, w_141_1476, w_141_1479, w_141_1481, w_141_1484, w_141_1487, w_141_1490, w_141_1491, w_141_1498, w_141_1499, w_141_1504, w_141_1505, w_141_1506, w_141_1509, w_141_1515, w_141_1517, w_141_1520, w_141_1522, w_141_1523, w_141_1527, w_141_1533, w_141_1534, w_141_1537, w_141_1541, w_141_1546, w_141_1547, w_141_1548, w_141_1551, w_141_1555, w_141_1556, w_141_1560, w_141_1561, w_141_1562, w_141_1565, w_141_1569, w_141_1570, w_141_1571, w_141_1575, w_141_1576, w_141_1577, w_141_1579, w_141_1581, w_141_1584, w_141_1588, w_141_1589, w_141_1591, w_141_1592, w_141_1594, w_141_1601, w_141_1602, w_141_1605, w_141_1608, w_141_1616, w_141_1617, w_141_1618, w_141_1623, w_141_1625, w_141_1627, w_141_1628, w_141_1631, w_141_1633, w_141_1636, w_141_1637, w_141_1639, w_141_1642, w_141_1645, w_141_1652, w_141_1657, w_141_1661, w_141_1662, w_141_1664, w_141_1665, w_141_1667, w_141_1668, w_141_1676, w_141_1683, w_141_1685, w_141_1690, w_141_1691, w_141_1694, w_141_1701, w_141_1702, w_141_1704, w_141_1708, w_141_1711, w_141_1713, w_141_1714, w_141_1715, w_141_1718, w_141_1723, w_141_1725, w_141_1729, w_141_1733, w_141_1734, w_141_1738, w_141_1739, w_141_1744, w_141_1745, w_141_1746, w_141_1748, w_141_1749, w_141_1750, w_141_1752, w_141_1754, w_141_1764, w_141_1766, w_141_1770, w_141_1772, w_141_1773, w_141_1775, w_141_1784, w_141_1786, w_141_1790, w_141_1792, w_141_1793, w_141_1794, w_141_1800, w_141_1803, w_141_1805, w_141_1808, w_141_1810, w_141_1811, w_141_1815, w_141_1816, w_141_1817, w_141_1818, w_141_1820, w_141_1822, w_141_1823, w_141_1824, w_141_1825, w_141_1826, w_141_1828;
  wire w_142_003, w_142_005, w_142_007, w_142_008, w_142_009, w_142_016, w_142_018, w_142_020, w_142_021, w_142_022, w_142_029, w_142_030, w_142_032, w_142_036, w_142_040, w_142_041, w_142_043, w_142_047, w_142_052, w_142_053, w_142_054, w_142_062, w_142_064, w_142_066, w_142_070, w_142_071, w_142_072, w_142_074, w_142_075, w_142_082, w_142_083, w_142_090, w_142_093, w_142_103, w_142_106, w_142_108, w_142_109, w_142_112, w_142_113, w_142_114, w_142_124, w_142_125, w_142_129, w_142_131, w_142_134, w_142_138, w_142_139, w_142_143, w_142_151, w_142_158, w_142_163, w_142_172, w_142_173, w_142_177, w_142_181, w_142_184, w_142_189, w_142_190, w_142_191, w_142_194, w_142_197, w_142_216, w_142_220, w_142_227, w_142_231, w_142_232, w_142_235, w_142_238, w_142_242, w_142_243, w_142_246, w_142_248, w_142_251, w_142_259, w_142_262, w_142_273, w_142_288, w_142_291, w_142_294, w_142_296, w_142_299, w_142_306, w_142_309, w_142_312, w_142_313, w_142_319, w_142_323, w_142_324, w_142_332, w_142_339, w_142_340, w_142_341, w_142_347, w_142_353, w_142_356, w_142_365, w_142_376, w_142_378, w_142_381, w_142_383, w_142_384, w_142_385, w_142_396, w_142_405, w_142_418, w_142_421, w_142_434, w_142_454, w_142_456, w_142_457, w_142_458, w_142_464, w_142_465, w_142_466, w_142_471, w_142_477, w_142_479, w_142_488, w_142_490, w_142_497, w_142_499, w_142_505, w_142_507, w_142_508, w_142_512, w_142_513, w_142_521, w_142_526, w_142_530, w_142_537, w_142_541, w_142_544, w_142_554, w_142_558, w_142_571, w_142_574, w_142_586, w_142_595, w_142_610, w_142_617, w_142_627, w_142_631, w_142_632, w_142_634, w_142_646, w_142_651, w_142_657, w_142_660, w_142_668, w_142_669, w_142_673, w_142_678, w_142_680, w_142_682, w_142_690, w_142_693, w_142_700, w_142_708, w_142_718, w_142_720, w_142_729, w_142_749, w_142_759, w_142_761, w_142_766, w_142_770, w_142_772, w_142_774, w_142_779, w_142_782, w_142_784, w_142_797, w_142_801, w_142_809, w_142_817, w_142_822, w_142_827, w_142_838, w_142_840, w_142_863, w_142_864, w_142_872, w_142_877, w_142_880, w_142_881, w_142_889, w_142_893, w_142_902, w_142_907, w_142_909, w_142_910, w_142_911, w_142_913, w_142_916, w_142_919, w_142_925, w_142_928, w_142_929, w_142_946, w_142_948, w_142_951, w_142_955, w_142_958, w_142_963, w_142_971, w_142_980, w_142_981, w_142_991, w_142_1006, w_142_1042, w_142_1044, w_142_1072, w_142_1077, w_142_1078, w_142_1082, w_142_1086, w_142_1087, w_142_1098, w_142_1101, w_142_1102, w_142_1103, w_142_1108, w_142_1110, w_142_1111, w_142_1115, w_142_1120, w_142_1121, w_142_1128, w_142_1130, w_142_1135, w_142_1138, w_142_1145, w_142_1152, w_142_1172, w_142_1173, w_142_1174, w_142_1177, w_142_1186, w_142_1188, w_142_1191, w_142_1208, w_142_1212, w_142_1218, w_142_1230, w_142_1234, w_142_1239, w_142_1243, w_142_1247, w_142_1248, w_142_1252, w_142_1269, w_142_1276, w_142_1280, w_142_1296, w_142_1297, w_142_1307, w_142_1309, w_142_1310, w_142_1314, w_142_1319, w_142_1322, w_142_1325, w_142_1337, w_142_1339, w_142_1342, w_142_1344, w_142_1351, w_142_1355, w_142_1357, w_142_1366, w_142_1372, w_142_1386, w_142_1392, w_142_1398, w_142_1405, w_142_1406, w_142_1410, w_142_1416, w_142_1427, w_142_1432, w_142_1434, w_142_1437, w_142_1441, w_142_1442, w_142_1448, w_142_1461, w_142_1463, w_142_1466, w_142_1475, w_142_1476, w_142_1480, w_142_1484, w_142_1497, w_142_1498, w_142_1499, w_142_1506, w_142_1517, w_142_1521, w_142_1524, w_142_1547, w_142_1555, w_142_1560, w_142_1562, w_142_1564, w_142_1566, w_142_1568, w_142_1574, w_142_1575, w_142_1579, w_142_1581, w_142_1592, w_142_1596, w_142_1608, w_142_1619, w_142_1623, w_142_1633, w_142_1640, w_142_1651, w_142_1664, w_142_1669, w_142_1678, w_142_1679, w_142_1680, w_142_1681, w_142_1685, w_142_1687, w_142_1692, w_142_1693, w_142_1694, w_142_1695, w_142_1710, w_142_1713, w_142_1718, w_142_1719, w_142_1720, w_142_1728, w_142_1737, w_142_1738, w_142_1741, w_142_1744, w_142_1749, w_142_1754, w_142_1759, w_142_1761, w_142_1775, w_142_1782, w_142_1788, w_142_1791, w_142_1794, w_142_1805, w_142_1811, w_142_1813, w_142_1814, w_142_1815, w_142_1816, w_142_1821, w_142_1822, w_142_1825, w_142_1830, w_142_1839, w_142_1847, w_142_1851, w_142_1867, w_142_1881, w_142_1890, w_142_1896, w_142_1897, w_142_1900, w_142_1901, w_142_1908, w_142_1910, w_142_1911, w_142_1913, w_142_1916, w_142_1918, w_142_1920, w_142_1925, w_142_1930, w_142_1932, w_142_1937, w_142_1940, w_142_1955, w_142_1965, w_142_1967, w_142_1972, w_142_1974, w_142_1980, w_142_1982, w_142_1983, w_142_1998, w_142_2004, w_142_2010, w_142_2016, w_142_2024, w_142_2029, w_142_2037, w_142_2041, w_142_2049, w_142_2060, w_142_2071, w_142_2078, w_142_2079, w_142_2080, w_142_2084, w_142_2087, w_142_2091, w_142_2092, w_142_2102, w_142_2106, w_142_2114, w_142_2117, w_142_2120, w_142_2126, w_142_2128, w_142_2130, w_142_2142, w_142_2145, w_142_2146, w_142_2150, w_142_2154, w_142_2158, w_142_2171, w_142_2174, w_142_2179, w_142_2180, w_142_2181, w_142_2184, w_142_2186, w_142_2187, w_142_2200, w_142_2204, w_142_2205, w_142_2207, w_142_2213, w_142_2217, w_142_2225, w_142_2226, w_142_2228, w_142_2235, w_142_2236, w_142_2238, w_142_2246, w_142_2265, w_142_2267, w_142_2268, w_142_2270, w_142_2289, w_142_2299, w_142_2304, w_142_2313, w_142_2315, w_142_2325, w_142_2328, w_142_2332, w_142_2351, w_142_2362, w_142_2368, w_142_2369, w_142_2377, w_142_2390, w_142_2408, w_142_2423, w_142_2424, w_142_2438, w_142_2448, w_142_2453, w_142_2456, w_142_2459, w_142_2472, w_142_2477, w_142_2480, w_142_2482, w_142_2483, w_142_2486, w_142_2491, w_142_2500, w_142_2503, w_142_2504, w_142_2523, w_142_2526, w_142_2534, w_142_2536, w_142_2540, w_142_2545, w_142_2548, w_142_2550, w_142_2551, w_142_2553, w_142_2565, w_142_2569, w_142_2570, w_142_2584, w_142_2585, w_142_2594, w_142_2598, w_142_2599, w_142_2603, w_142_2606, w_142_2620, w_142_2633, w_142_2636, w_142_2637, w_142_2644, w_142_2649, w_142_2651, w_142_2652, w_142_2663, w_142_2668, w_142_2673, w_142_2679, w_142_2681, w_142_2683, w_142_2684, w_142_2689, w_142_2690, w_142_2701, w_142_2706, w_142_2710, w_142_2711, w_142_2718, w_142_2720, w_142_2723, w_142_2726, w_142_2730, w_142_2733, w_142_2736, w_142_2743, w_142_2747, w_142_2766, w_142_2767, w_142_2769, w_142_2773, w_142_2774, w_142_2777, w_142_2781, w_142_2784, w_142_2792, w_142_2808, w_142_2812, w_142_2815, w_142_2816, w_142_2817, w_142_2820, w_142_2821, w_142_2827, w_142_2828, w_142_2830, w_142_2835, w_142_2837, w_142_2841, w_142_2845, w_142_2846, w_142_2848, w_142_2849, w_142_2852, w_142_2858, w_142_2865, w_142_2877, w_142_2880, w_142_2882, w_142_2883, w_142_2889, w_142_2897, w_142_2900, w_142_2918, w_142_2920, w_142_2935, w_142_2948, w_142_2949, w_142_2958, w_142_2959, w_142_2962, w_142_2963, w_142_2973, w_142_2982, w_142_2983, w_142_2987, w_142_2993, w_142_3002, w_142_3007, w_142_3009, w_142_3014, w_142_3015, w_142_3016, w_142_3037, w_142_3038, w_142_3039, w_142_3046, w_142_3050, w_142_3051, w_142_3055, w_142_3057, w_142_3060, w_142_3071, w_142_3072, w_142_3084, w_142_3089, w_142_3098, w_142_3106, w_142_3110, w_142_3112, w_142_3123, w_142_3124, w_142_3131, w_142_3136, w_142_3137, w_142_3140, w_142_3147, w_142_3151, w_142_3152, w_142_3164, w_142_3170, w_142_3171, w_142_3172, w_142_3174, w_142_3183, w_142_3188, w_142_3196, w_142_3202, w_142_3203, w_142_3204, w_142_3209, w_142_3211, w_142_3220, w_142_3221, w_142_3222, w_142_3226, w_142_3239, w_142_3245, w_142_3246, w_142_3250, w_142_3257, w_142_3265, w_142_3269, w_142_3270, w_142_3274, w_142_3275, w_142_3276, w_142_3282, w_142_3288, w_142_3289, w_142_3291, w_142_3294, w_142_3296, w_142_3297, w_142_3308, w_142_3309, w_142_3310, w_142_3315, w_142_3322, w_142_3324, w_142_3330, w_142_3342, w_142_3343, w_142_3346, w_142_3352, w_142_3353, w_142_3354, w_142_3355, w_142_3357, w_142_3359, w_142_3371, w_142_3375, w_142_3390, w_142_3393, w_142_3396, w_142_3398, w_142_3402, w_142_3403, w_142_3407, w_142_3419, w_142_3421, w_142_3422, w_142_3423, w_142_3435, w_142_3440, w_142_3452, w_142_3454, w_142_3455, w_142_3458, w_142_3464, w_142_3471, w_142_3476, w_142_3481, w_142_3482, w_142_3492, w_142_3513, w_142_3514, w_142_3516, w_142_3521, w_142_3522, w_142_3536, w_142_3539, w_142_3542, w_142_3548, w_142_3549, w_142_3550, w_142_3553, w_142_3560, w_142_3562, w_142_3583, w_142_3587, w_142_3592, w_142_3598, w_142_3599, w_142_3605, w_142_3624, w_142_3627, w_142_3636, w_142_3644, w_142_3647, w_142_3653, w_142_3657, w_142_3663, w_142_3668, w_142_3674, w_142_3677, w_142_3692, w_142_3707, w_142_3710, w_142_3715, w_142_3716, w_142_3717, w_142_3743, w_142_3754, w_142_3756, w_142_3773, w_142_3774, w_142_3778, w_142_3791, w_142_3792, w_142_3794, w_142_3801, w_142_3802, w_142_3810, w_142_3814, w_142_3821, w_142_3823, w_142_3824, w_142_3838, w_142_3839, w_142_3840, w_142_3841, w_142_3842, w_142_3852, w_142_3854, w_142_3856, w_142_3857, w_142_3858, w_142_3861, w_142_3864, w_142_3871, w_142_3879, w_142_3880, w_142_3889, w_142_3894, w_142_3901, w_142_3903, w_142_3907, w_142_3912, w_142_3913, w_142_3916, w_142_3923, w_142_3925, w_142_3927, w_142_3928, w_142_3933, w_142_3936, w_142_3941, w_142_3948, w_142_3962, w_142_3967, w_142_3989, w_142_3990, w_142_3994, w_142_4011, w_142_4022, w_142_4025, w_142_4031, w_142_4032, w_142_4035, w_142_4036, w_142_4039, w_142_4040, w_142_4043, w_142_4046, w_142_4051, w_142_4054, w_142_4058, w_142_4060, w_142_4080, w_142_4082, w_142_4087, w_142_4088, w_142_4097, w_142_4108, w_142_4112, w_142_4118, w_142_4128, w_142_4131, w_142_4133, w_142_4140, w_142_4145, w_142_4146, w_142_4158, w_142_4163, w_142_4168, w_142_4171, w_142_4176, w_142_4178, w_142_4195, w_142_4207, w_142_4211, w_142_4218, w_142_4224, w_142_4225, w_142_4231, w_142_4244, w_142_4250, w_142_4253, w_142_4255, w_142_4262, w_142_4266, w_142_4270, w_142_4273, w_142_4274, w_142_4275, w_142_4276, w_142_4288, w_142_4289, w_142_4297, w_142_4302, w_142_4306, w_142_4314, w_142_4318, w_142_4325, w_142_4326, w_142_4335, w_142_4337, w_142_4343, w_142_4369, w_142_4371, w_142_4378, w_142_4379, w_142_4380, w_142_4381, w_142_4388, w_142_4395, w_142_4398, w_142_4402, w_142_4405, w_142_4412, w_142_4415, w_142_4416, w_142_4421, w_142_4422, w_142_4424, w_142_4427, w_142_4432, w_142_4442, w_142_4443, w_142_4447, w_142_4449, w_142_4455, w_142_4456, w_142_4459, w_142_4463, w_142_4475, w_142_4478, w_142_4488, w_142_4490, w_142_4492, w_142_4494, w_142_4498, w_142_4505, w_142_4510, w_142_4516, w_142_4522, w_142_4534, w_142_4539, w_142_4541, w_142_4563, w_142_4564, w_142_4565, w_142_4575, w_142_4579, w_142_4580, w_142_4597, w_142_4598, w_142_4604, w_142_4605, w_142_4606, w_142_4612, w_142_4622, w_142_4626, w_142_4627, w_142_4630, w_142_4637, w_142_4638, w_142_4645, w_142_4648, w_142_4654, w_142_4688, w_142_4700, w_142_4704, w_142_4706, w_142_4707, w_142_4709, w_142_4717, w_142_4733, w_142_4740, w_142_4741, w_142_4748, w_142_4755, w_142_4762, w_142_4767, w_142_4769, w_142_4772, w_142_4775, w_142_4776, w_142_4779, w_142_4785, w_142_4789, w_142_4790, w_142_4791, w_142_4792, w_142_4793, w_142_4796, w_142_4797, w_142_4798, w_142_4808, w_142_4822, w_142_4835, w_142_4838, w_142_4848;
  wire w_143_000, w_143_001, w_143_002, w_143_003, w_143_004, w_143_005, w_143_006, w_143_007, w_143_009, w_143_010, w_143_011, w_143_012, w_143_013, w_143_015, w_143_017, w_143_018, w_143_020, w_143_021, w_143_022, w_143_023, w_143_025, w_143_026, w_143_027, w_143_028, w_143_030, w_143_032, w_143_033, w_143_034, w_143_036, w_143_038, w_143_039, w_143_041, w_143_042, w_143_043, w_143_044, w_143_045, w_143_046, w_143_048, w_143_049, w_143_051, w_143_052, w_143_053, w_143_054, w_143_055, w_143_056, w_143_057, w_143_058, w_143_060, w_143_061, w_143_062, w_143_063, w_143_064, w_143_065, w_143_068, w_143_069, w_143_072, w_143_073, w_143_074, w_143_075, w_143_076, w_143_078, w_143_079, w_143_080, w_143_082, w_143_083, w_143_085, w_143_086, w_143_088, w_143_089, w_143_091, w_143_092, w_143_095, w_143_096, w_143_097, w_143_098, w_143_099, w_143_100, w_143_101, w_143_102, w_143_104, w_143_105, w_143_106, w_143_108, w_143_112, w_143_113, w_143_114, w_143_116, w_143_117, w_143_118, w_143_120, w_143_121, w_143_123, w_143_125, w_143_126, w_143_132, w_143_135, w_143_136, w_143_137, w_143_140, w_143_142, w_143_143, w_143_145, w_143_146, w_143_147, w_143_150, w_143_151, w_143_152, w_143_153, w_143_154, w_143_155, w_143_156, w_143_158, w_143_159, w_143_160, w_143_163, w_143_164, w_143_165, w_143_166, w_143_167, w_143_168, w_143_171, w_143_172, w_143_173, w_143_174, w_143_177, w_143_178, w_143_179, w_143_181, w_143_183, w_143_185, w_143_186, w_143_187, w_143_190, w_143_191, w_143_192, w_143_194, w_143_195, w_143_196, w_143_197, w_143_198, w_143_200, w_143_201, w_143_202, w_143_203, w_143_204, w_143_206, w_143_207, w_143_208, w_143_209, w_143_210, w_143_211, w_143_212, w_143_213, w_143_214, w_143_217, w_143_218, w_143_222, w_143_225, w_143_229, w_143_230, w_143_235, w_143_236, w_143_237, w_143_238, w_143_239, w_143_240, w_143_241, w_143_244, w_143_245, w_143_246, w_143_247, w_143_248, w_143_249, w_143_250, w_143_251, w_143_253, w_143_254, w_143_255, w_143_256, w_143_257, w_143_260, w_143_261, w_143_264, w_143_265, w_143_266, w_143_267, w_143_270, w_143_271, w_143_274, w_143_276, w_143_277, w_143_278, w_143_280, w_143_289, w_143_290, w_143_291, w_143_292, w_143_294, w_143_296, w_143_298, w_143_299, w_143_300, w_143_306, w_143_308, w_143_309, w_143_310, w_143_311, w_143_313, w_143_314, w_143_315, w_143_316, w_143_317, w_143_318, w_143_322, w_143_325, w_143_328, w_143_329, w_143_331, w_143_332, w_143_334, w_143_337, w_143_338, w_143_339, w_143_341, w_143_342, w_143_343, w_143_344, w_143_345, w_143_347, w_143_349, w_143_350, w_143_352, w_143_353, w_143_354, w_143_355, w_143_356, w_143_357, w_143_359, w_143_360, w_143_364, w_143_365, w_143_367, w_143_369, w_143_370, w_143_373, w_143_375, w_143_379, w_143_380, w_143_381, w_143_384, w_143_385, w_143_386, w_143_387, w_143_391, w_143_392, w_143_393, w_143_394, w_143_395, w_143_399, w_143_401, w_143_403, w_143_404, w_143_405, w_143_406, w_143_408, w_143_410, w_143_411, w_143_412, w_143_414, w_143_415, w_143_416, w_143_419, w_143_420, w_143_421, w_143_422, w_143_423, w_143_424, w_143_427, w_143_428, w_143_429, w_143_432, w_143_434, w_143_435, w_143_436, w_143_437, w_143_438, w_143_439, w_143_440, w_143_444, w_143_445, w_143_446, w_143_447, w_143_448, w_143_450, w_143_451, w_143_453, w_143_454, w_143_455, w_143_457, w_143_460, w_143_461, w_143_462, w_143_463, w_143_466, w_143_467, w_143_469, w_143_470, w_143_471, w_143_474, w_143_476, w_143_477, w_143_478, w_143_479, w_143_480, w_143_481, w_143_482, w_143_483, w_143_484, w_143_488, w_143_491, w_143_492, w_143_493, w_143_494, w_143_496, w_143_497, w_143_498, w_143_499, w_143_500, w_143_501, w_143_502, w_143_503, w_143_504, w_143_505, w_143_507, w_143_508, w_143_510, w_143_511, w_143_512, w_143_513, w_143_514, w_143_516, w_143_519, w_143_522, w_143_523, w_143_525, w_143_526, w_143_528, w_143_530, w_143_532, w_143_533, w_143_534, w_143_536, w_143_537, w_143_539, w_143_540, w_143_541, w_143_543, w_143_544, w_143_545, w_143_546, w_143_547, w_143_549, w_143_550, w_143_551, w_143_552, w_143_554, w_143_556, w_143_558, w_143_561, w_143_562, w_143_563, w_143_565, w_143_566, w_143_567, w_143_569, w_143_571, w_143_573, w_143_576, w_143_580, w_143_582, w_143_583, w_143_584, w_143_585, w_143_586, w_143_587, w_143_591, w_143_593, w_143_595, w_143_597, w_143_598, w_143_599, w_143_600, w_143_602, w_143_603, w_143_604, w_143_605, w_143_607, w_143_611, w_143_612, w_143_614, w_143_615, w_143_616, w_143_618, w_143_620, w_143_621, w_143_622, w_143_627, w_143_628, w_143_629, w_143_630, w_143_632, w_143_633, w_143_635, w_143_638, w_143_643, w_143_646, w_143_648, w_143_650, w_143_651, w_143_654, w_143_655, w_143_657, w_143_660, w_143_663, w_143_664, w_143_665, w_143_666, w_143_667, w_143_669, w_143_671, w_143_672, w_143_673, w_143_674, w_143_676, w_143_677, w_143_678, w_143_682, w_143_683, w_143_684, w_143_685, w_143_687, w_143_688, w_143_689, w_143_690, w_143_691, w_143_694, w_143_695, w_143_696, w_143_698, w_143_699, w_143_700, w_143_702, w_143_703, w_143_706, w_143_709, w_143_710, w_143_711, w_143_713, w_143_715, w_143_716, w_143_718, w_143_719, w_143_721, w_143_722, w_143_725, w_143_726, w_143_729, w_143_731, w_143_733, w_143_734, w_143_735, w_143_736, w_143_738, w_143_740, w_143_742, w_143_743, w_143_744, w_143_745, w_143_746, w_143_747, w_143_750, w_143_751, w_143_753, w_143_757, w_143_759, w_143_760, w_143_765, w_143_766, w_143_767, w_143_770, w_143_771, w_143_772, w_143_773, w_143_775, w_143_776, w_143_777, w_143_779, w_143_780, w_143_782, w_143_783, w_143_786, w_143_787, w_143_788, w_143_789, w_143_790, w_143_792, w_143_793, w_143_794, w_143_795, w_143_797, w_143_800, w_143_801, w_143_802, w_143_805, w_143_806, w_143_810, w_143_812, w_143_814, w_143_815, w_143_816, w_143_818, w_143_819, w_143_820, w_143_821, w_143_823, w_143_825, w_143_826, w_143_828, w_143_829, w_143_830, w_143_831, w_143_832, w_143_834, w_143_835, w_143_837, w_143_841, w_143_843, w_143_844, w_143_846, w_143_847, w_143_848, w_143_849, w_143_852, w_143_855, w_143_856, w_143_858, w_143_859, w_143_860, w_143_861, w_143_862, w_143_864, w_143_866, w_143_867, w_143_869, w_143_870, w_143_872, w_143_875, w_143_878, w_143_880, w_143_881, w_143_882, w_143_883, w_143_884, w_143_885, w_143_886, w_143_888, w_143_890, w_143_894, w_143_896, w_143_897, w_143_898, w_143_899, w_143_900, w_143_901, w_143_902, w_143_903, w_143_905, w_143_906, w_143_907, w_143_908, w_143_909, w_143_911, w_143_912, w_143_915, w_143_916, w_143_921, w_143_927, w_143_928, w_143_929, w_143_930, w_143_931, w_143_932, w_143_933, w_143_935, w_143_937, w_143_938, w_143_939, w_143_940, w_143_942, w_143_945, w_143_946, w_143_947, w_143_949, w_143_950, w_143_951, w_143_953, w_143_954, w_143_955, w_143_956, w_143_957, w_143_959, w_143_960, w_143_961, w_143_962, w_143_963, w_143_964, w_143_965, w_143_967, w_143_968, w_143_969, w_143_970, w_143_971, w_143_975, w_143_976, w_143_977, w_143_978, w_143_979, w_143_984, w_143_985, w_143_986, w_143_987, w_143_988, w_143_989, w_143_990, w_143_991, w_143_992, w_143_994, w_143_996, w_143_997, w_143_998, w_143_999, w_143_1000, w_143_1001, w_143_1002, w_143_1003, w_143_1004, w_143_1005, w_143_1009, w_143_1010, w_143_1011, w_143_1012, w_143_1013, w_143_1014, w_143_1015, w_143_1016, w_143_1017, w_143_1018, w_143_1019, w_143_1021, w_143_1023, w_143_1024, w_143_1025, w_143_1026, w_143_1027, w_143_1029, w_143_1031, w_143_1032, w_143_1033, w_143_1034, w_143_1035, w_143_1036, w_143_1038;
  wire w_144_000, w_144_001, w_144_005, w_144_011, w_144_012, w_144_014, w_144_015, w_144_018, w_144_025, w_144_026, w_144_029, w_144_031, w_144_035, w_144_040, w_144_045, w_144_048, w_144_052, w_144_053, w_144_054, w_144_055, w_144_056, w_144_057, w_144_059, w_144_062, w_144_066, w_144_072, w_144_077, w_144_080, w_144_081, w_144_082, w_144_087, w_144_095, w_144_097, w_144_098, w_144_100, w_144_108, w_144_109, w_144_110, w_144_111, w_144_115, w_144_119, w_144_124, w_144_126, w_144_134, w_144_135, w_144_136, w_144_142, w_144_143, w_144_144, w_144_146, w_144_153, w_144_154, w_144_156, w_144_157, w_144_158, w_144_163, w_144_168, w_144_171, w_144_175, w_144_176, w_144_178, w_144_179, w_144_182, w_144_184, w_144_185, w_144_188, w_144_190, w_144_192, w_144_196, w_144_197, w_144_199, w_144_206, w_144_209, w_144_212, w_144_217, w_144_219, w_144_220, w_144_221, w_144_228, w_144_229, w_144_234, w_144_235, w_144_239, w_144_248, w_144_249, w_144_253, w_144_254, w_144_258, w_144_259, w_144_262, w_144_265, w_144_270, w_144_271, w_144_277, w_144_279, w_144_281, w_144_282, w_144_283, w_144_287, w_144_288, w_144_293, w_144_294, w_144_298, w_144_301, w_144_303, w_144_305, w_144_308, w_144_312, w_144_313, w_144_315, w_144_316, w_144_320, w_144_321, w_144_325, w_144_332, w_144_333, w_144_334, w_144_335, w_144_337, w_144_338, w_144_345, w_144_348, w_144_351, w_144_352, w_144_355, w_144_358, w_144_359, w_144_361, w_144_362, w_144_373, w_144_375, w_144_378, w_144_379, w_144_380, w_144_381, w_144_382, w_144_383, w_144_387, w_144_388, w_144_391, w_144_395, w_144_401, w_144_402, w_144_408, w_144_410, w_144_411, w_144_413, w_144_417, w_144_419, w_144_421, w_144_425, w_144_426, w_144_430, w_144_434, w_144_435, w_144_437, w_144_440, w_144_441, w_144_442, w_144_447, w_144_450, w_144_451, w_144_454, w_144_455, w_144_459, w_144_460, w_144_470, w_144_472, w_144_475, w_144_480, w_144_482, w_144_484, w_144_485, w_144_487, w_144_490, w_144_493, w_144_497, w_144_503, w_144_512, w_144_517, w_144_520, w_144_530, w_144_539, w_144_544, w_144_548, w_144_561, w_144_563, w_144_566, w_144_570, w_144_574, w_144_578, w_144_581, w_144_586, w_144_590, w_144_593, w_144_594, w_144_607, w_144_610, w_144_611, w_144_612, w_144_625, w_144_627, w_144_634, w_144_636, w_144_639, w_144_641, w_144_645, w_144_647, w_144_649, w_144_653, w_144_662, w_144_669, w_144_677, w_144_678, w_144_687, w_144_693, w_144_701, w_144_709, w_144_713, w_144_716, w_144_720, w_144_721, w_144_722, w_144_730, w_144_738, w_144_741, w_144_744, w_144_745, w_144_752, w_144_757, w_144_769, w_144_780, w_144_781, w_144_783, w_144_786, w_144_787, w_144_794, w_144_795, w_144_801, w_144_806, w_144_811, w_144_813, w_144_815, w_144_819, w_144_822, w_144_824, w_144_827, w_144_841, w_144_842, w_144_850, w_144_853, w_144_856, w_144_857, w_144_858, w_144_872, w_144_874, w_144_875, w_144_885, w_144_891, w_144_899, w_144_909, w_144_910, w_144_911, w_144_914, w_144_915, w_144_916, w_144_921, w_144_922, w_144_924, w_144_925, w_144_927, w_144_931, w_144_932, w_144_941, w_144_944, w_144_952, w_144_957, w_144_961, w_144_963, w_144_969, w_144_976, w_144_991, w_144_995, w_144_1002, w_144_1007, w_144_1013, w_144_1014, w_144_1039, w_144_1041, w_144_1047, w_144_1048, w_144_1049, w_144_1055, w_144_1058, w_144_1064, w_144_1072, w_144_1073, w_144_1092, w_144_1095, w_144_1098, w_144_1100, w_144_1109, w_144_1110, w_144_1116, w_144_1120, w_144_1122, w_144_1125, w_144_1126, w_144_1132, w_144_1140, w_144_1144, w_144_1153, w_144_1159, w_144_1163, w_144_1173, w_144_1175, w_144_1181, w_144_1196, w_144_1197, w_144_1199, w_144_1200, w_144_1203, w_144_1216, w_144_1236, w_144_1242, w_144_1245, w_144_1251, w_144_1254, w_144_1257, w_144_1262, w_144_1268, w_144_1274, w_144_1275, w_144_1287, w_144_1291, w_144_1299, w_144_1301, w_144_1312, w_144_1313, w_144_1324, w_144_1325, w_144_1334, w_144_1340, w_144_1356, w_144_1358, w_144_1362, w_144_1382, w_144_1387, w_144_1396, w_144_1398, w_144_1403, w_144_1404, w_144_1423, w_144_1431, w_144_1435, w_144_1437, w_144_1440, w_144_1445, w_144_1451, w_144_1455, w_144_1456, w_144_1466, w_144_1470, w_144_1473, w_144_1484, w_144_1487, w_144_1491, w_144_1503, w_144_1508, w_144_1512, w_144_1517, w_144_1524, w_144_1526, w_144_1527, w_144_1531, w_144_1537, w_144_1542, w_144_1544, w_144_1550, w_144_1557, w_144_1560, w_144_1580, w_144_1581, w_144_1591, w_144_1592, w_144_1600, w_144_1601, w_144_1607, w_144_1608, w_144_1619, w_144_1621, w_144_1645, w_144_1651, w_144_1656, w_144_1661, w_144_1668, w_144_1669, w_144_1676, w_144_1680, w_144_1685, w_144_1688, w_144_1692, w_144_1697, w_144_1707, w_144_1708, w_144_1718, w_144_1726, w_144_1732, w_144_1733, w_144_1736, w_144_1756, w_144_1759, w_144_1760, w_144_1774, w_144_1775, w_144_1776, w_144_1778, w_144_1786, w_144_1787, w_144_1794, w_144_1796, w_144_1803, w_144_1810, w_144_1814, w_144_1816, w_144_1818, w_144_1820, w_144_1825, w_144_1828, w_144_1829, w_144_1835, w_144_1841, w_144_1850, w_144_1853, w_144_1860, w_144_1861, w_144_1863, w_144_1872, w_144_1878, w_144_1884, w_144_1902, w_144_1907, w_144_1912, w_144_1927, w_144_1928, w_144_1931, w_144_1937, w_144_1944, w_144_1945, w_144_1948, w_144_1964, w_144_1969, w_144_1978, w_144_1979, w_144_1980, w_144_1984, w_144_1995, w_144_1996, w_144_2005, w_144_2009, w_144_2026, w_144_2033, w_144_2038, w_144_2041, w_144_2046, w_144_2047, w_144_2050, w_144_2067, w_144_2075, w_144_2077, w_144_2088, w_144_2090, w_144_2100, w_144_2115, w_144_2117, w_144_2121, w_144_2142, w_144_2147, w_144_2151, w_144_2160, w_144_2164, w_144_2174, w_144_2175, w_144_2179, w_144_2180, w_144_2185, w_144_2186, w_144_2193, w_144_2198, w_144_2200, w_144_2202, w_144_2203, w_144_2211, w_144_2213, w_144_2214, w_144_2217, w_144_2226, w_144_2235, w_144_2236, w_144_2239, w_144_2241, w_144_2245, w_144_2251, w_144_2252, w_144_2255, w_144_2273, w_144_2278, w_144_2284, w_144_2285, w_144_2288, w_144_2292, w_144_2294, w_144_2301, w_144_2303, w_144_2317, w_144_2318, w_144_2326, w_144_2331, w_144_2346, w_144_2356, w_144_2357, w_144_2358, w_144_2364, w_144_2373, w_144_2376, w_144_2377, w_144_2378, w_144_2379, w_144_2382, w_144_2384, w_144_2396, w_144_2401, w_144_2404, w_144_2417, w_144_2422, w_144_2427, w_144_2430, w_144_2441, w_144_2443, w_144_2446, w_144_2450, w_144_2454, w_144_2455, w_144_2458, w_144_2463, w_144_2468, w_144_2469, w_144_2473, w_144_2476, w_144_2478, w_144_2490, w_144_2492, w_144_2501, w_144_2504, w_144_2511, w_144_2515, w_144_2516, w_144_2521, w_144_2533, w_144_2542, w_144_2548, w_144_2550, w_144_2551, w_144_2555, w_144_2560, w_144_2561, w_144_2577, w_144_2582, w_144_2586, w_144_2601, w_144_2612, w_144_2627, w_144_2635, w_144_2636, w_144_2637, w_144_2641, w_144_2642, w_144_2646, w_144_2649, w_144_2655, w_144_2658, w_144_2667, w_144_2671, w_144_2672, w_144_2680, w_144_2684, w_144_2690, w_144_2696, w_144_2704, w_144_2722, w_144_2741, w_144_2745, w_144_2751, w_144_2755, w_144_2759, w_144_2762, w_144_2767, w_144_2773, w_144_2775, w_144_2790, w_144_2803, w_144_2805, w_144_2806, w_144_2813, w_144_2815, w_144_2820, w_144_2823, w_144_2827, w_144_2829, w_144_2833, w_144_2840, w_144_2841, w_144_2844, w_144_2849, w_144_2850, w_144_2865, w_144_2867, w_144_2872, w_144_2875, w_144_2887, w_144_2900, w_144_2902, w_144_2909, w_144_2917, w_144_2923, w_144_2926, w_144_2934, w_144_2936, w_144_2937, w_144_2941, w_144_2945, w_144_2946, w_144_2948, w_144_2949, w_144_2950, w_144_2958, w_144_2960, w_144_2962, w_144_2968, w_144_2973, w_144_2974, w_144_2975, w_144_2977, w_144_2985, w_144_2987, w_144_2996, w_144_3007, w_144_3014, w_144_3024, w_144_3035, w_144_3038, w_144_3046, w_144_3047, w_144_3048, w_144_3050, w_144_3059, w_144_3068, w_144_3074, w_144_3079, w_144_3085, w_144_3088, w_144_3093, w_144_3097, w_144_3098, w_144_3102, w_144_3106, w_144_3107, w_144_3114, w_144_3117, w_144_3133, w_144_3146, w_144_3152, w_144_3154, w_144_3157, w_144_3160, w_144_3161, w_144_3162, w_144_3169, w_144_3170, w_144_3184, w_144_3188, w_144_3189, w_144_3190, w_144_3202, w_144_3210, w_144_3211, w_144_3216, w_144_3218, w_144_3231, w_144_3239, w_144_3240, w_144_3241, w_144_3245, w_144_3269, w_144_3270, w_144_3281, w_144_3283, w_144_3290, w_144_3296, w_144_3297, w_144_3300, w_144_3305, w_144_3312, w_144_3313, w_144_3318, w_144_3322, w_144_3325, w_144_3335, w_144_3339, w_144_3349, w_144_3353, w_144_3355, w_144_3356, w_144_3372, w_144_3377, w_144_3388, w_144_3393, w_144_3395, w_144_3402, w_144_3416, w_144_3418, w_144_3421, w_144_3422, w_144_3431, w_144_3433, w_144_3434, w_144_3437, w_144_3441, w_144_3445, w_144_3453, w_144_3454, w_144_3455, w_144_3458, w_144_3462, w_144_3465, w_144_3466, w_144_3471, w_144_3477, w_144_3481, w_144_3487, w_144_3489, w_144_3496, w_144_3498, w_144_3499, w_144_3500, w_144_3504, w_144_3506, w_144_3514, w_144_3522, w_144_3523, w_144_3535, w_144_3546, w_144_3552, w_144_3557, w_144_3559, w_144_3560, w_144_3562, w_144_3567, w_144_3568, w_144_3579, w_144_3581, w_144_3582, w_144_3585, w_144_3594, w_144_3596, w_144_3597, w_144_3600, w_144_3602, w_144_3605, w_144_3606, w_144_3608, w_144_3615, w_144_3618, w_144_3619, w_144_3620, w_144_3623, w_144_3629, w_144_3635, w_144_3636, w_144_3645, w_144_3647, w_144_3649, w_144_3652, w_144_3654, w_144_3659, w_144_3667, w_144_3672, w_144_3676, w_144_3683, w_144_3684, w_144_3686, w_144_3697, w_144_3701, w_144_3704, w_144_3709, w_144_3711, w_144_3717, w_144_3719, w_144_3720, w_144_3730, w_144_3735, w_144_3739, w_144_3745, w_144_3746, w_144_3756, w_144_3757, w_144_3763, w_144_3766, w_144_3778, w_144_3780, w_144_3784, w_144_3787, w_144_3795, w_144_3797, w_144_3804, w_144_3811, w_144_3814, w_144_3822, w_144_3834, w_144_3836, w_144_3854, w_144_3856, w_144_3861, w_144_3863, w_144_3864, w_144_3871, w_144_3872, w_144_3873, w_144_3879, w_144_3896, w_144_3897, w_144_3906, w_144_3907, w_144_3911, w_144_3922, w_144_3925, w_144_3929, w_144_3932, w_144_3937, w_144_3942, w_144_3946, w_144_3949, w_144_3955, w_144_3963, w_144_3966, w_144_3983, w_144_3985, w_144_3991, w_144_4007, w_144_4020, w_144_4025, w_144_4038, w_144_4045, w_144_4046, w_144_4047, w_144_4060, w_144_4068, w_144_4075, w_144_4078, w_144_4085, w_144_4095, w_144_4108, w_144_4112, w_144_4113, w_144_4128, w_144_4132, w_144_4138, w_144_4156, w_144_4159, w_144_4161, w_144_4163, w_144_4164, w_144_4168, w_144_4174, w_144_4176, w_144_4178, w_144_4184, w_144_4186, w_144_4193, w_144_4194, w_144_4195, w_144_4198, w_144_4216, w_144_4217, w_144_4222, w_144_4225, w_144_4230, w_144_4232, w_144_4236, w_144_4243, w_144_4244, w_144_4252, w_144_4258, w_144_4269, w_144_4273, w_144_4275, w_144_4278, w_144_4279, w_144_4290, w_144_4291, w_144_4297, w_144_4309, w_144_4313, w_144_4315, w_144_4322, w_144_4326, w_144_4329, w_144_4336, w_144_4342, w_144_4345, w_144_4356, w_144_4389, w_144_4397, w_144_4409, w_144_4413, w_144_4414, w_144_4419, w_144_4424, w_144_4428, w_144_4429, w_144_4430, w_144_4435, w_144_4436, w_144_4453, w_144_4455, w_144_4459, w_144_4460, w_144_4462, w_144_4470, w_144_4473, w_144_4478, w_144_4479, w_144_4480, w_144_4482;
  wire w_145_004, w_145_005, w_145_010, w_145_011, w_145_012, w_145_016, w_145_028, w_145_030, w_145_031, w_145_033, w_145_034, w_145_041, w_145_048, w_145_050, w_145_051, w_145_062, w_145_064, w_145_066, w_145_067, w_145_071, w_145_072, w_145_073, w_145_075, w_145_077, w_145_079, w_145_081, w_145_085, w_145_089, w_145_091, w_145_092, w_145_094, w_145_095, w_145_099, w_145_102, w_145_103, w_145_105, w_145_106, w_145_111, w_145_118, w_145_119, w_145_122, w_145_128, w_145_129, w_145_130, w_145_132, w_145_133, w_145_135, w_145_140, w_145_141, w_145_146, w_145_148, w_145_152, w_145_155, w_145_156, w_145_157, w_145_159, w_145_161, w_145_164, w_145_165, w_145_166, w_145_174, w_145_179, w_145_182, w_145_183, w_145_187, w_145_189, w_145_193, w_145_195, w_145_196, w_145_200, w_145_201, w_145_207, w_145_219, w_145_222, w_145_224, w_145_226, w_145_227, w_145_232, w_145_234, w_145_241, w_145_250, w_145_252, w_145_256, w_145_259, w_145_267, w_145_270, w_145_271, w_145_274, w_145_281, w_145_285, w_145_288, w_145_293, w_145_296, w_145_297, w_145_298, w_145_299, w_145_301, w_145_303, w_145_305, w_145_306, w_145_307, w_145_308, w_145_309, w_145_316, w_145_327, w_145_328, w_145_332, w_145_333, w_145_335, w_145_340, w_145_342, w_145_348, w_145_350, w_145_354, w_145_356, w_145_359, w_145_360, w_145_363, w_145_367, w_145_376, w_145_377, w_145_379, w_145_380, w_145_382, w_145_385, w_145_388, w_145_391, w_145_392, w_145_393, w_145_395, w_145_400, w_145_404, w_145_405, w_145_407, w_145_409, w_145_417, w_145_418, w_145_426, w_145_427, w_145_429, w_145_438, w_145_440, w_145_441, w_145_443, w_145_448, w_145_451, w_145_454, w_145_457, w_145_458, w_145_461, w_145_462, w_145_470, w_145_475, w_145_477, w_145_479, w_145_483, w_145_484, w_145_486, w_145_489, w_145_490, w_145_492, w_145_497, w_145_498, w_145_501, w_145_506, w_145_509, w_145_512, w_145_513, w_145_517, w_145_523, w_145_524, w_145_528, w_145_531, w_145_534, w_145_535, w_145_543, w_145_544, w_145_545, w_145_546, w_145_552, w_145_555, w_145_556, w_145_557, w_145_559, w_145_564, w_145_566, w_145_567, w_145_568, w_145_570, w_145_580, w_145_582, w_145_587, w_145_588, w_145_593, w_145_594, w_145_597, w_145_603, w_145_612, w_145_613, w_145_614, w_145_616, w_145_618, w_145_621, w_145_624, w_145_625, w_145_626, w_145_631, w_145_632, w_145_634, w_145_635, w_145_636, w_145_637, w_145_638, w_145_640, w_145_644, w_145_645, w_145_648, w_145_649, w_145_650, w_145_653, w_145_655, w_145_656, w_145_661, w_145_662, w_145_665, w_145_667, w_145_668, w_145_670, w_145_674, w_145_676, w_145_678, w_145_682, w_145_684, w_145_688, w_145_690, w_145_696, w_145_698, w_145_704, w_145_708, w_145_711, w_145_714, w_145_716, w_145_720, w_145_726, w_145_727, w_145_731, w_145_734, w_145_736, w_145_740, w_145_744, w_145_745, w_145_747, w_145_748, w_145_749, w_145_750, w_145_754, w_145_755, w_145_760, w_145_763, w_145_765, w_145_766, w_145_767, w_145_768, w_145_772, w_145_773, w_145_774, w_145_783, w_145_784, w_145_787, w_145_788, w_145_789, w_145_792, w_145_794, w_145_796, w_145_798, w_145_803, w_145_806, w_145_811, w_145_815, w_145_824, w_145_829, w_145_834, w_145_837, w_145_838, w_145_840, w_145_843, w_145_845, w_145_847, w_145_848, w_145_849, w_145_850, w_145_854, w_145_862, w_145_867, w_145_869, w_145_872, w_145_879, w_145_885, w_145_888, w_145_889, w_145_892, w_145_893, w_145_895, w_145_898, w_145_900, w_145_902, w_145_903, w_145_906, w_145_908, w_145_909, w_145_911, w_145_913, w_145_914, w_145_916, w_145_917, w_145_918, w_145_922, w_145_927, w_145_928, w_145_940, w_145_941, w_145_943, w_145_950, w_145_954, w_145_959, w_145_960, w_145_964, w_145_978, w_145_980, w_145_981, w_145_988, w_145_990, w_145_992, w_145_993, w_145_996, w_145_1003, w_145_1007, w_145_1010, w_145_1011, w_145_1012, w_145_1020, w_145_1023, w_145_1026, w_145_1027, w_145_1030, w_145_1033, w_145_1035, w_145_1037, w_145_1038, w_145_1039, w_145_1040, w_145_1042, w_145_1048, w_145_1049, w_145_1050, w_145_1051, w_145_1053, w_145_1065, w_145_1070, w_145_1077, w_145_1078, w_145_1080, w_145_1089, w_145_1098, w_145_1100, w_145_1103, w_145_1105, w_145_1108, w_145_1112, w_145_1115, w_145_1132, w_145_1133, w_145_1137, w_145_1145, w_145_1148, w_145_1153, w_145_1161, w_145_1162, w_145_1166, w_145_1169, w_145_1170, w_145_1172, w_145_1175, w_145_1176, w_145_1177, w_145_1181, w_145_1186, w_145_1193, w_145_1194, w_145_1195, w_145_1197, w_145_1204, w_145_1206, w_145_1209, w_145_1212, w_145_1215, w_145_1219, w_145_1221, w_145_1222, w_145_1224, w_145_1225, w_145_1227, w_145_1238, w_145_1239, w_145_1240, w_145_1241, w_145_1242, w_145_1245, w_145_1249, w_145_1254, w_145_1255, w_145_1257, w_145_1258, w_145_1261, w_145_1262, w_145_1263, w_145_1268, w_145_1271, w_145_1273, w_145_1280, w_145_1281, w_145_1297, w_145_1298, w_145_1302, w_145_1303, w_145_1304, w_145_1305, w_145_1308, w_145_1310, w_145_1314, w_145_1320, w_145_1323, w_145_1326, w_145_1327, w_145_1346, w_145_1348, w_145_1349, w_145_1350, w_145_1352, w_145_1354, w_145_1358, w_145_1359, w_145_1361, w_145_1362, w_145_1367, w_145_1372, w_145_1373, w_145_1374, w_145_1375, w_145_1377, w_145_1379, w_145_1380, w_145_1381, w_145_1382, w_145_1384, w_145_1386, w_145_1387, w_145_1389, w_145_1390, w_145_1391, w_145_1392, w_145_1395, w_145_1402, w_145_1406, w_145_1407, w_145_1410, w_145_1412, w_145_1416, w_145_1419, w_145_1420, w_145_1422, w_145_1427, w_145_1430, w_145_1432, w_145_1435, w_145_1436, w_145_1438, w_145_1446, w_145_1449, w_145_1458, w_145_1459, w_145_1461, w_145_1462, w_145_1467, w_145_1468, w_145_1471, w_145_1477, w_145_1482, w_145_1484, w_145_1487, w_145_1490, w_145_1492, w_145_1501, w_145_1503, w_145_1504, w_145_1511, w_145_1512, w_145_1513, w_145_1516, w_145_1518, w_145_1521, w_145_1523, w_145_1527, w_145_1529, w_145_1530, w_145_1531, w_145_1534, w_145_1542, w_145_1544, w_145_1549, w_145_1553, w_145_1559, w_145_1565, w_145_1566, w_145_1576, w_145_1578, w_145_1581, w_145_1584, w_145_1585, w_145_1589, w_145_1590, w_145_1595, w_145_1596, w_145_1601, w_145_1603, w_145_1624, w_145_1626, w_145_1630, w_145_1634, w_145_1635, w_145_1640, w_145_1649, w_145_1650, w_145_1653, w_145_1654, w_145_1655, w_145_1656, w_145_1657, w_145_1658, w_145_1660, w_145_1661, w_145_1663, w_145_1664, w_145_1673, w_145_1674, w_145_1676, w_145_1681, w_145_1683, w_145_1684, w_145_1686, w_145_1687, w_145_1693, w_145_1696, w_145_1697, w_145_1700, w_145_1701, w_145_1704, w_145_1705, w_145_1706, w_145_1707, w_145_1708, w_145_1709, w_145_1712, w_145_1714, w_145_1718, w_145_1724, w_145_1725, w_145_1727, w_145_1728, w_145_1731, w_145_1736, w_145_1740, w_145_1741, w_145_1746, w_145_1748, w_145_1753, w_145_1756, w_145_1757, w_145_1762, w_145_1765, w_145_1768, w_145_1769, w_145_1770, w_145_1771, w_145_1774, w_145_1778, w_145_1780, w_145_1781, w_145_1782, w_145_1783, w_145_1784, w_145_1785, w_145_1786, w_145_1788, w_145_1790, w_145_1792, w_145_1793, w_145_1795, w_145_1799, w_145_1801, w_145_1809, w_145_1810, w_145_1811, w_145_1816, w_145_1817, w_145_1821, w_145_1824, w_145_1828, w_145_1832, w_145_1836, w_145_1837, w_145_1841, w_145_1843, w_145_1848, w_145_1850, w_145_1856, w_145_1859, w_145_1863, w_145_1866, w_145_1870, w_145_1874, w_145_1877, w_145_1883, w_145_1888, w_145_1891, w_145_1893, w_145_1897, w_145_1903, w_145_1907, w_145_1910, w_145_1914, w_145_1915, w_145_1923, w_145_1926, w_145_1936, w_145_1937, w_145_1938, w_145_1939, w_145_1941, w_145_1943, w_145_1946, w_145_1947, w_145_1948, w_145_1950, w_145_1959, w_145_1960, w_145_1962, w_145_1964, w_145_1968, w_145_1969, w_145_1973, w_145_1975, w_145_1977, w_145_1979, w_145_1981, w_145_1983, w_145_1986, w_145_1987, w_145_1994, w_145_1995, w_145_1996, w_145_1998, w_145_2000, w_145_2001, w_145_2011, w_145_2017, w_145_2018, w_145_2022, w_145_2024, w_145_2026, w_145_2036, w_145_2037, w_145_2038, w_145_2041, w_145_2045, w_145_2052, w_145_2054, w_145_2055, w_145_2058, w_145_2060, w_145_2065, w_145_2066, w_145_2068, w_145_2071, w_145_2074, w_145_2076, w_145_2077, w_145_2079, w_145_2081, w_145_2082, w_145_2083, w_145_2084, w_145_2085, w_145_2089, w_145_2091, w_145_2095, w_145_2096, w_145_2100, w_145_2103, w_145_2106, w_145_2111, w_145_2114, w_145_2116, w_145_2122, w_145_2128, w_145_2130, w_145_2131, w_145_2133, w_145_2134, w_145_2142, w_145_2143, w_145_2146, w_145_2151, w_145_2152, w_145_2159, w_145_2163, w_145_2164, w_145_2165, w_145_2166, w_145_2170, w_145_2171, w_145_2177, w_145_2179, w_145_2187, w_145_2189, w_145_2193, w_145_2194, w_145_2199, w_145_2200, w_145_2201, w_145_2202, w_145_2210, w_145_2213, w_145_2214, w_145_2215, w_145_2218, w_145_2224, w_145_2225, w_145_2230, w_145_2231, w_145_2240, w_145_2241, w_145_2242, w_145_2243, w_145_2246, w_145_2250, w_145_2252, w_145_2255, w_145_2256, w_145_2257, w_145_2259, w_145_2266, w_145_2268, w_145_2270, w_145_2272, w_145_2279, w_145_2281, w_145_2284, w_145_2287, w_145_2289, w_145_2291, w_145_2295, w_145_2296, w_145_2297, w_145_2300, w_145_2304, w_145_2306, w_145_2308, w_145_2310, w_145_2316, w_145_2320, w_145_2332, w_145_2333, w_145_2334, w_145_2336, w_145_2338, w_145_2344, w_145_2350, w_145_2353, w_145_2354, w_145_2356, w_145_2360, w_145_2361, w_145_2364, w_145_2368, w_145_2371, w_145_2372, w_145_2373, w_145_2374, w_145_2375, w_145_2376, w_145_2379, w_145_2380, w_145_2383, w_145_2386, w_145_2387, w_145_2388, w_145_2390, w_145_2391, w_145_2392, w_145_2395, w_145_2396, w_145_2401, w_145_2402, w_145_2406, w_145_2407, w_145_2408, w_145_2409, w_145_2410, w_145_2414, w_145_2421, w_145_2426, w_145_2427, w_145_2428, w_145_2436, w_145_2438, w_145_2440, w_145_2444, w_145_2449, w_145_2453, w_145_2458, w_145_2459, w_145_2460, w_145_2463, w_145_2464, w_145_2466, w_145_2469, w_145_2474, w_145_2478, w_145_2479, w_145_2480, w_145_2481, w_145_2483, w_145_2490, w_145_2491;
  wire w_146_000, w_146_001, w_146_005, w_146_006, w_146_007, w_146_009, w_146_010, w_146_011, w_146_013, w_146_014, w_146_015, w_146_016, w_146_017, w_146_018, w_146_020, w_146_021, w_146_022, w_146_023, w_146_024, w_146_025, w_146_027, w_146_028, w_146_029, w_146_030, w_146_032, w_146_033, w_146_034, w_146_038, w_146_040, w_146_041, w_146_043, w_146_045, w_146_047, w_146_048, w_146_049, w_146_055, w_146_058, w_146_062, w_146_063, w_146_065, w_146_066, w_146_067, w_146_069, w_146_070, w_146_072, w_146_073, w_146_074, w_146_075, w_146_077, w_146_080, w_146_081, w_146_084, w_146_085, w_146_087, w_146_088, w_146_089, w_146_091, w_146_095, w_146_096, w_146_097, w_146_098, w_146_100, w_146_103, w_146_104, w_146_105, w_146_106, w_146_111, w_146_112, w_146_115, w_146_118, w_146_122, w_146_124, w_146_125, w_146_127, w_146_128, w_146_129, w_146_130, w_146_134, w_146_135, w_146_136, w_146_137, w_146_138, w_146_139, w_146_140, w_146_141, w_146_142, w_146_143, w_146_145, w_146_146, w_146_147, w_146_148, w_146_150, w_146_154, w_146_155, w_146_156, w_146_157, w_146_159, w_146_160, w_146_161, w_146_162, w_146_163, w_146_164, w_146_167, w_146_169, w_146_170, w_146_171, w_146_172, w_146_173, w_146_174, w_146_177, w_146_178, w_146_179, w_146_181, w_146_182, w_146_183, w_146_187, w_146_189, w_146_190, w_146_193, w_146_194, w_146_197, w_146_198, w_146_199, w_146_200, w_146_202, w_146_203, w_146_205, w_146_206, w_146_207, w_146_209, w_146_210, w_146_211, w_146_212, w_146_217, w_146_219, w_146_220, w_146_222, w_146_223, w_146_224, w_146_227, w_146_230, w_146_232, w_146_233, w_146_235, w_146_237, w_146_238, w_146_239, w_146_241, w_146_243, w_146_244, w_146_245, w_146_246, w_146_247, w_146_250, w_146_251, w_146_252, w_146_253, w_146_254, w_146_255, w_146_256, w_146_258, w_146_259, w_146_261, w_146_262, w_146_263, w_146_267, w_146_268, w_146_269, w_146_270, w_146_271, w_146_272, w_146_273, w_146_274, w_146_275, w_146_276, w_146_279, w_146_280, w_146_282, w_146_283, w_146_285, w_146_286, w_146_288, w_146_289, w_146_293, w_146_296, w_146_297, w_146_298, w_146_299, w_146_300, w_146_302, w_146_305, w_146_306, w_146_308, w_146_309, w_146_310, w_146_312, w_146_316, w_146_317, w_146_319, w_146_320, w_146_321, w_146_322, w_146_323, w_146_325, w_146_330, w_146_331, w_146_333, w_146_334, w_146_336, w_146_340, w_146_341, w_146_342, w_146_343, w_146_347, w_146_350, w_146_352, w_146_353, w_146_355, w_146_356, w_146_357, w_146_360, w_146_361, w_146_362, w_146_363, w_146_364, w_146_365, w_146_370, w_146_371, w_146_372, w_146_374, w_146_376, w_146_377, w_146_379, w_146_380, w_146_381, w_146_383, w_146_385, w_146_390, w_146_391, w_146_393, w_146_394, w_146_395, w_146_397, w_146_399, w_146_400, w_146_402, w_146_404, w_146_405, w_146_407, w_146_408, w_146_410, w_146_411, w_146_412, w_146_413, w_146_414, w_146_421, w_146_422, w_146_427, w_146_428, w_146_429, w_146_430, w_146_431, w_146_437, w_146_439, w_146_440, w_146_443, w_146_444, w_146_445, w_146_446, w_146_447, w_146_448, w_146_450, w_146_451, w_146_452, w_146_453, w_146_454, w_146_455, w_146_456, w_146_457, w_146_460, w_146_465, w_146_466, w_146_469, w_146_471, w_146_473, w_146_474, w_146_475, w_146_476, w_146_481, w_146_485, w_146_489, w_146_490, w_146_491, w_146_493, w_146_495, w_146_501, w_146_504, w_146_505, w_146_507, w_146_508, w_146_511, w_146_516, w_146_517, w_146_520, w_146_522, w_146_523, w_146_526, w_146_527, w_146_529, w_146_530, w_146_531, w_146_532, w_146_533, w_146_537, w_146_539, w_146_540, w_146_541, w_146_546, w_146_547, w_146_548, w_146_549, w_146_553, w_146_557, w_146_560, w_146_561, w_146_562, w_146_565, w_146_566, w_146_567, w_146_568, w_146_569, w_146_572, w_146_576, w_146_577, w_146_579, w_146_582, w_146_584, w_146_586, w_146_587, w_146_588, w_146_589, w_146_590, w_146_591, w_146_593, w_146_596, w_146_598, w_146_599, w_146_600, w_146_601, w_146_602, w_146_603, w_146_604, w_146_610, w_146_612, w_146_613, w_146_614, w_146_615, w_146_616, w_146_618, w_146_620, w_146_621, w_146_622, w_146_629, w_146_631, w_146_632, w_146_635, w_146_638, w_146_639, w_146_642, w_146_643, w_146_646, w_146_650, w_146_651, w_146_652, w_146_653, w_146_654, w_146_655, w_146_656, w_146_657, w_146_658, w_146_659, w_146_660, w_146_661, w_146_664, w_146_665, w_146_667, w_146_669, w_146_672, w_146_673, w_146_674, w_146_677, w_146_678, w_146_680, w_146_687, w_146_688, w_146_689, w_146_690, w_146_691, w_146_692, w_146_694, w_146_696, w_146_702, w_146_705, w_146_707, w_146_719, w_146_720, w_146_722, w_146_723, w_146_724, w_146_725, w_146_729, w_146_730, w_146_731, w_146_732, w_146_733, w_146_737, w_146_738, w_146_739, w_146_740, w_146_743, w_146_744, w_146_746, w_146_747, w_146_750, w_146_753, w_146_754, w_146_755, w_146_756, w_146_757, w_146_758, w_146_761, w_146_766, w_146_767, w_146_770, w_146_773, w_146_774, w_146_776, w_146_778, w_146_782, w_146_783, w_146_787, w_146_788, w_146_791, w_146_793, w_146_794, w_146_795, w_146_796, w_146_797, w_146_799, w_146_800, w_146_805, w_146_806, w_146_807, w_146_812, w_146_813, w_146_815, w_146_816, w_146_817, w_146_818, w_146_820, w_146_821, w_146_823, w_146_826, w_146_829, w_146_830, w_146_831, w_146_832, w_146_834, w_146_836, w_146_837, w_146_838, w_146_839, w_146_840, w_146_844, w_146_845, w_146_846, w_146_848, w_146_849, w_146_850, w_146_851, w_146_853, w_146_856, w_146_857, w_146_859, w_146_860, w_146_861, w_146_863, w_146_864, w_146_866, w_146_869, w_146_870, w_146_871, w_146_880, w_146_883, w_146_884, w_146_886, w_146_887, w_146_888, w_146_889, w_146_890, w_146_891, w_146_893, w_146_894, w_146_896, w_146_898, w_146_899, w_146_900, w_146_902, w_146_903, w_146_904, w_146_905, w_146_907, w_146_912, w_146_916, w_146_917, w_146_918, w_146_921, w_146_922, w_146_923, w_146_924, w_146_926, w_146_927, w_146_928, w_146_931, w_146_933, w_146_934, w_146_935, w_146_936, w_146_937, w_146_938, w_146_940, w_146_944, w_146_945, w_146_952, w_146_953, w_146_954, w_146_955, w_146_958, w_146_961, w_146_962, w_146_963, w_146_967, w_146_968, w_146_969, w_146_972, w_146_973, w_146_975, w_146_977, w_146_978, w_146_983, w_146_984, w_146_985, w_146_987, w_146_988, w_146_990, w_146_992, w_146_993, w_146_994, w_146_995, w_146_997, w_146_998, w_146_999, w_146_1000, w_146_1001, w_146_1002, w_146_1003, w_146_1005, w_146_1006, w_146_1008, w_146_1010, w_146_1013, w_146_1014, w_146_1017, w_146_1018, w_146_1019, w_146_1020, w_146_1022, w_146_1023, w_146_1025, w_146_1026, w_146_1028, w_146_1029, w_146_1035, w_146_1036, w_146_1037, w_146_1038, w_146_1039, w_146_1041, w_146_1047, w_146_1051, w_146_1054, w_146_1059, w_146_1061, w_146_1062, w_146_1065, w_146_1067, w_146_1069, w_146_1072, w_146_1074, w_146_1075, w_146_1077, w_146_1079, w_146_1080, w_146_1082, w_146_1083, w_146_1084, w_146_1087, w_146_1089, w_146_1090, w_146_1092, w_146_1093, w_146_1096, w_146_1097, w_146_1098, w_146_1099, w_146_1100, w_146_1101, w_146_1102, w_146_1103, w_146_1105, w_146_1107, w_146_1108, w_146_1109, w_146_1113, w_146_1115, w_146_1116, w_146_1117, w_146_1120, w_146_1121, w_146_1123, w_146_1124, w_146_1125, w_146_1126, w_146_1128, w_146_1130, w_146_1131, w_146_1133, w_146_1134, w_146_1136, w_146_1138, w_146_1139, w_146_1140, w_146_1141, w_146_1142, w_146_1143, w_146_1144, w_146_1145, w_146_1149, w_146_1151, w_146_1152, w_146_1154, w_146_1156, w_146_1159, w_146_1160, w_146_1162, w_146_1164, w_146_1167, w_146_1168, w_146_1170, w_146_1171, w_146_1172, w_146_1173, w_146_1174, w_146_1175, w_146_1184, w_146_1185, w_146_1189, w_146_1191, w_146_1193, w_146_1195, w_146_1196, w_146_1198, w_146_1199, w_146_1200, w_146_1201, w_146_1203, w_146_1205, w_146_1206, w_146_1207, w_146_1208, w_146_1216, w_146_1217, w_146_1218, w_146_1221, w_146_1223, w_146_1227, w_146_1232;
  wire w_147_009, w_147_013, w_147_014, w_147_018, w_147_024, w_147_026, w_147_032, w_147_033, w_147_035, w_147_037, w_147_040, w_147_041, w_147_042, w_147_048, w_147_049, w_147_050, w_147_053, w_147_056, w_147_058, w_147_059, w_147_065, w_147_067, w_147_070, w_147_071, w_147_074, w_147_080, w_147_082, w_147_083, w_147_084, w_147_085, w_147_086, w_147_094, w_147_096, w_147_102, w_147_104, w_147_108, w_147_111, w_147_112, w_147_113, w_147_116, w_147_117, w_147_118, w_147_119, w_147_120, w_147_123, w_147_126, w_147_127, w_147_131, w_147_133, w_147_138, w_147_142, w_147_143, w_147_147, w_147_148, w_147_151, w_147_152, w_147_156, w_147_157, w_147_158, w_147_159, w_147_161, w_147_162, w_147_165, w_147_168, w_147_183, w_147_184, w_147_187, w_147_189, w_147_190, w_147_194, w_147_199, w_147_201, w_147_202, w_147_209, w_147_210, w_147_211, w_147_216, w_147_217, w_147_222, w_147_225, w_147_229, w_147_230, w_147_232, w_147_237, w_147_238, w_147_239, w_147_246, w_147_250, w_147_255, w_147_256, w_147_257, w_147_260, w_147_262, w_147_263, w_147_265, w_147_268, w_147_275, w_147_277, w_147_279, w_147_282, w_147_283, w_147_285, w_147_287, w_147_288, w_147_291, w_147_292, w_147_302, w_147_306, w_147_307, w_147_310, w_147_315, w_147_316, w_147_319, w_147_323, w_147_324, w_147_325, w_147_328, w_147_330, w_147_335, w_147_337, w_147_339, w_147_341, w_147_351, w_147_354, w_147_355, w_147_358, w_147_360, w_147_362, w_147_364, w_147_365, w_147_368, w_147_374, w_147_379, w_147_382, w_147_384, w_147_395, w_147_396, w_147_398, w_147_405, w_147_406, w_147_409, w_147_414, w_147_415, w_147_417, w_147_418, w_147_422, w_147_426, w_147_434, w_147_436, w_147_437, w_147_438, w_147_440, w_147_443, w_147_445, w_147_451, w_147_452, w_147_453, w_147_461, w_147_462, w_147_463, w_147_464, w_147_469, w_147_470, w_147_473, w_147_475, w_147_479, w_147_484, w_147_485, w_147_488, w_147_494, w_147_497, w_147_504, w_147_506, w_147_513, w_147_516, w_147_517, w_147_523, w_147_524, w_147_526, w_147_527, w_147_531, w_147_534, w_147_537, w_147_540, w_147_541, w_147_545, w_147_546, w_147_553, w_147_554, w_147_555, w_147_561, w_147_563, w_147_564, w_147_566, w_147_569, w_147_577, w_147_579, w_147_580, w_147_582, w_147_584, w_147_592, w_147_594, w_147_595, w_147_597, w_147_598, w_147_599, w_147_603, w_147_604, w_147_606, w_147_611, w_147_613, w_147_617, w_147_618, w_147_619, w_147_620, w_147_622, w_147_624, w_147_625, w_147_641, w_147_645, w_147_647, w_147_648, w_147_656, w_147_657, w_147_660, w_147_665, w_147_668, w_147_671, w_147_673, w_147_676, w_147_679, w_147_680, w_147_697, w_147_700, w_147_701, w_147_703, w_147_704, w_147_708, w_147_720, w_147_721, w_147_724, w_147_725, w_147_727, w_147_732, w_147_745, w_147_753, w_147_754, w_147_756, w_147_757, w_147_764, w_147_768, w_147_769, w_147_771, w_147_773, w_147_776, w_147_778, w_147_780, w_147_782, w_147_783, w_147_790, w_147_791, w_147_800, w_147_803, w_147_807, w_147_808, w_147_809, w_147_813, w_147_817, w_147_821, w_147_824, w_147_828, w_147_831, w_147_834, w_147_839, w_147_842, w_147_843, w_147_848, w_147_855, w_147_858, w_147_860, w_147_862, w_147_863, w_147_866, w_147_868, w_147_870, w_147_874, w_147_876, w_147_878, w_147_880, w_147_884, w_147_886, w_147_888, w_147_892, w_147_895, w_147_900, w_147_903, w_147_909, w_147_911, w_147_912, w_147_914, w_147_916, w_147_919, w_147_924, w_147_928, w_147_930, w_147_932, w_147_934, w_147_937, w_147_939, w_147_943, w_147_944, w_147_947, w_147_951, w_147_952, w_147_959, w_147_962, w_147_963, w_147_966, w_147_970, w_147_975, w_147_976, w_147_985, w_147_993, w_147_996, w_147_998, w_147_999, w_147_1001, w_147_1002, w_147_1013, w_147_1014, w_147_1020, w_147_1022, w_147_1024, w_147_1025, w_147_1027, w_147_1028, w_147_1032, w_147_1034, w_147_1036, w_147_1040, w_147_1046, w_147_1047, w_147_1055, w_147_1061, w_147_1062, w_147_1064, w_147_1067, w_147_1073, w_147_1075, w_147_1084, w_147_1096, w_147_1098, w_147_1100, w_147_1101, w_147_1102, w_147_1103, w_147_1105, w_147_1116, w_147_1119, w_147_1125, w_147_1126, w_147_1129, w_147_1130, w_147_1135, w_147_1136, w_147_1137, w_147_1138, w_147_1143, w_147_1145, w_147_1149, w_147_1150, w_147_1152, w_147_1157, w_147_1158, w_147_1159, w_147_1161, w_147_1162, w_147_1166, w_147_1168, w_147_1182, w_147_1185, w_147_1188, w_147_1190, w_147_1191, w_147_1195, w_147_1196, w_147_1197, w_147_1199, w_147_1200, w_147_1210, w_147_1214, w_147_1218, w_147_1225, w_147_1226, w_147_1228, w_147_1229, w_147_1234, w_147_1236, w_147_1238, w_147_1239, w_147_1243, w_147_1248, w_147_1249, w_147_1250, w_147_1251, w_147_1254, w_147_1255, w_147_1256, w_147_1262, w_147_1267, w_147_1271, w_147_1279, w_147_1280, w_147_1282, w_147_1285, w_147_1287, w_147_1296, w_147_1297, w_147_1300, w_147_1305, w_147_1306, w_147_1307, w_147_1311, w_147_1313, w_147_1314, w_147_1327, w_147_1329, w_147_1331, w_147_1332, w_147_1339, w_147_1342, w_147_1349, w_147_1351, w_147_1356, w_147_1362, w_147_1363, w_147_1366, w_147_1367, w_147_1368, w_147_1375, w_147_1377, w_147_1388, w_147_1394, w_147_1401, w_147_1404, w_147_1405, w_147_1409, w_147_1410, w_147_1417, w_147_1418, w_147_1419, w_147_1421, w_147_1429, w_147_1430, w_147_1431, w_147_1432, w_147_1435, w_147_1436, w_147_1442, w_147_1445, w_147_1450, w_147_1452, w_147_1453, w_147_1455, w_147_1456, w_147_1458, w_147_1459, w_147_1460, w_147_1465, w_147_1466, w_147_1467, w_147_1470, w_147_1471, w_147_1473, w_147_1478, w_147_1479, w_147_1481, w_147_1482, w_147_1483, w_147_1484, w_147_1485, w_147_1489, w_147_1490, w_147_1492, w_147_1494, w_147_1500, w_147_1503, w_147_1508, w_147_1511, w_147_1513, w_147_1515, w_147_1516, w_147_1519, w_147_1524, w_147_1529, w_147_1530, w_147_1534, w_147_1536, w_147_1539, w_147_1540, w_147_1541, w_147_1543, w_147_1545, w_147_1550, w_147_1554, w_147_1555, w_147_1556, w_147_1557, w_147_1567, w_147_1569, w_147_1574, w_147_1576, w_147_1577, w_147_1578, w_147_1584, w_147_1589, w_147_1592, w_147_1593, w_147_1594, w_147_1595, w_147_1599, w_147_1600, w_147_1601, w_147_1604, w_147_1612, w_147_1613, w_147_1614, w_147_1619, w_147_1622, w_147_1623, w_147_1628, w_147_1629, w_147_1632, w_147_1634, w_147_1635, w_147_1637, w_147_1639, w_147_1643, w_147_1644, w_147_1646, w_147_1648, w_147_1649, w_147_1650, w_147_1652, w_147_1654, w_147_1655, w_147_1658, w_147_1659, w_147_1663, w_147_1664, w_147_1665, w_147_1669, w_147_1670, w_147_1671, w_147_1672, w_147_1674, w_147_1681, w_147_1684, w_147_1689, w_147_1692, w_147_1694, w_147_1704, w_147_1709, w_147_1713, w_147_1715, w_147_1717, w_147_1719, w_147_1720, w_147_1722, w_147_1724, w_147_1726, w_147_1727, w_147_1731, w_147_1735, w_147_1743, w_147_1744, w_147_1747, w_147_1749, w_147_1763, w_147_1776, w_147_1781, w_147_1782, w_147_1787, w_147_1796, w_147_1797, w_147_1803, w_147_1804, w_147_1816, w_147_1839, w_147_1844, w_147_1845, w_147_1855, w_147_1857, w_147_1863, w_147_1877, w_147_1880, w_147_1883, w_147_1887, w_147_1888, w_147_1897, w_147_1898, w_147_1902, w_147_1904, w_147_1923, w_147_1929, w_147_1932, w_147_1933, w_147_1936, w_147_1940, w_147_1950, w_147_1954, w_147_1956, w_147_1959, w_147_1968, w_147_1986, w_147_1988, w_147_1990, w_147_1999, w_147_2004, w_147_2006, w_147_2010, w_147_2012, w_147_2013, w_147_2014, w_147_2016, w_147_2023, w_147_2038, w_147_2039, w_147_2041, w_147_2044, w_147_2060, w_147_2070, w_147_2075, w_147_2080, w_147_2092, w_147_2096, w_147_2097, w_147_2108, w_147_2109, w_147_2114, w_147_2116, w_147_2134, w_147_2144, w_147_2150, w_147_2161, w_147_2162, w_147_2168, w_147_2179, w_147_2183, w_147_2191, w_147_2195, w_147_2204, w_147_2214, w_147_2229, w_147_2230, w_147_2241, w_147_2246, w_147_2247, w_147_2257, w_147_2274, w_147_2284, w_147_2310, w_147_2315, w_147_2330, w_147_2338, w_147_2347, w_147_2350, w_147_2355, w_147_2368, w_147_2371, w_147_2386, w_147_2388, w_147_2392, w_147_2405, w_147_2408, w_147_2413, w_147_2421, w_147_2425, w_147_2445, w_147_2446, w_147_2466, w_147_2500, w_147_2504, w_147_2514, w_147_2519, w_147_2521, w_147_2523, w_147_2525, w_147_2527, w_147_2534, w_147_2539, w_147_2544, w_147_2545, w_147_2556, w_147_2557, w_147_2561, w_147_2562, w_147_2568, w_147_2573, w_147_2578, w_147_2595, w_147_2596, w_147_2600, w_147_2604, w_147_2614, w_147_2620, w_147_2623, w_147_2635, w_147_2637, w_147_2638, w_147_2639, w_147_2642, w_147_2653, w_147_2655, w_147_2659, w_147_2660, w_147_2666, w_147_2669, w_147_2677, w_147_2682, w_147_2684, w_147_2689, w_147_2693, w_147_2700, w_147_2703, w_147_2711, w_147_2712, w_147_2716, w_147_2726, w_147_2728, w_147_2729, w_147_2735, w_147_2751, w_147_2753, w_147_2755, w_147_2768, w_147_2776, w_147_2781, w_147_2786, w_147_2789, w_147_2795, w_147_2800, w_147_2802, w_147_2817, w_147_2834, w_147_2837, w_147_2851, w_147_2862, w_147_2868, w_147_2871, w_147_2873, w_147_2874, w_147_2883, w_147_2886, w_147_2890, w_147_2891, w_147_2894, w_147_2898, w_147_2901, w_147_2905, w_147_2910, w_147_2913, w_147_2914, w_147_2916, w_147_2919, w_147_2923, w_147_2924, w_147_2934, w_147_2945, w_147_2955, w_147_2961, w_147_2967, w_147_2973, w_147_2975, w_147_2976, w_147_2989, w_147_2992, w_147_2995, w_147_3000, w_147_3012, w_147_3019, w_147_3024, w_147_3025, w_147_3040, w_147_3044, w_147_3050, w_147_3052, w_147_3054, w_147_3056, w_147_3059, w_147_3061, w_147_3077, w_147_3097, w_147_3121, w_147_3133, w_147_3141, w_147_3152, w_147_3157, w_147_3162, w_147_3163, w_147_3168, w_147_3171, w_147_3172, w_147_3174, w_147_3176, w_147_3181, w_147_3184, w_147_3189, w_147_3190, w_147_3191, w_147_3197, w_147_3204, w_147_3205, w_147_3222, w_147_3224, w_147_3226, w_147_3233, w_147_3234, w_147_3242;
  wire w_148_000, w_148_001, w_148_004, w_148_005, w_148_008, w_148_009, w_148_010, w_148_013, w_148_015, w_148_018, w_148_020, w_148_026, w_148_029, w_148_032, w_148_036, w_148_037, w_148_039, w_148_048, w_148_049, w_148_053, w_148_054, w_148_058, w_148_067, w_148_073, w_148_074, w_148_078, w_148_079, w_148_083, w_148_097, w_148_099, w_148_101, w_148_104, w_148_107, w_148_110, w_148_111, w_148_114, w_148_116, w_148_118, w_148_123, w_148_124, w_148_133, w_148_136, w_148_138, w_148_147, w_148_149, w_148_154, w_148_159, w_148_161, w_148_163, w_148_164, w_148_167, w_148_169, w_148_170, w_148_182, w_148_184, w_148_186, w_148_191, w_148_192, w_148_194, w_148_195, w_148_197, w_148_198, w_148_205, w_148_206, w_148_208, w_148_211, w_148_214, w_148_215, w_148_219, w_148_220, w_148_223, w_148_224, w_148_225, w_148_229, w_148_230, w_148_234, w_148_243, w_148_244, w_148_247, w_148_251, w_148_255, w_148_263, w_148_267, w_148_268, w_148_269, w_148_271, w_148_272, w_148_273, w_148_274, w_148_275, w_148_280, w_148_282, w_148_283, w_148_286, w_148_293, w_148_295, w_148_296, w_148_297, w_148_298, w_148_299, w_148_303, w_148_304, w_148_305, w_148_307, w_148_310, w_148_315, w_148_319, w_148_320, w_148_321, w_148_325, w_148_328, w_148_332, w_148_334, w_148_340, w_148_342, w_148_349, w_148_353, w_148_354, w_148_364, w_148_366, w_148_368, w_148_370, w_148_373, w_148_378, w_148_382, w_148_383, w_148_386, w_148_388, w_148_390, w_148_392, w_148_397, w_148_398, w_148_399, w_148_403, w_148_404, w_148_412, w_148_416, w_148_417, w_148_418, w_148_420, w_148_423, w_148_429, w_148_430, w_148_434, w_148_437, w_148_443, w_148_447, w_148_461, w_148_464, w_148_473, w_148_474, w_148_475, w_148_476, w_148_479, w_148_480, w_148_484, w_148_485, w_148_486, w_148_489, w_148_491, w_148_492, w_148_495, w_148_504, w_148_507, w_148_511, w_148_512, w_148_515, w_148_517, w_148_519, w_148_522, w_148_524, w_148_525, w_148_534, w_148_535, w_148_539, w_148_540, w_148_542, w_148_545, w_148_548, w_148_549, w_148_550, w_148_551, w_148_553, w_148_555, w_148_564, w_148_570, w_148_574, w_148_577, w_148_585, w_148_588, w_148_589, w_148_593, w_148_594, w_148_597, w_148_603, w_148_604, w_148_605, w_148_609, w_148_612, w_148_614, w_148_615, w_148_618, w_148_621, w_148_622, w_148_623, w_148_624, w_148_629, w_148_631, w_148_632, w_148_633, w_148_635, w_148_636, w_148_638, w_148_639, w_148_646, w_148_655, w_148_664, w_148_666, w_148_667, w_148_668, w_148_675, w_148_676, w_148_679, w_148_680, w_148_682, w_148_683, w_148_684, w_148_686, w_148_687, w_148_689, w_148_691, w_148_692, w_148_697, w_148_705, w_148_706, w_148_707, w_148_711, w_148_712, w_148_713, w_148_716, w_148_720, w_148_721, w_148_724, w_148_728, w_148_732, w_148_737, w_148_742, w_148_744, w_148_746, w_148_748, w_148_749, w_148_755, w_148_756, w_148_762, w_148_763, w_148_767, w_148_769, w_148_773, w_148_777, w_148_783, w_148_784, w_148_795, w_148_798, w_148_800, w_148_803, w_148_804, w_148_812, w_148_819, w_148_824, w_148_825, w_148_826, w_148_829, w_148_832, w_148_833, w_148_834, w_148_835, w_148_836, w_148_839, w_148_844, w_148_850, w_148_851, w_148_854, w_148_856, w_148_857, w_148_860, w_148_865, w_148_873, w_148_877, w_148_878, w_148_879, w_148_882, w_148_883, w_148_884, w_148_886, w_148_887, w_148_894, w_148_895, w_148_898, w_148_899, w_148_900, w_148_905, w_148_907, w_148_910, w_148_916, w_148_927, w_148_928, w_148_929, w_148_933, w_148_934, w_148_949, w_148_951, w_148_952, w_148_958, w_148_959, w_148_960, w_148_963, w_148_964, w_148_965, w_148_967, w_148_970, w_148_972, w_148_976, w_148_985, w_148_987, w_148_994, w_148_997, w_148_1003, w_148_1005, w_148_1007, w_148_1010, w_148_1011, w_148_1014, w_148_1017, w_148_1025, w_148_1027, w_148_1029, w_148_1031, w_148_1035, w_148_1038, w_148_1044, w_148_1049, w_148_1050, w_148_1052, w_148_1053, w_148_1055, w_148_1059, w_148_1073, w_148_1084, w_148_1098, w_148_1099, w_148_1103, w_148_1104, w_148_1107, w_148_1112, w_148_1113, w_148_1114, w_148_1115, w_148_1118, w_148_1121, w_148_1129, w_148_1134, w_148_1135, w_148_1137, w_148_1141, w_148_1152, w_148_1166, w_148_1171, w_148_1173, w_148_1177, w_148_1180, w_148_1185, w_148_1186, w_148_1187, w_148_1203, w_148_1204, w_148_1208, w_148_1219, w_148_1221, w_148_1223, w_148_1232, w_148_1237, w_148_1251, w_148_1261, w_148_1274, w_148_1277, w_148_1286, w_148_1293, w_148_1301, w_148_1302, w_148_1304, w_148_1309, w_148_1311, w_148_1313, w_148_1324, w_148_1331, w_148_1334, w_148_1335, w_148_1338, w_148_1360, w_148_1361, w_148_1370, w_148_1371, w_148_1372, w_148_1376, w_148_1385, w_148_1390, w_148_1399, w_148_1407, w_148_1408, w_148_1431, w_148_1438, w_148_1443, w_148_1452, w_148_1454, w_148_1461, w_148_1463, w_148_1465, w_148_1472, w_148_1479, w_148_1480, w_148_1483, w_148_1493, w_148_1495, w_148_1505, w_148_1515, w_148_1516, w_148_1517, w_148_1520, w_148_1523, w_148_1524, w_148_1527, w_148_1528, w_148_1534, w_148_1542, w_148_1544, w_148_1550, w_148_1554, w_148_1559, w_148_1561, w_148_1562, w_148_1567, w_148_1591, w_148_1596, w_148_1598, w_148_1620, w_148_1629, w_148_1631, w_148_1633, w_148_1634, w_148_1639, w_148_1646, w_148_1647, w_148_1664, w_148_1667, w_148_1669, w_148_1672, w_148_1675, w_148_1681, w_148_1689, w_148_1694, w_148_1698, w_148_1710, w_148_1719, w_148_1727, w_148_1729, w_148_1730, w_148_1732, w_148_1733, w_148_1739, w_148_1741, w_148_1742, w_148_1747, w_148_1748, w_148_1751, w_148_1754, w_148_1756, w_148_1758, w_148_1760, w_148_1761, w_148_1762, w_148_1763, w_148_1774, w_148_1777, w_148_1779, w_148_1784, w_148_1786, w_148_1791, w_148_1795, w_148_1801, w_148_1805, w_148_1810, w_148_1811, w_148_1812, w_148_1814, w_148_1822, w_148_1824, w_148_1836, w_148_1852, w_148_1853, w_148_1859, w_148_1867, w_148_1868, w_148_1869, w_148_1870, w_148_1871, w_148_1873, w_148_1882, w_148_1888, w_148_1890, w_148_1902, w_148_1920, w_148_1924, w_148_1925, w_148_1929, w_148_1948, w_148_1957, w_148_1960, w_148_1961, w_148_1967, w_148_1968, w_148_1969, w_148_1970, w_148_1975, w_148_1986, w_148_1988, w_148_1996, w_148_1997, w_148_2002, w_148_2013, w_148_2016, w_148_2017, w_148_2022, w_148_2036, w_148_2045, w_148_2048, w_148_2054, w_148_2060, w_148_2089, w_148_2091, w_148_2095, w_148_2104, w_148_2127, w_148_2128, w_148_2134, w_148_2136, w_148_2139, w_148_2148, w_148_2160, w_148_2163, w_148_2164, w_148_2174, w_148_2203, w_148_2206, w_148_2209, w_148_2219, w_148_2221, w_148_2226, w_148_2232, w_148_2234, w_148_2244, w_148_2247, w_148_2254, w_148_2255, w_148_2258, w_148_2264, w_148_2265, w_148_2272, w_148_2280, w_148_2291, w_148_2299, w_148_2302, w_148_2312, w_148_2318, w_148_2323, w_148_2325, w_148_2332, w_148_2341, w_148_2353, w_148_2354, w_148_2357, w_148_2360, w_148_2364, w_148_2370, w_148_2374, w_148_2377, w_148_2382, w_148_2395, w_148_2396, w_148_2403, w_148_2415, w_148_2417, w_148_2418, w_148_2419, w_148_2429, w_148_2432, w_148_2437, w_148_2438, w_148_2440, w_148_2448, w_148_2451, w_148_2470, w_148_2472, w_148_2474, w_148_2477, w_148_2479, w_148_2481, w_148_2482, w_148_2487, w_148_2499, w_148_2503, w_148_2513, w_148_2518, w_148_2521, w_148_2523, w_148_2538, w_148_2550, w_148_2563, w_148_2565, w_148_2571, w_148_2575, w_148_2576, w_148_2585, w_148_2596, w_148_2598, w_148_2600, w_148_2629, w_148_2635, w_148_2642, w_148_2651, w_148_2658, w_148_2677, w_148_2686, w_148_2687, w_148_2693, w_148_2695, w_148_2696, w_148_2705, w_148_2706, w_148_2708, w_148_2709, w_148_2713, w_148_2717, w_148_2718, w_148_2719, w_148_2723, w_148_2725, w_148_2733, w_148_2734, w_148_2739, w_148_2742, w_148_2744, w_148_2746, w_148_2749, w_148_2754, w_148_2756, w_148_2771, w_148_2773, w_148_2775, w_148_2776, w_148_2779, w_148_2788, w_148_2793, w_148_2801, w_148_2808, w_148_2813, w_148_2834, w_148_2853, w_148_2857, w_148_2864, w_148_2876, w_148_2879, w_148_2880, w_148_2906, w_148_2914, w_148_2929, w_148_2933, w_148_2945, w_148_2985, w_148_2997, w_148_3004, w_148_3009, w_148_3013, w_148_3015, w_148_3019, w_148_3032, w_148_3034, w_148_3044, w_148_3045, w_148_3050, w_148_3056, w_148_3058, w_148_3065, w_148_3069, w_148_3070, w_148_3075, w_148_3080, w_148_3083, w_148_3091, w_148_3092, w_148_3096, w_148_3107, w_148_3114, w_148_3120, w_148_3123, w_148_3124, w_148_3132, w_148_3137, w_148_3138, w_148_3139, w_148_3143, w_148_3150, w_148_3154, w_148_3169, w_148_3171, w_148_3183, w_148_3195, w_148_3197, w_148_3198, w_148_3199, w_148_3202, w_148_3208, w_148_3213, w_148_3218, w_148_3219, w_148_3220, w_148_3223, w_148_3227, w_148_3229, w_148_3236, w_148_3254, w_148_3255, w_148_3256, w_148_3262, w_148_3264, w_148_3267, w_148_3269, w_148_3278, w_148_3281, w_148_3287, w_148_3288, w_148_3312, w_148_3315, w_148_3323, w_148_3325, w_148_3327, w_148_3335, w_148_3338, w_148_3343, w_148_3348, w_148_3352, w_148_3353, w_148_3354, w_148_3360, w_148_3363, w_148_3365, w_148_3370, w_148_3371, w_148_3380, w_148_3382, w_148_3386, w_148_3392, w_148_3393, w_148_3397, w_148_3398, w_148_3400, w_148_3407, w_148_3417, w_148_3420, w_148_3430, w_148_3433, w_148_3434, w_148_3443, w_148_3444, w_148_3446, w_148_3447, w_148_3449, w_148_3450, w_148_3457, w_148_3470, w_148_3472, w_148_3473, w_148_3483, w_148_3495, w_148_3503, w_148_3515, w_148_3519, w_148_3528, w_148_3532, w_148_3537, w_148_3539, w_148_3542, w_148_3562, w_148_3564, w_148_3571, w_148_3577, w_148_3583, w_148_3584, w_148_3598, w_148_3607, w_148_3610, w_148_3622, w_148_3626, w_148_3627, w_148_3630, w_148_3635, w_148_3640, w_148_3644, w_148_3645, w_148_3665, w_148_3667, w_148_3672, w_148_3674, w_148_3677, w_148_3691, w_148_3701, w_148_3709, w_148_3713, w_148_3717, w_148_3720, w_148_3722, w_148_3747, w_148_3752, w_148_3757, w_148_3758, w_148_3769, w_148_3772, w_148_3775, w_148_3776, w_148_3786, w_148_3788, w_148_3801, w_148_3803, w_148_3808, w_148_3809, w_148_3810, w_148_3811, w_148_3827, w_148_3836, w_148_3842, w_148_3844, w_148_3859, w_148_3868, w_148_3870, w_148_3878, w_148_3894, w_148_3906, w_148_3909, w_148_3915, w_148_3918, w_148_3921, w_148_3938, w_148_3939;
  wire w_149_000, w_149_001, w_149_002, w_149_003, w_149_006, w_149_007, w_149_008, w_149_009, w_149_010, w_149_011, w_149_012, w_149_013, w_149_014, w_149_015, w_149_016, w_149_018, w_149_019, w_149_021, w_149_023, w_149_024, w_149_025, w_149_026, w_149_027, w_149_028, w_149_030, w_149_031, w_149_032, w_149_033, w_149_035, w_149_036, w_149_037, w_149_039, w_149_040, w_149_041, w_149_042, w_149_043, w_149_046, w_149_047, w_149_049, w_149_050, w_149_051, w_149_052, w_149_053, w_149_054, w_149_055, w_149_056, w_149_057, w_149_058, w_149_059, w_149_060, w_149_061, w_149_062, w_149_064, w_149_065, w_149_066, w_149_068, w_149_069, w_149_070, w_149_071, w_149_072, w_149_073, w_149_074, w_149_075, w_149_076, w_149_078, w_149_079, w_149_080, w_149_083, w_149_085, w_149_086, w_149_087, w_149_088, w_149_089, w_149_090, w_149_091, w_149_092, w_149_093, w_149_094, w_149_095, w_149_096, w_149_097, w_149_098, w_149_099, w_149_100, w_149_101, w_149_102, w_149_103, w_149_104, w_149_105, w_149_106, w_149_107, w_149_108, w_149_109, w_149_110, w_149_111, w_149_112, w_149_113, w_149_115, w_149_116, w_149_117, w_149_118, w_149_119, w_149_120, w_149_121, w_149_122, w_149_124, w_149_126, w_149_127, w_149_128, w_149_129, w_149_132, w_149_133, w_149_134, w_149_135, w_149_136, w_149_137, w_149_138, w_149_139, w_149_140, w_149_142, w_149_143, w_149_145, w_149_147, w_149_148, w_149_151, w_149_152, w_149_153, w_149_154, w_149_155, w_149_157, w_149_158, w_149_159, w_149_160, w_149_161, w_149_162, w_149_163, w_149_164, w_149_165, w_149_166, w_149_167, w_149_168, w_149_169, w_149_170, w_149_171, w_149_172, w_149_173, w_149_174, w_149_175, w_149_176, w_149_177, w_149_178, w_149_179, w_149_180, w_149_181, w_149_182, w_149_183, w_149_184, w_149_185, w_149_186, w_149_187, w_149_188, w_149_189, w_149_190, w_149_193, w_149_194, w_149_195, w_149_196, w_149_197, w_149_198, w_149_199, w_149_200, w_149_201, w_149_202, w_149_203, w_149_204, w_149_205, w_149_206, w_149_207, w_149_208, w_149_209, w_149_210, w_149_211, w_149_213, w_149_214, w_149_216, w_149_217, w_149_218, w_149_219, w_149_222, w_149_223, w_149_224, w_149_225, w_149_227, w_149_228, w_149_229, w_149_230, w_149_231, w_149_232, w_149_233, w_149_234, w_149_236, w_149_238, w_149_240, w_149_242, w_149_243, w_149_245, w_149_246, w_149_247, w_149_248, w_149_249, w_149_250, w_149_251, w_149_253, w_149_256, w_149_257, w_149_258, w_149_262, w_149_263, w_149_264, w_149_266, w_149_267, w_149_270, w_149_271, w_149_272, w_149_273, w_149_274, w_149_275, w_149_276, w_149_277, w_149_278, w_149_279, w_149_280, w_149_281, w_149_282, w_149_284, w_149_285, w_149_286, w_149_287, w_149_288, w_149_289, w_149_290, w_149_291, w_149_292, w_149_293, w_149_294, w_149_295, w_149_297, w_149_298, w_149_299, w_149_300, w_149_301, w_149_302, w_149_303, w_149_304, w_149_308, w_149_309, w_149_310, w_149_311, w_149_312, w_149_313, w_149_314, w_149_315, w_149_316, w_149_317, w_149_318, w_149_319, w_149_320, w_149_321, w_149_322, w_149_323, w_149_324, w_149_326, w_149_328, w_149_329, w_149_330, w_149_331, w_149_332, w_149_333, w_149_334, w_149_335, w_149_336, w_149_337, w_149_338, w_149_339, w_149_340, w_149_341, w_149_342, w_149_344, w_149_345, w_149_347, w_149_348, w_149_349, w_149_350, w_149_351, w_149_352, w_149_353, w_149_355, w_149_356, w_149_357, w_149_358, w_149_359, w_149_360, w_149_361, w_149_362, w_149_363, w_149_364, w_149_365, w_149_366, w_149_367, w_149_368, w_149_369, w_149_370, w_149_371, w_149_372, w_149_373, w_149_374, w_149_375, w_149_376, w_149_377, w_149_378, w_149_379, w_149_380, w_149_381, w_149_382, w_149_385, w_149_386, w_149_387, w_149_388, w_149_390, w_149_391, w_149_392, w_149_393, w_149_394, w_149_395, w_149_396, w_149_397, w_149_399, w_149_401, w_149_402, w_149_403, w_149_406, w_149_407, w_149_409, w_149_410, w_149_411, w_149_412, w_149_413, w_149_415, w_149_416, w_149_417, w_149_419, w_149_420, w_149_421, w_149_422, w_149_423, w_149_425, w_149_427, w_149_429, w_149_431, w_149_432, w_149_433, w_149_434, w_149_435, w_149_436, w_149_437, w_149_438, w_149_440, w_149_441, w_149_442, w_149_444, w_149_445, w_149_446, w_149_448, w_149_450, w_149_452, w_149_453, w_149_454, w_149_455, w_149_456, w_149_457, w_149_458, w_149_459, w_149_462, w_149_463, w_149_464, w_149_465, w_149_466, w_149_467, w_149_468, w_149_469, w_149_471, w_149_475, w_149_476, w_149_477, w_149_478, w_149_479, w_149_480, w_149_482, w_149_483, w_149_484, w_149_486, w_149_487, w_149_489, w_149_490, w_149_491, w_149_492, w_149_493, w_149_495, w_149_496, w_149_497, w_149_498, w_149_499, w_149_500, w_149_501, w_149_502, w_149_503, w_149_504, w_149_505, w_149_506, w_149_508, w_149_509, w_149_510, w_149_511, w_149_512, w_149_513, w_149_514, w_149_515, w_149_516, w_149_519, w_149_520, w_149_521, w_149_522, w_149_525, w_149_526, w_149_527, w_149_528, w_149_530, w_149_532, w_149_533, w_149_536, w_149_538, w_149_539, w_149_541, w_149_543, w_149_544, w_149_546, w_149_547, w_149_548, w_149_549, w_149_550, w_149_551, w_149_552, w_149_553, w_149_554, w_149_555, w_149_556, w_149_557, w_149_558, w_149_559, w_149_560, w_149_562, w_149_563, w_149_564, w_149_565, w_149_566, w_149_567, w_149_568, w_149_569, w_149_570, w_149_573, w_149_574, w_149_577, w_149_578, w_149_579, w_149_580, w_149_581, w_149_582, w_149_584, w_149_585, w_149_586, w_149_588, w_149_589, w_149_590, w_149_591, w_149_592, w_149_593;
  wire w_150_000, w_150_001, w_150_002, w_150_003, w_150_004, w_150_005, w_150_006, w_150_007, w_150_008, w_150_009, w_150_010, w_150_011, w_150_012, w_150_013, w_150_014, w_150_015, w_150_016, w_150_017, w_150_018, w_150_019, w_150_020, w_150_021, w_150_022, w_150_023, w_150_024, w_150_025, w_150_026, w_150_027, w_150_028, w_150_029, w_150_030, w_150_031, w_150_032, w_150_033, w_150_034, w_150_035, w_150_036, w_150_037, w_150_038, w_150_039, w_150_040, w_150_041, w_150_042, w_150_043, w_150_044, w_150_045, w_150_046, w_150_047, w_150_048, w_150_049, w_150_050, w_150_051, w_150_052, w_150_053, w_150_054, w_150_055, w_150_056, w_150_057, w_150_058, w_150_059, w_150_060, w_150_061, w_150_062, w_150_063, w_150_064, w_150_065, w_150_066, w_150_067, w_150_068, w_150_069, w_150_071, w_150_072, w_150_073, w_150_074, w_150_075, w_150_076, w_150_077, w_150_078, w_150_080, w_150_081, w_150_082, w_150_083, w_150_084, w_150_085, w_150_086, w_150_087, w_150_088, w_150_089, w_150_090, w_150_091, w_150_093, w_150_094, w_150_095, w_150_096, w_150_097, w_150_098, w_150_099, w_150_100, w_150_101, w_150_102, w_150_103, w_150_104, w_150_105, w_150_106, w_150_107, w_150_108, w_150_109, w_150_110, w_150_111, w_150_112, w_150_113, w_150_114, w_150_115, w_150_116, w_150_117, w_150_118, w_150_119, w_150_120, w_150_121, w_150_122, w_150_123, w_150_124, w_150_125, w_150_126, w_150_127, w_150_128, w_150_129, w_150_130, w_150_131, w_150_132, w_150_133, w_150_134, w_150_135, w_150_136, w_150_137, w_150_138, w_150_139, w_150_140, w_150_141, w_150_142, w_150_143, w_150_144, w_150_145, w_150_146, w_150_147, w_150_148, w_150_149, w_150_150, w_150_151, w_150_153, w_150_154, w_150_155, w_150_156, w_150_157, w_150_158, w_150_159, w_150_160, w_150_161, w_150_162, w_150_163, w_150_164, w_150_165, w_150_166, w_150_167, w_150_168, w_150_169, w_150_170, w_150_171, w_150_172, w_150_173, w_150_174, w_150_175, w_150_176, w_150_177, w_150_178, w_150_179, w_150_180, w_150_181, w_150_182, w_150_183, w_150_184, w_150_185, w_150_186, w_150_187, w_150_188, w_150_189, w_150_190, w_150_191, w_150_192, w_150_193, w_150_194, w_150_195, w_150_196, w_150_197, w_150_198, w_150_199, w_150_200, w_150_201, w_150_202, w_150_203, w_150_204, w_150_205, w_150_206, w_150_207, w_150_208, w_150_209, w_150_210, w_150_211, w_150_212, w_150_213, w_150_214, w_150_215, w_150_216, w_150_217, w_150_218, w_150_219, w_150_220, w_150_222, w_150_223, w_150_224, w_150_225, w_150_226, w_150_227, w_150_228, w_150_229, w_150_230, w_150_231, w_150_232, w_150_233, w_150_234, w_150_235, w_150_236, w_150_237, w_150_238, w_150_239, w_150_240, w_150_241, w_150_242, w_150_243, w_150_244, w_150_245, w_150_246, w_150_247, w_150_248, w_150_249, w_150_250, w_150_251, w_150_252, w_150_253, w_150_254, w_150_255, w_150_256, w_150_257, w_150_258, w_150_259, w_150_260, w_150_261, w_150_262, w_150_263, w_150_264, w_150_265, w_150_266, w_150_267, w_150_268, w_150_269, w_150_270, w_150_272, w_150_273, w_150_274, w_150_275, w_150_276, w_150_277, w_150_278, w_150_279, w_150_280, w_150_281, w_150_282, w_150_283, w_150_284, w_150_287, w_150_288, w_150_289, w_150_290, w_150_294, w_150_295, w_150_296, w_150_297, w_150_298, w_150_299, w_150_301;
  wire w_151_004, w_151_005, w_151_006, w_151_007, w_151_013, w_151_015, w_151_019, w_151_024, w_151_030, w_151_032, w_151_035, w_151_037, w_151_043, w_151_046, w_151_047, w_151_048, w_151_052, w_151_060, w_151_061, w_151_062, w_151_065, w_151_068, w_151_075, w_151_076, w_151_078, w_151_080, w_151_082, w_151_085, w_151_093, w_151_098, w_151_112, w_151_113, w_151_116, w_151_117, w_151_120, w_151_121, w_151_123, w_151_124, w_151_129, w_151_133, w_151_136, w_151_137, w_151_138, w_151_142, w_151_145, w_151_147, w_151_151, w_151_152, w_151_153, w_151_156, w_151_157, w_151_159, w_151_166, w_151_172, w_151_173, w_151_176, w_151_179, w_151_180, w_151_185, w_151_186, w_151_191, w_151_193, w_151_196, w_151_199, w_151_206, w_151_207, w_151_208, w_151_214, w_151_217, w_151_231, w_151_232, w_151_233, w_151_234, w_151_237, w_151_238, w_151_239, w_151_244, w_151_245, w_151_247, w_151_251, w_151_252, w_151_254, w_151_260, w_151_264, w_151_266, w_151_271, w_151_273, w_151_275, w_151_282, w_151_283, w_151_287, w_151_291, w_151_294, w_151_295, w_151_297, w_151_298, w_151_300, w_151_303, w_151_305, w_151_309, w_151_310, w_151_311, w_151_314, w_151_317, w_151_321, w_151_322, w_151_328, w_151_338, w_151_339, w_151_346, w_151_348, w_151_350, w_151_352, w_151_357, w_151_358, w_151_359, w_151_362, w_151_363, w_151_369, w_151_380, w_151_383, w_151_388, w_151_390, w_151_394, w_151_397, w_151_403, w_151_404, w_151_406, w_151_408, w_151_410, w_151_411, w_151_412, w_151_418, w_151_424, w_151_429, w_151_431, w_151_432, w_151_439, w_151_440, w_151_446, w_151_448, w_151_450, w_151_455, w_151_459, w_151_460, w_151_461, w_151_462, w_151_464, w_151_466, w_151_469, w_151_471, w_151_473, w_151_477, w_151_479, w_151_492, w_151_503, w_151_505, w_151_507, w_151_521, w_151_527, w_151_535, w_151_541, w_151_548, w_151_549, w_151_557, w_151_558, w_151_563, w_151_567, w_151_568, w_151_571, w_151_573, w_151_574, w_151_580, w_151_582, w_151_585, w_151_596, w_151_599, w_151_602, w_151_605, w_151_608, w_151_613, w_151_621, w_151_622, w_151_625, w_151_629, w_151_631, w_151_632, w_151_634, w_151_646, w_151_648, w_151_649, w_151_653, w_151_656, w_151_662, w_151_669, w_151_671, w_151_674, w_151_679, w_151_681, w_151_683, w_151_692, w_151_694, w_151_695, w_151_703, w_151_706, w_151_718, w_151_722, w_151_724, w_151_726, w_151_732, w_151_735, w_151_736, w_151_739, w_151_741, w_151_747, w_151_754, w_151_755, w_151_760, w_151_763, w_151_765, w_151_770, w_151_776, w_151_784, w_151_790, w_151_794, w_151_795, w_151_796, w_151_799, w_151_801, w_151_808, w_151_811, w_151_812, w_151_814, w_151_815, w_151_821, w_151_822, w_151_824, w_151_827, w_151_831, w_151_835, w_151_836, w_151_837, w_151_842, w_151_851, w_151_854, w_151_862, w_151_863, w_151_869, w_151_871, w_151_874, w_151_875, w_151_876, w_151_879, w_151_890, w_151_894, w_151_898, w_151_901, w_151_905, w_151_914, w_151_916, w_151_919, w_151_922, w_151_923, w_151_926, w_151_928, w_151_929, w_151_937, w_151_941, w_151_942, w_151_943, w_151_947, w_151_953, w_151_954, w_151_955, w_151_957, w_151_959, w_151_961, w_151_962, w_151_971, w_151_978, w_151_986, w_151_987, w_151_990, w_151_998, w_151_1003, w_151_1008, w_151_1009, w_151_1010, w_151_1011, w_151_1019, w_151_1021, w_151_1026, w_151_1027, w_151_1028, w_151_1030, w_151_1032, w_151_1033, w_151_1037, w_151_1040, w_151_1041, w_151_1042, w_151_1043, w_151_1049, w_151_1053, w_151_1058, w_151_1060, w_151_1063, w_151_1068, w_151_1070, w_151_1073, w_151_1074, w_151_1077, w_151_1084, w_151_1086, w_151_1088, w_151_1092, w_151_1096, w_151_1098, w_151_1103, w_151_1105, w_151_1106, w_151_1109, w_151_1110, w_151_1114, w_151_1115, w_151_1116, w_151_1123, w_151_1124, w_151_1126, w_151_1127, w_151_1129, w_151_1132, w_151_1141, w_151_1142, w_151_1143, w_151_1150, w_151_1153, w_151_1156, w_151_1165, w_151_1168, w_151_1171, w_151_1173, w_151_1174, w_151_1175, w_151_1177, w_151_1179, w_151_1183, w_151_1187, w_151_1189, w_151_1190, w_151_1191, w_151_1194, w_151_1195, w_151_1196, w_151_1198, w_151_1202, w_151_1204, w_151_1206, w_151_1207, w_151_1211, w_151_1212, w_151_1213, w_151_1215, w_151_1216, w_151_1218, w_151_1221, w_151_1224, w_151_1225, w_151_1226, w_151_1228, w_151_1232, w_151_1235, w_151_1242, w_151_1244, w_151_1246, w_151_1248, w_151_1249, w_151_1253, w_151_1255, w_151_1259, w_151_1260, w_151_1264, w_151_1265, w_151_1266, w_151_1267, w_151_1271, w_151_1273, w_151_1274, w_151_1281, w_151_1286, w_151_1289, w_151_1291, w_151_1292, w_151_1293, w_151_1297, w_151_1299, w_151_1300, w_151_1304, w_151_1307, w_151_1312, w_151_1313, w_151_1316, w_151_1322, w_151_1324, w_151_1325, w_151_1329, w_151_1332, w_151_1333, w_151_1342, w_151_1343, w_151_1346, w_151_1352, w_151_1358, w_151_1359, w_151_1360, w_151_1364, w_151_1366, w_151_1367, w_151_1372, w_151_1376, w_151_1378, w_151_1382, w_151_1384, w_151_1385, w_151_1386, w_151_1387, w_151_1388, w_151_1394, w_151_1395, w_151_1397, w_151_1403, w_151_1404, w_151_1410, w_151_1411, w_151_1412, w_151_1415, w_151_1417, w_151_1420, w_151_1423, w_151_1425, w_151_1429, w_151_1431, w_151_1432, w_151_1434, w_151_1435, w_151_1437, w_151_1438, w_151_1442, w_151_1443, w_151_1445, w_151_1446, w_151_1449, w_151_1456, w_151_1457, w_151_1464, w_151_1466, w_151_1472, w_151_1473, w_151_1475, w_151_1477, w_151_1479, w_151_1480, w_151_1482, w_151_1484, w_151_1489, w_151_1494, w_151_1496, w_151_1497, w_151_1498, w_151_1501, w_151_1505, w_151_1510, w_151_1516, w_151_1522, w_151_1526, w_151_1528, w_151_1533, w_151_1536, w_151_1537, w_151_1542, w_151_1558, w_151_1560, w_151_1562, w_151_1564, w_151_1565, w_151_1570, w_151_1575, w_151_1576, w_151_1578, w_151_1579, w_151_1582, w_151_1583, w_151_1591, w_151_1592, w_151_1595, w_151_1596, w_151_1597, w_151_1599, w_151_1600, w_151_1601, w_151_1603, w_151_1615, w_151_1620, w_151_1633, w_151_1634, w_151_1638, w_151_1641, w_151_1647, w_151_1648, w_151_1649, w_151_1652, w_151_1653, w_151_1655, w_151_1659, w_151_1662, w_151_1664, w_151_1668, w_151_1672, w_151_1674, w_151_1676, w_151_1677, w_151_1681, w_151_1682, w_151_1689, w_151_1693, w_151_1697, w_151_1700, w_151_1701, w_151_1708, w_151_1713, w_151_1718, w_151_1719, w_151_1726, w_151_1729, w_151_1730, w_151_1731, w_151_1735, w_151_1740, w_151_1752, w_151_1753, w_151_1756, w_151_1759, w_151_1760, w_151_1763, w_151_1765, w_151_1766, w_151_1768, w_151_1770, w_151_1773, w_151_1774, w_151_1776, w_151_1781, w_151_1785, w_151_1787, w_151_1788, w_151_1789, w_151_1793, w_151_1795, w_151_1801, w_151_1806, w_151_1809, w_151_1812, w_151_1813, w_151_1816, w_151_1820, w_151_1822, w_151_1823, w_151_1826, w_151_1832, w_151_1834, w_151_1836, w_151_1838, w_151_1839, w_151_1846, w_151_1852, w_151_1855, w_151_1856, w_151_1866, w_151_1867, w_151_1868, w_151_1871, w_151_1876, w_151_1879, w_151_1881, w_151_1891, w_151_1897, w_151_1899, w_151_1906, w_151_1913, w_151_1915, w_151_1920, w_151_1923, w_151_1924, w_151_1928, w_151_1930, w_151_1934, w_151_1937, w_151_1942, w_151_1945, w_151_1946, w_151_1948, w_151_1950, w_151_1959, w_151_1960, w_151_1962, w_151_1963, w_151_1964, w_151_1965, w_151_1966, w_151_1977, w_151_1979, w_151_1981, w_151_1984, w_151_1991, w_151_1992, w_151_1995, w_151_1996, w_151_1997, w_151_1999, w_151_2002, w_151_2004, w_151_2005, w_151_2007, w_151_2008, w_151_2009, w_151_2011, w_151_2012, w_151_2014, w_151_2015, w_151_2021, w_151_2025, w_151_2030, w_151_2031, w_151_2032, w_151_2033, w_151_2040, w_151_2041, w_151_2044, w_151_2047, w_151_2048, w_151_2058, w_151_2063, w_151_2068, w_151_2069, w_151_2073, w_151_2074, w_151_2078, w_151_2083, w_151_2084, w_151_2086, w_151_2095, w_151_2103, w_151_2126, w_151_2129, w_151_2138, w_151_2151, w_151_2157, w_151_2158, w_151_2165, w_151_2172, w_151_2182, w_151_2187, w_151_2199, w_151_2207, w_151_2212, w_151_2218, w_151_2228, w_151_2229, w_151_2236, w_151_2240, w_151_2243, w_151_2251, w_151_2255, w_151_2259, w_151_2261, w_151_2265, w_151_2276, w_151_2277, w_151_2279, w_151_2283, w_151_2288, w_151_2297, w_151_2300, w_151_2307, w_151_2309, w_151_2310, w_151_2319, w_151_2320, w_151_2322, w_151_2323, w_151_2324, w_151_2336, w_151_2340, w_151_2344, w_151_2346, w_151_2348, w_151_2355, w_151_2358, w_151_2364, w_151_2366, w_151_2367, w_151_2372, w_151_2373, w_151_2378, w_151_2380, w_151_2383, w_151_2405, w_151_2410, w_151_2413, w_151_2415, w_151_2416, w_151_2418, w_151_2419, w_151_2441, w_151_2463, w_151_2468, w_151_2469, w_151_2471, w_151_2479, w_151_2483, w_151_2486, w_151_2490, w_151_2493, w_151_2495, w_151_2498, w_151_2500, w_151_2506, w_151_2508, w_151_2530, w_151_2538, w_151_2543, w_151_2548, w_151_2549, w_151_2553, w_151_2557, w_151_2563, w_151_2568, w_151_2578, w_151_2582, w_151_2591, w_151_2593, w_151_2596, w_151_2609, w_151_2619, w_151_2621, w_151_2631, w_151_2632, w_151_2636, w_151_2638, w_151_2645, w_151_2656, w_151_2665, w_151_2672, w_151_2674, w_151_2680, w_151_2686, w_151_2690, w_151_2692, w_151_2695, w_151_2701, w_151_2702, w_151_2710, w_151_2711, w_151_2714, w_151_2717, w_151_2722, w_151_2726, w_151_2727, w_151_2729, w_151_2758, w_151_2772, w_151_2774, w_151_2776, w_151_2780, w_151_2782, w_151_2789, w_151_2790, w_151_2793, w_151_2809, w_151_2821, w_151_2824, w_151_2834, w_151_2840, w_151_2845, w_151_2860, w_151_2862, w_151_2864, w_151_2872, w_151_2874, w_151_2883, w_151_2886, w_151_2894, w_151_2899, w_151_2908, w_151_2909, w_151_2913;
  wire w_152_002, w_152_003, w_152_004, w_152_006, w_152_009, w_152_010, w_152_016, w_152_017, w_152_019, w_152_026, w_152_030, w_152_037, w_152_038, w_152_039, w_152_041, w_152_046, w_152_049, w_152_053, w_152_054, w_152_056, w_152_059, w_152_062, w_152_066, w_152_070, w_152_076, w_152_078, w_152_079, w_152_080, w_152_081, w_152_083, w_152_087, w_152_092, w_152_093, w_152_095, w_152_096, w_152_100, w_152_104, w_152_105, w_152_109, w_152_110, w_152_112, w_152_119, w_152_121, w_152_122, w_152_124, w_152_134, w_152_144, w_152_148, w_152_149, w_152_150, w_152_151, w_152_157, w_152_158, w_152_160, w_152_161, w_152_163, w_152_165, w_152_166, w_152_167, w_152_170, w_152_174, w_152_175, w_152_179, w_152_181, w_152_183, w_152_184, w_152_187, w_152_189, w_152_191, w_152_192, w_152_194, w_152_198, w_152_204, w_152_213, w_152_215, w_152_219, w_152_220, w_152_225, w_152_229, w_152_235, w_152_237, w_152_238, w_152_239, w_152_240, w_152_244, w_152_245, w_152_247, w_152_251, w_152_255, w_152_256, w_152_257, w_152_259, w_152_264, w_152_266, w_152_267, w_152_271, w_152_276, w_152_277, w_152_281, w_152_286, w_152_287, w_152_290, w_152_293, w_152_299, w_152_300, w_152_302, w_152_305, w_152_306, w_152_307, w_152_310, w_152_311, w_152_313, w_152_316, w_152_317, w_152_319, w_152_320, w_152_321, w_152_322, w_152_325, w_152_327, w_152_329, w_152_331, w_152_332, w_152_343, w_152_344, w_152_346, w_152_347, w_152_351, w_152_353, w_152_354, w_152_362, w_152_372, w_152_378, w_152_380, w_152_381, w_152_382, w_152_385, w_152_386, w_152_388, w_152_389, w_152_395, w_152_398, w_152_402, w_152_404, w_152_409, w_152_410, w_152_412, w_152_413, w_152_416, w_152_419, w_152_423, w_152_430, w_152_431, w_152_434, w_152_436, w_152_438, w_152_440, w_152_444, w_152_448, w_152_454, w_152_456, w_152_459, w_152_461, w_152_462, w_152_468, w_152_470, w_152_471, w_152_474, w_152_475, w_152_476, w_152_483, w_152_484, w_152_486, w_152_490, w_152_496, w_152_498, w_152_504, w_152_505, w_152_510, w_152_514, w_152_515, w_152_519, w_152_521, w_152_523, w_152_529, w_152_530, w_152_532, w_152_535, w_152_536, w_152_538, w_152_539, w_152_544, w_152_548, w_152_555, w_152_556, w_152_560, w_152_562, w_152_569, w_152_571, w_152_572, w_152_574, w_152_575, w_152_578, w_152_580, w_152_583, w_152_590, w_152_591, w_152_592, w_152_597, w_152_600, w_152_602, w_152_603, w_152_608, w_152_610, w_152_615, w_152_617, w_152_619, w_152_625, w_152_626, w_152_629, w_152_630, w_152_632, w_152_634, w_152_638, w_152_640, w_152_641, w_152_642, w_152_643, w_152_644, w_152_645, w_152_647, w_152_648, w_152_650, w_152_652, w_152_653, w_152_656, w_152_657, w_152_665, w_152_666, w_152_668, w_152_669, w_152_673, w_152_674, w_152_680, w_152_693, w_152_695, w_152_696, w_152_699, w_152_701, w_152_702, w_152_705, w_152_710, w_152_711, w_152_714, w_152_718, w_152_719, w_152_727, w_152_729, w_152_730, w_152_735, w_152_741, w_152_742, w_152_754, w_152_756, w_152_757, w_152_763, w_152_765, w_152_768, w_152_769, w_152_772, w_152_773, w_152_775, w_152_776, w_152_779, w_152_782, w_152_788, w_152_795, w_152_801, w_152_802, w_152_803, w_152_807, w_152_813, w_152_814, w_152_816, w_152_820, w_152_825, w_152_829, w_152_831, w_152_832, w_152_837, w_152_839, w_152_847, w_152_849, w_152_850, w_152_854, w_152_855, w_152_856, w_152_862, w_152_864, w_152_865, w_152_871, w_152_874, w_152_876, w_152_877, w_152_878, w_152_880, w_152_884, w_152_901, w_152_902, w_152_905, w_152_908, w_152_909, w_152_910, w_152_912, w_152_917, w_152_926, w_152_934, w_152_941, w_152_942, w_152_944, w_152_946, w_152_952, w_152_958, w_152_959, w_152_968, w_152_970, w_152_972, w_152_974, w_152_977, w_152_979, w_152_983, w_152_984, w_152_987, w_152_988, w_152_992, w_152_993, w_152_994, w_152_997, w_152_1001, w_152_1002, w_152_1004, w_152_1011, w_152_1014, w_152_1016, w_152_1018, w_152_1021, w_152_1026, w_152_1029, w_152_1031, w_152_1032, w_152_1037, w_152_1038, w_152_1041, w_152_1049, w_152_1067, w_152_1068, w_152_1069, w_152_1072, w_152_1074, w_152_1078, w_152_1093, w_152_1106, w_152_1109, w_152_1110, w_152_1112, w_152_1117, w_152_1118, w_152_1119, w_152_1123, w_152_1136, w_152_1137, w_152_1142, w_152_1145, w_152_1147, w_152_1150, w_152_1153, w_152_1158, w_152_1159, w_152_1160, w_152_1163, w_152_1164, w_152_1167, w_152_1168, w_152_1171, w_152_1176, w_152_1177, w_152_1179, w_152_1182, w_152_1183, w_152_1187, w_152_1190, w_152_1192, w_152_1194, w_152_1195, w_152_1197, w_152_1201, w_152_1209, w_152_1212, w_152_1216, w_152_1217, w_152_1221, w_152_1222, w_152_1231, w_152_1233, w_152_1236, w_152_1243, w_152_1247, w_152_1248, w_152_1249, w_152_1253, w_152_1258, w_152_1262, w_152_1266, w_152_1268, w_152_1269, w_152_1270, w_152_1274, w_152_1284, w_152_1285, w_152_1288, w_152_1292, w_152_1293, w_152_1297, w_152_1298, w_152_1301, w_152_1305, w_152_1315, w_152_1316, w_152_1317, w_152_1318, w_152_1321, w_152_1322, w_152_1327, w_152_1328, w_152_1329, w_152_1336, w_152_1342, w_152_1344, w_152_1346, w_152_1349, w_152_1350, w_152_1354, w_152_1359, w_152_1368, w_152_1383, w_152_1386, w_152_1388, w_152_1390, w_152_1391, w_152_1396, w_152_1398, w_152_1399, w_152_1406, w_152_1410, w_152_1415, w_152_1418, w_152_1419, w_152_1426, w_152_1427, w_152_1428, w_152_1432, w_152_1437, w_152_1438, w_152_1441, w_152_1442, w_152_1445, w_152_1451, w_152_1460, w_152_1461, w_152_1463, w_152_1472, w_152_1473, w_152_1475, w_152_1476, w_152_1479, w_152_1482, w_152_1483, w_152_1484, w_152_1488, w_152_1497, w_152_1499, w_152_1501, w_152_1510, w_152_1515, w_152_1519, w_152_1520, w_152_1523, w_152_1524, w_152_1527, w_152_1531, w_152_1535, w_152_1538, w_152_1542, w_152_1544, w_152_1545, w_152_1547, w_152_1549, w_152_1551, w_152_1552, w_152_1556, w_152_1564, w_152_1566, w_152_1575, w_152_1579, w_152_1580, w_152_1582, w_152_1587, w_152_1590, w_152_1591, w_152_1599, w_152_1601, w_152_1608, w_152_1610, w_152_1614, w_152_1618, w_152_1623, w_152_1627, w_152_1628, w_152_1630, w_152_1631, w_152_1635, w_152_1637, w_152_1643, w_152_1648, w_152_1652, w_152_1654, w_152_1656, w_152_1663, w_152_1665, w_152_1670, w_152_1671, w_152_1673, w_152_1674, w_152_1678, w_152_1680, w_152_1685, w_152_1686, w_152_1688, w_152_1691, w_152_1693, w_152_1697, w_152_1698, w_152_1701, w_152_1707, w_152_1708, w_152_1709, w_152_1711, w_152_1716, w_152_1717, w_152_1720, w_152_1723, w_152_1724, w_152_1725, w_152_1729, w_152_1734, w_152_1735, w_152_1738, w_152_1741, w_152_1745, w_152_1750, w_152_1751, w_152_1753, w_152_1754, w_152_1755, w_152_1770, w_152_1771, w_152_1773, w_152_1775, w_152_1776, w_152_1778, w_152_1780, w_152_1784, w_152_1786, w_152_1787, w_152_1788, w_152_1790, w_152_1791, w_152_1793, w_152_1794, w_152_1795, w_152_1796, w_152_1801, w_152_1804, w_152_1807, w_152_1811, w_152_1813, w_152_1814, w_152_1823, w_152_1827, w_152_1831, w_152_1833, w_152_1834, w_152_1835, w_152_1837, w_152_1842, w_152_1845, w_152_1851, w_152_1852, w_152_1859, w_152_1861, w_152_1862, w_152_1867, w_152_1868, w_152_1870, w_152_1873, w_152_1874, w_152_1875, w_152_1878, w_152_1880, w_152_1882, w_152_1883, w_152_1885, w_152_1887, w_152_1893, w_152_1895, w_152_1897, w_152_1912, w_152_1913, w_152_1923, w_152_1925, w_152_1931, w_152_1937, w_152_1940, w_152_1941, w_152_1950, w_152_1954, w_152_1956, w_152_1971, w_152_1978, w_152_1984, w_152_1994, w_152_1998, w_152_2002, w_152_2006, w_152_2014, w_152_2017, w_152_2018, w_152_2033, w_152_2046, w_152_2058, w_152_2067, w_152_2068, w_152_2069, w_152_2074, w_152_2086, w_152_2088, w_152_2096, w_152_2101, w_152_2104, w_152_2113, w_152_2115, w_152_2124, w_152_2133, w_152_2145, w_152_2146, w_152_2152, w_152_2158, w_152_2169, w_152_2171, w_152_2178, w_152_2196, w_152_2199, w_152_2207, w_152_2234, w_152_2252, w_152_2258, w_152_2259, w_152_2263, w_152_2278, w_152_2295, w_152_2299, w_152_2311, w_152_2312, w_152_2321, w_152_2325, w_152_2335, w_152_2338, w_152_2340, w_152_2342, w_152_2352, w_152_2356, w_152_2357, w_152_2367, w_152_2376, w_152_2380, w_152_2382, w_152_2390, w_152_2393, w_152_2395, w_152_2397, w_152_2401, w_152_2402, w_152_2411, w_152_2413, w_152_2420, w_152_2426, w_152_2440, w_152_2441, w_152_2444, w_152_2446, w_152_2448, w_152_2452, w_152_2461, w_152_2462, w_152_2467, w_152_2471, w_152_2479, w_152_2482, w_152_2484, w_152_2490, w_152_2495, w_152_2496, w_152_2498, w_152_2505, w_152_2531, w_152_2547, w_152_2551, w_152_2556, w_152_2571, w_152_2581, w_152_2582, w_152_2593, w_152_2595, w_152_2596, w_152_2601, w_152_2605, w_152_2613, w_152_2615, w_152_2633, w_152_2657, w_152_2663, w_152_2665, w_152_2674, w_152_2682, w_152_2689, w_152_2690, w_152_2700, w_152_2701, w_152_2705, w_152_2707, w_152_2721, w_152_2724, w_152_2729, w_152_2730, w_152_2750, w_152_2751, w_152_2755, w_152_2765, w_152_2775, w_152_2776, w_152_2781, w_152_2789, w_152_2806, w_152_2826, w_152_2841, w_152_2844, w_152_2858, w_152_2859, w_152_2869, w_152_2876, w_152_2877, w_152_2883, w_152_2907, w_152_2919, w_152_2922, w_152_2931, w_152_2937, w_152_2942, w_152_2951, w_152_2955, w_152_2958, w_152_2975, w_152_2990, w_152_2996, w_152_3007, w_152_3023, w_152_3024, w_152_3035, w_152_3038, w_152_3046, w_152_3047, w_152_3055, w_152_3056, w_152_3057, w_152_3058, w_152_3059, w_152_3060, w_152_3061, w_152_3062, w_152_3063, w_152_3065, w_152_3067, w_152_3068, w_152_3069, w_152_3070, w_152_3071, w_152_3072, w_152_3073, w_152_3074, w_152_3075, w_152_3076, w_152_3077, w_152_3078;
  wire w_153_000, w_153_006, w_153_008, w_153_010, w_153_013, w_153_015, w_153_016, w_153_018, w_153_019, w_153_023, w_153_024, w_153_032, w_153_033, w_153_037, w_153_039, w_153_040, w_153_041, w_153_042, w_153_043, w_153_049, w_153_052, w_153_053, w_153_064, w_153_067, w_153_069, w_153_071, w_153_074, w_153_086, w_153_093, w_153_122, w_153_126, w_153_131, w_153_136, w_153_145, w_153_157, w_153_174, w_153_183, w_153_185, w_153_196, w_153_200, w_153_201, w_153_203, w_153_205, w_153_208, w_153_215, w_153_217, w_153_223, w_153_224, w_153_228, w_153_232, w_153_233, w_153_236, w_153_246, w_153_251, w_153_260, w_153_263, w_153_264, w_153_265, w_153_266, w_153_270, w_153_276, w_153_286, w_153_290, w_153_306, w_153_311, w_153_312, w_153_313, w_153_321, w_153_335, w_153_337, w_153_338, w_153_339, w_153_341, w_153_343, w_153_346, w_153_347, w_153_350, w_153_352, w_153_357, w_153_364, w_153_375, w_153_381, w_153_383, w_153_388, w_153_393, w_153_394, w_153_399, w_153_413, w_153_420, w_153_425, w_153_431, w_153_432, w_153_434, w_153_465, w_153_467, w_153_484, w_153_493, w_153_494, w_153_502, w_153_511, w_153_512, w_153_518, w_153_531, w_153_534, w_153_543, w_153_546, w_153_551, w_153_556, w_153_557, w_153_561, w_153_565, w_153_568, w_153_580, w_153_582, w_153_592, w_153_597, w_153_598, w_153_601, w_153_604, w_153_610, w_153_621, w_153_627, w_153_633, w_153_638, w_153_650, w_153_651, w_153_663, w_153_666, w_153_667, w_153_670, w_153_684, w_153_686, w_153_692, w_153_699, w_153_706, w_153_714, w_153_715, w_153_716, w_153_717, w_153_718, w_153_727, w_153_733, w_153_735, w_153_752, w_153_774, w_153_779, w_153_787, w_153_789, w_153_791, w_153_792, w_153_793, w_153_794, w_153_798, w_153_804, w_153_806, w_153_816, w_153_819, w_153_823, w_153_825, w_153_828, w_153_832, w_153_836, w_153_839, w_153_840, w_153_852, w_153_873, w_153_875, w_153_881, w_153_886, w_153_896, w_153_899, w_153_915, w_153_917, w_153_919, w_153_920, w_153_926, w_153_929, w_153_956, w_153_972, w_153_977, w_153_980, w_153_988, w_153_991, w_153_994, w_153_997, w_153_998, w_153_1000, w_153_1003, w_153_1019, w_153_1025, w_153_1031, w_153_1034, w_153_1035, w_153_1039, w_153_1043, w_153_1045, w_153_1057, w_153_1063, w_153_1065, w_153_1067, w_153_1068, w_153_1075, w_153_1084, w_153_1088, w_153_1089, w_153_1094, w_153_1100, w_153_1106, w_153_1113, w_153_1120, w_153_1121, w_153_1125, w_153_1131, w_153_1133, w_153_1138, w_153_1139, w_153_1140, w_153_1147, w_153_1155, w_153_1160, w_153_1175, w_153_1179, w_153_1200, w_153_1204, w_153_1207, w_153_1215, w_153_1216, w_153_1220, w_153_1227, w_153_1230, w_153_1231, w_153_1232, w_153_1235, w_153_1238, w_153_1241, w_153_1251, w_153_1264, w_153_1265, w_153_1266, w_153_1267, w_153_1269, w_153_1277, w_153_1285, w_153_1286, w_153_1289, w_153_1291, w_153_1292, w_153_1298, w_153_1299, w_153_1302, w_153_1303, w_153_1305, w_153_1315, w_153_1317, w_153_1334, w_153_1337, w_153_1341, w_153_1342, w_153_1346, w_153_1354, w_153_1358, w_153_1367, w_153_1368, w_153_1371, w_153_1372, w_153_1392, w_153_1394, w_153_1400, w_153_1401, w_153_1402, w_153_1406, w_153_1410, w_153_1416, w_153_1423, w_153_1437, w_153_1443, w_153_1447, w_153_1448, w_153_1451, w_153_1457, w_153_1462, w_153_1469, w_153_1483, w_153_1485, w_153_1496, w_153_1497, w_153_1507, w_153_1520, w_153_1521, w_153_1525, w_153_1526, w_153_1531, w_153_1539, w_153_1540, w_153_1542, w_153_1550, w_153_1556, w_153_1564, w_153_1569, w_153_1571, w_153_1578, w_153_1580, w_153_1623, w_153_1641, w_153_1644, w_153_1653, w_153_1654, w_153_1657, w_153_1671, w_153_1676, w_153_1694, w_153_1704, w_153_1705, w_153_1706, w_153_1707, w_153_1713, w_153_1719, w_153_1720, w_153_1725, w_153_1727, w_153_1743, w_153_1746, w_153_1754, w_153_1758, w_153_1760, w_153_1769, w_153_1772, w_153_1778, w_153_1797, w_153_1800, w_153_1802, w_153_1804, w_153_1825, w_153_1826, w_153_1829, w_153_1830, w_153_1837, w_153_1839, w_153_1841, w_153_1842, w_153_1844, w_153_1846, w_153_1849, w_153_1852, w_153_1854, w_153_1856, w_153_1863, w_153_1868, w_153_1869, w_153_1870, w_153_1873, w_153_1874, w_153_1876, w_153_1878, w_153_1893, w_153_1906, w_153_1910, w_153_1917, w_153_1921, w_153_1925, w_153_1926, w_153_1935, w_153_1937, w_153_1949, w_153_1951, w_153_1959, w_153_1976, w_153_1978, w_153_1983, w_153_1987, w_153_1988, w_153_2001, w_153_2013, w_153_2016, w_153_2022, w_153_2023, w_153_2031, w_153_2032, w_153_2037, w_153_2045, w_153_2057, w_153_2060, w_153_2066, w_153_2079, w_153_2089, w_153_2093, w_153_2098, w_153_2107, w_153_2109, w_153_2110, w_153_2120, w_153_2125, w_153_2129, w_153_2132, w_153_2134, w_153_2142, w_153_2143, w_153_2145, w_153_2154, w_153_2162, w_153_2173, w_153_2175, w_153_2177, w_153_2181, w_153_2188, w_153_2189, w_153_2194, w_153_2195, w_153_2196, w_153_2218, w_153_2226, w_153_2228, w_153_2235, w_153_2243, w_153_2248, w_153_2251, w_153_2257, w_153_2265, w_153_2266, w_153_2272, w_153_2280, w_153_2296, w_153_2300, w_153_2313, w_153_2325, w_153_2326, w_153_2327, w_153_2337, w_153_2352, w_153_2354, w_153_2366, w_153_2369, w_153_2386, w_153_2399, w_153_2402, w_153_2404, w_153_2406, w_153_2408, w_153_2409, w_153_2417, w_153_2432, w_153_2451, w_153_2456, w_153_2461, w_153_2469, w_153_2475, w_153_2476, w_153_2486, w_153_2488, w_153_2499, w_153_2501, w_153_2504, w_153_2507, w_153_2515, w_153_2518, w_153_2522, w_153_2526, w_153_2530, w_153_2532, w_153_2533, w_153_2542, w_153_2544, w_153_2550, w_153_2568, w_153_2570, w_153_2581, w_153_2593, w_153_2604, w_153_2613, w_153_2618, w_153_2621, w_153_2624, w_153_2637, w_153_2639, w_153_2640, w_153_2668, w_153_2686, w_153_2697, w_153_2704, w_153_2705, w_153_2708, w_153_2712, w_153_2716, w_153_2722, w_153_2727, w_153_2749, w_153_2751, w_153_2756, w_153_2765, w_153_2767, w_153_2770, w_153_2786, w_153_2791, w_153_2794, w_153_2805, w_153_2807, w_153_2811, w_153_2812, w_153_2822, w_153_2823, w_153_2835, w_153_2845, w_153_2847, w_153_2848, w_153_2854, w_153_2857, w_153_2876, w_153_2886, w_153_2889, w_153_2891, w_153_2892, w_153_2895, w_153_2898, w_153_2903, w_153_2910, w_153_2923, w_153_2946, w_153_2950, w_153_2952, w_153_2960, w_153_2965, w_153_2968, w_153_2970, w_153_2982, w_153_2984, w_153_2985, w_153_2986, w_153_2995, w_153_3006, w_153_3007, w_153_3008, w_153_3010, w_153_3014, w_153_3015, w_153_3024, w_153_3041, w_153_3053, w_153_3054, w_153_3067, w_153_3069, w_153_3074, w_153_3080, w_153_3081, w_153_3090, w_153_3093, w_153_3114, w_153_3117, w_153_3122, w_153_3124, w_153_3126, w_153_3127, w_153_3128, w_153_3132, w_153_3135, w_153_3137, w_153_3138, w_153_3141, w_153_3152, w_153_3154, w_153_3156, w_153_3157, w_153_3163, w_153_3182, w_153_3183, w_153_3188, w_153_3195, w_153_3197, w_153_3198, w_153_3203, w_153_3205, w_153_3211, w_153_3220, w_153_3221, w_153_3225, w_153_3234, w_153_3240, w_153_3247, w_153_3248, w_153_3262, w_153_3263, w_153_3266, w_153_3267, w_153_3272, w_153_3274, w_153_3277, w_153_3279, w_153_3281, w_153_3282, w_153_3283, w_153_3285, w_153_3294, w_153_3297, w_153_3301, w_153_3304, w_153_3313, w_153_3318, w_153_3319, w_153_3325, w_153_3328, w_153_3352, w_153_3362, w_153_3375, w_153_3377, w_153_3385, w_153_3389, w_153_3415, w_153_3426, w_153_3432, w_153_3452, w_153_3454, w_153_3455, w_153_3462, w_153_3465, w_153_3472, w_153_3483, w_153_3489, w_153_3492, w_153_3493, w_153_3494, w_153_3496, w_153_3497, w_153_3499, w_153_3500, w_153_3503, w_153_3504, w_153_3511, w_153_3517, w_153_3520, w_153_3521, w_153_3527, w_153_3530, w_153_3533, w_153_3534, w_153_3539, w_153_3557, w_153_3566, w_153_3582, w_153_3588, w_153_3589, w_153_3590, w_153_3596, w_153_3599, w_153_3602, w_153_3607, w_153_3609, w_153_3621, w_153_3622, w_153_3623, w_153_3625, w_153_3626, w_153_3629, w_153_3638, w_153_3639, w_153_3657, w_153_3659, w_153_3660, w_153_3661, w_153_3662, w_153_3667, w_153_3674, w_153_3677, w_153_3681, w_153_3686, w_153_3690, w_153_3705, w_153_3710, w_153_3711, w_153_3720, w_153_3729, w_153_3737, w_153_3745, w_153_3756, w_153_3765, w_153_3776, w_153_3783, w_153_3786, w_153_3790, w_153_3794, w_153_3797, w_153_3801, w_153_3806, w_153_3818, w_153_3819, w_153_3821, w_153_3826, w_153_3834, w_153_3835, w_153_3836, w_153_3846, w_153_3847, w_153_3851, w_153_3853, w_153_3862, w_153_3884, w_153_3894, w_153_3898, w_153_3899, w_153_3901, w_153_3905, w_153_3908, w_153_3919, w_153_3922, w_153_3925, w_153_3930, w_153_3935, w_153_3939, w_153_3945, w_153_3950, w_153_3957, w_153_3962, w_153_3969, w_153_3970, w_153_3974, w_153_3979, w_153_3981, w_153_3984, w_153_3990, w_153_3992, w_153_3994, w_153_4000, w_153_4003, w_153_4010, w_153_4011, w_153_4014, w_153_4016, w_153_4022, w_153_4028, w_153_4031, w_153_4036, w_153_4041, w_153_4042, w_153_4045, w_153_4047, w_153_4056, w_153_4064, w_153_4069, w_153_4077, w_153_4080, w_153_4082, w_153_4093, w_153_4101, w_153_4102, w_153_4105, w_153_4113, w_153_4115, w_153_4121, w_153_4125, w_153_4132, w_153_4138, w_153_4145, w_153_4155, w_153_4169, w_153_4173, w_153_4182, w_153_4195, w_153_4198, w_153_4210, w_153_4213, w_153_4214, w_153_4218, w_153_4222, w_153_4230, w_153_4237, w_153_4238, w_153_4240, w_153_4246, w_153_4247, w_153_4263, w_153_4286, w_153_4289, w_153_4290, w_153_4291, w_153_4294, w_153_4298, w_153_4300, w_153_4303, w_153_4317, w_153_4318, w_153_4321, w_153_4322, w_153_4326, w_153_4335, w_153_4354, w_153_4359, w_153_4365, w_153_4367, w_153_4369, w_153_4370, w_153_4371, w_153_4375, w_153_4382, w_153_4386, w_153_4390, w_153_4398, w_153_4400, w_153_4415, w_153_4417, w_153_4421, w_153_4432, w_153_4434, w_153_4435, w_153_4444, w_153_4447, w_153_4454, w_153_4458, w_153_4467, w_153_4469, w_153_4476, w_153_4482, w_153_4485, w_153_4487, w_153_4496, w_153_4505, w_153_4516, w_153_4518, w_153_4522, w_153_4528, w_153_4534, w_153_4539, w_153_4540, w_153_4565, w_153_4566, w_153_4571, w_153_4574, w_153_4575, w_153_4589, w_153_4591, w_153_4600, w_153_4606, w_153_4610, w_153_4611, w_153_4615, w_153_4628, w_153_4632, w_153_4635, w_153_4638, w_153_4640, w_153_4641, w_153_4645, w_153_4647, w_153_4650, w_153_4661, w_153_4664, w_153_4668, w_153_4671, w_153_4675, w_153_4680, w_153_4686, w_153_4702, w_153_4706, w_153_4709, w_153_4712, w_153_4713, w_153_4722, w_153_4723, w_153_4727, w_153_4730, w_153_4732, w_153_4755, w_153_4764, w_153_4765, w_153_4766, w_153_4768, w_153_4775, w_153_4776, w_153_4792, w_153_4806, w_153_4814, w_153_4817, w_153_4818, w_153_4819, w_153_4821, w_153_4822, w_153_4826, w_153_4831, w_153_4842, w_153_4843, w_153_4861, w_153_4862, w_153_4878, w_153_4880, w_153_4886, w_153_4895, w_153_4896, w_153_4920, w_153_4926, w_153_4935;
  wire w_154_002, w_154_005, w_154_007, w_154_013, w_154_014, w_154_016, w_154_020, w_154_025, w_154_027, w_154_032, w_154_034, w_154_035, w_154_036, w_154_037, w_154_038, w_154_039, w_154_040, w_154_044, w_154_045, w_154_047, w_154_048, w_154_049, w_154_051, w_154_061, w_154_067, w_154_070, w_154_071, w_154_072, w_154_073, w_154_074, w_154_077, w_154_078, w_154_079, w_154_080, w_154_081, w_154_084, w_154_085, w_154_088, w_154_089, w_154_090, w_154_094, w_154_095, w_154_096, w_154_097, w_154_102, w_154_104, w_154_105, w_154_106, w_154_109, w_154_110, w_154_113, w_154_118, w_154_120, w_154_122, w_154_125, w_154_127, w_154_128, w_154_129, w_154_132, w_154_135, w_154_136, w_154_139, w_154_140, w_154_142, w_154_144, w_154_145, w_154_146, w_154_148, w_154_150, w_154_151, w_154_152, w_154_153, w_154_154, w_154_157, w_154_158, w_154_159, w_154_164, w_154_168, w_154_170, w_154_172, w_154_174, w_154_177, w_154_179, w_154_181, w_154_182, w_154_184, w_154_185, w_154_186, w_154_187, w_154_188, w_154_190, w_154_193, w_154_195, w_154_197, w_154_200, w_154_201, w_154_202, w_154_203, w_154_204, w_154_209, w_154_213, w_154_215, w_154_218, w_154_219, w_154_222, w_154_223, w_154_224, w_154_225, w_154_228, w_154_229, w_154_230, w_154_232, w_154_234, w_154_236, w_154_237, w_154_242, w_154_251, w_154_252, w_154_254, w_154_256, w_154_258, w_154_260, w_154_262, w_154_263, w_154_264, w_154_265, w_154_266, w_154_267, w_154_268, w_154_269, w_154_272, w_154_274, w_154_278, w_154_279, w_154_285, w_154_289, w_154_291, w_154_297, w_154_302, w_154_303, w_154_305, w_154_308, w_154_311, w_154_313, w_154_317, w_154_321, w_154_323, w_154_324, w_154_326, w_154_327, w_154_333, w_154_338, w_154_342, w_154_343, w_154_345, w_154_350, w_154_352, w_154_354, w_154_356, w_154_357, w_154_360, w_154_362, w_154_365, w_154_368, w_154_370, w_154_373, w_154_374, w_154_375, w_154_377, w_154_378, w_154_380, w_154_382, w_154_385, w_154_386, w_154_394, w_154_395, w_154_397, w_154_398, w_154_400, w_154_402, w_154_405, w_154_407, w_154_409, w_154_413, w_154_414, w_154_415, w_154_417, w_154_419, w_154_422, w_154_423, w_154_425, w_154_426, w_154_428, w_154_429, w_154_430, w_154_434, w_154_435, w_154_436, w_154_438, w_154_439, w_154_440, w_154_444, w_154_447, w_154_448, w_154_451, w_154_452, w_154_458, w_154_462, w_154_463, w_154_464, w_154_466, w_154_467, w_154_469, w_154_471, w_154_472, w_154_473, w_154_474, w_154_475, w_154_477, w_154_478, w_154_481, w_154_482, w_154_483, w_154_491, w_154_494, w_154_495, w_154_496, w_154_498, w_154_499, w_154_501, w_154_504, w_154_506, w_154_508, w_154_509, w_154_513, w_154_514, w_154_516, w_154_517, w_154_519, w_154_521, w_154_523, w_154_525, w_154_526, w_154_533, w_154_537, w_154_538, w_154_540, w_154_543, w_154_546, w_154_548, w_154_551, w_154_556, w_154_558, w_154_562, w_154_563, w_154_567, w_154_568, w_154_569, w_154_573, w_154_574, w_154_575, w_154_579, w_154_580, w_154_581, w_154_582, w_154_583, w_154_584, w_154_588, w_154_590, w_154_591, w_154_593, w_154_597, w_154_598, w_154_601, w_154_603, w_154_605, w_154_607, w_154_608, w_154_609, w_154_617, w_154_618, w_154_619, w_154_622, w_154_623, w_154_626, w_154_631, w_154_632, w_154_634, w_154_637, w_154_639, w_154_642, w_154_643, w_154_648, w_154_649, w_154_654, w_154_658, w_154_660, w_154_661, w_154_662, w_154_663, w_154_664, w_154_667, w_154_668, w_154_669, w_154_675, w_154_677, w_154_678, w_154_679, w_154_683, w_154_688, w_154_696, w_154_697, w_154_700, w_154_702, w_154_705, w_154_706, w_154_709, w_154_711, w_154_712, w_154_713, w_154_716, w_154_719, w_154_721, w_154_724, w_154_725, w_154_729, w_154_730, w_154_731, w_154_733, w_154_734, w_154_735, w_154_737, w_154_739, w_154_740, w_154_741, w_154_742, w_154_743, w_154_744, w_154_745, w_154_746, w_154_753, w_154_756, w_154_757, w_154_758, w_154_759, w_154_760, w_154_762, w_154_764, w_154_765, w_154_766, w_154_768, w_154_771, w_154_772, w_154_775, w_154_781, w_154_782, w_154_784, w_154_787, w_154_788, w_154_789, w_154_790, w_154_796, w_154_798, w_154_800, w_154_801, w_154_804, w_154_807, w_154_808, w_154_809, w_154_810, w_154_811, w_154_812, w_154_813, w_154_815, w_154_816, w_154_818, w_154_823, w_154_824, w_154_825, w_154_829, w_154_836, w_154_842, w_154_849, w_154_850, w_154_853, w_154_855, w_154_856, w_154_858, w_154_860, w_154_862, w_154_866, w_154_867, w_154_869, w_154_871, w_154_874, w_154_878, w_154_880, w_154_882, w_154_885, w_154_886, w_154_887, w_154_888, w_154_892, w_154_893, w_154_897, w_154_898, w_154_900, w_154_902, w_154_904, w_154_909, w_154_911, w_154_913, w_154_914, w_154_915, w_154_917, w_154_918, w_154_924, w_154_930, w_154_932, w_154_934, w_154_935, w_154_938, w_154_939, w_154_942, w_154_943, w_154_946, w_154_952, w_154_957, w_154_962, w_154_963, w_154_964, w_154_968, w_154_975, w_154_976, w_154_979, w_154_989, w_154_990, w_154_992, w_154_993, w_154_994, w_154_998, w_154_1000, w_154_1003, w_154_1006, w_154_1011, w_154_1016, w_154_1017, w_154_1018, w_154_1019, w_154_1022, w_154_1023, w_154_1025, w_154_1026, w_154_1028, w_154_1029, w_154_1030, w_154_1032, w_154_1037, w_154_1043, w_154_1046, w_154_1047, w_154_1050, w_154_1051, w_154_1053, w_154_1054, w_154_1056, w_154_1061, w_154_1063, w_154_1065, w_154_1066, w_154_1069, w_154_1071, w_154_1072, w_154_1073, w_154_1076, w_154_1081, w_154_1082, w_154_1085, w_154_1088, w_154_1093, w_154_1098, w_154_1099, w_154_1102, w_154_1104, w_154_1106, w_154_1107, w_154_1112, w_154_1114, w_154_1115, w_154_1116, w_154_1124, w_154_1126, w_154_1127, w_154_1128, w_154_1131, w_154_1132, w_154_1133, w_154_1134, w_154_1135, w_154_1139, w_154_1141, w_154_1143, w_154_1144, w_154_1147, w_154_1150, w_154_1152, w_154_1153, w_154_1158, w_154_1159, w_154_1160, w_154_1161, w_154_1163, w_154_1165, w_154_1167, w_154_1168, w_154_1169, w_154_1171, w_154_1177, w_154_1178, w_154_1179, w_154_1180, w_154_1184, w_154_1185, w_154_1190, w_154_1191, w_154_1195, w_154_1202, w_154_1205, w_154_1207, w_154_1208, w_154_1210, w_154_1212, w_154_1213, w_154_1220, w_154_1231, w_154_1232, w_154_1236, w_154_1240, w_154_1244, w_154_1248, w_154_1249, w_154_1254, w_154_1258, w_154_1259, w_154_1260, w_154_1261, w_154_1266, w_154_1268, w_154_1269, w_154_1275, w_154_1277, w_154_1279, w_154_1283, w_154_1284, w_154_1293, w_154_1297, w_154_1300, w_154_1302, w_154_1306, w_154_1310, w_154_1311, w_154_1312, w_154_1313, w_154_1316, w_154_1319, w_154_1320, w_154_1322, w_154_1323, w_154_1327, w_154_1330, w_154_1335, w_154_1337, w_154_1343, w_154_1345, w_154_1348, w_154_1350, w_154_1351, w_154_1354, w_154_1360, w_154_1362, w_154_1364, w_154_1365, w_154_1367, w_154_1368, w_154_1369, w_154_1370, w_154_1372, w_154_1374, w_154_1376, w_154_1377, w_154_1379, w_154_1381, w_154_1384, w_154_1388, w_154_1391, w_154_1392, w_154_1396, w_154_1398, w_154_1399, w_154_1403, w_154_1404, w_154_1408, w_154_1411, w_154_1414, w_154_1415, w_154_1416, w_154_1418, w_154_1422, w_154_1424, w_154_1426, w_154_1430, w_154_1431, w_154_1436, w_154_1437, w_154_1438, w_154_1439, w_154_1445, w_154_1449, w_154_1452, w_154_1454, w_154_1457, w_154_1458, w_154_1459, w_154_1461, w_154_1463, w_154_1465, w_154_1466, w_154_1469, w_154_1471, w_154_1475, w_154_1476, w_154_1477, w_154_1482, w_154_1487, w_154_1490, w_154_1503, w_154_1504, w_154_1505, w_154_1507, w_154_1511, w_154_1512, w_154_1519, w_154_1520, w_154_1522, w_154_1532, w_154_1533, w_154_1536, w_154_1541, w_154_1542, w_154_1544, w_154_1546, w_154_1550, w_154_1551, w_154_1552, w_154_1553, w_154_1558, w_154_1564, w_154_1566, w_154_1569, w_154_1572, w_154_1574, w_154_1575, w_154_1577, w_154_1578, w_154_1581, w_154_1583, w_154_1585, w_154_1589, w_154_1590, w_154_1591, w_154_1592, w_154_1595, w_154_1601, w_154_1606, w_154_1610, w_154_1612, w_154_1615, w_154_1617, w_154_1620, w_154_1621, w_154_1624, w_154_1627, w_154_1631, w_154_1638, w_154_1640, w_154_1645, w_154_1646, w_154_1648, w_154_1649, w_154_1656, w_154_1660, w_154_1662, w_154_1666, w_154_1673, w_154_1676, w_154_1677, w_154_1680, w_154_1682, w_154_1683, w_154_1685, w_154_1686, w_154_1693, w_154_1696, w_154_1700, w_154_1707, w_154_1710, w_154_1711, w_154_1712, w_154_1713, w_154_1714, w_154_1716, w_154_1720, w_154_1724, w_154_1725, w_154_1726, w_154_1730, w_154_1737, w_154_1738, w_154_1741, w_154_1744, w_154_1745, w_154_1750, w_154_1753, w_154_1760, w_154_1766, w_154_1770, w_154_1771, w_154_1774, w_154_1777, w_154_1786, w_154_1793, w_154_1797, w_154_1800, w_154_1802, w_154_1804, w_154_1806, w_154_1808, w_154_1816, w_154_1819, w_154_1823, w_154_1827, w_154_1829, w_154_1832, w_154_1835, w_154_1836, w_154_1838, w_154_1841, w_154_1842, w_154_1844, w_154_1847, w_154_1850, w_154_1851, w_154_1852, w_154_1853, w_154_1855, w_154_1856, w_154_1861, w_154_1862, w_154_1869, w_154_1870, w_154_1873, w_154_1876, w_154_1879, w_154_1888, w_154_1890;
  wire w_155_000, w_155_001, w_155_002, w_155_003, w_155_004, w_155_005, w_155_006;
  wire w_156_000, w_156_001, w_156_002, w_156_003, w_156_005, w_156_006, w_156_007, w_156_010, w_156_012, w_156_014, w_156_016, w_156_017, w_156_019, w_156_020, w_156_021, w_156_023, w_156_024, w_156_027, w_156_029, w_156_031, w_156_036, w_156_039, w_156_040, w_156_042, w_156_045, w_156_046, w_156_047, w_156_048, w_156_049, w_156_056, w_156_057, w_156_060, w_156_062, w_156_063, w_156_065, w_156_066, w_156_067, w_156_068, w_156_070, w_156_071, w_156_073, w_156_079, w_156_080, w_156_084, w_156_086, w_156_088, w_156_089, w_156_090, w_156_092, w_156_094, w_156_095, w_156_097, w_156_098, w_156_100, w_156_101, w_156_102, w_156_103, w_156_104, w_156_105, w_156_109, w_156_111, w_156_112, w_156_113, w_156_116, w_156_118, w_156_120, w_156_121, w_156_123, w_156_124, w_156_126, w_156_127, w_156_128, w_156_129, w_156_130, w_156_131, w_156_134, w_156_135, w_156_136, w_156_138, w_156_142, w_156_144, w_156_145, w_156_146, w_156_148, w_156_149, w_156_151, w_156_152, w_156_155, w_156_156, w_156_157, w_156_158, w_156_164, w_156_165, w_156_166, w_156_167, w_156_170, w_156_171, w_156_172, w_156_174, w_156_177, w_156_178, w_156_181, w_156_183, w_156_184, w_156_186, w_156_187, w_156_190, w_156_191, w_156_193, w_156_196, w_156_197, w_156_198, w_156_201, w_156_203, w_156_204, w_156_205, w_156_206, w_156_210, w_156_211, w_156_212, w_156_215, w_156_219, w_156_221, w_156_222, w_156_223, w_156_226, w_156_230, w_156_234, w_156_235, w_156_242, w_156_244, w_156_245, w_156_247, w_156_256, w_156_257, w_156_258, w_156_261, w_156_262, w_156_263, w_156_264, w_156_265, w_156_266, w_156_267, w_156_270, w_156_273, w_156_276, w_156_277, w_156_279, w_156_280, w_156_281, w_156_282, w_156_283, w_156_284, w_156_285, w_156_287, w_156_289, w_156_291, w_156_294, w_156_296, w_156_297, w_156_299, w_156_300, w_156_301, w_156_307, w_156_308, w_156_309, w_156_313, w_156_318, w_156_320, w_156_321, w_156_322, w_156_325, w_156_327, w_156_328, w_156_329, w_156_333, w_156_334, w_156_336, w_156_338, w_156_340, w_156_341, w_156_343, w_156_344, w_156_345, w_156_346, w_156_348, w_156_349, w_156_350, w_156_351, w_156_352, w_156_354, w_156_355, w_156_356, w_156_359, w_156_361, w_156_362, w_156_366, w_156_367, w_156_369, w_156_370, w_156_373, w_156_374, w_156_375, w_156_377, w_156_378, w_156_379, w_156_381, w_156_383, w_156_384, w_156_385, w_156_386, w_156_388, w_156_390, w_156_393, w_156_394, w_156_395, w_156_398, w_156_402, w_156_403, w_156_404, w_156_406, w_156_409, w_156_410, w_156_412, w_156_417, w_156_420, w_156_421, w_156_422, w_156_423, w_156_426, w_156_427, w_156_428, w_156_429, w_156_430, w_156_434, w_156_439, w_156_440, w_156_441, w_156_443, w_156_444, w_156_448, w_156_450, w_156_451, w_156_454, w_156_455, w_156_457, w_156_458, w_156_459, w_156_460, w_156_461, w_156_465, w_156_467, w_156_468, w_156_469, w_156_471, w_156_475, w_156_476, w_156_477, w_156_478, w_156_480, w_156_481, w_156_483, w_156_484, w_156_486, w_156_487, w_156_488, w_156_491, w_156_492, w_156_493, w_156_499, w_156_503, w_156_504, w_156_506, w_156_509, w_156_511, w_156_512, w_156_513, w_156_518, w_156_521, w_156_523, w_156_524, w_156_527, w_156_528, w_156_529, w_156_533, w_156_534, w_156_535, w_156_536, w_156_538, w_156_540, w_156_541, w_156_544, w_156_552, w_156_553, w_156_555, w_156_559, w_156_561, w_156_563, w_156_564, w_156_565, w_156_566, w_156_567, w_156_570, w_156_571, w_156_572, w_156_573, w_156_574, w_156_575, w_156_576, w_156_577, w_156_578, w_156_579, w_156_585, w_156_588, w_156_589, w_156_590, w_156_591, w_156_592, w_156_597, w_156_599, w_156_601, w_156_605, w_156_611, w_156_613, w_156_615, w_156_617, w_156_621, w_156_622, w_156_623, w_156_624, w_156_625, w_156_628, w_156_629, w_156_631, w_156_632, w_156_633, w_156_634, w_156_638, w_156_640, w_156_641, w_156_642, w_156_646, w_156_647, w_156_651, w_156_652, w_156_653, w_156_654, w_156_657, w_156_659, w_156_660, w_156_661, w_156_662, w_156_663, w_156_664, w_156_665, w_156_666, w_156_667, w_156_669, w_156_671, w_156_672, w_156_673, w_156_674, w_156_677, w_156_678, w_156_679, w_156_681, w_156_682, w_156_684, w_156_685, w_156_686, w_156_687, w_156_690, w_156_692, w_156_693, w_156_694, w_156_695, w_156_696, w_156_697, w_156_698, w_156_699, w_156_700, w_156_703, w_156_705, w_156_707, w_156_709, w_156_710, w_156_711, w_156_712, w_156_714, w_156_715, w_156_717, w_156_718, w_156_719, w_156_720, w_156_721, w_156_726, w_156_728, w_156_732, w_156_734, w_156_735, w_156_736, w_156_737, w_156_740, w_156_745, w_156_747, w_156_748, w_156_749, w_156_750, w_156_752, w_156_753, w_156_755, w_156_756, w_156_757, w_156_758, w_156_759, w_156_761, w_156_765, w_156_767, w_156_768, w_156_769, w_156_770, w_156_775, w_156_777, w_156_778, w_156_781, w_156_784, w_156_785, w_156_786, w_156_787, w_156_788, w_156_789, w_156_792, w_156_793, w_156_794, w_156_797, w_156_799, w_156_800, w_156_801, w_156_802, w_156_803, w_156_804, w_156_806, w_156_807, w_156_809, w_156_815, w_156_816, w_156_817, w_156_818, w_156_820, w_156_821, w_156_822, w_156_823, w_156_826, w_156_827, w_156_830, w_156_834, w_156_837, w_156_840, w_156_842, w_156_843, w_156_845, w_156_848, w_156_850, w_156_853, w_156_855, w_156_862, w_156_863, w_156_869, w_156_870, w_156_872, w_156_874, w_156_877, w_156_878, w_156_883, w_156_886, w_156_887, w_156_888, w_156_889, w_156_890, w_156_891, w_156_893, w_156_894, w_156_896, w_156_897, w_156_899, w_156_900, w_156_901, w_156_902, w_156_903, w_156_905, w_156_907, w_156_908, w_156_913, w_156_916, w_156_918, w_156_921, w_156_931, w_156_933, w_156_940, w_156_941, w_156_943, w_156_944, w_156_945, w_156_948, w_156_951, w_156_953, w_156_954, w_156_961, w_156_968, w_156_970, w_156_971, w_156_972, w_156_973, w_156_976, w_156_977, w_156_978, w_156_979, w_156_980, w_156_981, w_156_982, w_156_983, w_156_987, w_156_989, w_156_992, w_156_993, w_156_995, w_156_996, w_156_999, w_156_1000, w_156_1004, w_156_1007, w_156_1008, w_156_1011, w_156_1014, w_156_1015, w_156_1016, w_156_1019, w_156_1022, w_156_1026, w_156_1028, w_156_1029, w_156_1031, w_156_1033, w_156_1034, w_156_1039, w_156_1040, w_156_1043, w_156_1044, w_156_1045, w_156_1047, w_156_1049, w_156_1050, w_156_1052, w_156_1053, w_156_1055, w_156_1057, w_156_1059, w_156_1060, w_156_1061, w_156_1062, w_156_1064, w_156_1071, w_156_1074, w_156_1075, w_156_1076, w_156_1078, w_156_1079, w_156_1080, w_156_1083, w_156_1084, w_156_1087, w_156_1088, w_156_1089, w_156_1091, w_156_1092, w_156_1093, w_156_1094, w_156_1096, w_156_1098, w_156_1100, w_156_1101, w_156_1103, w_156_1104, w_156_1105, w_156_1107, w_156_1115, w_156_1116, w_156_1118, w_156_1120, w_156_1122, w_156_1125, w_156_1127, w_156_1129, w_156_1132, w_156_1133, w_156_1134, w_156_1137, w_156_1139, w_156_1140, w_156_1143, w_156_1148, w_156_1149, w_156_1156, w_156_1157, w_156_1165, w_156_1166, w_156_1167, w_156_1168, w_156_1172, w_156_1173, w_156_1174, w_156_1175, w_156_1181, w_156_1182, w_156_1184, w_156_1188, w_156_1190, w_156_1192, w_156_1193, w_156_1200, w_156_1206, w_156_1207, w_156_1210, w_156_1215, w_156_1218, w_156_1220, w_156_1222, w_156_1224, w_156_1229, w_156_1231, w_156_1236, w_156_1237, w_156_1238, w_156_1239, w_156_1241, w_156_1242, w_156_1244, w_156_1248, w_156_1250, w_156_1252, w_156_1254, w_156_1255, w_156_1256, w_156_1257, w_156_1258, w_156_1259, w_156_1261, w_156_1265, w_156_1268, w_156_1270, w_156_1271, w_156_1273, w_156_1274, w_156_1278, w_156_1282, w_156_1285, w_156_1289, w_156_1290, w_156_1295, w_156_1296, w_156_1297, w_156_1299, w_156_1307, w_156_1308, w_156_1313, w_156_1315, w_156_1316, w_156_1317, w_156_1319, w_156_1325, w_156_1327, w_156_1328, w_156_1329, w_156_1330, w_156_1332, w_156_1333, w_156_1335, w_156_1342, w_156_1343, w_156_1344, w_156_1345, w_156_1346, w_156_1351, w_156_1352, w_156_1353, w_156_1354, w_156_1356, w_156_1358, w_156_1361;
  wire w_157_000, w_157_003, w_157_004, w_157_005, w_157_008, w_157_009, w_157_012, w_157_014, w_157_015, w_157_016, w_157_017, w_157_022, w_157_023, w_157_024, w_157_025, w_157_026, w_157_028, w_157_034, w_157_038, w_157_039, w_157_040, w_157_043, w_157_046, w_157_048, w_157_049, w_157_050, w_157_051, w_157_053, w_157_054, w_157_055, w_157_056, w_157_059, w_157_060, w_157_061, w_157_062, w_157_064, w_157_067, w_157_068, w_157_071, w_157_074, w_157_077, w_157_081, w_157_082, w_157_087, w_157_089, w_157_091, w_157_093, w_157_097, w_157_100, w_157_101, w_157_105, w_157_106, w_157_107, w_157_109, w_157_110, w_157_114, w_157_115, w_157_116, w_157_117, w_157_122, w_157_123, w_157_124, w_157_125, w_157_126, w_157_128, w_157_129, w_157_131, w_157_132, w_157_133, w_157_134, w_157_136, w_157_138, w_157_140, w_157_141, w_157_142, w_157_147, w_157_149, w_157_150, w_157_152, w_157_153, w_157_154, w_157_155, w_157_159, w_157_161, w_157_162, w_157_163, w_157_164, w_157_165, w_157_166, w_157_167, w_157_169, w_157_171, w_157_172, w_157_174, w_157_176, w_157_177, w_157_178, w_157_180, w_157_181, w_157_182, w_157_184, w_157_186, w_157_187, w_157_189, w_157_190, w_157_193, w_157_194, w_157_198, w_157_199, w_157_200, w_157_201, w_157_204, w_157_205, w_157_206, w_157_209, w_157_213, w_157_214, w_157_215, w_157_216, w_157_218, w_157_221, w_157_223, w_157_225, w_157_228, w_157_230, w_157_232, w_157_234, w_157_236, w_157_237, w_157_239, w_157_240, w_157_243, w_157_244, w_157_245, w_157_246, w_157_248, w_157_250, w_157_251, w_157_254, w_157_256, w_157_259, w_157_260, w_157_261, w_157_264, w_157_265, w_157_267, w_157_268, w_157_272, w_157_274, w_157_277, w_157_280, w_157_281, w_157_285, w_157_286, w_157_287, w_157_288, w_157_289, w_157_290, w_157_293, w_157_294, w_157_295, w_157_302, w_157_305, w_157_307, w_157_308, w_157_313, w_157_314, w_157_317, w_157_318, w_157_320, w_157_321, w_157_322, w_157_328, w_157_330, w_157_331, w_157_332, w_157_333, w_157_339, w_157_341, w_157_342, w_157_343, w_157_344, w_157_346, w_157_347, w_157_348, w_157_350, w_157_351, w_157_355, w_157_356, w_157_357, w_157_359, w_157_360, w_157_361, w_157_363, w_157_365, w_157_367, w_157_368, w_157_369, w_157_374, w_157_375, w_157_376, w_157_378, w_157_380, w_157_381, w_157_383, w_157_384, w_157_385, w_157_387, w_157_388, w_157_389, w_157_390, w_157_392, w_157_394, w_157_396, w_157_399, w_157_401, w_157_402, w_157_403, w_157_405, w_157_407, w_157_409, w_157_411, w_157_412, w_157_413, w_157_414, w_157_417, w_157_420, w_157_421, w_157_423, w_157_424, w_157_425, w_157_426, w_157_428, w_157_430, w_157_431, w_157_432, w_157_433, w_157_434, w_157_435, w_157_436, w_157_437, w_157_440, w_157_442, w_157_444, w_157_445, w_157_446, w_157_447, w_157_452, w_157_457, w_157_459, w_157_460, w_157_461, w_157_463, w_157_468, w_157_469, w_157_470, w_157_471, w_157_474, w_157_475, w_157_476, w_157_477, w_157_478, w_157_479, w_157_481, w_157_483, w_157_488, w_157_489, w_157_491, w_157_492, w_157_494, w_157_497, w_157_498, w_157_500, w_157_501, w_157_502, w_157_504, w_157_505, w_157_507, w_157_510, w_157_511, w_157_512, w_157_517, w_157_524, w_157_526, w_157_527, w_157_528, w_157_531, w_157_532, w_157_534, w_157_536, w_157_537, w_157_539, w_157_540, w_157_542, w_157_544, w_157_546, w_157_548, w_157_549, w_157_550, w_157_552, w_157_553, w_157_554, w_157_555, w_157_556, w_157_560, w_157_562, w_157_565, w_157_572, w_157_573, w_157_574, w_157_575, w_157_576, w_157_578, w_157_580, w_157_582, w_157_584, w_157_585, w_157_589, w_157_590, w_157_591, w_157_595, w_157_596, w_157_597, w_157_600, w_157_603, w_157_605, w_157_606, w_157_610, w_157_613, w_157_617, w_157_618, w_157_619, w_157_621, w_157_622, w_157_623, w_157_624, w_157_627, w_157_629, w_157_630, w_157_632, w_157_636, w_157_637, w_157_638, w_157_642, w_157_643, w_157_645, w_157_646, w_157_650, w_157_654, w_157_655, w_157_657, w_157_661, w_157_662, w_157_663, w_157_664, w_157_669, w_157_670, w_157_671, w_157_672, w_157_674, w_157_675, w_157_676, w_157_680, w_157_682, w_157_683, w_157_684, w_157_687, w_157_689, w_157_690, w_157_691, w_157_693, w_157_694, w_157_698, w_157_699, w_157_700, w_157_703, w_157_704, w_157_707, w_157_708, w_157_709, w_157_711, w_157_712, w_157_716, w_157_717, w_157_719, w_157_720, w_157_724, w_157_725, w_157_726, w_157_729, w_157_731, w_157_732, w_157_738, w_157_739, w_157_740, w_157_741, w_157_742, w_157_743, w_157_744, w_157_745, w_157_748, w_157_749, w_157_750, w_157_751, w_157_753, w_157_755, w_157_756, w_157_757, w_157_759, w_157_760, w_157_761, w_157_762, w_157_763, w_157_765, w_157_771, w_157_772, w_157_774, w_157_776, w_157_780, w_157_783, w_157_786, w_157_788, w_157_795, w_157_799, w_157_801, w_157_803, w_157_804, w_157_806, w_157_807, w_157_808, w_157_809, w_157_811, w_157_817, w_157_818, w_157_820, w_157_821, w_157_824, w_157_825, w_157_827, w_157_828, w_157_829, w_157_830, w_157_832, w_157_834, w_157_836, w_157_839, w_157_840, w_157_842, w_157_843, w_157_844, w_157_847, w_157_849, w_157_850, w_157_853, w_157_854, w_157_855, w_157_860, w_157_861, w_157_864, w_157_866, w_157_868, w_157_870, w_157_872, w_157_879, w_157_880, w_157_881, w_157_882, w_157_884, w_157_885, w_157_889, w_157_891, w_157_893, w_157_894, w_157_896, w_157_897, w_157_898, w_157_899, w_157_901, w_157_903, w_157_905, w_157_906, w_157_907, w_157_908, w_157_912, w_157_913, w_157_916, w_157_917, w_157_918, w_157_925, w_157_928, w_157_930, w_157_931, w_157_932, w_157_933, w_157_937, w_157_938, w_157_939, w_157_942, w_157_943, w_157_945, w_157_949, w_157_950, w_157_953, w_157_960, w_157_961, w_157_962, w_157_964, w_157_965, w_157_972, w_157_973, w_157_974, w_157_975, w_157_980, w_157_981, w_157_982, w_157_983, w_157_985, w_157_986, w_157_987, w_157_991, w_157_994, w_157_995, w_157_998, w_157_999, w_157_1000, w_157_1003, w_157_1004, w_157_1006, w_157_1012, w_157_1016, w_157_1021, w_157_1027, w_157_1028, w_157_1029, w_157_1031, w_157_1034, w_157_1037, w_157_1039, w_157_1040, w_157_1041, w_157_1042, w_157_1043, w_157_1044, w_157_1045, w_157_1046, w_157_1049, w_157_1053, w_157_1056, w_157_1057, w_157_1061, w_157_1062, w_157_1065, w_157_1068, w_157_1069, w_157_1070, w_157_1071, w_157_1072, w_157_1073, w_157_1074, w_157_1078, w_157_1079, w_157_1083, w_157_1084, w_157_1088, w_157_1090, w_157_1091, w_157_1093, w_157_1094, w_157_1095, w_157_1099, w_157_1100, w_157_1101, w_157_1102, w_157_1105, w_157_1108, w_157_1109, w_157_1112, w_157_1114, w_157_1117, w_157_1119, w_157_1120, w_157_1121, w_157_1125, w_157_1127, w_157_1129, w_157_1131, w_157_1135, w_157_1137, w_157_1139, w_157_1140, w_157_1145, w_157_1147, w_157_1148, w_157_1149, w_157_1150, w_157_1152, w_157_1154, w_157_1156, w_157_1157, w_157_1163, w_157_1167, w_157_1171, w_157_1173, w_157_1175, w_157_1176, w_157_1177, w_157_1178, w_157_1179, w_157_1184, w_157_1186, w_157_1187, w_157_1189, w_157_1192, w_157_1194, w_157_1195, w_157_1198, w_157_1199, w_157_1200, w_157_1207, w_157_1211, w_157_1212, w_157_1214, w_157_1215, w_157_1217, w_157_1218, w_157_1219, w_157_1220, w_157_1221, w_157_1222, w_157_1228, w_157_1229, w_157_1231, w_157_1232, w_157_1235, w_157_1243, w_157_1245, w_157_1249, w_157_1253, w_157_1254, w_157_1258, w_157_1263, w_157_1266, w_157_1269, w_157_1273, w_157_1274, w_157_1275, w_157_1277, w_157_1278, w_157_1279, w_157_1280, w_157_1281, w_157_1284, w_157_1285, w_157_1287, w_157_1290, w_157_1294, w_157_1296, w_157_1297, w_157_1298, w_157_1301, w_157_1302, w_157_1304, w_157_1307, w_157_1311, w_157_1312, w_157_1313, w_157_1314, w_157_1316, w_157_1317, w_157_1318, w_157_1319, w_157_1324, w_157_1326, w_157_1329, w_157_1330, w_157_1331, w_157_1336, w_157_1340, w_157_1341, w_157_1342, w_157_1344, w_157_1345, w_157_1346, w_157_1350, w_157_1353, w_157_1357, w_157_1358, w_157_1359, w_157_1360, w_157_1361, w_157_1366, w_157_1370, w_157_1371;
  wire w_158_001, w_158_004, w_158_005, w_158_007, w_158_008, w_158_009, w_158_010, w_158_011, w_158_013, w_158_014, w_158_016, w_158_018, w_158_022, w_158_023, w_158_025, w_158_030, w_158_034, w_158_035, w_158_036, w_158_037, w_158_038, w_158_039, w_158_040, w_158_041, w_158_043, w_158_045, w_158_047, w_158_048, w_158_053, w_158_054, w_158_055, w_158_056, w_158_057, w_158_059, w_158_060, w_158_061, w_158_063, w_158_064, w_158_065, w_158_066, w_158_067, w_158_068, w_158_069, w_158_070, w_158_071, w_158_072, w_158_074, w_158_076, w_158_081, w_158_083, w_158_087, w_158_088, w_158_090, w_158_091, w_158_095, w_158_097, w_158_098, w_158_099, w_158_100, w_158_106, w_158_107, w_158_109, w_158_110, w_158_112, w_158_114, w_158_116, w_158_118, w_158_122, w_158_124, w_158_128, w_158_129, w_158_130, w_158_131, w_158_134, w_158_138, w_158_140, w_158_142, w_158_143, w_158_144, w_158_145, w_158_146, w_158_147, w_158_148, w_158_151, w_158_153, w_158_154, w_158_157, w_158_162, w_158_164, w_158_168, w_158_171, w_158_173, w_158_174, w_158_176, w_158_177, w_158_178, w_158_182, w_158_186, w_158_187, w_158_188, w_158_191, w_158_194, w_158_195, w_158_197, w_158_198, w_158_200, w_158_203, w_158_205, w_158_208, w_158_211, w_158_214, w_158_215, w_158_218, w_158_219, w_158_221, w_158_222, w_158_223, w_158_226, w_158_227, w_158_229, w_158_230, w_158_231, w_158_232, w_158_233, w_158_243, w_158_244, w_158_246, w_158_248, w_158_250, w_158_253, w_158_255, w_158_258, w_158_260, w_158_261, w_158_262, w_158_271, w_158_272, w_158_273, w_158_277, w_158_280, w_158_283, w_158_284, w_158_285, w_158_286, w_158_287, w_158_289, w_158_291, w_158_293, w_158_297, w_158_298, w_158_299, w_158_302, w_158_304, w_158_306, w_158_307, w_158_308, w_158_312, w_158_317, w_158_318, w_158_319, w_158_320, w_158_323, w_158_327, w_158_329, w_158_330, w_158_331, w_158_335, w_158_336, w_158_338, w_158_339, w_158_341, w_158_342, w_158_347, w_158_350, w_158_352, w_158_353, w_158_355, w_158_357, w_158_359, w_158_360, w_158_362, w_158_364, w_158_365, w_158_367, w_158_369, w_158_372, w_158_375, w_158_378, w_158_379, w_158_383, w_158_384, w_158_385, w_158_386, w_158_387, w_158_390, w_158_391, w_158_395, w_158_396, w_158_398, w_158_399, w_158_400, w_158_402, w_158_405, w_158_408, w_158_409, w_158_411, w_158_412, w_158_413, w_158_417, w_158_420, w_158_421, w_158_426, w_158_427, w_158_428, w_158_433, w_158_434, w_158_436, w_158_437, w_158_439, w_158_440, w_158_441, w_158_442, w_158_443, w_158_444, w_158_448, w_158_450, w_158_451, w_158_456, w_158_457, w_158_458, w_158_459, w_158_460, w_158_461, w_158_462, w_158_464, w_158_468, w_158_471, w_158_472, w_158_478, w_158_482, w_158_484, w_158_486, w_158_492, w_158_495, w_158_496, w_158_497, w_158_499, w_158_503, w_158_504, w_158_507, w_158_508, w_158_511, w_158_512, w_158_513, w_158_516, w_158_517, w_158_520, w_158_527, w_158_529, w_158_533, w_158_535, w_158_536, w_158_537, w_158_543, w_158_548, w_158_549, w_158_551, w_158_552, w_158_554, w_158_555, w_158_557, w_158_560, w_158_562, w_158_563, w_158_568, w_158_569, w_158_573, w_158_574, w_158_577, w_158_578, w_158_579, w_158_580, w_158_582, w_158_583, w_158_591, w_158_593, w_158_594, w_158_595, w_158_596, w_158_598, w_158_602, w_158_603, w_158_604, w_158_610, w_158_614, w_158_617, w_158_619, w_158_620, w_158_622, w_158_623, w_158_627, w_158_628, w_158_631, w_158_634, w_158_637, w_158_639, w_158_642, w_158_644, w_158_645, w_158_646, w_158_648, w_158_651, w_158_656, w_158_657, w_158_658, w_158_661, w_158_662, w_158_663, w_158_665, w_158_676, w_158_677, w_158_678, w_158_679, w_158_682, w_158_684, w_158_686, w_158_689, w_158_690, w_158_692, w_158_700, w_158_701, w_158_702, w_158_705, w_158_706, w_158_709, w_158_710, w_158_715, w_158_722, w_158_729, w_158_731, w_158_734, w_158_735, w_158_737, w_158_738, w_158_742, w_158_746, w_158_748, w_158_750, w_158_751, w_158_756, w_158_757, w_158_759, w_158_760, w_158_761, w_158_762, w_158_766, w_158_768, w_158_769, w_158_775, w_158_776, w_158_777, w_158_779, w_158_780, w_158_782, w_158_785, w_158_787, w_158_790, w_158_792, w_158_794, w_158_796, w_158_800, w_158_803, w_158_804, w_158_805, w_158_806, w_158_808, w_158_809, w_158_810, w_158_812, w_158_813, w_158_814, w_158_815, w_158_816, w_158_818, w_158_819, w_158_821, w_158_822, w_158_823, w_158_824, w_158_828, w_158_829, w_158_833, w_158_835, w_158_838, w_158_840, w_158_841, w_158_844, w_158_845, w_158_849, w_158_852, w_158_859, w_158_860, w_158_867, w_158_870, w_158_871, w_158_872, w_158_875, w_158_876, w_158_877, w_158_878, w_158_879, w_158_884, w_158_886, w_158_888, w_158_890, w_158_896, w_158_897, w_158_899, w_158_900, w_158_903, w_158_908, w_158_910, w_158_911, w_158_912, w_158_915, w_158_917, w_158_930, w_158_931, w_158_934, w_158_935, w_158_937, w_158_939, w_158_942, w_158_943, w_158_945, w_158_946, w_158_947, w_158_950, w_158_951, w_158_955, w_158_958, w_158_965, w_158_968, w_158_970, w_158_971, w_158_974, w_158_977, w_158_981, w_158_982, w_158_985, w_158_986, w_158_990, w_158_996, w_158_997, w_158_998, w_158_999, w_158_1002, w_158_1004, w_158_1007, w_158_1011, w_158_1012, w_158_1015, w_158_1020, w_158_1021, w_158_1025, w_158_1027, w_158_1031, w_158_1033, w_158_1034, w_158_1035, w_158_1036, w_158_1038, w_158_1043, w_158_1044, w_158_1046, w_158_1047, w_158_1050, w_158_1051, w_158_1053, w_158_1054, w_158_1055, w_158_1058, w_158_1059, w_158_1063, w_158_1064, w_158_1066, w_158_1068, w_158_1069, w_158_1070, w_158_1073, w_158_1076, w_158_1077, w_158_1079, w_158_1081, w_158_1085, w_158_1086, w_158_1088, w_158_1089, w_158_1093, w_158_1095, w_158_1096, w_158_1098, w_158_1099, w_158_1103, w_158_1105, w_158_1106, w_158_1119, w_158_1122, w_158_1123, w_158_1127, w_158_1129, w_158_1130, w_158_1133, w_158_1134, w_158_1136, w_158_1137, w_158_1138, w_158_1139, w_158_1141, w_158_1142, w_158_1147, w_158_1150, w_158_1154, w_158_1155, w_158_1157, w_158_1158, w_158_1159, w_158_1160, w_158_1162, w_158_1166, w_158_1167, w_158_1173, w_158_1177, w_158_1179, w_158_1180, w_158_1186, w_158_1187, w_158_1190, w_158_1191, w_158_1192, w_158_1197, w_158_1198, w_158_1199, w_158_1200, w_158_1203, w_158_1204, w_158_1206, w_158_1209, w_158_1211, w_158_1215, w_158_1216, w_158_1217, w_158_1219, w_158_1222, w_158_1224, w_158_1225, w_158_1226, w_158_1227, w_158_1230, w_158_1238, w_158_1241, w_158_1242, w_158_1243, w_158_1244, w_158_1250, w_158_1253, w_158_1258, w_158_1259, w_158_1260, w_158_1261, w_158_1265, w_158_1266, w_158_1267, w_158_1269, w_158_1274, w_158_1277, w_158_1278, w_158_1282, w_158_1286, w_158_1287, w_158_1288, w_158_1291, w_158_1293, w_158_1294, w_158_1296, w_158_1298, w_158_1300, w_158_1304, w_158_1306, w_158_1307, w_158_1310, w_158_1311, w_158_1314, w_158_1315, w_158_1316, w_158_1318, w_158_1319, w_158_1322, w_158_1328, w_158_1330, w_158_1331, w_158_1332, w_158_1333, w_158_1339, w_158_1344, w_158_1345, w_158_1346, w_158_1347, w_158_1348, w_158_1351, w_158_1358, w_158_1360, w_158_1362, w_158_1366, w_158_1367, w_158_1370, w_158_1371, w_158_1372, w_158_1374, w_158_1375, w_158_1376, w_158_1380, w_158_1382, w_158_1383, w_158_1384, w_158_1385, w_158_1388, w_158_1391, w_158_1397, w_158_1398, w_158_1400, w_158_1401, w_158_1402, w_158_1403, w_158_1404, w_158_1407, w_158_1408, w_158_1409, w_158_1410, w_158_1412, w_158_1413, w_158_1415, w_158_1420, w_158_1421, w_158_1422, w_158_1423, w_158_1424, w_158_1425, w_158_1429, w_158_1430, w_158_1432, w_158_1433, w_158_1440, w_158_1445, w_158_1451, w_158_1456, w_158_1457, w_158_1458, w_158_1463, w_158_1464, w_158_1465, w_158_1471, w_158_1474, w_158_1480, w_158_1483, w_158_1485, w_158_1486, w_158_1488, w_158_1493, w_158_1494, w_158_1495, w_158_1500, w_158_1501, w_158_1502, w_158_1505, w_158_1506, w_158_1508, w_158_1509, w_158_1510, w_158_1512, w_158_1518, w_158_1519, w_158_1521, w_158_1522, w_158_1524, w_158_1527, w_158_1528, w_158_1531, w_158_1533, w_158_1538, w_158_1539, w_158_1540, w_158_1541, w_158_1544, w_158_1546, w_158_1547, w_158_1550, w_158_1551, w_158_1552, w_158_1553, w_158_1555, w_158_1556, w_158_1558, w_158_1561, w_158_1563, w_158_1564, w_158_1565, w_158_1573, w_158_1574, w_158_1579, w_158_1581, w_158_1583, w_158_1588, w_158_1590, w_158_1596, w_158_1598, w_158_1599, w_158_1601, w_158_1602, w_158_1610, w_158_1612, w_158_1615, w_158_1616, w_158_1617, w_158_1623, w_158_1624, w_158_1630, w_158_1632, w_158_1636;
  wire w_159_000, w_159_001, w_159_010, w_159_011, w_159_013, w_159_015, w_159_016, w_159_018, w_159_019, w_159_020, w_159_021, w_159_022, w_159_025, w_159_029, w_159_030, w_159_032, w_159_033, w_159_034, w_159_035, w_159_036, w_159_037, w_159_039, w_159_041, w_159_042, w_159_043, w_159_044, w_159_045, w_159_046, w_159_049, w_159_055, w_159_057, w_159_058, w_159_059, w_159_060, w_159_061, w_159_064, w_159_066, w_159_067, w_159_068, w_159_069, w_159_070, w_159_071, w_159_074, w_159_076, w_159_077, w_159_080, w_159_084, w_159_086, w_159_088, w_159_089, w_159_090, w_159_093, w_159_096, w_159_099, w_159_101, w_159_102, w_159_104, w_159_105, w_159_110, w_159_114, w_159_116, w_159_117, w_159_118, w_159_119, w_159_120, w_159_121, w_159_123, w_159_125, w_159_127, w_159_128, w_159_129, w_159_130, w_159_137, w_159_141, w_159_142, w_159_144, w_159_145, w_159_146, w_159_147, w_159_148, w_159_150, w_159_152, w_159_155, w_159_156, w_159_157, w_159_160, w_159_167, w_159_169, w_159_170, w_159_171, w_159_172, w_159_176, w_159_178, w_159_180, w_159_184, w_159_189, w_159_191, w_159_193, w_159_194, w_159_195, w_159_196, w_159_197, w_159_199, w_159_202, w_159_203, w_159_204, w_159_207, w_159_208, w_159_209, w_159_211, w_159_212, w_159_214, w_159_215, w_159_216, w_159_219, w_159_222, w_159_225, w_159_226, w_159_229, w_159_230, w_159_233, w_159_236, w_159_240, w_159_245, w_159_247, w_159_250, w_159_254, w_159_256, w_159_257, w_159_260, w_159_262, w_159_266, w_159_270, w_159_272, w_159_274, w_159_276, w_159_279, w_159_282, w_159_283, w_159_284, w_159_285, w_159_286, w_159_287, w_159_290, w_159_291, w_159_295, w_159_297, w_159_301, w_159_304, w_159_305, w_159_307, w_159_308, w_159_312, w_159_314, w_159_315, w_159_317, w_159_320, w_159_322, w_159_324, w_159_325, w_159_329, w_159_330, w_159_335, w_159_336, w_159_342, w_159_345, w_159_346, w_159_348, w_159_352, w_159_355, w_159_356, w_159_357, w_159_362, w_159_367, w_159_370, w_159_371, w_159_373, w_159_381, w_159_385, w_159_389, w_159_390, w_159_391, w_159_392, w_159_395, w_159_399, w_159_400, w_159_404, w_159_409, w_159_410, w_159_416, w_159_417, w_159_419, w_159_420, w_159_426, w_159_428, w_159_432, w_159_433, w_159_439, w_159_447, w_159_448, w_159_449, w_159_450, w_159_452, w_159_454, w_159_455, w_159_456, w_159_461, w_159_462, w_159_464, w_159_467, w_159_471, w_159_476, w_159_478, w_159_479, w_159_481, w_159_482, w_159_483, w_159_484, w_159_486, w_159_487, w_159_492, w_159_494, w_159_495, w_159_499, w_159_500, w_159_501, w_159_504, w_159_505, w_159_506, w_159_509, w_159_511, w_159_517, w_159_519, w_159_520, w_159_521, w_159_524, w_159_525, w_159_527, w_159_528, w_159_530, w_159_531, w_159_532, w_159_533, w_159_536, w_159_539, w_159_540, w_159_543, w_159_545, w_159_546, w_159_548, w_159_551, w_159_552, w_159_553, w_159_554, w_159_555, w_159_558, w_159_559, w_159_561, w_159_563, w_159_566, w_159_568, w_159_572, w_159_575, w_159_578, w_159_579, w_159_580, w_159_581, w_159_583, w_159_585, w_159_587, w_159_588, w_159_590, w_159_592, w_159_594, w_159_595, w_159_598, w_159_600, w_159_601, w_159_603, w_159_604, w_159_608, w_159_613, w_159_616, w_159_622, w_159_624, w_159_626, w_159_628, w_159_629, w_159_637, w_159_640, w_159_644, w_159_645, w_159_646, w_159_647, w_159_648, w_159_651, w_159_653, w_159_658, w_159_659, w_159_665, w_159_666, w_159_670, w_159_674, w_159_675, w_159_677, w_159_679, w_159_680, w_159_681, w_159_683, w_159_684, w_159_688, w_159_689, w_159_693, w_159_694, w_159_696, w_159_700, w_159_701, w_159_702, w_159_705, w_159_708, w_159_710, w_159_711, w_159_712, w_159_713, w_159_714, w_159_715, w_159_717, w_159_719, w_159_722, w_159_725, w_159_726, w_159_730, w_159_731, w_159_734, w_159_736, w_159_739, w_159_743, w_159_748, w_159_749, w_159_750, w_159_751, w_159_758, w_159_759, w_159_760, w_159_763, w_159_764, w_159_769, w_159_770, w_159_771, w_159_772, w_159_774, w_159_777, w_159_778, w_159_779, w_159_781, w_159_783, w_159_784, w_159_787, w_159_788, w_159_789, w_159_790, w_159_797, w_159_801, w_159_803, w_159_804, w_159_809, w_159_811, w_159_812, w_159_814, w_159_816, w_159_817, w_159_820, w_159_822, w_159_825, w_159_826, w_159_830, w_159_832, w_159_835, w_159_842, w_159_843, w_159_844, w_159_845, w_159_849, w_159_854, w_159_855, w_159_856, w_159_859, w_159_860, w_159_862, w_159_864, w_159_865, w_159_867, w_159_872, w_159_874, w_159_876, w_159_878, w_159_879, w_159_881, w_159_883, w_159_887, w_159_888, w_159_890, w_159_891, w_159_895, w_159_897, w_159_898, w_159_899, w_159_908, w_159_911, w_159_913, w_159_914, w_159_918, w_159_920, w_159_921, w_159_922, w_159_923, w_159_925, w_159_931, w_159_934, w_159_935, w_159_936, w_159_939, w_159_941, w_159_942, w_159_950, w_159_951, w_159_952, w_159_953, w_159_954, w_159_955, w_159_957, w_159_958, w_159_959, w_159_961, w_159_963, w_159_968, w_159_970, w_159_972, w_159_975, w_159_980, w_159_981, w_159_983, w_159_985, w_159_986, w_159_987, w_159_988, w_159_991, w_159_996, w_159_997, w_159_1002, w_159_1006, w_159_1015, w_159_1017, w_159_1018, w_159_1019, w_159_1020, w_159_1021, w_159_1022, w_159_1023, w_159_1027, w_159_1028, w_159_1029, w_159_1031, w_159_1032, w_159_1034, w_159_1038, w_159_1040, w_159_1044, w_159_1045, w_159_1047, w_159_1050, w_159_1051, w_159_1052, w_159_1054, w_159_1057, w_159_1058, w_159_1062, w_159_1068, w_159_1069, w_159_1070, w_159_1073, w_159_1082, w_159_1085, w_159_1087, w_159_1090, w_159_1093, w_159_1097, w_159_1100, w_159_1105, w_159_1106, w_159_1107, w_159_1108, w_159_1112, w_159_1116, w_159_1118, w_159_1119, w_159_1120, w_159_1121, w_159_1123, w_159_1127, w_159_1128, w_159_1130, w_159_1131, w_159_1135, w_159_1137, w_159_1138, w_159_1145, w_159_1147, w_159_1148, w_159_1149, w_159_1150, w_159_1156, w_159_1157, w_159_1160, w_159_1163, w_159_1166, w_159_1167, w_159_1168, w_159_1171, w_159_1176, w_159_1178, w_159_1181, w_159_1183, w_159_1184, w_159_1186, w_159_1190, w_159_1194, w_159_1196, w_159_1197, w_159_1199, w_159_1200, w_159_1204, w_159_1205, w_159_1207, w_159_1209, w_159_1211, w_159_1212, w_159_1213, w_159_1214, w_159_1215, w_159_1217, w_159_1219, w_159_1221, w_159_1222, w_159_1223, w_159_1224, w_159_1226, w_159_1227, w_159_1228, w_159_1229, w_159_1230, w_159_1231, w_159_1232, w_159_1233, w_159_1237, w_159_1240, w_159_1241, w_159_1248, w_159_1250, w_159_1259, w_159_1260, w_159_1262, w_159_1265, w_159_1266, w_159_1267, w_159_1269, w_159_1270, w_159_1271, w_159_1273, w_159_1274, w_159_1275, w_159_1277, w_159_1280, w_159_1282, w_159_1284, w_159_1285, w_159_1287, w_159_1290, w_159_1292, w_159_1295, w_159_1297, w_159_1301, w_159_1302, w_159_1309, w_159_1310, w_159_1314, w_159_1317, w_159_1319, w_159_1321, w_159_1322, w_159_1325, w_159_1328, w_159_1330, w_159_1331, w_159_1334, w_159_1338, w_159_1340, w_159_1344, w_159_1347, w_159_1352, w_159_1359, w_159_1360, w_159_1363, w_159_1365, w_159_1366, w_159_1368, w_159_1369, w_159_1375, w_159_1378, w_159_1379, w_159_1381, w_159_1382, w_159_1383, w_159_1385, w_159_1387, w_159_1391, w_159_1396, w_159_1399, w_159_1400, w_159_1409, w_159_1410, w_159_1412, w_159_1416, w_159_1417, w_159_1418, w_159_1419, w_159_1422, w_159_1423, w_159_1425, w_159_1426, w_159_1428, w_159_1429, w_159_1430, w_159_1433, w_159_1434, w_159_1436, w_159_1437, w_159_1438, w_159_1441, w_159_1443, w_159_1447, w_159_1450, w_159_1452, w_159_1453, w_159_1454, w_159_1455, w_159_1458, w_159_1460, w_159_1462, w_159_1464, w_159_1467, w_159_1469, w_159_1471, w_159_1473, w_159_1474, w_159_1477, w_159_1482, w_159_1483, w_159_1484, w_159_1486, w_159_1491, w_159_1493, w_159_1496, w_159_1497, w_159_1501, w_159_1503, w_159_1506, w_159_1513, w_159_1514, w_159_1515, w_159_1516, w_159_1517, w_159_1524, w_159_1528, w_159_1529, w_159_1534, w_159_1535, w_159_1537, w_159_1538, w_159_1539, w_159_1542, w_159_1545, w_159_1549, w_159_1550, w_159_1552, w_159_1553, w_159_1554, w_159_1555, w_159_1556, w_159_1562, w_159_1563, w_159_1564, w_159_1565, w_159_1566, w_159_1569, w_159_1570, w_159_1573, w_159_1576, w_159_1577, w_159_1586, w_159_1590, w_159_1591, w_159_1592, w_159_1593, w_159_1594, w_159_1595, w_159_1598, w_159_1600, w_159_1601, w_159_1604, w_159_1605, w_159_1609, w_159_1610, w_159_1612, w_159_1616, w_159_1618, w_159_1620;
  wire w_160_002, w_160_004, w_160_006, w_160_007, w_160_009, w_160_010, w_160_011, w_160_012, w_160_013, w_160_015, w_160_016, w_160_017, w_160_019, w_160_021, w_160_025, w_160_026, w_160_030, w_160_031, w_160_032, w_160_038, w_160_039, w_160_040, w_160_042, w_160_044, w_160_045, w_160_046, w_160_047, w_160_048, w_160_049, w_160_051, w_160_055, w_160_056, w_160_062, w_160_065, w_160_066, w_160_067, w_160_069, w_160_070, w_160_071, w_160_073, w_160_076, w_160_077, w_160_078, w_160_082, w_160_084, w_160_086, w_160_087, w_160_088, w_160_089, w_160_091, w_160_092, w_160_094, w_160_095, w_160_097, w_160_098, w_160_099, w_160_100, w_160_101, w_160_103, w_160_104, w_160_106, w_160_107, w_160_109, w_160_111, w_160_113, w_160_114, w_160_115, w_160_116, w_160_119, w_160_122, w_160_124, w_160_126, w_160_128, w_160_131, w_160_132, w_160_133, w_160_136, w_160_138, w_160_139, w_160_140, w_160_142, w_160_144, w_160_145, w_160_148, w_160_149, w_160_153, w_160_159, w_160_160, w_160_161, w_160_162, w_160_163, w_160_164, w_160_165, w_160_166, w_160_168, w_160_169, w_160_170, w_160_171, w_160_173, w_160_175, w_160_176, w_160_177, w_160_178, w_160_179, w_160_180, w_160_181, w_160_182, w_160_184, w_160_185, w_160_186, w_160_187, w_160_188, w_160_189, w_160_192, w_160_195, w_160_197, w_160_199, w_160_201, w_160_202, w_160_203, w_160_205, w_160_206, w_160_207, w_160_208, w_160_209, w_160_211, w_160_212, w_160_217, w_160_219, w_160_220, w_160_222, w_160_223, w_160_224, w_160_225, w_160_226, w_160_227, w_160_228, w_160_229, w_160_230, w_160_231, w_160_235, w_160_237, w_160_238, w_160_239, w_160_241, w_160_243, w_160_244, w_160_248, w_160_250, w_160_252, w_160_254, w_160_256, w_160_258, w_160_264, w_160_266, w_160_268, w_160_270, w_160_271, w_160_272, w_160_273, w_160_274, w_160_277, w_160_279, w_160_280, w_160_282, w_160_283, w_160_284, w_160_289, w_160_290, w_160_292, w_160_294, w_160_295, w_160_299, w_160_300, w_160_301, w_160_302, w_160_303, w_160_304, w_160_307, w_160_310, w_160_312, w_160_315, w_160_321, w_160_322, w_160_325, w_160_332, w_160_333, w_160_334, w_160_337, w_160_338, w_160_339, w_160_340, w_160_341, w_160_342, w_160_344, w_160_346, w_160_348, w_160_351, w_160_355, w_160_358, w_160_359, w_160_360, w_160_361, w_160_362, w_160_363, w_160_364, w_160_365, w_160_366, w_160_367, w_160_368, w_160_369, w_160_370, w_160_372, w_160_373, w_160_374, w_160_377, w_160_381, w_160_382, w_160_383, w_160_384, w_160_388, w_160_389, w_160_390, w_160_395, w_160_396, w_160_397, w_160_399, w_160_400, w_160_401, w_160_403, w_160_404, w_160_405, w_160_408, w_160_409, w_160_410, w_160_415, w_160_416, w_160_417, w_160_420, w_160_422, w_160_423, w_160_424, w_160_425, w_160_426, w_160_427, w_160_430, w_160_431, w_160_432, w_160_433, w_160_434, w_160_437, w_160_440, w_160_442, w_160_443, w_160_444, w_160_445, w_160_448, w_160_451, w_160_454, w_160_455, w_160_456, w_160_457, w_160_459, w_160_461, w_160_464, w_160_465, w_160_468, w_160_469, w_160_471, w_160_472, w_160_476, w_160_477, w_160_479, w_160_481, w_160_482, w_160_483, w_160_485, w_160_486, w_160_488, w_160_489, w_160_490, w_160_492, w_160_493, w_160_497, w_160_499, w_160_501, w_160_502, w_160_504, w_160_506, w_160_507, w_160_511, w_160_514, w_160_515, w_160_516, w_160_517, w_160_518, w_160_520, w_160_522, w_160_524, w_160_525, w_160_526, w_160_528, w_160_529, w_160_533, w_160_538, w_160_539, w_160_540, w_160_541, w_160_542, w_160_545, w_160_547, w_160_549, w_160_550, w_160_555, w_160_556, w_160_558, w_160_559, w_160_567, w_160_568, w_160_569, w_160_571, w_160_572, w_160_573, w_160_574, w_160_575, w_160_576, w_160_577, w_160_578, w_160_582, w_160_584, w_160_585, w_160_586, w_160_587, w_160_588, w_160_589, w_160_591, w_160_594, w_160_597, w_160_600, w_160_603, w_160_605, w_160_606, w_160_609, w_160_610, w_160_614, w_160_615, w_160_616, w_160_618, w_160_619, w_160_620, w_160_621, w_160_623, w_160_625, w_160_626, w_160_629, w_160_630, w_160_631, w_160_632, w_160_633, w_160_634, w_160_638, w_160_639, w_160_641, w_160_643, w_160_644, w_160_645, w_160_647, w_160_649, w_160_650, w_160_651, w_160_652, w_160_653, w_160_654, w_160_655, w_160_659, w_160_662, w_160_663, w_160_664, w_160_665, w_160_668, w_160_670, w_160_671, w_160_672, w_160_673, w_160_674, w_160_677, w_160_680, w_160_682, w_160_683, w_160_684, w_160_685, w_160_686, w_160_687, w_160_688, w_160_694, w_160_695, w_160_697, w_160_699, w_160_701, w_160_703, w_160_705, w_160_706, w_160_707, w_160_710, w_160_712, w_160_713, w_160_715, w_160_723, w_160_727, w_160_730, w_160_731, w_160_733, w_160_734, w_160_735, w_160_738, w_160_739, w_160_742, w_160_743, w_160_744, w_160_745, w_160_746, w_160_747, w_160_750, w_160_756, w_160_757, w_160_758, w_160_759, w_160_761, w_160_762, w_160_763, w_160_764, w_160_765, w_160_767, w_160_769, w_160_774, w_160_777, w_160_778, w_160_780, w_160_781, w_160_782, w_160_784, w_160_787, w_160_788, w_160_790, w_160_794, w_160_796, w_160_797, w_160_798, w_160_799, w_160_800, w_160_802, w_160_804, w_160_805, w_160_808, w_160_813, w_160_814, w_160_815, w_160_816, w_160_818, w_160_819, w_160_823, w_160_824, w_160_826, w_160_828, w_160_829, w_160_831, w_160_832, w_160_833, w_160_836, w_160_839, w_160_840, w_160_841, w_160_852, w_160_854, w_160_860, w_160_861, w_160_863, w_160_866, w_160_867, w_160_868, w_160_869, w_160_874, w_160_875, w_160_876, w_160_877, w_160_879, w_160_881, w_160_882, w_160_883, w_160_884, w_160_886, w_160_889, w_160_891, w_160_892, w_160_893, w_160_894, w_160_895, w_160_896, w_160_900, w_160_902, w_160_903, w_160_904, w_160_908, w_160_909, w_160_910, w_160_913, w_160_915, w_160_918, w_160_919, w_160_920, w_160_923, w_160_924, w_160_926, w_160_927, w_160_928, w_160_930, w_160_932, w_160_933, w_160_935, w_160_936, w_160_938, w_160_940, w_160_942, w_160_943, w_160_944, w_160_946, w_160_948, w_160_949, w_160_951, w_160_959, w_160_960, w_160_962, w_160_965, w_160_967, w_160_971, w_160_972, w_160_973, w_160_977, w_160_980, w_160_983, w_160_984, w_160_985, w_160_989, w_160_992, w_160_994, w_160_995, w_160_998, w_160_999, w_160_1001, w_160_1010, w_160_1013, w_160_1021, w_160_1024, w_160_1026, w_160_1029, w_160_1039, w_160_1040, w_160_1041, w_160_1042, w_160_1045, w_160_1047, w_160_1049, w_160_1051, w_160_1055, w_160_1059, w_160_1060, w_160_1062, w_160_1064, w_160_1066, w_160_1069, w_160_1076, w_160_1079, w_160_1081, w_160_1082, w_160_1087, w_160_1088, w_160_1089, w_160_1094, w_160_1095, w_160_1100, w_160_1101, w_160_1102, w_160_1105, w_160_1106, w_160_1110, w_160_1113, w_160_1114, w_160_1115, w_160_1118, w_160_1119, w_160_1121, w_160_1123, w_160_1128, w_160_1129, w_160_1130, w_160_1135, w_160_1136, w_160_1142, w_160_1147, w_160_1148, w_160_1149, w_160_1150, w_160_1154, w_160_1159, w_160_1164, w_160_1168, w_160_1172, w_160_1174, w_160_1179, w_160_1180, w_160_1184, w_160_1185, w_160_1187, w_160_1190, w_160_1192, w_160_1193, w_160_1194, w_160_1196, w_160_1197, w_160_1198, w_160_1200, w_160_1204, w_160_1208, w_160_1212, w_160_1219, w_160_1220, w_160_1221, w_160_1228, w_160_1229, w_160_1230, w_160_1231, w_160_1232, w_160_1235, w_160_1236, w_160_1238, w_160_1240, w_160_1241, w_160_1242, w_160_1246, w_160_1247, w_160_1249, w_160_1250, w_160_1251, w_160_1258, w_160_1261, w_160_1262, w_160_1263, w_160_1264, w_160_1271, w_160_1272, w_160_1274, w_160_1276, w_160_1279, w_160_1285, w_160_1286, w_160_1290, w_160_1291, w_160_1292, w_160_1294, w_160_1298, w_160_1302, w_160_1309, w_160_1311, w_160_1314, w_160_1315, w_160_1317, w_160_1318, w_160_1321, w_160_1323, w_160_1324, w_160_1325, w_160_1327, w_160_1329, w_160_1332, w_160_1337, w_160_1340, w_160_1342, w_160_1343, w_160_1345, w_160_1346, w_160_1347, w_160_1349, w_160_1351, w_160_1352;
  wire w_161_000, w_161_001, w_161_003, w_161_005, w_161_006, w_161_008, w_161_009, w_161_010, w_161_011, w_161_012, w_161_013, w_161_014, w_161_016, w_161_018, w_161_019, w_161_020, w_161_021, w_161_022, w_161_024, w_161_026, w_161_027, w_161_029, w_161_030, w_161_031, w_161_032, w_161_033, w_161_034, w_161_035, w_161_036, w_161_037, w_161_038, w_161_039, w_161_040, w_161_041, w_161_042, w_161_043, w_161_044, w_161_045, w_161_046, w_161_047, w_161_048, w_161_049, w_161_051, w_161_052, w_161_054, w_161_057, w_161_059, w_161_060, w_161_061, w_161_062, w_161_063, w_161_064, w_161_065, w_161_066, w_161_067, w_161_068, w_161_069, w_161_071, w_161_072, w_161_073, w_161_074, w_161_075, w_161_076, w_161_078, w_161_079, w_161_081, w_161_083, w_161_084, w_161_085, w_161_086, w_161_090, w_161_091, w_161_092, w_161_095, w_161_096, w_161_097, w_161_098, w_161_099, w_161_100, w_161_101, w_161_102, w_161_103, w_161_104, w_161_105, w_161_106, w_161_107, w_161_108, w_161_109, w_161_110, w_161_111, w_161_112, w_161_113, w_161_114, w_161_116, w_161_117, w_161_118, w_161_119, w_161_120, w_161_121, w_161_122, w_161_123, w_161_124, w_161_125, w_161_126, w_161_127, w_161_128, w_161_129, w_161_130, w_161_133, w_161_134, w_161_135, w_161_136, w_161_137, w_161_138, w_161_140, w_161_141, w_161_142, w_161_143, w_161_144, w_161_145, w_161_146, w_161_148, w_161_150, w_161_151, w_161_152, w_161_153, w_161_155, w_161_156, w_161_157, w_161_159, w_161_160, w_161_161, w_161_162, w_161_165, w_161_166, w_161_168, w_161_171, w_161_172, w_161_173, w_161_174, w_161_175, w_161_176, w_161_177, w_161_178, w_161_179, w_161_180, w_161_181, w_161_182, w_161_184, w_161_185, w_161_186, w_161_187, w_161_188, w_161_189, w_161_190, w_161_191, w_161_193, w_161_194, w_161_195, w_161_196, w_161_197, w_161_198, w_161_199, w_161_201, w_161_202, w_161_205, w_161_207, w_161_208, w_161_209, w_161_210, w_161_211, w_161_212, w_161_213, w_161_214, w_161_215, w_161_216, w_161_217, w_161_218, w_161_219, w_161_220, w_161_222, w_161_223, w_161_224, w_161_226, w_161_227, w_161_228, w_161_229, w_161_231, w_161_232, w_161_233, w_161_234, w_161_235, w_161_236, w_161_237, w_161_238, w_161_239, w_161_240, w_161_241, w_161_242, w_161_243, w_161_244, w_161_245, w_161_247, w_161_248, w_161_249, w_161_251, w_161_252, w_161_253, w_161_255, w_161_256, w_161_257, w_161_258, w_161_259, w_161_261, w_161_262, w_161_263, w_161_264, w_161_265, w_161_269, w_161_270, w_161_273, w_161_274, w_161_275, w_161_276, w_161_277, w_161_278, w_161_279, w_161_281, w_161_283, w_161_284, w_161_285, w_161_286, w_161_287, w_161_288, w_161_289, w_161_290, w_161_291, w_161_293, w_161_294, w_161_295, w_161_296, w_161_297, w_161_299, w_161_300, w_161_301, w_161_302, w_161_304, w_161_306, w_161_307, w_161_308, w_161_309, w_161_310, w_161_311, w_161_313, w_161_314, w_161_315, w_161_316, w_161_317, w_161_318, w_161_319, w_161_320, w_161_321, w_161_323, w_161_324, w_161_325, w_161_326, w_161_328, w_161_329, w_161_330, w_161_336, w_161_337, w_161_338, w_161_339, w_161_342, w_161_343, w_161_344, w_161_345, w_161_346, w_161_347, w_161_348, w_161_349, w_161_351, w_161_352, w_161_353, w_161_354, w_161_356, w_161_357, w_161_359, w_161_362, w_161_364, w_161_365, w_161_366, w_161_367, w_161_369, w_161_370, w_161_371, w_161_372, w_161_373, w_161_375, w_161_377, w_161_380, w_161_384, w_161_385, w_161_387, w_161_388, w_161_389, w_161_390, w_161_391, w_161_392, w_161_394, w_161_396, w_161_397, w_161_398, w_161_399, w_161_401, w_161_402, w_161_404, w_161_406, w_161_407, w_161_408, w_161_409, w_161_411, w_161_412, w_161_413, w_161_414, w_161_418, w_161_419, w_161_420, w_161_421, w_161_422, w_161_423, w_161_424, w_161_425, w_161_426, w_161_427, w_161_428, w_161_430, w_161_431, w_161_432, w_161_434, w_161_435, w_161_437, w_161_439, w_161_440, w_161_441, w_161_442, w_161_443, w_161_444, w_161_446, w_161_447, w_161_448, w_161_449, w_161_450, w_161_454, w_161_455, w_161_460, w_161_461, w_161_467, w_161_468, w_161_469, w_161_471, w_161_473, w_161_474, w_161_475, w_161_476, w_161_477, w_161_478, w_161_479, w_161_480, w_161_484, w_161_486, w_161_489, w_161_491, w_161_492, w_161_493, w_161_494, w_161_495, w_161_498, w_161_499, w_161_500, w_161_502, w_161_503, w_161_504, w_161_505, w_161_506, w_161_507, w_161_508, w_161_509, w_161_510, w_161_511, w_161_512, w_161_516, w_161_517, w_161_518, w_161_520, w_161_521, w_161_522, w_161_523, w_161_524, w_161_528, w_161_529, w_161_530, w_161_531, w_161_533, w_161_535, w_161_536, w_161_539, w_161_540, w_161_541, w_161_542, w_161_543, w_161_544, w_161_546, w_161_547, w_161_548, w_161_549, w_161_550, w_161_552, w_161_554, w_161_555, w_161_556, w_161_559, w_161_560, w_161_561, w_161_562, w_161_563, w_161_564, w_161_565, w_161_566, w_161_567, w_161_568, w_161_569, w_161_570, w_161_572, w_161_573, w_161_574, w_161_575, w_161_576, w_161_577, w_161_580, w_161_581, w_161_582, w_161_584, w_161_586, w_161_588, w_161_589, w_161_591, w_161_592, w_161_595, w_161_596, w_161_598, w_161_599, w_161_600;
  wire w_162_006, w_162_012, w_162_014, w_162_019, w_162_025, w_162_031, w_162_035, w_162_040, w_162_041, w_162_048, w_162_055, w_162_056, w_162_061, w_162_068, w_162_071, w_162_084, w_162_085, w_162_089, w_162_095, w_162_096, w_162_097, w_162_098, w_162_103, w_162_107, w_162_109, w_162_113, w_162_117, w_162_118, w_162_120, w_162_130, w_162_131, w_162_137, w_162_141, w_162_142, w_162_143, w_162_144, w_162_148, w_162_153, w_162_156, w_162_161, w_162_164, w_162_167, w_162_169, w_162_171, w_162_173, w_162_176, w_162_180, w_162_188, w_162_193, w_162_194, w_162_195, w_162_196, w_162_197, w_162_198, w_162_201, w_162_204, w_162_205, w_162_209, w_162_210, w_162_211, w_162_215, w_162_218, w_162_223, w_162_230, w_162_231, w_162_234, w_162_238, w_162_241, w_162_242, w_162_246, w_162_249, w_162_254, w_162_256, w_162_260, w_162_268, w_162_269, w_162_270, w_162_273, w_162_274, w_162_275, w_162_276, w_162_277, w_162_282, w_162_284, w_162_294, w_162_296, w_162_297, w_162_298, w_162_299, w_162_300, w_162_313, w_162_315, w_162_317, w_162_322, w_162_324, w_162_325, w_162_327, w_162_328, w_162_329, w_162_335, w_162_338, w_162_339, w_162_340, w_162_341, w_162_343, w_162_345, w_162_347, w_162_349, w_162_352, w_162_353, w_162_358, w_162_367, w_162_374, w_162_376, w_162_379, w_162_380, w_162_386, w_162_387, w_162_393, w_162_400, w_162_401, w_162_404, w_162_405, w_162_413, w_162_418, w_162_420, w_162_430, w_162_435, w_162_436, w_162_437, w_162_438, w_162_443, w_162_446, w_162_453, w_162_455, w_162_459, w_162_460, w_162_461, w_162_465, w_162_466, w_162_469, w_162_470, w_162_473, w_162_477, w_162_479, w_162_480, w_162_486, w_162_490, w_162_492, w_162_496, w_162_500, w_162_503, w_162_504, w_162_506, w_162_508, w_162_512, w_162_515, w_162_519, w_162_521, w_162_524, w_162_527, w_162_530, w_162_532, w_162_534, w_162_536, w_162_542, w_162_551, w_162_552, w_162_562, w_162_564, w_162_565, w_162_566, w_162_569, w_162_570, w_162_571, w_162_574, w_162_575, w_162_580, w_162_586, w_162_587, w_162_588, w_162_590, w_162_591, w_162_595, w_162_596, w_162_597, w_162_599, w_162_600, w_162_601, w_162_603, w_162_609, w_162_614, w_162_617, w_162_619, w_162_623, w_162_624, w_162_634, w_162_636, w_162_637, w_162_639, w_162_647, w_162_648, w_162_658, w_162_664, w_162_667, w_162_672, w_162_673, w_162_674, w_162_678, w_162_679, w_162_682, w_162_683, w_162_685, w_162_686, w_162_691, w_162_693, w_162_699, w_162_700, w_162_702, w_162_703, w_162_704, w_162_710, w_162_712, w_162_713, w_162_714, w_162_715, w_162_718, w_162_720, w_162_722, w_162_723, w_162_727, w_162_733, w_162_737, w_162_741, w_162_745, w_162_750, w_162_755, w_162_770, w_162_771, w_162_773, w_162_775, w_162_776, w_162_777, w_162_782, w_162_786, w_162_788, w_162_791, w_162_792, w_162_793, w_162_798, w_162_801, w_162_802, w_162_804, w_162_810, w_162_812, w_162_820, w_162_826, w_162_828, w_162_830, w_162_837, w_162_840, w_162_843, w_162_846, w_162_848, w_162_849, w_162_853, w_162_857, w_162_858, w_162_862, w_162_874, w_162_877, w_162_887, w_162_894, w_162_900, w_162_902, w_162_904, w_162_908, w_162_912, w_162_913, w_162_916, w_162_919, w_162_923, w_162_924, w_162_925, w_162_926, w_162_931, w_162_932, w_162_933, w_162_940, w_162_941, w_162_942, w_162_948, w_162_950, w_162_952, w_162_955, w_162_956, w_162_964, w_162_966, w_162_968, w_162_969, w_162_971, w_162_977, w_162_984, w_162_987, w_162_989, w_162_993, w_162_996, w_162_998, w_162_1008, w_162_1009, w_162_1015, w_162_1016, w_162_1017, w_162_1023, w_162_1026, w_162_1028, w_162_1033, w_162_1047, w_162_1051, w_162_1052, w_162_1056, w_162_1058, w_162_1060, w_162_1062, w_162_1065, w_162_1069, w_162_1072, w_162_1073, w_162_1076, w_162_1081, w_162_1088, w_162_1092, w_162_1094, w_162_1095, w_162_1101, w_162_1110, w_162_1112, w_162_1114, w_162_1118, w_162_1119, w_162_1126, w_162_1128, w_162_1129, w_162_1131, w_162_1137, w_162_1138, w_162_1141, w_162_1149, w_162_1150, w_162_1154, w_162_1156, w_162_1161, w_162_1167, w_162_1168, w_162_1170, w_162_1173, w_162_1174, w_162_1175, w_162_1177, w_162_1178, w_162_1179, w_162_1187, w_162_1188, w_162_1189, w_162_1193, w_162_1196, w_162_1197, w_162_1199, w_162_1200, w_162_1203, w_162_1210, w_162_1212, w_162_1213, w_162_1216, w_162_1220, w_162_1222, w_162_1224, w_162_1227, w_162_1229, w_162_1230, w_162_1231, w_162_1233, w_162_1234, w_162_1237, w_162_1238, w_162_1242, w_162_1244, w_162_1247, w_162_1248, w_162_1250, w_162_1254, w_162_1257, w_162_1262, w_162_1264, w_162_1266, w_162_1269, w_162_1270, w_162_1273, w_162_1276, w_162_1279, w_162_1283, w_162_1287, w_162_1294, w_162_1296, w_162_1298, w_162_1300, w_162_1304, w_162_1307, w_162_1310, w_162_1317, w_162_1321, w_162_1324, w_162_1330, w_162_1331, w_162_1332, w_162_1339, w_162_1340, w_162_1353, w_162_1357, w_162_1359, w_162_1361, w_162_1363, w_162_1365, w_162_1367, w_162_1368, w_162_1369, w_162_1378, w_162_1381, w_162_1383, w_162_1389, w_162_1400, w_162_1402, w_162_1404, w_162_1405, w_162_1406, w_162_1408, w_162_1410, w_162_1415, w_162_1419, w_162_1424, w_162_1425, w_162_1427, w_162_1436, w_162_1437, w_162_1439, w_162_1440, w_162_1444, w_162_1445, w_162_1452, w_162_1453, w_162_1454, w_162_1455, w_162_1456, w_162_1457, w_162_1463, w_162_1464, w_162_1467, w_162_1473, w_162_1474, w_162_1481, w_162_1485, w_162_1494, w_162_1512, w_162_1518, w_162_1526, w_162_1531, w_162_1534, w_162_1541, w_162_1545, w_162_1546, w_162_1548, w_162_1549, w_162_1560, w_162_1563, w_162_1566, w_162_1567, w_162_1569, w_162_1577, w_162_1578, w_162_1582, w_162_1593, w_162_1595, w_162_1596, w_162_1597, w_162_1601, w_162_1603, w_162_1607, w_162_1619, w_162_1620, w_162_1622, w_162_1625, w_162_1626, w_162_1627, w_162_1632, w_162_1633, w_162_1635, w_162_1654, w_162_1661, w_162_1677, w_162_1679, w_162_1681, w_162_1682, w_162_1683, w_162_1686, w_162_1688, w_162_1694, w_162_1705, w_162_1711, w_162_1713, w_162_1718, w_162_1745, w_162_1747, w_162_1750, w_162_1755, w_162_1765, w_162_1767, w_162_1773, w_162_1809, w_162_1810, w_162_1824, w_162_1836, w_162_1845, w_162_1853, w_162_1865, w_162_1870, w_162_1871, w_162_1874, w_162_1875, w_162_1877, w_162_1882, w_162_1886, w_162_1905, w_162_1906, w_162_1912, w_162_1920, w_162_1925, w_162_1927, w_162_1931, w_162_1936, w_162_1946, w_162_1954, w_162_1956, w_162_1958, w_162_1965, w_162_1968, w_162_1983, w_162_1985, w_162_1992, w_162_1993, w_162_2002, w_162_2020, w_162_2037, w_162_2043, w_162_2047, w_162_2057, w_162_2060, w_162_2064, w_162_2065, w_162_2066, w_162_2079, w_162_2081, w_162_2093, w_162_2096, w_162_2107, w_162_2110, w_162_2117, w_162_2126, w_162_2133, w_162_2138, w_162_2142, w_162_2159, w_162_2173, w_162_2175, w_162_2176, w_162_2179, w_162_2183, w_162_2189, w_162_2190, w_162_2194, w_162_2195, w_162_2201, w_162_2215, w_162_2216, w_162_2222, w_162_2227, w_162_2228, w_162_2230, w_162_2232, w_162_2257, w_162_2265, w_162_2266, w_162_2270, w_162_2283, w_162_2284, w_162_2287, w_162_2290, w_162_2292, w_162_2296, w_162_2302, w_162_2304, w_162_2305, w_162_2307, w_162_2308, w_162_2316, w_162_2320, w_162_2331, w_162_2352, w_162_2356, w_162_2360, w_162_2361, w_162_2365, w_162_2368, w_162_2375, w_162_2379, w_162_2384, w_162_2392, w_162_2401, w_162_2405, w_162_2413, w_162_2417, w_162_2418, w_162_2433, w_162_2442, w_162_2444, w_162_2462, w_162_2476, w_162_2486, w_162_2496, w_162_2503, w_162_2505, w_162_2522, w_162_2542, w_162_2543, w_162_2545, w_162_2550, w_162_2552, w_162_2563, w_162_2564, w_162_2589, w_162_2590, w_162_2591, w_162_2598, w_162_2603, w_162_2604, w_162_2616, w_162_2619, w_162_2624, w_162_2630, w_162_2649, w_162_2651, w_162_2652, w_162_2660, w_162_2661, w_162_2666, w_162_2689, w_162_2699, w_162_2711, w_162_2712, w_162_2724, w_162_2727, w_162_2730, w_162_2734, w_162_2736, w_162_2743, w_162_2746, w_162_2752, w_162_2772, w_162_2777, w_162_2779, w_162_2792, w_162_2795, w_162_2797, w_162_2800, w_162_2802, w_162_2805, w_162_2806, w_162_2813, w_162_2819, w_162_2828, w_162_2834, w_162_2836, w_162_2841, w_162_2845, w_162_2852, w_162_2856, w_162_2861, w_162_2870, w_162_2871, w_162_2883, w_162_2890, w_162_2892, w_162_2893, w_162_2895, w_162_2897, w_162_2900, w_162_2903, w_162_2913, w_162_2914, w_162_2921, w_162_2922, w_162_2940, w_162_2951, w_162_2953, w_162_2963, w_162_2964, w_162_2968, w_162_2980, w_162_2981, w_162_2995, w_162_3004, w_162_3005, w_162_3015, w_162_3016, w_162_3020, w_162_3022, w_162_3024, w_162_3031, w_162_3044, w_162_3046, w_162_3050, w_162_3052, w_162_3065, w_162_3068, w_162_3076, w_162_3078, w_162_3080, w_162_3082, w_162_3083, w_162_3088, w_162_3089, w_162_3090, w_162_3109, w_162_3110, w_162_3116, w_162_3122, w_162_3123, w_162_3127, w_162_3134, w_162_3146, w_162_3149, w_162_3154, w_162_3159, w_162_3163, w_162_3170, w_162_3173, w_162_3176, w_162_3181, w_162_3183, w_162_3185, w_162_3190, w_162_3206, w_162_3210, w_162_3212, w_162_3219, w_162_3220, w_162_3228, w_162_3235, w_162_3240, w_162_3253, w_162_3262, w_162_3263, w_162_3276, w_162_3278, w_162_3279, w_162_3284, w_162_3286, w_162_3291, w_162_3299, w_162_3300, w_162_3316, w_162_3320, w_162_3321, w_162_3323, w_162_3332, w_162_3334, w_162_3335, w_162_3338, w_162_3341, w_162_3354, w_162_3355, w_162_3364, w_162_3376, w_162_3381, w_162_3386, w_162_3387, w_162_3389, w_162_3398, w_162_3400, w_162_3403, w_162_3409, w_162_3414, w_162_3419, w_162_3423, w_162_3426, w_162_3428, w_162_3436, w_162_3450, w_162_3453, w_162_3457, w_162_3462, w_162_3466, w_162_3468, w_162_3484, w_162_3490, w_162_3498, w_162_3502, w_162_3507, w_162_3513, w_162_3517, w_162_3520, w_162_3521, w_162_3523;
  wire w_163_002, w_163_005, w_163_008, w_163_011, w_163_015, w_163_018, w_163_025, w_163_028, w_163_029, w_163_032, w_163_044, w_163_051, w_163_053, w_163_054, w_163_056, w_163_065, w_163_066, w_163_067, w_163_073, w_163_074, w_163_075, w_163_080, w_163_083, w_163_087, w_163_088, w_163_090, w_163_091, w_163_097, w_163_098, w_163_099, w_163_105, w_163_109, w_163_110, w_163_111, w_163_112, w_163_114, w_163_118, w_163_120, w_163_124, w_163_128, w_163_129, w_163_130, w_163_136, w_163_138, w_163_140, w_163_141, w_163_147, w_163_148, w_163_151, w_163_154, w_163_156, w_163_157, w_163_158, w_163_159, w_163_160, w_163_163, w_163_165, w_163_166, w_163_167, w_163_170, w_163_177, w_163_178, w_163_185, w_163_186, w_163_187, w_163_194, w_163_202, w_163_203, w_163_209, w_163_210, w_163_212, w_163_213, w_163_214, w_163_215, w_163_216, w_163_218, w_163_219, w_163_220, w_163_221, w_163_222, w_163_223, w_163_225, w_163_226, w_163_227, w_163_230, w_163_236, w_163_245, w_163_247, w_163_248, w_163_249, w_163_252, w_163_256, w_163_258, w_163_261, w_163_263, w_163_264, w_163_265, w_163_266, w_163_270, w_163_275, w_163_280, w_163_283, w_163_284, w_163_286, w_163_287, w_163_289, w_163_291, w_163_292, w_163_295, w_163_296, w_163_297, w_163_302, w_163_303, w_163_305, w_163_306, w_163_307, w_163_308, w_163_309, w_163_313, w_163_316, w_163_317, w_163_319, w_163_320, w_163_321, w_163_322, w_163_325, w_163_330, w_163_331, w_163_338, w_163_339, w_163_340, w_163_344, w_163_346, w_163_348, w_163_356, w_163_360, w_163_361, w_163_362, w_163_366, w_163_371, w_163_383, w_163_385, w_163_390, w_163_393, w_163_394, w_163_399, w_163_400, w_163_405, w_163_408, w_163_409, w_163_411, w_163_413, w_163_420, w_163_425, w_163_436, w_163_437, w_163_439, w_163_446, w_163_447, w_163_449, w_163_451, w_163_456, w_163_457, w_163_459, w_163_464, w_163_467, w_163_469, w_163_476, w_163_477, w_163_479, w_163_480, w_163_483, w_163_484, w_163_488, w_163_489, w_163_490, w_163_491, w_163_492, w_163_497, w_163_499, w_163_506, w_163_508, w_163_511, w_163_513, w_163_515, w_163_527, w_163_532, w_163_537, w_163_538, w_163_542, w_163_543, w_163_544, w_163_552, w_163_553, w_163_554, w_163_555, w_163_556, w_163_557, w_163_559, w_163_561, w_163_565, w_163_567, w_163_569, w_163_571, w_163_573, w_163_576, w_163_578, w_163_580, w_163_583, w_163_586, w_163_596, w_163_598, w_163_600, w_163_603, w_163_607, w_163_609, w_163_611, w_163_614, w_163_616, w_163_617, w_163_618, w_163_619, w_163_628, w_163_629, w_163_632, w_163_636, w_163_639, w_163_640, w_163_642, w_163_647, w_163_648, w_163_650, w_163_651, w_163_655, w_163_656, w_163_657, w_163_660, w_163_661, w_163_663, w_163_664, w_163_670, w_163_671, w_163_672, w_163_675, w_163_676, w_163_678, w_163_679, w_163_682, w_163_683, w_163_685, w_163_686, w_163_687, w_163_688, w_163_690, w_163_692, w_163_693, w_163_697, w_163_698, w_163_699, w_163_703, w_163_704, w_163_705, w_163_708, w_163_710, w_163_712, w_163_714, w_163_719, w_163_725, w_163_726, w_163_729, w_163_731, w_163_732, w_163_735, w_163_742, w_163_744, w_163_747, w_163_748, w_163_749, w_163_751, w_163_753, w_163_754, w_163_759, w_163_761, w_163_763, w_163_766, w_163_772, w_163_773, w_163_775, w_163_776, w_163_778, w_163_782, w_163_783, w_163_786, w_163_789, w_163_790, w_163_796, w_163_800, w_163_801, w_163_803, w_163_804, w_163_805, w_163_809, w_163_811, w_163_812, w_163_813, w_163_814, w_163_815, w_163_822, w_163_823, w_163_828, w_163_829, w_163_830, w_163_833, w_163_834, w_163_836, w_163_837, w_163_839, w_163_840, w_163_843, w_163_850, w_163_851, w_163_852, w_163_853, w_163_854, w_163_855, w_163_859, w_163_860, w_163_862, w_163_863, w_163_865, w_163_866, w_163_868, w_163_871, w_163_872, w_163_875, w_163_879, w_163_883, w_163_884, w_163_887, w_163_888, w_163_889, w_163_891, w_163_893, w_163_894, w_163_895, w_163_897, w_163_900, w_163_905, w_163_906, w_163_907, w_163_910, w_163_913, w_163_915, w_163_919, w_163_923, w_163_925, w_163_926, w_163_927, w_163_928, w_163_931, w_163_934, w_163_935, w_163_938, w_163_941, w_163_945, w_163_946, w_163_947, w_163_948, w_163_950, w_163_951, w_163_952, w_163_954, w_163_955, w_163_958, w_163_963, w_163_964, w_163_965, w_163_966, w_163_968, w_163_969, w_163_970, w_163_971, w_163_974, w_163_976, w_163_978, w_163_986, w_163_987, w_163_989, w_163_990, w_163_992, w_163_995, w_163_996, w_163_1001, w_163_1004, w_163_1005, w_163_1007, w_163_1008, w_163_1011, w_163_1014, w_163_1017, w_163_1019, w_163_1021, w_163_1024, w_163_1025, w_163_1026, w_163_1029, w_163_1033, w_163_1037, w_163_1044, w_163_1045, w_163_1046, w_163_1047, w_163_1048, w_163_1049, w_163_1051, w_163_1052, w_163_1054, w_163_1055, w_163_1059, w_163_1062, w_163_1066, w_163_1068, w_163_1073, w_163_1076, w_163_1082, w_163_1085, w_163_1086, w_163_1090, w_163_1095, w_163_1098, w_163_1107, w_163_1108, w_163_1111, w_163_1114, w_163_1115, w_163_1116, w_163_1120, w_163_1125, w_163_1126, w_163_1133, w_163_1134, w_163_1136, w_163_1139, w_163_1144, w_163_1145, w_163_1149, w_163_1156, w_163_1158, w_163_1163, w_163_1164, w_163_1167, w_163_1170, w_163_1173, w_163_1176, w_163_1184, w_163_1186, w_163_1188, w_163_1189, w_163_1192, w_163_1195, w_163_1197, w_163_1198, w_163_1204, w_163_1210, w_163_1212, w_163_1213, w_163_1216, w_163_1219, w_163_1220, w_163_1221, w_163_1225, w_163_1227, w_163_1229, w_163_1230, w_163_1232, w_163_1234, w_163_1235, w_163_1236, w_163_1237, w_163_1239, w_163_1242, w_163_1244, w_163_1249, w_163_1251, w_163_1253, w_163_1255, w_163_1259, w_163_1262, w_163_1263, w_163_1264, w_163_1266, w_163_1267, w_163_1272, w_163_1273, w_163_1278, w_163_1281, w_163_1282, w_163_1284, w_163_1285, w_163_1287, w_163_1290, w_163_1303, w_163_1305, w_163_1313, w_163_1314, w_163_1316, w_163_1318, w_163_1324, w_163_1326, w_163_1330, w_163_1332, w_163_1336, w_163_1339, w_163_1340, w_163_1341, w_163_1353, w_163_1354, w_163_1356, w_163_1357, w_163_1369, w_163_1370, w_163_1373, w_163_1377, w_163_1378, w_163_1388, w_163_1389, w_163_1396, w_163_1398, w_163_1400, w_163_1408, w_163_1412, w_163_1417, w_163_1418, w_163_1425, w_163_1427, w_163_1431, w_163_1433, w_163_1436, w_163_1438, w_163_1442, w_163_1447, w_163_1448, w_163_1449, w_163_1453, w_163_1454, w_163_1457, w_163_1458, w_163_1464, w_163_1465, w_163_1467, w_163_1470, w_163_1473, w_163_1475, w_163_1478, w_163_1479, w_163_1485, w_163_1490, w_163_1496, w_163_1498, w_163_1499, w_163_1500, w_163_1508, w_163_1512, w_163_1514, w_163_1519, w_163_1521, w_163_1525, w_163_1526, w_163_1531, w_163_1533, w_163_1537, w_163_1543, w_163_1545, w_163_1546, w_163_1550, w_163_1553, w_163_1554, w_163_1558, w_163_1563, w_163_1564, w_163_1567, w_163_1572, w_163_1574, w_163_1583, w_163_1584, w_163_1585, w_163_1588, w_163_1590, w_163_1597, w_163_1598, w_163_1600, w_163_1602, w_163_1605, w_163_1606, w_163_1607, w_163_1610, w_163_1620, w_163_1630, w_163_1640, w_163_1645, w_163_1646, w_163_1653, w_163_1658, w_163_1659, w_163_1661, w_163_1663, w_163_1670, w_163_1671, w_163_1673, w_163_1676, w_163_1678, w_163_1679, w_163_1687, w_163_1688, w_163_1690, w_163_1692, w_163_1695, w_163_1696, w_163_1699, w_163_1701, w_163_1705, w_163_1710, w_163_1712, w_163_1716, w_163_1726, w_163_1728, w_163_1731, w_163_1732, w_163_1736, w_163_1740, w_163_1747, w_163_1757, w_163_1760, w_163_1761, w_163_1765, w_163_1772, w_163_1774, w_163_1775, w_163_1779, w_163_1787, w_163_1798, w_163_1803, w_163_1805, w_163_1806, w_163_1808, w_163_1818, w_163_1820, w_163_1826, w_163_1835, w_163_1836, w_163_1838, w_163_1840, w_163_1842, w_163_1846, w_163_1852, w_163_1854, w_163_1857, w_163_1858, w_163_1859, w_163_1862;
  wire w_164_000, w_164_001, w_164_002, w_164_003, w_164_004, w_164_005, w_164_006, w_164_007, w_164_008, w_164_009, w_164_010, w_164_011, w_164_012, w_164_013;
  wire w_165_000, w_165_002, w_165_004, w_165_006, w_165_007, w_165_010, w_165_011, w_165_016, w_165_018, w_165_019, w_165_020, w_165_022, w_165_024, w_165_025, w_165_026, w_165_029, w_165_038, w_165_040, w_165_041, w_165_043, w_165_044, w_165_045, w_165_046, w_165_048, w_165_051, w_165_052, w_165_054, w_165_055, w_165_056, w_165_057, w_165_058, w_165_059, w_165_061, w_165_062, w_165_063, w_165_069, w_165_071, w_165_077, w_165_079, w_165_080, w_165_082, w_165_086, w_165_089, w_165_090, w_165_097, w_165_099, w_165_100, w_165_103, w_165_104, w_165_107, w_165_108, w_165_109, w_165_110, w_165_112, w_165_120, w_165_121, w_165_125, w_165_127, w_165_128, w_165_134, w_165_137, w_165_139, w_165_142, w_165_143, w_165_144, w_165_147, w_165_148, w_165_149, w_165_150, w_165_152, w_165_156, w_165_160, w_165_162, w_165_163, w_165_164, w_165_165, w_165_170, w_165_173, w_165_174, w_165_176, w_165_177, w_165_179, w_165_180, w_165_183, w_165_184, w_165_186, w_165_192, w_165_196, w_165_200, w_165_204, w_165_207, w_165_208, w_165_212, w_165_216, w_165_218, w_165_219, w_165_221, w_165_222, w_165_223, w_165_229, w_165_232, w_165_237, w_165_239, w_165_242, w_165_249, w_165_251, w_165_253, w_165_254, w_165_255, w_165_256, w_165_258, w_165_262, w_165_266, w_165_267, w_165_268, w_165_271, w_165_276, w_165_277, w_165_279, w_165_281, w_165_286, w_165_292, w_165_294, w_165_295, w_165_298, w_165_299, w_165_300, w_165_303, w_165_304, w_165_305, w_165_310, w_165_311, w_165_314, w_165_316, w_165_318, w_165_321, w_165_323, w_165_324, w_165_325, w_165_327, w_165_329, w_165_331, w_165_332, w_165_333, w_165_336, w_165_337, w_165_340, w_165_343, w_165_348, w_165_350, w_165_351, w_165_361, w_165_362, w_165_364, w_165_365, w_165_367, w_165_368, w_165_369, w_165_370, w_165_371, w_165_374, w_165_375, w_165_376, w_165_377, w_165_378, w_165_381, w_165_382, w_165_387, w_165_390, w_165_396, w_165_397, w_165_398, w_165_399, w_165_403, w_165_404, w_165_406, w_165_408, w_165_409, w_165_411, w_165_415, w_165_416, w_165_419, w_165_422, w_165_424, w_165_427, w_165_430, w_165_433, w_165_435, w_165_445, w_165_446, w_165_447, w_165_453, w_165_454, w_165_456, w_165_457, w_165_458, w_165_459, w_165_461, w_165_468, w_165_473, w_165_476, w_165_481, w_165_483, w_165_488, w_165_491, w_165_492, w_165_494, w_165_497, w_165_500, w_165_502, w_165_504, w_165_505, w_165_506, w_165_513, w_165_519, w_165_521, w_165_523, w_165_524, w_165_527, w_165_531, w_165_534, w_165_537, w_165_540, w_165_543, w_165_546, w_165_550, w_165_560, w_165_569, w_165_572, w_165_574, w_165_577, w_165_578, w_165_582, w_165_586, w_165_587, w_165_588, w_165_590, w_165_601, w_165_604, w_165_605, w_165_608, w_165_610, w_165_614, w_165_615, w_165_618, w_165_619, w_165_621, w_165_622, w_165_623, w_165_633, w_165_642, w_165_644, w_165_645, w_165_650, w_165_654, w_165_662, w_165_663, w_165_664, w_165_665, w_165_666, w_165_667, w_165_670, w_165_671, w_165_674, w_165_675, w_165_679, w_165_680, w_165_682, w_165_687, w_165_688, w_165_690, w_165_693, w_165_701, w_165_703, w_165_705, w_165_707, w_165_713, w_165_714, w_165_715, w_165_721, w_165_722, w_165_724, w_165_730, w_165_731, w_165_733, w_165_737, w_165_739, w_165_742, w_165_751, w_165_758, w_165_760, w_165_761, w_165_766, w_165_767, w_165_768, w_165_769, w_165_772, w_165_776, w_165_789, w_165_790, w_165_796, w_165_797, w_165_801, w_165_802, w_165_808, w_165_817, w_165_818, w_165_823, w_165_824, w_165_825, w_165_828, w_165_835, w_165_838, w_165_839, w_165_842, w_165_843, w_165_844, w_165_848, w_165_853, w_165_855, w_165_860, w_165_861, w_165_872, w_165_873, w_165_874, w_165_883, w_165_885, w_165_894, w_165_899, w_165_906, w_165_912, w_165_914, w_165_922, w_165_923, w_165_924, w_165_930, w_165_931, w_165_934, w_165_935, w_165_937, w_165_938, w_165_939, w_165_947, w_165_948, w_165_952, w_165_953, w_165_954, w_165_955, w_165_958, w_165_959, w_165_960, w_165_962, w_165_965, w_165_967, w_165_971, w_165_972, w_165_975, w_165_977, w_165_987, w_165_988, w_165_989, w_165_990, w_165_996, w_165_1001, w_165_1002, w_165_1003, w_165_1006, w_165_1007, w_165_1009, w_165_1010, w_165_1012, w_165_1013, w_165_1014, w_165_1015, w_165_1019, w_165_1020, w_165_1021, w_165_1023, w_165_1024, w_165_1029, w_165_1030, w_165_1031, w_165_1036, w_165_1040, w_165_1041, w_165_1042, w_165_1043, w_165_1046, w_165_1047, w_165_1048, w_165_1050, w_165_1051, w_165_1055, w_165_1057, w_165_1061, w_165_1068, w_165_1074, w_165_1077, w_165_1081, w_165_1092, w_165_1093, w_165_1095, w_165_1097, w_165_1099, w_165_1102, w_165_1103, w_165_1109, w_165_1110, w_165_1113, w_165_1118, w_165_1119, w_165_1125, w_165_1132, w_165_1133, w_165_1134, w_165_1136, w_165_1139, w_165_1140, w_165_1143, w_165_1144, w_165_1150, w_165_1153, w_165_1155, w_165_1156, w_165_1161, w_165_1163, w_165_1164, w_165_1167, w_165_1177, w_165_1186, w_165_1188, w_165_1192, w_165_1194, w_165_1195, w_165_1202, w_165_1205, w_165_1209, w_165_1211, w_165_1219, w_165_1221, w_165_1224, w_165_1227, w_165_1233, w_165_1235, w_165_1236, w_165_1237, w_165_1239, w_165_1241, w_165_1244, w_165_1248, w_165_1251, w_165_1258, w_165_1262, w_165_1264, w_165_1267, w_165_1278, w_165_1281, w_165_1296, w_165_1297, w_165_1308, w_165_1309, w_165_1312, w_165_1313, w_165_1318, w_165_1326, w_165_1327, w_165_1328, w_165_1333, w_165_1334, w_165_1337, w_165_1340, w_165_1342, w_165_1348, w_165_1349, w_165_1350, w_165_1351, w_165_1352, w_165_1359, w_165_1360, w_165_1370, w_165_1372, w_165_1373, w_165_1375, w_165_1383, w_165_1385, w_165_1392, w_165_1393, w_165_1399, w_165_1400, w_165_1402, w_165_1405, w_165_1407, w_165_1408, w_165_1409, w_165_1410, w_165_1414, w_165_1416, w_165_1420, w_165_1424, w_165_1426, w_165_1428, w_165_1431, w_165_1436, w_165_1440, w_165_1441, w_165_1448, w_165_1450, w_165_1452, w_165_1454, w_165_1465, w_165_1466, w_165_1467, w_165_1468, w_165_1475, w_165_1479, w_165_1482, w_165_1483, w_165_1487, w_165_1490, w_165_1492, w_165_1496, w_165_1502, w_165_1504, w_165_1506, w_165_1514, w_165_1517, w_165_1519, w_165_1526, w_165_1527, w_165_1530, w_165_1534, w_165_1536, w_165_1542, w_165_1543, w_165_1550, w_165_1551, w_165_1552, w_165_1555, w_165_1556, w_165_1561, w_165_1562, w_165_1566, w_165_1568, w_165_1569, w_165_1570, w_165_1573, w_165_1575, w_165_1576, w_165_1579, w_165_1583, w_165_1591, w_165_1593, w_165_1594, w_165_1597, w_165_1598, w_165_1600, w_165_1601, w_165_1606, w_165_1608, w_165_1609, w_165_1611, w_165_1612, w_165_1622, w_165_1623, w_165_1624, w_165_1625, w_165_1628, w_165_1636, w_165_1639, w_165_1640, w_165_1642, w_165_1645, w_165_1650, w_165_1651, w_165_1661, w_165_1662, w_165_1663, w_165_1665, w_165_1673, w_165_1678, w_165_1680, w_165_1683, w_165_1684, w_165_1688, w_165_1693, w_165_1707, w_165_1708, w_165_1709, w_165_1715, w_165_1717, w_165_1724, w_165_1727, w_165_1732, w_165_1741, w_165_1752, w_165_1760, w_165_1763, w_165_1767, w_165_1768, w_165_1769, w_165_1772, w_165_1775, w_165_1776, w_165_1777, w_165_1778, w_165_1779, w_165_1780, w_165_1782, w_165_1786, w_165_1795, w_165_1798, w_165_1805, w_165_1809, w_165_1812, w_165_1813, w_165_1814, w_165_1817, w_165_1825, w_165_1827, w_165_1828, w_165_1834, w_165_1839, w_165_1841, w_165_1844, w_165_1852, w_165_1855, w_165_1857, w_165_1860, w_165_1861, w_165_1864, w_165_1868, w_165_1872, w_165_1890, w_165_1892, w_165_1893, w_165_1894, w_165_1895, w_165_1898, w_165_1908, w_165_1914, w_165_1918, w_165_1920, w_165_1922, w_165_1924, w_165_1928, w_165_1930, w_165_1931, w_165_1932, w_165_1941, w_165_1955, w_165_1963, w_165_1973, w_165_1974, w_165_1978, w_165_1984, w_165_1988, w_165_1989, w_165_1990, w_165_1991, w_165_1992, w_165_1995, w_165_1997, w_165_1999, w_165_2000, w_165_2002, w_165_2004, w_165_2005, w_165_2009, w_165_2025, w_165_2026, w_165_2028, w_165_2030, w_165_2031, w_165_2036, w_165_2038, w_165_2039, w_165_2042, w_165_2044, w_165_2048, w_165_2050, w_165_2052, w_165_2054, w_165_2055, w_165_2056, w_165_2057, w_165_2058, w_165_2059, w_165_2061, w_165_2067, w_165_2068, w_165_2075, w_165_2080, w_165_2083, w_165_2089, w_165_2092, w_165_2102, w_165_2104, w_165_2107, w_165_2112, w_165_2117, w_165_2118, w_165_2121, w_165_2124, w_165_2125, w_165_2130, w_165_2131, w_165_2132, w_165_2135, w_165_2136, w_165_2137, w_165_2144, w_165_2146, w_165_2149, w_165_2150, w_165_2154, w_165_2155, w_165_2160, w_165_2163, w_165_2165, w_165_2173, w_165_2174, w_165_2191, w_165_2192, w_165_2193, w_165_2195, w_165_2197, w_165_2199, w_165_2209, w_165_2211, w_165_2215, w_165_2216, w_165_2219, w_165_2222, w_165_2225, w_165_2226, w_165_2229, w_165_2230, w_165_2233, w_165_2236, w_165_2239, w_165_2246, w_165_2250, w_165_2252, w_165_2253, w_165_2254, w_165_2255, w_165_2256, w_165_2260, w_165_2261, w_165_2262, w_165_2263, w_165_2264, w_165_2265, w_165_2267, w_165_2269, w_165_2270, w_165_2271, w_165_2272, w_165_2273, w_165_2274, w_165_2275, w_165_2277, w_165_2279, w_165_2280, w_165_2281, w_165_2282, w_165_2283, w_165_2284, w_165_2286, w_165_2288, w_165_2289, w_165_2290, w_165_2291, w_165_2292, w_165_2293, w_165_2294, w_165_2295, w_165_2296, w_165_2297, w_165_2299, w_165_2301, w_165_2302, w_165_2303, w_165_2304, w_165_2305, w_165_2306, w_165_2307, w_165_2308, w_165_2309, w_165_2310, w_165_2312;
  wire w_166_000, w_166_004, w_166_005, w_166_006, w_166_007, w_166_008, w_166_011, w_166_014, w_166_016, w_166_017, w_166_025, w_166_027, w_166_033, w_166_035, w_166_038, w_166_042, w_166_047, w_166_051, w_166_060, w_166_061, w_166_064, w_166_069, w_166_071, w_166_082, w_166_086, w_166_093, w_166_096, w_166_110, w_166_111, w_166_112, w_166_117, w_166_118, w_166_120, w_166_129, w_166_132, w_166_134, w_166_140, w_166_142, w_166_144, w_166_149, w_166_152, w_166_153, w_166_164, w_166_165, w_166_168, w_166_169, w_166_170, w_166_172, w_166_177, w_166_188, w_166_189, w_166_190, w_166_193, w_166_212, w_166_213, w_166_219, w_166_222, w_166_223, w_166_226, w_166_229, w_166_235, w_166_245, w_166_253, w_166_257, w_166_259, w_166_260, w_166_261, w_166_264, w_166_267, w_166_273, w_166_280, w_166_283, w_166_290, w_166_291, w_166_292, w_166_294, w_166_295, w_166_298, w_166_301, w_166_310, w_166_316, w_166_323, w_166_332, w_166_335, w_166_341, w_166_345, w_166_349, w_166_351, w_166_357, w_166_358, w_166_359, w_166_361, w_166_362, w_166_371, w_166_377, w_166_379, w_166_381, w_166_382, w_166_384, w_166_387, w_166_389, w_166_393, w_166_394, w_166_398, w_166_399, w_166_403, w_166_406, w_166_415, w_166_421, w_166_438, w_166_439, w_166_441, w_166_446, w_166_447, w_166_448, w_166_449, w_166_451, w_166_452, w_166_460, w_166_463, w_166_469, w_166_470, w_166_472, w_166_473, w_166_476, w_166_481, w_166_483, w_166_487, w_166_489, w_166_490, w_166_492, w_166_498, w_166_499, w_166_501, w_166_502, w_166_506, w_166_509, w_166_515, w_166_522, w_166_527, w_166_529, w_166_532, w_166_540, w_166_547, w_166_550, w_166_553, w_166_558, w_166_559, w_166_564, w_166_565, w_166_568, w_166_569, w_166_570, w_166_572, w_166_579, w_166_580, w_166_583, w_166_587, w_166_593, w_166_594, w_166_599, w_166_602, w_166_603, w_166_607, w_166_609, w_166_611, w_166_612, w_166_613, w_166_614, w_166_615, w_166_629, w_166_631, w_166_634, w_166_636, w_166_639, w_166_642, w_166_646, w_166_651, w_166_660, w_166_661, w_166_662, w_166_671, w_166_673, w_166_677, w_166_681, w_166_682, w_166_683, w_166_688, w_166_691, w_166_693, w_166_695, w_166_697, w_166_700, w_166_702, w_166_711, w_166_712, w_166_714, w_166_729, w_166_736, w_166_740, w_166_741, w_166_742, w_166_745, w_166_749, w_166_755, w_166_756, w_166_757, w_166_758, w_166_760, w_166_764, w_166_765, w_166_771, w_166_774, w_166_775, w_166_781, w_166_790, w_166_801, w_166_818, w_166_823, w_166_824, w_166_826, w_166_828, w_166_829, w_166_833, w_166_834, w_166_835, w_166_836, w_166_847, w_166_850, w_166_851, w_166_852, w_166_853, w_166_854, w_166_855, w_166_859, w_166_860, w_166_861, w_166_866, w_166_871, w_166_874, w_166_884, w_166_887, w_166_892, w_166_896, w_166_897, w_166_905, w_166_908, w_166_911, w_166_912, w_166_913, w_166_914, w_166_921, w_166_927, w_166_928, w_166_929, w_166_930, w_166_934, w_166_937, w_166_943, w_166_945, w_166_948, w_166_951, w_166_955, w_166_960, w_166_963, w_166_966, w_166_969, w_166_970, w_166_973, w_166_976, w_166_977, w_166_980, w_166_984, w_166_988, w_166_989, w_166_991, w_166_996, w_166_1003, w_166_1012, w_166_1013, w_166_1014, w_166_1018, w_166_1020, w_166_1025, w_166_1035, w_166_1038, w_166_1043, w_166_1048, w_166_1056, w_166_1058, w_166_1066, w_166_1078, w_166_1081, w_166_1082, w_166_1083, w_166_1084, w_166_1089, w_166_1090, w_166_1100, w_166_1102, w_166_1105, w_166_1107, w_166_1108, w_166_1111, w_166_1117, w_166_1120, w_166_1127, w_166_1133, w_166_1141, w_166_1142, w_166_1143, w_166_1145, w_166_1148, w_166_1151, w_166_1152, w_166_1155, w_166_1158, w_166_1159, w_166_1163, w_166_1164, w_166_1165, w_166_1166, w_166_1173, w_166_1178, w_166_1182, w_166_1185, w_166_1187, w_166_1190, w_166_1194, w_166_1197, w_166_1198, w_166_1199, w_166_1202, w_166_1203, w_166_1205, w_166_1206, w_166_1208, w_166_1212, w_166_1213, w_166_1214, w_166_1215, w_166_1223, w_166_1225, w_166_1227, w_166_1229, w_166_1230, w_166_1234, w_166_1235, w_166_1236, w_166_1241, w_166_1247, w_166_1249, w_166_1251, w_166_1259, w_166_1271, w_166_1277, w_166_1278, w_166_1281, w_166_1283, w_166_1284, w_166_1285, w_166_1287, w_166_1290, w_166_1291, w_166_1293, w_166_1294, w_166_1295, w_166_1297, w_166_1298, w_166_1299, w_166_1301, w_166_1302, w_166_1303, w_166_1306, w_166_1309, w_166_1310, w_166_1318, w_166_1322, w_166_1332, w_166_1335, w_166_1344, w_166_1348, w_166_1351, w_166_1353, w_166_1370, w_166_1373, w_166_1378, w_166_1380, w_166_1386, w_166_1387, w_166_1392, w_166_1395, w_166_1396, w_166_1397, w_166_1399, w_166_1400, w_166_1401, w_166_1404, w_166_1405, w_166_1407, w_166_1411, w_166_1414, w_166_1417, w_166_1419, w_166_1420, w_166_1422, w_166_1423, w_166_1425, w_166_1426, w_166_1427, w_166_1428, w_166_1429, w_166_1430, w_166_1433, w_166_1434, w_166_1435, w_166_1436, w_166_1439, w_166_1441, w_166_1448, w_166_1449, w_166_1457, w_166_1458, w_166_1460, w_166_1461, w_166_1462, w_166_1464, w_166_1466, w_166_1472, w_166_1473, w_166_1474, w_166_1479, w_166_1481, w_166_1482, w_166_1484, w_166_1493, w_166_1497, w_166_1501, w_166_1502, w_166_1504, w_166_1508, w_166_1511, w_166_1515, w_166_1516, w_166_1518, w_166_1519, w_166_1522, w_166_1530, w_166_1531, w_166_1533, w_166_1534, w_166_1542, w_166_1543, w_166_1546, w_166_1554, w_166_1559, w_166_1565, w_166_1566, w_166_1569, w_166_1572, w_166_1573, w_166_1574, w_166_1577, w_166_1585, w_166_1589, w_166_1594, w_166_1596, w_166_1599, w_166_1600, w_166_1611, w_166_1612, w_166_1613, w_166_1614, w_166_1616, w_166_1619, w_166_1620, w_166_1622, w_166_1623, w_166_1625, w_166_1632, w_166_1635, w_166_1641, w_166_1642, w_166_1650, w_166_1651, w_166_1652, w_166_1658, w_166_1660, w_166_1663, w_166_1664, w_166_1667, w_166_1674, w_166_1676, w_166_1679, w_166_1680, w_166_1681, w_166_1682, w_166_1683, w_166_1685, w_166_1689, w_166_1690, w_166_1692, w_166_1695, w_166_1700, w_166_1702, w_166_1703, w_166_1714, w_166_1725, w_166_1729, w_166_1734, w_166_1741, w_166_1742, w_166_1746, w_166_1756, w_166_1767, w_166_1773, w_166_1780, w_166_1784, w_166_1786, w_166_1793, w_166_1795, w_166_1798, w_166_1803, w_166_1804, w_166_1805, w_166_1815, w_166_1819, w_166_1821, w_166_1827, w_166_1828, w_166_1833, w_166_1836, w_166_1842, w_166_1847, w_166_1848, w_166_1850, w_166_1851, w_166_1859, w_166_1860, w_166_1864, w_166_1873, w_166_1874, w_166_1879, w_166_1881, w_166_1886, w_166_1888, w_166_1899, w_166_1909, w_166_1910, w_166_1912, w_166_1913, w_166_1915, w_166_1917, w_166_1919, w_166_1920, w_166_1925, w_166_1927, w_166_1931, w_166_1933, w_166_1934, w_166_1935, w_166_1941, w_166_1943, w_166_1944, w_166_1948, w_166_1952, w_166_1961, w_166_1962, w_166_1969, w_166_1973, w_166_1976, w_166_1978, w_166_1981, w_166_1982, w_166_1983, w_166_1984, w_166_1986, w_166_1996, w_166_1998, w_166_2009, w_166_2019, w_166_2021, w_166_2024, w_166_2026, w_166_2029, w_166_2032, w_166_2033, w_166_2035, w_166_2043, w_166_2045, w_166_2047, w_166_2049, w_166_2053, w_166_2054, w_166_2056, w_166_2057, w_166_2058, w_166_2067, w_166_2074, w_166_2085, w_166_2088, w_166_2092, w_166_2093, w_166_2096, w_166_2098, w_166_2099, w_166_2107, w_166_2123, w_166_2128, w_166_2135, w_166_2137, w_166_2142, w_166_2145, w_166_2147, w_166_2148, w_166_2155, w_166_2163, w_166_2164, w_166_2172, w_166_2173, w_166_2175, w_166_2187, w_166_2191, w_166_2207, w_166_2208, w_166_2211, w_166_2230, w_166_2240, w_166_2242, w_166_2244, w_166_2248, w_166_2257, w_166_2265, w_166_2268, w_166_2281, w_166_2285, w_166_2288, w_166_2290, w_166_2297, w_166_2302, w_166_2305, w_166_2309, w_166_2311, w_166_2314, w_166_2318, w_166_2320, w_166_2324, w_166_2326, w_166_2330, w_166_2332, w_166_2333, w_166_2335, w_166_2338, w_166_2339, w_166_2343, w_166_2347, w_166_2357, w_166_2372, w_166_2383, w_166_2391, w_166_2392, w_166_2402, w_166_2414, w_166_2425, w_166_2437, w_166_2439, w_166_2440, w_166_2444, w_166_2448, w_166_2458, w_166_2466, w_166_2470, w_166_2474, w_166_2477, w_166_2484, w_166_2488, w_166_2494, w_166_2498, w_166_2499, w_166_2500, w_166_2507, w_166_2514, w_166_2515, w_166_2518, w_166_2528, w_166_2533, w_166_2542, w_166_2552, w_166_2563, w_166_2565, w_166_2570, w_166_2571, w_166_2574, w_166_2575, w_166_2587, w_166_2609, w_166_2612, w_166_2613, w_166_2620, w_166_2622, w_166_2629, w_166_2637, w_166_2643, w_166_2647, w_166_2649, w_166_2665, w_166_2666, w_166_2674, w_166_2682, w_166_2725, w_166_2730, w_166_2734, w_166_2736, w_166_2739, w_166_2775, w_166_2779, w_166_2785, w_166_2787, w_166_2791, w_166_2797, w_166_2799, w_166_2802, w_166_2805, w_166_2815, w_166_2816, w_166_2830, w_166_2834, w_166_2840, w_166_2844, w_166_2845, w_166_2847, w_166_2850, w_166_2856, w_166_2867, w_166_2871, w_166_2872, w_166_2876, w_166_2878, w_166_2885, w_166_2887, w_166_2899, w_166_2910, w_166_2913, w_166_2915, w_166_2918, w_166_2920, w_166_2921, w_166_2928, w_166_2937, w_166_2938, w_166_2939, w_166_2942, w_166_2943, w_166_2944, w_166_2945, w_166_2946, w_166_2947, w_166_2948, w_166_2949, w_166_2950;
  wire w_167_001, w_167_003, w_167_004, w_167_005, w_167_006, w_167_009, w_167_012, w_167_014, w_167_016, w_167_017, w_167_018, w_167_021, w_167_023, w_167_025, w_167_026, w_167_028, w_167_029, w_167_031, w_167_033, w_167_035, w_167_036, w_167_037, w_167_038, w_167_039, w_167_041, w_167_042, w_167_044, w_167_045, w_167_048, w_167_050, w_167_054, w_167_056, w_167_057, w_167_058, w_167_060, w_167_061, w_167_062, w_167_063, w_167_064, w_167_067, w_167_068, w_167_069, w_167_070, w_167_071, w_167_073, w_167_077, w_167_078, w_167_080, w_167_085, w_167_087, w_167_088, w_167_090, w_167_094, w_167_095, w_167_096, w_167_099, w_167_100, w_167_101, w_167_102, w_167_106, w_167_107, w_167_108, w_167_112, w_167_114, w_167_116, w_167_117, w_167_118, w_167_119, w_167_120, w_167_123, w_167_124, w_167_126, w_167_131, w_167_132, w_167_133, w_167_134, w_167_135, w_167_137, w_167_139, w_167_140, w_167_141, w_167_142, w_167_143, w_167_144, w_167_145, w_167_146, w_167_149, w_167_152, w_167_153, w_167_154, w_167_155, w_167_157, w_167_162, w_167_163, w_167_164, w_167_166, w_167_167, w_167_168, w_167_169, w_167_171, w_167_172, w_167_176, w_167_179, w_167_180, w_167_182, w_167_183, w_167_185, w_167_186, w_167_187, w_167_188, w_167_189, w_167_191, w_167_192, w_167_193, w_167_194, w_167_195, w_167_196, w_167_199, w_167_200, w_167_203, w_167_204, w_167_206, w_167_209, w_167_210, w_167_211, w_167_212, w_167_213, w_167_215, w_167_217, w_167_218, w_167_219, w_167_222, w_167_224, w_167_225, w_167_226, w_167_227, w_167_228, w_167_234, w_167_235, w_167_236, w_167_237, w_167_238, w_167_240, w_167_241, w_167_242, w_167_244, w_167_245, w_167_246, w_167_247, w_167_248, w_167_250, w_167_252, w_167_256, w_167_258, w_167_260, w_167_262, w_167_263, w_167_266, w_167_267, w_167_269, w_167_270, w_167_273, w_167_276, w_167_277, w_167_281, w_167_284, w_167_285, w_167_286, w_167_288, w_167_292, w_167_293, w_167_294, w_167_295, w_167_296, w_167_297, w_167_299, w_167_300, w_167_301, w_167_302, w_167_304, w_167_305, w_167_309, w_167_310, w_167_311, w_167_314, w_167_315, w_167_317, w_167_318, w_167_319, w_167_320, w_167_321, w_167_322, w_167_323, w_167_325, w_167_326, w_167_328, w_167_329, w_167_331, w_167_333, w_167_336, w_167_337, w_167_339, w_167_341, w_167_343, w_167_345, w_167_346, w_167_348, w_167_349, w_167_350, w_167_351, w_167_353, w_167_356, w_167_357, w_167_359, w_167_360, w_167_362, w_167_364, w_167_366, w_167_368, w_167_370, w_167_372, w_167_373, w_167_377, w_167_379, w_167_380, w_167_381, w_167_382, w_167_384, w_167_385, w_167_387, w_167_389, w_167_390, w_167_392, w_167_394, w_167_397, w_167_399, w_167_400, w_167_402, w_167_403, w_167_405, w_167_406, w_167_409, w_167_410, w_167_411, w_167_412, w_167_413, w_167_414, w_167_415, w_167_416, w_167_418, w_167_419, w_167_426, w_167_427, w_167_428, w_167_429, w_167_430, w_167_432, w_167_433, w_167_434, w_167_438, w_167_439, w_167_440, w_167_441, w_167_444, w_167_445, w_167_446, w_167_447, w_167_448, w_167_449, w_167_452, w_167_454, w_167_456, w_167_458, w_167_459, w_167_461, w_167_462, w_167_465, w_167_468, w_167_469, w_167_470, w_167_471, w_167_472, w_167_474, w_167_475, w_167_476, w_167_481, w_167_484, w_167_485, w_167_488, w_167_489, w_167_490, w_167_492, w_167_495, w_167_497, w_167_499, w_167_500, w_167_501, w_167_502, w_167_503, w_167_506, w_167_507, w_167_508, w_167_513, w_167_519, w_167_520, w_167_522, w_167_523, w_167_524, w_167_525, w_167_526, w_167_529, w_167_531, w_167_532, w_167_534, w_167_538, w_167_539, w_167_543, w_167_546, w_167_547, w_167_549, w_167_551, w_167_553, w_167_555, w_167_557, w_167_558, w_167_559, w_167_561, w_167_564, w_167_566, w_167_567, w_167_568, w_167_571, w_167_572, w_167_575, w_167_577, w_167_578, w_167_580, w_167_584, w_167_586, w_167_587, w_167_589, w_167_591, w_167_596, w_167_599, w_167_600, w_167_602, w_167_604, w_167_608, w_167_611, w_167_613, w_167_614, w_167_616, w_167_617, w_167_621, w_167_622, w_167_625, w_167_626, w_167_628, w_167_629, w_167_632, w_167_635, w_167_638, w_167_640, w_167_641, w_167_644, w_167_646, w_167_648, w_167_649, w_167_653, w_167_656, w_167_657, w_167_659, w_167_660, w_167_661, w_167_662, w_167_663, w_167_665, w_167_666, w_167_669, w_167_672, w_167_675, w_167_676, w_167_680, w_167_681, w_167_683, w_167_687, w_167_689, w_167_693, w_167_694, w_167_695, w_167_696, w_167_697, w_167_698, w_167_699, w_167_700, w_167_702, w_167_703, w_167_704, w_167_706, w_167_708, w_167_712, w_167_713, w_167_714, w_167_715, w_167_717, w_167_719, w_167_720, w_167_721, w_167_723, w_167_727, w_167_728, w_167_730, w_167_733, w_167_734, w_167_735, w_167_736, w_167_739, w_167_741, w_167_742, w_167_743, w_167_744, w_167_747, w_167_748, w_167_749, w_167_750, w_167_751, w_167_752, w_167_753, w_167_754, w_167_758, w_167_760, w_167_761, w_167_762, w_167_764, w_167_765, w_167_766, w_167_767, w_167_768, w_167_771, w_167_772, w_167_773, w_167_777, w_167_779, w_167_784, w_167_785, w_167_790, w_167_793, w_167_797, w_167_798, w_167_799, w_167_800, w_167_802, w_167_804, w_167_805, w_167_806, w_167_807, w_167_809, w_167_810, w_167_812, w_167_814, w_167_815, w_167_816, w_167_817, w_167_818, w_167_819, w_167_820, w_167_824, w_167_827, w_167_829, w_167_830, w_167_832, w_167_833, w_167_834, w_167_835, w_167_838, w_167_839, w_167_843, w_167_845, w_167_847, w_167_848, w_167_849, w_167_850, w_167_852, w_167_855, w_167_857, w_167_859, w_167_860, w_167_861, w_167_864, w_167_868, w_167_869, w_167_871, w_167_872, w_167_873, w_167_874, w_167_875, w_167_876, w_167_879, w_167_880, w_167_881, w_167_886, w_167_890, w_167_893, w_167_896, w_167_900, w_167_903, w_167_904, w_167_906, w_167_908, w_167_911, w_167_912, w_167_913, w_167_916, w_167_917, w_167_918, w_167_919, w_167_922, w_167_923, w_167_924, w_167_925, w_167_926, w_167_927, w_167_928, w_167_934, w_167_937, w_167_938, w_167_939, w_167_940, w_167_941, w_167_942, w_167_943, w_167_944, w_167_945, w_167_946, w_167_949, w_167_954, w_167_957, w_167_958, w_167_960, w_167_961, w_167_962, w_167_963, w_167_964, w_167_966, w_167_968, w_167_970, w_167_975, w_167_977, w_167_978, w_167_980, w_167_981, w_167_982, w_167_983, w_167_984, w_167_985, w_167_986, w_167_987, w_167_988, w_167_990, w_167_991, w_167_992, w_167_995, w_167_997, w_167_1000, w_167_1003, w_167_1004, w_167_1005, w_167_1007, w_167_1009, w_167_1014, w_167_1017, w_167_1019, w_167_1023, w_167_1024, w_167_1025, w_167_1027, w_167_1029, w_167_1030, w_167_1033, w_167_1034, w_167_1039, w_167_1040, w_167_1041, w_167_1046, w_167_1049, w_167_1050, w_167_1052, w_167_1053, w_167_1059, w_167_1060, w_167_1064, w_167_1066, w_167_1067, w_167_1069, w_167_1070, w_167_1073, w_167_1077, w_167_1078, w_167_1079, w_167_1081, w_167_1082, w_167_1083, w_167_1085, w_167_1088, w_167_1092, w_167_1093, w_167_1094, w_167_1096, w_167_1098, w_167_1106, w_167_1107, w_167_1108, w_167_1111, w_167_1115, w_167_1116, w_167_1118, w_167_1122, w_167_1125, w_167_1126, w_167_1127, w_167_1128, w_167_1129, w_167_1130, w_167_1132;
  wire w_168_000, w_168_004, w_168_008, w_168_012, w_168_013, w_168_015, w_168_016, w_168_018, w_168_019, w_168_024, w_168_026, w_168_027, w_168_031, w_168_038, w_168_043, w_168_044, w_168_047, w_168_049, w_168_051, w_168_053, w_168_055, w_168_057, w_168_060, w_168_063, w_168_065, w_168_068, w_168_069, w_168_073, w_168_074, w_168_076, w_168_077, w_168_078, w_168_080, w_168_083, w_168_084, w_168_085, w_168_087, w_168_088, w_168_091, w_168_092, w_168_098, w_168_101, w_168_102, w_168_105, w_168_110, w_168_111, w_168_113, w_168_118, w_168_119, w_168_122, w_168_123, w_168_124, w_168_125, w_168_127, w_168_129, w_168_131, w_168_132, w_168_133, w_168_134, w_168_135, w_168_136, w_168_137, w_168_138, w_168_139, w_168_141, w_168_142, w_168_143, w_168_145, w_168_147, w_168_148, w_168_149, w_168_151, w_168_152, w_168_154, w_168_157, w_168_158, w_168_160, w_168_162, w_168_166, w_168_167, w_168_168, w_168_170, w_168_173, w_168_176, w_168_178, w_168_181, w_168_187, w_168_188, w_168_189, w_168_191, w_168_192, w_168_194, w_168_195, w_168_196, w_168_197, w_168_200, w_168_201, w_168_204, w_168_206, w_168_207, w_168_211, w_168_219, w_168_228, w_168_233, w_168_238, w_168_241, w_168_242, w_168_245, w_168_247, w_168_251, w_168_252, w_168_256, w_168_262, w_168_264, w_168_265, w_168_270, w_168_272, w_168_275, w_168_276, w_168_277, w_168_280, w_168_281, w_168_283, w_168_289, w_168_292, w_168_296, w_168_298, w_168_299, w_168_300, w_168_301, w_168_308, w_168_309, w_168_310, w_168_314, w_168_317, w_168_318, w_168_319, w_168_321, w_168_322, w_168_324, w_168_327, w_168_328, w_168_330, w_168_332, w_168_335, w_168_343, w_168_344, w_168_345, w_168_346, w_168_348, w_168_349, w_168_356, w_168_360, w_168_362, w_168_363, w_168_365, w_168_367, w_168_368, w_168_369, w_168_372, w_168_376, w_168_381, w_168_383, w_168_393, w_168_403, w_168_404, w_168_408, w_168_410, w_168_413, w_168_415, w_168_416, w_168_417, w_168_419, w_168_421, w_168_423, w_168_431, w_168_433, w_168_435, w_168_436, w_168_437, w_168_438, w_168_439, w_168_446, w_168_451, w_168_452, w_168_457, w_168_458, w_168_460, w_168_462, w_168_463, w_168_466, w_168_468, w_168_469, w_168_470, w_168_473, w_168_474, w_168_477, w_168_478, w_168_479, w_168_481, w_168_483, w_168_486, w_168_487, w_168_489, w_168_490, w_168_491, w_168_492, w_168_496, w_168_498, w_168_502, w_168_506, w_168_507, w_168_510, w_168_512, w_168_513, w_168_514, w_168_515, w_168_518, w_168_520, w_168_523, w_168_524, w_168_526, w_168_534, w_168_536, w_168_538, w_168_541, w_168_542, w_168_543, w_168_549, w_168_551, w_168_552, w_168_555, w_168_556, w_168_557, w_168_558, w_168_561, w_168_564, w_168_565, w_168_567, w_168_568, w_168_570, w_168_571, w_168_582, w_168_585, w_168_588, w_168_592, w_168_593, w_168_597, w_168_598, w_168_601, w_168_603, w_168_605, w_168_607, w_168_611, w_168_612, w_168_615, w_168_616, w_168_621, w_168_624, w_168_626, w_168_627, w_168_628, w_168_630, w_168_631, w_168_632, w_168_635, w_168_637, w_168_638, w_168_640, w_168_641, w_168_644, w_168_645, w_168_648, w_168_649, w_168_651, w_168_654, w_168_658, w_168_660, w_168_661, w_168_663, w_168_664, w_168_669, w_168_671, w_168_678, w_168_681, w_168_682, w_168_684, w_168_689, w_168_691, w_168_695, w_168_698, w_168_699, w_168_700, w_168_704, w_168_707, w_168_709, w_168_711, w_168_712, w_168_714, w_168_717, w_168_720, w_168_721, w_168_723, w_168_726, w_168_728, w_168_729, w_168_731, w_168_732, w_168_733, w_168_735, w_168_736, w_168_739, w_168_741, w_168_743, w_168_744, w_168_747, w_168_748, w_168_750, w_168_751, w_168_752, w_168_753, w_168_754, w_168_755, w_168_756, w_168_758, w_168_759, w_168_760, w_168_761, w_168_762, w_168_765, w_168_766, w_168_770, w_168_774, w_168_779, w_168_788, w_168_792, w_168_794, w_168_797, w_168_798, w_168_799, w_168_808, w_168_810, w_168_813, w_168_820, w_168_821, w_168_824, w_168_825, w_168_827, w_168_829, w_168_830, w_168_834, w_168_835, w_168_836, w_168_845, w_168_846, w_168_847, w_168_848, w_168_853, w_168_861, w_168_866, w_168_868, w_168_875, w_168_881, w_168_885, w_168_889, w_168_895, w_168_901, w_168_904, w_168_906, w_168_911, w_168_916, w_168_926, w_168_931, w_168_932, w_168_934, w_168_938, w_168_943, w_168_944, w_168_945, w_168_946, w_168_951, w_168_958, w_168_963, w_168_965, w_168_975, w_168_976, w_168_978, w_168_979, w_168_983, w_168_985, w_168_986, w_168_989, w_168_991, w_168_992, w_168_993, w_168_995, w_168_996, w_168_997, w_168_998, w_168_1004, w_168_1006, w_168_1008, w_168_1010, w_168_1013, w_168_1014, w_168_1019, w_168_1029, w_168_1033, w_168_1036, w_168_1041, w_168_1043, w_168_1045, w_168_1050, w_168_1051, w_168_1052, w_168_1055, w_168_1057, w_168_1060, w_168_1065, w_168_1071, w_168_1072, w_168_1074, w_168_1075, w_168_1079, w_168_1081, w_168_1082, w_168_1084, w_168_1091, w_168_1093, w_168_1099, w_168_1106, w_168_1107, w_168_1111, w_168_1112, w_168_1113, w_168_1114, w_168_1119, w_168_1124, w_168_1125, w_168_1127, w_168_1130, w_168_1131, w_168_1137, w_168_1146, w_168_1149, w_168_1151, w_168_1152, w_168_1156, w_168_1163, w_168_1165, w_168_1167, w_168_1172, w_168_1179, w_168_1183, w_168_1184, w_168_1190, w_168_1192, w_168_1203, w_168_1204, w_168_1205, w_168_1210, w_168_1212, w_168_1213, w_168_1218, w_168_1220, w_168_1224, w_168_1230, w_168_1231, w_168_1232, w_168_1234, w_168_1239, w_168_1242, w_168_1243, w_168_1248, w_168_1252, w_168_1257, w_168_1263, w_168_1266, w_168_1272, w_168_1274, w_168_1276, w_168_1277, w_168_1278, w_168_1282, w_168_1285, w_168_1287, w_168_1290, w_168_1294, w_168_1303, w_168_1304, w_168_1305, w_168_1307, w_168_1309, w_168_1312, w_168_1315, w_168_1320, w_168_1321, w_168_1322, w_168_1327, w_168_1328, w_168_1329, w_168_1332, w_168_1333, w_168_1344, w_168_1345, w_168_1352, w_168_1353, w_168_1354, w_168_1360, w_168_1364, w_168_1370, w_168_1374, w_168_1375, w_168_1376, w_168_1380, w_168_1383, w_168_1384, w_168_1385, w_168_1386, w_168_1387, w_168_1388, w_168_1390, w_168_1392, w_168_1395, w_168_1398, w_168_1399, w_168_1404, w_168_1407, w_168_1417, w_168_1418, w_168_1426, w_168_1431, w_168_1432, w_168_1435, w_168_1436, w_168_1440, w_168_1443, w_168_1446, w_168_1447, w_168_1451, w_168_1452, w_168_1453, w_168_1456, w_168_1460, w_168_1462, w_168_1469, w_168_1470, w_168_1479, w_168_1488, w_168_1494, w_168_1498, w_168_1500, w_168_1503, w_168_1508, w_168_1517, w_168_1520, w_168_1529, w_168_1542, w_168_1544, w_168_1545, w_168_1547, w_168_1552, w_168_1554, w_168_1558, w_168_1563, w_168_1564, w_168_1565, w_168_1577, w_168_1578, w_168_1580, w_168_1581, w_168_1582, w_168_1587, w_168_1588, w_168_1594, w_168_1600, w_168_1602, w_168_1605, w_168_1606, w_168_1609, w_168_1610, w_168_1616, w_168_1617, w_168_1618, w_168_1621, w_168_1625, w_168_1627, w_168_1632, w_168_1640, w_168_1646, w_168_1649, w_168_1651, w_168_1652, w_168_1653, w_168_1655, w_168_1656, w_168_1659, w_168_1664, w_168_1665, w_168_1669, w_168_1678, w_168_1681, w_168_1682, w_168_1683, w_168_1686, w_168_1687, w_168_1688, w_168_1690, w_168_1692, w_168_1693, w_168_1712, w_168_1713, w_168_1718, w_168_1722, w_168_1726, w_168_1729, w_168_1731, w_168_1743, w_168_1750, w_168_1755, w_168_1757, w_168_1758, w_168_1763, w_168_1768, w_168_1771, w_168_1772, w_168_1777, w_168_1781, w_168_1782, w_168_1786, w_168_1787, w_168_1791, w_168_1793, w_168_1796, w_168_1800, w_168_1802, w_168_1810, w_168_1814, w_168_1823, w_168_1828, w_168_1831, w_168_1836, w_168_1837, w_168_1840, w_168_1841, w_168_1844, w_168_1857, w_168_1860, w_168_1861, w_168_1862, w_168_1866, w_168_1869, w_168_1873, w_168_1878, w_168_1880, w_168_1885, w_168_1896, w_168_1900, w_168_1901, w_168_1905, w_168_1922, w_168_1923, w_168_1927, w_168_1937, w_168_1941, w_168_1946, w_168_1948, w_168_1950, w_168_1952, w_168_1955, w_168_1957, w_168_1958, w_168_1961, w_168_1963, w_168_1965, w_168_1970, w_168_1972, w_168_1975, w_168_1976, w_168_1980, w_168_1983, w_168_1987, w_168_1988, w_168_1992, w_168_2000, w_168_2003, w_168_2004, w_168_2005, w_168_2007, w_168_2008, w_168_2009, w_168_2019, w_168_2021, w_168_2022, w_168_2024, w_168_2029, w_168_2032, w_168_2034, w_168_2039, w_168_2044, w_168_2060, w_168_2065, w_168_2067, w_168_2068, w_168_2069, w_168_2070, w_168_2074, w_168_2076, w_168_2080, w_168_2086, w_168_2087, w_168_2089, w_168_2090, w_168_2094;
  wire w_169_001, w_169_007, w_169_009, w_169_010, w_169_013, w_169_015, w_169_023, w_169_027, w_169_029, w_169_037, w_169_038, w_169_040, w_169_041, w_169_044, w_169_046, w_169_048, w_169_051, w_169_053, w_169_058, w_169_067, w_169_068, w_169_070, w_169_073, w_169_074, w_169_075, w_169_081, w_169_085, w_169_098, w_169_099, w_169_100, w_169_101, w_169_102, w_169_103, w_169_104, w_169_109, w_169_111, w_169_120, w_169_121, w_169_122, w_169_123, w_169_129, w_169_130, w_169_132, w_169_133, w_169_138, w_169_142, w_169_144, w_169_154, w_169_155, w_169_166, w_169_168, w_169_170, w_169_171, w_169_175, w_169_178, w_169_179, w_169_187, w_169_188, w_169_189, w_169_201, w_169_202, w_169_203, w_169_206, w_169_210, w_169_219, w_169_221, w_169_225, w_169_226, w_169_233, w_169_234, w_169_238, w_169_240, w_169_241, w_169_246, w_169_251, w_169_252, w_169_265, w_169_272, w_169_275, w_169_279, w_169_285, w_169_288, w_169_291, w_169_292, w_169_299, w_169_300, w_169_302, w_169_303, w_169_307, w_169_313, w_169_316, w_169_318, w_169_320, w_169_322, w_169_326, w_169_331, w_169_335, w_169_336, w_169_340, w_169_341, w_169_342, w_169_346, w_169_347, w_169_352, w_169_358, w_169_359, w_169_360, w_169_362, w_169_363, w_169_369, w_169_370, w_169_371, w_169_373, w_169_376, w_169_392, w_169_393, w_169_396, w_169_398, w_169_399, w_169_403, w_169_405, w_169_409, w_169_411, w_169_413, w_169_416, w_169_419, w_169_427, w_169_433, w_169_434, w_169_438, w_169_441, w_169_448, w_169_452, w_169_454, w_169_460, w_169_462, w_169_467, w_169_471, w_169_474, w_169_475, w_169_476, w_169_477, w_169_489, w_169_492, w_169_493, w_169_494, w_169_496, w_169_498, w_169_506, w_169_509, w_169_513, w_169_521, w_169_524, w_169_525, w_169_527, w_169_531, w_169_536, w_169_539, w_169_542, w_169_543, w_169_544, w_169_545, w_169_548, w_169_552, w_169_554, w_169_555, w_169_556, w_169_563, w_169_566, w_169_573, w_169_576, w_169_580, w_169_582, w_169_583, w_169_585, w_169_587, w_169_596, w_169_599, w_169_602, w_169_604, w_169_609, w_169_611, w_169_613, w_169_627, w_169_631, w_169_632, w_169_642, w_169_643, w_169_645, w_169_649, w_169_655, w_169_657, w_169_658, w_169_660, w_169_662, w_169_664, w_169_671, w_169_677, w_169_680, w_169_687, w_169_688, w_169_692, w_169_693, w_169_694, w_169_695, w_169_701, w_169_702, w_169_703, w_169_704, w_169_714, w_169_719, w_169_723, w_169_726, w_169_728, w_169_736, w_169_745, w_169_747, w_169_748, w_169_751, w_169_756, w_169_760, w_169_761, w_169_762, w_169_763, w_169_773, w_169_776, w_169_783, w_169_785, w_169_786, w_169_793, w_169_798, w_169_799, w_169_802, w_169_808, w_169_814, w_169_816, w_169_822, w_169_829, w_169_834, w_169_841, w_169_842, w_169_846, w_169_849, w_169_852, w_169_853, w_169_868, w_169_877, w_169_879, w_169_882, w_169_898, w_169_901, w_169_906, w_169_908, w_169_910, w_169_911, w_169_912, w_169_916, w_169_924, w_169_927, w_169_934, w_169_938, w_169_944, w_169_946, w_169_952, w_169_959, w_169_960, w_169_962, w_169_963, w_169_964, w_169_965, w_169_972, w_169_973, w_169_977, w_169_979, w_169_981, w_169_982, w_169_990, w_169_991, w_169_995, w_169_996, w_169_1005, w_169_1006, w_169_1007, w_169_1009, w_169_1010, w_169_1011, w_169_1013, w_169_1015, w_169_1016, w_169_1017, w_169_1026, w_169_1027, w_169_1030, w_169_1031, w_169_1032, w_169_1033, w_169_1037, w_169_1054, w_169_1056, w_169_1059, w_169_1062, w_169_1065, w_169_1066, w_169_1074, w_169_1091, w_169_1092, w_169_1094, w_169_1098, w_169_1101, w_169_1103, w_169_1109, w_169_1110, w_169_1112, w_169_1114, w_169_1121, w_169_1127, w_169_1130, w_169_1131, w_169_1134, w_169_1135, w_169_1137, w_169_1139, w_169_1143, w_169_1148, w_169_1149, w_169_1151, w_169_1156, w_169_1158, w_169_1162, w_169_1168, w_169_1169, w_169_1177, w_169_1178, w_169_1180, w_169_1181, w_169_1182, w_169_1185, w_169_1192, w_169_1193, w_169_1199, w_169_1206, w_169_1207, w_169_1209, w_169_1210, w_169_1222, w_169_1228, w_169_1234, w_169_1236, w_169_1238, w_169_1240, w_169_1242, w_169_1246, w_169_1249, w_169_1251, w_169_1252, w_169_1253, w_169_1254, w_169_1256, w_169_1258, w_169_1259, w_169_1260, w_169_1261, w_169_1269, w_169_1270, w_169_1273, w_169_1274, w_169_1276, w_169_1279, w_169_1281, w_169_1286, w_169_1290, w_169_1294, w_169_1295, w_169_1297, w_169_1299, w_169_1306, w_169_1311, w_169_1315, w_169_1316, w_169_1318, w_169_1321, w_169_1322, w_169_1325, w_169_1330, w_169_1331, w_169_1338, w_169_1339, w_169_1341, w_169_1351, w_169_1360, w_169_1363, w_169_1366, w_169_1367, w_169_1368, w_169_1377, w_169_1384, w_169_1389, w_169_1392, w_169_1393, w_169_1402, w_169_1403, w_169_1406, w_169_1410, w_169_1412, w_169_1413, w_169_1415, w_169_1416, w_169_1417, w_169_1423, w_169_1425, w_169_1426, w_169_1435, w_169_1436, w_169_1437, w_169_1438, w_169_1446, w_169_1451, w_169_1454, w_169_1455, w_169_1463, w_169_1465, w_169_1467, w_169_1468, w_169_1472, w_169_1474, w_169_1475, w_169_1478, w_169_1482, w_169_1483, w_169_1484, w_169_1485, w_169_1489, w_169_1491, w_169_1494, w_169_1501, w_169_1503, w_169_1505, w_169_1507, w_169_1510, w_169_1513, w_169_1514, w_169_1519, w_169_1524, w_169_1525, w_169_1529, w_169_1532, w_169_1539, w_169_1541, w_169_1549, w_169_1550, w_169_1551, w_169_1561, w_169_1562, w_169_1563, w_169_1568, w_169_1573, w_169_1576, w_169_1580, w_169_1582, w_169_1585, w_169_1588, w_169_1594, w_169_1603, w_169_1605, w_169_1616, w_169_1617, w_169_1618, w_169_1623, w_169_1635, w_169_1639, w_169_1646, w_169_1647, w_169_1657, w_169_1660, w_169_1662, w_169_1669, w_169_1670, w_169_1672, w_169_1675, w_169_1677, w_169_1679, w_169_1680, w_169_1681, w_169_1683, w_169_1691, w_169_1692, w_169_1699, w_169_1704, w_169_1705, w_169_1710, w_169_1712, w_169_1715, w_169_1716, w_169_1722, w_169_1723, w_169_1729, w_169_1734, w_169_1738, w_169_1744, w_169_1751, w_169_1756, w_169_1760, w_169_1763, w_169_1767, w_169_1768, w_169_1769, w_169_1770, w_169_1774, w_169_1779, w_169_1780, w_169_1788, w_169_1789, w_169_1790, w_169_1795, w_169_1797, w_169_1798, w_169_1809, w_169_1814, w_169_1817, w_169_1819, w_169_1828, w_169_1829, w_169_1832, w_169_1836, w_169_1838, w_169_1842, w_169_1843, w_169_1846, w_169_1848, w_169_1852, w_169_1853, w_169_1855, w_169_1859, w_169_1863, w_169_1868, w_169_1876, w_169_1877, w_169_1878, w_169_1893, w_169_1896, w_169_1898, w_169_1906, w_169_1907, w_169_1908, w_169_1914, w_169_1917, w_169_1918, w_169_1919, w_169_1920, w_169_1921, w_169_1925, w_169_1926, w_169_1929, w_169_1931, w_169_1932, w_169_1933, w_169_1935, w_169_1939, w_169_1941, w_169_1945, w_169_1949, w_169_1952, w_169_1953, w_169_1954, w_169_1958, w_169_1961, w_169_1963, w_169_1966, w_169_1967, w_169_1972, w_169_1977, w_169_1987, w_169_1991, w_169_1993, w_169_2005, w_169_2011, w_169_2015, w_169_2020, w_169_2026, w_169_2028, w_169_2029, w_169_2032, w_169_2033, w_169_2034, w_169_2035, w_169_2040, w_169_2041, w_169_2046, w_169_2051, w_169_2053, w_169_2054, w_169_2056, w_169_2059, w_169_2064, w_169_2070, w_169_2071, w_169_2073, w_169_2075, w_169_2077, w_169_2078, w_169_2080, w_169_2081, w_169_2082, w_169_2083, w_169_2085, w_169_2087, w_169_2089, w_169_2091, w_169_2094, w_169_2098, w_169_2099, w_169_2100, w_169_2107, w_169_2109, w_169_2111, w_169_2115, w_169_2117, w_169_2123, w_169_2124, w_169_2129, w_169_2131, w_169_2141, w_169_2143, w_169_2148, w_169_2149, w_169_2150, w_169_2151, w_169_2153, w_169_2155, w_169_2157, w_169_2158, w_169_2160, w_169_2166, w_169_2167, w_169_2172, w_169_2175, w_169_2176, w_169_2182, w_169_2189, w_169_2191, w_169_2192, w_169_2197, w_169_2212, w_169_2218, w_169_2220, w_169_2232, w_169_2233, w_169_2236, w_169_2237, w_169_2240, w_169_2247, w_169_2250, w_169_2253, w_169_2254, w_169_2257, w_169_2264, w_169_2278, w_169_2279, w_169_2287, w_169_2300, w_169_2302, w_169_2303, w_169_2313, w_169_2315, w_169_2316, w_169_2322, w_169_2329, w_169_2344, w_169_2346, w_169_2348, w_169_2351, w_169_2357, w_169_2372, w_169_2376, w_169_2380, w_169_2383, w_169_2389, w_169_2392, w_169_2396, w_169_2400, w_169_2407, w_169_2426, w_169_2428, w_169_2451, w_169_2461, w_169_2462, w_169_2464, w_169_2467, w_169_2469, w_169_2477, w_169_2488, w_169_2494, w_169_2501, w_169_2502, w_169_2506, w_169_2508, w_169_2512, w_169_2522, w_169_2531, w_169_2543, w_169_2557, w_169_2561, w_169_2572, w_169_2576, w_169_2581, w_169_2583, w_169_2595, w_169_2606, w_169_2607, w_169_2621, w_169_2624, w_169_2631, w_169_2632, w_169_2633, w_169_2636, w_169_2643, w_169_2663, w_169_2669, w_169_2671, w_169_2672, w_169_2687, w_169_2691, w_169_2707, w_169_2712, w_169_2715, w_169_2717, w_169_2723, w_169_2750, w_169_2753, w_169_2758, w_169_2762, w_169_2770, w_169_2796, w_169_2798;
  wire w_170_000, w_170_001, w_170_003, w_170_004, w_170_006, w_170_007, w_170_008, w_170_009, w_170_010, w_170_013, w_170_014, w_170_015, w_170_017, w_170_018, w_170_019, w_170_020, w_170_021, w_170_022, w_170_023, w_170_024, w_170_025, w_170_027, w_170_028, w_170_029, w_170_030, w_170_031, w_170_033, w_170_036, w_170_037, w_170_038, w_170_039, w_170_040, w_170_043, w_170_044, w_170_045, w_170_046, w_170_047, w_170_048, w_170_049, w_170_050, w_170_051, w_170_052, w_170_053, w_170_054, w_170_055, w_170_056, w_170_057, w_170_058, w_170_059, w_170_060, w_170_062, w_170_065, w_170_066, w_170_067, w_170_069, w_170_070, w_170_071, w_170_072, w_170_073, w_170_074, w_170_075, w_170_076, w_170_077, w_170_078, w_170_079, w_170_080, w_170_083, w_170_084, w_170_085, w_170_086, w_170_087, w_170_088, w_170_089, w_170_090, w_170_091, w_170_093, w_170_094, w_170_095, w_170_096, w_170_098, w_170_099, w_170_100, w_170_102, w_170_103, w_170_104, w_170_105, w_170_106, w_170_107, w_170_108, w_170_109, w_170_110, w_170_111, w_170_112, w_170_113, w_170_115, w_170_116, w_170_117, w_170_118, w_170_119, w_170_125, w_170_126, w_170_127, w_170_128, w_170_129, w_170_131, w_170_132, w_170_133, w_170_134, w_170_136, w_170_137, w_170_138, w_170_139, w_170_140, w_170_141, w_170_142, w_170_143, w_170_144, w_170_145, w_170_146, w_170_147, w_170_149, w_170_150, w_170_151, w_170_152, w_170_153, w_170_155, w_170_157, w_170_158, w_170_159, w_170_160, w_170_161, w_170_162, w_170_163, w_170_164, w_170_165, w_170_167, w_170_168, w_170_169, w_170_170, w_170_172, w_170_173, w_170_174, w_170_175, w_170_176, w_170_177, w_170_178, w_170_179, w_170_180, w_170_181, w_170_184, w_170_188, w_170_189, w_170_190, w_170_191, w_170_192, w_170_194, w_170_195, w_170_197, w_170_198, w_170_200, w_170_201, w_170_202, w_170_203, w_170_204, w_170_205, w_170_206, w_170_208, w_170_209, w_170_210, w_170_212, w_170_213, w_170_214, w_170_215, w_170_216, w_170_218, w_170_219, w_170_220, w_170_221, w_170_222, w_170_223, w_170_224, w_170_225, w_170_226, w_170_227, w_170_228, w_170_230, w_170_231, w_170_232, w_170_233, w_170_234, w_170_235, w_170_236, w_170_239, w_170_240, w_170_241, w_170_242, w_170_243, w_170_244, w_170_245, w_170_247, w_170_248, w_170_249, w_170_251, w_170_252, w_170_253, w_170_254, w_170_255, w_170_256, w_170_257, w_170_258, w_170_259, w_170_260, w_170_263, w_170_264, w_170_265, w_170_266, w_170_267, w_170_269, w_170_271, w_170_272, w_170_273, w_170_276, w_170_277, w_170_279, w_170_280, w_170_281, w_170_282, w_170_283, w_170_284, w_170_286, w_170_287, w_170_288, w_170_289, w_170_290, w_170_293, w_170_294, w_170_296, w_170_299, w_170_301, w_170_302, w_170_303, w_170_304, w_170_305, w_170_307, w_170_308, w_170_309, w_170_310, w_170_311, w_170_312, w_170_313, w_170_314, w_170_315, w_170_316, w_170_317, w_170_318, w_170_319, w_170_320, w_170_321, w_170_322, w_170_323, w_170_324, w_170_325, w_170_327, w_170_330, w_170_331, w_170_332, w_170_334, w_170_335, w_170_337, w_170_338, w_170_339, w_170_340, w_170_341, w_170_342, w_170_343, w_170_344, w_170_345, w_170_346, w_170_347, w_170_348, w_170_349, w_170_351, w_170_352, w_170_353, w_170_354, w_170_355, w_170_356, w_170_357, w_170_358, w_170_360, w_170_361, w_170_362, w_170_363, w_170_364, w_170_365, w_170_367, w_170_368, w_170_370, w_170_373, w_170_374, w_170_375, w_170_376, w_170_377, w_170_381, w_170_382, w_170_383, w_170_384, w_170_385, w_170_386, w_170_387, w_170_388, w_170_389, w_170_390, w_170_391, w_170_394, w_170_395, w_170_396, w_170_397, w_170_398, w_170_399, w_170_400, w_170_403, w_170_404, w_170_407, w_170_408, w_170_409, w_170_410, w_170_412, w_170_413, w_170_414, w_170_415, w_170_416, w_170_418, w_170_419, w_170_420, w_170_421, w_170_422, w_170_423, w_170_424, w_170_425, w_170_426, w_170_428, w_170_430, w_170_432, w_170_434, w_170_435, w_170_436, w_170_438, w_170_439, w_170_441, w_170_442, w_170_443, w_170_445, w_170_446, w_170_447, w_170_449, w_170_451, w_170_453, w_170_454, w_170_455, w_170_457, w_170_458, w_170_459, w_170_463, w_170_464, w_170_465, w_170_466, w_170_468, w_170_469, w_170_473, w_170_474, w_170_475, w_170_476, w_170_477, w_170_478, w_170_481, w_170_482, w_170_483, w_170_484, w_170_488, w_170_489, w_170_490, w_170_494, w_170_495, w_170_497, w_170_498, w_170_499, w_170_500, w_170_501, w_170_502, w_170_503, w_170_504, w_170_505, w_170_507, w_170_510, w_170_511, w_170_512, w_170_513, w_170_514, w_170_515, w_170_517, w_170_519, w_170_520, w_170_521, w_170_522, w_170_523, w_170_524, w_170_525, w_170_526, w_170_527, w_170_529, w_170_531, w_170_533, w_170_534, w_170_535, w_170_536, w_170_538, w_170_539, w_170_540, w_170_541, w_170_542, w_170_543, w_170_544, w_170_546, w_170_548, w_170_549, w_170_550, w_170_552, w_170_554, w_170_555, w_170_557, w_170_558, w_170_559, w_170_563, w_170_565, w_170_567, w_170_570, w_170_571, w_170_572, w_170_573, w_170_574, w_170_576, w_170_577, w_170_578, w_170_581, w_170_582, w_170_583, w_170_585, w_170_587, w_170_588, w_170_589, w_170_593, w_170_594, w_170_595, w_170_596, w_170_597, w_170_598, w_170_600;
  wire w_171_003, w_171_006, w_171_008, w_171_012, w_171_013, w_171_014, w_171_016, w_171_018, w_171_024, w_171_025, w_171_028, w_171_034, w_171_035, w_171_037, w_171_045, w_171_047, w_171_048, w_171_052, w_171_054, w_171_055, w_171_056, w_171_061, w_171_062, w_171_065, w_171_066, w_171_068, w_171_071, w_171_072, w_171_080, w_171_084, w_171_091, w_171_092, w_171_097, w_171_108, w_171_109, w_171_110, w_171_117, w_171_118, w_171_123, w_171_124, w_171_128, w_171_129, w_171_134, w_171_138, w_171_139, w_171_140, w_171_148, w_171_154, w_171_156, w_171_158, w_171_161, w_171_162, w_171_166, w_171_168, w_171_169, w_171_171, w_171_174, w_171_181, w_171_186, w_171_190, w_171_194, w_171_195, w_171_197, w_171_198, w_171_203, w_171_206, w_171_216, w_171_218, w_171_230, w_171_234, w_171_238, w_171_248, w_171_249, w_171_258, w_171_259, w_171_261, w_171_262, w_171_266, w_171_267, w_171_270, w_171_273, w_171_276, w_171_281, w_171_283, w_171_284, w_171_289, w_171_290, w_171_295, w_171_302, w_171_309, w_171_319, w_171_325, w_171_327, w_171_332, w_171_333, w_171_335, w_171_337, w_171_339, w_171_341, w_171_347, w_171_349, w_171_350, w_171_352, w_171_353, w_171_354, w_171_367, w_171_368, w_171_370, w_171_372, w_171_373, w_171_378, w_171_379, w_171_383, w_171_384, w_171_387, w_171_388, w_171_389, w_171_390, w_171_392, w_171_393, w_171_397, w_171_401, w_171_406, w_171_410, w_171_415, w_171_422, w_171_423, w_171_426, w_171_428, w_171_431, w_171_438, w_171_443, w_171_444, w_171_445, w_171_450, w_171_453, w_171_454, w_171_461, w_171_462, w_171_464, w_171_466, w_171_471, w_171_472, w_171_475, w_171_477, w_171_484, w_171_491, w_171_495, w_171_498, w_171_499, w_171_504, w_171_505, w_171_506, w_171_512, w_171_515, w_171_516, w_171_521, w_171_530, w_171_534, w_171_535, w_171_536, w_171_542, w_171_547, w_171_552, w_171_555, w_171_566, w_171_567, w_171_569, w_171_571, w_171_573, w_171_574, w_171_581, w_171_582, w_171_588, w_171_590, w_171_594, w_171_601, w_171_605, w_171_619, w_171_620, w_171_623, w_171_628, w_171_629, w_171_635, w_171_636, w_171_637, w_171_639, w_171_640, w_171_643, w_171_650, w_171_653, w_171_655, w_171_662, w_171_663, w_171_665, w_171_671, w_171_673, w_171_676, w_171_679, w_171_681, w_171_682, w_171_687, w_171_690, w_171_691, w_171_699, w_171_704, w_171_709, w_171_714, w_171_716, w_171_717, w_171_722, w_171_723, w_171_724, w_171_728, w_171_730, w_171_734, w_171_735, w_171_737, w_171_741, w_171_743, w_171_748, w_171_749, w_171_751, w_171_753, w_171_758, w_171_759, w_171_763, w_171_768, w_171_770, w_171_771, w_171_775, w_171_777, w_171_779, w_171_782, w_171_784, w_171_786, w_171_788, w_171_793, w_171_797, w_171_804, w_171_809, w_171_812, w_171_813, w_171_816, w_171_820, w_171_825, w_171_829, w_171_832, w_171_835, w_171_846, w_171_850, w_171_851, w_171_853, w_171_855, w_171_856, w_171_863, w_171_864, w_171_866, w_171_869, w_171_882, w_171_888, w_171_898, w_171_902, w_171_904, w_171_906, w_171_912, w_171_914, w_171_920, w_171_921, w_171_922, w_171_926, w_171_928, w_171_929, w_171_931, w_171_934, w_171_938, w_171_939, w_171_944, w_171_947, w_171_950, w_171_951, w_171_952, w_171_955, w_171_960, w_171_964, w_171_969, w_171_975, w_171_976, w_171_977, w_171_979, w_171_984, w_171_989, w_171_991, w_171_992, w_171_994, w_171_997, w_171_1007, w_171_1017, w_171_1024, w_171_1030, w_171_1031, w_171_1033, w_171_1036, w_171_1037, w_171_1041, w_171_1042, w_171_1046, w_171_1047, w_171_1053, w_171_1072, w_171_1073, w_171_1080, w_171_1082, w_171_1084, w_171_1085, w_171_1086, w_171_1091, w_171_1095, w_171_1098, w_171_1099, w_171_1112, w_171_1113, w_171_1131, w_171_1132, w_171_1137, w_171_1144, w_171_1146, w_171_1150, w_171_1154, w_171_1159, w_171_1161, w_171_1166, w_171_1183, w_171_1185, w_171_1189, w_171_1195, w_171_1199, w_171_1214, w_171_1217, w_171_1218, w_171_1220, w_171_1225, w_171_1232, w_171_1239, w_171_1241, w_171_1245, w_171_1250, w_171_1253, w_171_1258, w_171_1266, w_171_1268, w_171_1271, w_171_1275, w_171_1287, w_171_1302, w_171_1306, w_171_1313, w_171_1317, w_171_1319, w_171_1332, w_171_1335, w_171_1337, w_171_1344, w_171_1347, w_171_1352, w_171_1360, w_171_1362, w_171_1369, w_171_1374, w_171_1384, w_171_1393, w_171_1402, w_171_1403, w_171_1405, w_171_1410, w_171_1412, w_171_1422, w_171_1430, w_171_1431, w_171_1434, w_171_1443, w_171_1458, w_171_1485, w_171_1486, w_171_1496, w_171_1499, w_171_1508, w_171_1532, w_171_1538, w_171_1541, w_171_1556, w_171_1572, w_171_1573, w_171_1578, w_171_1584, w_171_1589, w_171_1610, w_171_1617, w_171_1618, w_171_1630, w_171_1637, w_171_1641, w_171_1643, w_171_1656, w_171_1658, w_171_1671, w_171_1677, w_171_1680, w_171_1681, w_171_1687, w_171_1688, w_171_1690, w_171_1691, w_171_1692, w_171_1693, w_171_1695, w_171_1696, w_171_1722, w_171_1731, w_171_1734, w_171_1740, w_171_1745, w_171_1762, w_171_1783, w_171_1790, w_171_1792, w_171_1793, w_171_1795, w_171_1796, w_171_1798, w_171_1804, w_171_1810, w_171_1813, w_171_1820, w_171_1829, w_171_1832, w_171_1849, w_171_1857, w_171_1863, w_171_1874, w_171_1890, w_171_1893, w_171_1914, w_171_1931, w_171_1938, w_171_1941, w_171_1945, w_171_1947, w_171_1954, w_171_1963, w_171_1975, w_171_1987, w_171_2006, w_171_2007, w_171_2022, w_171_2023, w_171_2026, w_171_2034, w_171_2035, w_171_2043, w_171_2056, w_171_2072, w_171_2082, w_171_2092, w_171_2093, w_171_2098, w_171_2113, w_171_2136, w_171_2137, w_171_2143, w_171_2144, w_171_2153, w_171_2163, w_171_2174, w_171_2180, w_171_2189, w_171_2196, w_171_2213, w_171_2220, w_171_2227, w_171_2232, w_171_2236, w_171_2239, w_171_2242, w_171_2253, w_171_2256, w_171_2260, w_171_2269, w_171_2270, w_171_2273, w_171_2277, w_171_2283, w_171_2290, w_171_2298, w_171_2308, w_171_2316, w_171_2331, w_171_2332, w_171_2335, w_171_2343, w_171_2348, w_171_2352, w_171_2354, w_171_2361, w_171_2378, w_171_2399, w_171_2432, w_171_2434, w_171_2445, w_171_2450, w_171_2451, w_171_2461, w_171_2462, w_171_2463, w_171_2464, w_171_2468, w_171_2474, w_171_2487, w_171_2488, w_171_2511, w_171_2513, w_171_2524, w_171_2527, w_171_2541, w_171_2557, w_171_2560, w_171_2562, w_171_2575, w_171_2590, w_171_2592, w_171_2595, w_171_2607, w_171_2609, w_171_2610, w_171_2626, w_171_2628, w_171_2631, w_171_2648, w_171_2649, w_171_2679, w_171_2687, w_171_2688, w_171_2699, w_171_2702, w_171_2706, w_171_2721, w_171_2733, w_171_2736, w_171_2739, w_171_2740, w_171_2743, w_171_2747, w_171_2751, w_171_2753, w_171_2772, w_171_2787, w_171_2794, w_171_2795, w_171_2796, w_171_2818, w_171_2828, w_171_2830, w_171_2834, w_171_2848, w_171_2853, w_171_2875, w_171_2876, w_171_2885, w_171_2892, w_171_2893, w_171_2895, w_171_2897, w_171_2901, w_171_2907, w_171_2913, w_171_2914, w_171_2916, w_171_2918, w_171_2922, w_171_2927, w_171_2932, w_171_2934, w_171_2945, w_171_2949, w_171_2952, w_171_2962, w_171_2975, w_171_2982, w_171_2996, w_171_2997, w_171_3003, w_171_3036, w_171_3038, w_171_3051, w_171_3052, w_171_3059, w_171_3070, w_171_3077, w_171_3085, w_171_3087, w_171_3093, w_171_3104, w_171_3108, w_171_3111, w_171_3116, w_171_3120, w_171_3130, w_171_3132, w_171_3145, w_171_3148, w_171_3149, w_171_3150, w_171_3167, w_171_3177, w_171_3180, w_171_3184, w_171_3188, w_171_3189, w_171_3190, w_171_3191, w_171_3194, w_171_3195, w_171_3201, w_171_3207, w_171_3217, w_171_3226, w_171_3238, w_171_3239, w_171_3249, w_171_3256, w_171_3263, w_171_3282, w_171_3288, w_171_3293, w_171_3296, w_171_3305, w_171_3308, w_171_3321, w_171_3328, w_171_3342, w_171_3351, w_171_3353, w_171_3355, w_171_3359, w_171_3361, w_171_3362, w_171_3367, w_171_3369, w_171_3371, w_171_3373, w_171_3376, w_171_3379, w_171_3381, w_171_3398, w_171_3402, w_171_3404, w_171_3409, w_171_3424, w_171_3427, w_171_3432, w_171_3440, w_171_3454, w_171_3459, w_171_3496, w_171_3508, w_171_3517, w_171_3518, w_171_3524, w_171_3531, w_171_3536, w_171_3540, w_171_3550, w_171_3566, w_171_3567, w_171_3568, w_171_3569, w_171_3570, w_171_3582, w_171_3583, w_171_3585, w_171_3587, w_171_3595, w_171_3599, w_171_3605, w_171_3610, w_171_3613, w_171_3630, w_171_3640, w_171_3645, w_171_3649, w_171_3650, w_171_3654, w_171_3667, w_171_3669, w_171_3675, w_171_3683, w_171_3689, w_171_3695, w_171_3696, w_171_3699, w_171_3701, w_171_3704, w_171_3710, w_171_3725, w_171_3742, w_171_3751, w_171_3756, w_171_3768, w_171_3777, w_171_3790, w_171_3794, w_171_3795, w_171_3800, w_171_3802, w_171_3813, w_171_3827, w_171_3832, w_171_3844, w_171_3855, w_171_3861, w_171_3862, w_171_3863, w_171_3865, w_171_3867, w_171_3868, w_171_3869, w_171_3870, w_171_3872;
  wire w_172_002, w_172_004, w_172_010, w_172_015, w_172_024, w_172_025, w_172_028, w_172_035, w_172_037, w_172_038, w_172_040, w_172_042, w_172_043, w_172_044, w_172_047, w_172_055, w_172_058, w_172_060, w_172_062, w_172_064, w_172_066, w_172_068, w_172_069, w_172_070, w_172_074, w_172_076, w_172_083, w_172_086, w_172_093, w_172_096, w_172_098, w_172_099, w_172_102, w_172_103, w_172_107, w_172_123, w_172_126, w_172_127, w_172_130, w_172_131, w_172_132, w_172_133, w_172_140, w_172_143, w_172_150, w_172_152, w_172_154, w_172_155, w_172_156, w_172_163, w_172_168, w_172_171, w_172_172, w_172_178, w_172_179, w_172_185, w_172_198, w_172_199, w_172_200, w_172_205, w_172_206, w_172_207, w_172_209, w_172_211, w_172_219, w_172_225, w_172_227, w_172_229, w_172_233, w_172_237, w_172_239, w_172_245, w_172_246, w_172_255, w_172_257, w_172_263, w_172_264, w_172_271, w_172_284, w_172_287, w_172_289, w_172_290, w_172_293, w_172_295, w_172_299, w_172_301, w_172_302, w_172_308, w_172_313, w_172_317, w_172_319, w_172_321, w_172_322, w_172_325, w_172_327, w_172_328, w_172_334, w_172_335, w_172_336, w_172_338, w_172_339, w_172_340, w_172_341, w_172_343, w_172_345, w_172_349, w_172_350, w_172_357, w_172_360, w_172_364, w_172_365, w_172_366, w_172_372, w_172_374, w_172_377, w_172_379, w_172_384, w_172_385, w_172_391, w_172_399, w_172_400, w_172_407, w_172_408, w_172_412, w_172_413, w_172_428, w_172_432, w_172_452, w_172_453, w_172_458, w_172_459, w_172_460, w_172_466, w_172_467, w_172_468, w_172_473, w_172_475, w_172_478, w_172_483, w_172_486, w_172_490, w_172_492, w_172_498, w_172_503, w_172_505, w_172_522, w_172_524, w_172_525, w_172_526, w_172_531, w_172_532, w_172_533, w_172_538, w_172_544, w_172_549, w_172_556, w_172_559, w_172_562, w_172_567, w_172_577, w_172_584, w_172_587, w_172_589, w_172_591, w_172_600, w_172_601, w_172_608, w_172_609, w_172_612, w_172_614, w_172_620, w_172_628, w_172_642, w_172_646, w_172_649, w_172_664, w_172_666, w_172_671, w_172_676, w_172_678, w_172_679, w_172_680, w_172_694, w_172_700, w_172_708, w_172_714, w_172_717, w_172_725, w_172_735, w_172_737, w_172_748, w_172_753, w_172_760, w_172_762, w_172_765, w_172_766, w_172_774, w_172_785, w_172_792, w_172_818, w_172_827, w_172_833, w_172_843, w_172_846, w_172_851, w_172_865, w_172_872, w_172_882, w_172_884, w_172_891, w_172_896, w_172_910, w_172_916, w_172_927, w_172_932, w_172_933, w_172_935, w_172_939, w_172_941, w_172_942, w_172_945, w_172_971, w_172_978, w_172_979, w_172_990, w_172_1013, w_172_1016, w_172_1017, w_172_1022, w_172_1027, w_172_1034, w_172_1043, w_172_1044, w_172_1045, w_172_1053, w_172_1054, w_172_1056, w_172_1059, w_172_1060, w_172_1065, w_172_1066, w_172_1072, w_172_1083, w_172_1085, w_172_1095, w_172_1099, w_172_1106, w_172_1112, w_172_1117, w_172_1119, w_172_1124, w_172_1127, w_172_1140, w_172_1143, w_172_1144, w_172_1151, w_172_1155, w_172_1164, w_172_1175, w_172_1176, w_172_1178, w_172_1184, w_172_1198, w_172_1233, w_172_1237, w_172_1244, w_172_1249, w_172_1252, w_172_1253, w_172_1264, w_172_1280, w_172_1284, w_172_1287, w_172_1291, w_172_1294, w_172_1306, w_172_1315, w_172_1321, w_172_1323, w_172_1325, w_172_1336, w_172_1343, w_172_1345, w_172_1351, w_172_1352, w_172_1355, w_172_1356, w_172_1360, w_172_1364, w_172_1379, w_172_1381, w_172_1385, w_172_1390, w_172_1399, w_172_1400, w_172_1413, w_172_1421, w_172_1423, w_172_1429, w_172_1430, w_172_1436, w_172_1441, w_172_1463, w_172_1466, w_172_1469, w_172_1475, w_172_1481, w_172_1494, w_172_1505, w_172_1508, w_172_1510, w_172_1512, w_172_1523, w_172_1524, w_172_1533, w_172_1538, w_172_1545, w_172_1568, w_172_1571, w_172_1574, w_172_1578, w_172_1583, w_172_1594, w_172_1596, w_172_1600, w_172_1617, w_172_1623, w_172_1633, w_172_1639, w_172_1645, w_172_1646, w_172_1666, w_172_1670, w_172_1680, w_172_1684, w_172_1694, w_172_1695, w_172_1709, w_172_1722, w_172_1727, w_172_1734, w_172_1737, w_172_1739, w_172_1744, w_172_1749, w_172_1774, w_172_1778, w_172_1794, w_172_1797, w_172_1815, w_172_1817, w_172_1826, w_172_1840, w_172_1843, w_172_1850, w_172_1856, w_172_1862, w_172_1864, w_172_1871, w_172_1880, w_172_1881, w_172_1882, w_172_1884, w_172_1894, w_172_1895, w_172_1907, w_172_1912, w_172_1914, w_172_1915, w_172_1922, w_172_1933, w_172_1948, w_172_1950, w_172_1953, w_172_1956, w_172_1957, w_172_1965, w_172_1967, w_172_1968, w_172_1973, w_172_1976, w_172_1999, w_172_2004, w_172_2011, w_172_2018, w_172_2037, w_172_2038, w_172_2040, w_172_2046, w_172_2048, w_172_2049, w_172_2053, w_172_2054, w_172_2056, w_172_2080, w_172_2090, w_172_2091, w_172_2094, w_172_2104, w_172_2122, w_172_2138, w_172_2142, w_172_2154, w_172_2155, w_172_2172, w_172_2181, w_172_2188, w_172_2192, w_172_2193, w_172_2202, w_172_2203, w_172_2223, w_172_2224, w_172_2242, w_172_2249, w_172_2256, w_172_2267, w_172_2270, w_172_2273, w_172_2276, w_172_2279, w_172_2282, w_172_2284, w_172_2289, w_172_2293, w_172_2294, w_172_2299, w_172_2306, w_172_2312, w_172_2326, w_172_2329, w_172_2335, w_172_2338, w_172_2340, w_172_2342, w_172_2343, w_172_2352, w_172_2353, w_172_2354, w_172_2356, w_172_2366, w_172_2368, w_172_2370, w_172_2380, w_172_2383, w_172_2393, w_172_2397, w_172_2411, w_172_2421, w_172_2441, w_172_2444, w_172_2459, w_172_2468, w_172_2475, w_172_2482, w_172_2485, w_172_2486, w_172_2494, w_172_2496, w_172_2501, w_172_2503, w_172_2512, w_172_2528, w_172_2545, w_172_2552, w_172_2553, w_172_2562, w_172_2571, w_172_2576, w_172_2581, w_172_2584, w_172_2597, w_172_2599, w_172_2601, w_172_2603, w_172_2605, w_172_2606, w_172_2607, w_172_2610, w_172_2619, w_172_2628, w_172_2648, w_172_2672, w_172_2675, w_172_2678, w_172_2682, w_172_2699, w_172_2705, w_172_2722, w_172_2730, w_172_2731, w_172_2737, w_172_2744, w_172_2745, w_172_2752, w_172_2753, w_172_2757, w_172_2763, w_172_2771, w_172_2772, w_172_2787, w_172_2793, w_172_2798, w_172_2806, w_172_2816, w_172_2822, w_172_2837, w_172_2839, w_172_2841, w_172_2842, w_172_2852, w_172_2857, w_172_2858, w_172_2865, w_172_2873, w_172_2921, w_172_2924, w_172_2925, w_172_2930, w_172_2932, w_172_2935, w_172_2937, w_172_2944, w_172_2947, w_172_2948, w_172_2950, w_172_2952, w_172_2954, w_172_2956, w_172_2963, w_172_2973, w_172_2975, w_172_2977, w_172_2996, w_172_2997, w_172_2999, w_172_3032, w_172_3044, w_172_3049, w_172_3080, w_172_3090, w_172_3095, w_172_3096, w_172_3113, w_172_3118, w_172_3126, w_172_3136, w_172_3142, w_172_3146, w_172_3175, w_172_3187, w_172_3188, w_172_3201, w_172_3211, w_172_3215, w_172_3226, w_172_3236, w_172_3238, w_172_3243, w_172_3248, w_172_3249, w_172_3256, w_172_3260, w_172_3272, w_172_3280, w_172_3282, w_172_3283, w_172_3299, w_172_3309, w_172_3318, w_172_3320, w_172_3335, w_172_3342, w_172_3345, w_172_3368, w_172_3371, w_172_3372, w_172_3374, w_172_3377, w_172_3406, w_172_3410, w_172_3425, w_172_3426, w_172_3430, w_172_3431, w_172_3434, w_172_3437, w_172_3438, w_172_3458, w_172_3459, w_172_3460, w_172_3466, w_172_3467, w_172_3468, w_172_3474, w_172_3480, w_172_3485, w_172_3486, w_172_3497, w_172_3501, w_172_3502, w_172_3507, w_172_3511, w_172_3520, w_172_3524, w_172_3527, w_172_3530, w_172_3537, w_172_3538, w_172_3539, w_172_3541, w_172_3543, w_172_3547, w_172_3552, w_172_3565, w_172_3571, w_172_3572, w_172_3586, w_172_3587, w_172_3590, w_172_3602, w_172_3617, w_172_3619, w_172_3625, w_172_3633, w_172_3636, w_172_3646, w_172_3654, w_172_3667, w_172_3675, w_172_3679, w_172_3681, w_172_3688, w_172_3693, w_172_3700, w_172_3713, w_172_3725, w_172_3756, w_172_3762, w_172_3766, w_172_3771, w_172_3775, w_172_3782, w_172_3803, w_172_3805, w_172_3816, w_172_3820, w_172_3821, w_172_3825, w_172_3837, w_172_3838, w_172_3839, w_172_3851, w_172_3860, w_172_3862, w_172_3880, w_172_3885, w_172_3891, w_172_3895, w_172_3896, w_172_3898, w_172_3906, w_172_3909, w_172_3912, w_172_3914, w_172_3915, w_172_3922, w_172_3934, w_172_3936, w_172_3946, w_172_3961, w_172_3971, w_172_3996, w_172_3999, w_172_4008, w_172_4009, w_172_4016, w_172_4024, w_172_4032, w_172_4035, w_172_4043, w_172_4045, w_172_4054, w_172_4055, w_172_4062, w_172_4067, w_172_4070, w_172_4078, w_172_4079, w_172_4088, w_172_4094, w_172_4095, w_172_4102, w_172_4103, w_172_4106, w_172_4114, w_172_4116, w_172_4124, w_172_4127, w_172_4140, w_172_4142, w_172_4148, w_172_4164, w_172_4168, w_172_4171, w_172_4173, w_172_4174, w_172_4195, w_172_4201, w_172_4207, w_172_4208, w_172_4209, w_172_4221, w_172_4225, w_172_4227, w_172_4230, w_172_4237, w_172_4241, w_172_4251, w_172_4258, w_172_4261, w_172_4262, w_172_4263, w_172_4266, w_172_4282, w_172_4286, w_172_4291, w_172_4296, w_172_4301, w_172_4302, w_172_4309, w_172_4312, w_172_4313, w_172_4315, w_172_4329, w_172_4344, w_172_4345, w_172_4348, w_172_4350, w_172_4351;
  wire w_173_000, w_173_003, w_173_005, w_173_009, w_173_013, w_173_014, w_173_017, w_173_019, w_173_023, w_173_025, w_173_027, w_173_031, w_173_033, w_173_035, w_173_036, w_173_045, w_173_056, w_173_062, w_173_066, w_173_069, w_173_072, w_173_074, w_173_075, w_173_076, w_173_083, w_173_084, w_173_096, w_173_097, w_173_099, w_173_104, w_173_108, w_173_112, w_173_116, w_173_122, w_173_124, w_173_125, w_173_126, w_173_127, w_173_129, w_173_130, w_173_131, w_173_140, w_173_144, w_173_149, w_173_152, w_173_159, w_173_161, w_173_168, w_173_170, w_173_171, w_173_173, w_173_176, w_173_179, w_173_181, w_173_185, w_173_186, w_173_192, w_173_195, w_173_196, w_173_199, w_173_203, w_173_205, w_173_214, w_173_217, w_173_219, w_173_221, w_173_223, w_173_235, w_173_237, w_173_240, w_173_246, w_173_253, w_173_257, w_173_260, w_173_262, w_173_263, w_173_265, w_173_273, w_173_275, w_173_276, w_173_282, w_173_291, w_173_303, w_173_305, w_173_316, w_173_320, w_173_328, w_173_336, w_173_341, w_173_346, w_173_348, w_173_355, w_173_356, w_173_360, w_173_363, w_173_373, w_173_380, w_173_381, w_173_383, w_173_384, w_173_386, w_173_387, w_173_395, w_173_398, w_173_401, w_173_403, w_173_405, w_173_408, w_173_409, w_173_411, w_173_415, w_173_420, w_173_424, w_173_425, w_173_438, w_173_447, w_173_450, w_173_452, w_173_455, w_173_456, w_173_459, w_173_461, w_173_463, w_173_465, w_173_470, w_173_472, w_173_474, w_173_482, w_173_484, w_173_485, w_173_486, w_173_490, w_173_491, w_173_493, w_173_498, w_173_500, w_173_501, w_173_502, w_173_505, w_173_509, w_173_512, w_173_519, w_173_520, w_173_521, w_173_527, w_173_538, w_173_546, w_173_548, w_173_549, w_173_554, w_173_558, w_173_562, w_173_563, w_173_567, w_173_568, w_173_575, w_173_577, w_173_585, w_173_602, w_173_604, w_173_606, w_173_615, w_173_626, w_173_627, w_173_628, w_173_632, w_173_637, w_173_638, w_173_641, w_173_643, w_173_645, w_173_648, w_173_651, w_173_653, w_173_654, w_173_656, w_173_659, w_173_662, w_173_664, w_173_669, w_173_672, w_173_675, w_173_678, w_173_687, w_173_689, w_173_690, w_173_691, w_173_692, w_173_694, w_173_696, w_173_698, w_173_700, w_173_701, w_173_706, w_173_710, w_173_713, w_173_715, w_173_716, w_173_717, w_173_720, w_173_721, w_173_732, w_173_737, w_173_740, w_173_746, w_173_749, w_173_760, w_173_763, w_173_766, w_173_769, w_173_770, w_173_772, w_173_774, w_173_781, w_173_784, w_173_786, w_173_793, w_173_798, w_173_805, w_173_806, w_173_810, w_173_813, w_173_815, w_173_819, w_173_822, w_173_826, w_173_828, w_173_833, w_173_835, w_173_836, w_173_843, w_173_844, w_173_845, w_173_848, w_173_849, w_173_855, w_173_856, w_173_862, w_173_870, w_173_880, w_173_883, w_173_884, w_173_886, w_173_888, w_173_909, w_173_912, w_173_913, w_173_917, w_173_918, w_173_919, w_173_920, w_173_922, w_173_924, w_173_925, w_173_926, w_173_927, w_173_931, w_173_932, w_173_936, w_173_937, w_173_947, w_173_951, w_173_957, w_173_958, w_173_961, w_173_963, w_173_964, w_173_966, w_173_973, w_173_974, w_173_976, w_173_979, w_173_981, w_173_985, w_173_988, w_173_993, w_173_995, w_173_1002, w_173_1005, w_173_1010, w_173_1016, w_173_1020, w_173_1027, w_173_1028, w_173_1029, w_173_1035, w_173_1036, w_173_1037, w_173_1039, w_173_1041, w_173_1043, w_173_1050, w_173_1051, w_173_1053, w_173_1065, w_173_1071, w_173_1079, w_173_1080, w_173_1081, w_173_1087, w_173_1088, w_173_1097, w_173_1103, w_173_1107, w_173_1110, w_173_1118, w_173_1120, w_173_1123, w_173_1128, w_173_1129, w_173_1137, w_173_1139, w_173_1145, w_173_1148, w_173_1158, w_173_1159, w_173_1160, w_173_1162, w_173_1164, w_173_1167, w_173_1168, w_173_1169, w_173_1172, w_173_1177, w_173_1178, w_173_1179, w_173_1180, w_173_1187, w_173_1193, w_173_1195, w_173_1202, w_173_1203, w_173_1204, w_173_1208, w_173_1210, w_173_1214, w_173_1215, w_173_1217, w_173_1219, w_173_1223, w_173_1225, w_173_1226, w_173_1227, w_173_1237, w_173_1242, w_173_1246, w_173_1251, w_173_1252, w_173_1253, w_173_1260, w_173_1261, w_173_1263, w_173_1271, w_173_1273, w_173_1274, w_173_1276, w_173_1282, w_173_1291, w_173_1305, w_173_1306, w_173_1307, w_173_1308, w_173_1312, w_173_1313, w_173_1315, w_173_1316, w_173_1318, w_173_1322, w_173_1325, w_173_1332, w_173_1333, w_173_1334, w_173_1335, w_173_1360, w_173_1361, w_173_1362, w_173_1363, w_173_1367, w_173_1368, w_173_1379, w_173_1388, w_173_1392, w_173_1399, w_173_1401, w_173_1407, w_173_1415, w_173_1416, w_173_1421, w_173_1422, w_173_1426, w_173_1428, w_173_1431, w_173_1432, w_173_1433, w_173_1435, w_173_1436, w_173_1439, w_173_1448, w_173_1464, w_173_1469, w_173_1471, w_173_1478, w_173_1481, w_173_1482, w_173_1483, w_173_1484, w_173_1485, w_173_1488, w_173_1489, w_173_1493, w_173_1496, w_173_1497, w_173_1499, w_173_1500, w_173_1503, w_173_1504, w_173_1506, w_173_1507, w_173_1515, w_173_1520, w_173_1528, w_173_1529, w_173_1532, w_173_1535, w_173_1540, w_173_1542, w_173_1543, w_173_1545, w_173_1546, w_173_1558, w_173_1559, w_173_1560, w_173_1571, w_173_1572, w_173_1574, w_173_1587, w_173_1594, w_173_1596, w_173_1603, w_173_1606, w_173_1609, w_173_1616, w_173_1619, w_173_1622, w_173_1634, w_173_1646, w_173_1647, w_173_1650, w_173_1655, w_173_1664, w_173_1667, w_173_1675, w_173_1676, w_173_1690, w_173_1710, w_173_1727, w_173_1728, w_173_1730, w_173_1734, w_173_1738, w_173_1752, w_173_1754, w_173_1757, w_173_1768, w_173_1769, w_173_1775, w_173_1777, w_173_1779, w_173_1788, w_173_1789, w_173_1792, w_173_1801, w_173_1804, w_173_1806, w_173_1808, w_173_1809, w_173_1810, w_173_1812, w_173_1817, w_173_1821, w_173_1845, w_173_1848, w_173_1860, w_173_1863, w_173_1867, w_173_1875, w_173_1880, w_173_1891, w_173_1893, w_173_1895, w_173_1900, w_173_1902, w_173_1904, w_173_1909, w_173_1918, w_173_1919, w_173_1920, w_173_1921, w_173_1934, w_173_1936, w_173_1940, w_173_1944, w_173_1951, w_173_1952, w_173_1975, w_173_1978, w_173_1994, w_173_1997, w_173_1999, w_173_2010, w_173_2019, w_173_2021, w_173_2023, w_173_2030, w_173_2049, w_173_2050, w_173_2054, w_173_2056, w_173_2062, w_173_2079, w_173_2089, w_173_2093, w_173_2094, w_173_2100, w_173_2112, w_173_2120, w_173_2135, w_173_2139, w_173_2140, w_173_2146, w_173_2152, w_173_2154, w_173_2157, w_173_2167, w_173_2169, w_173_2172, w_173_2174, w_173_2175, w_173_2186, w_173_2206, w_173_2207, w_173_2209, w_173_2216, w_173_2225, w_173_2237, w_173_2248, w_173_2259, w_173_2265, w_173_2269, w_173_2274, w_173_2275, w_173_2285, w_173_2288, w_173_2289, w_173_2311, w_173_2312, w_173_2321, w_173_2326, w_173_2330, w_173_2332, w_173_2333, w_173_2334, w_173_2337, w_173_2370, w_173_2379, w_173_2381, w_173_2386, w_173_2395, w_173_2396, w_173_2403, w_173_2422, w_173_2425, w_173_2431, w_173_2433, w_173_2438, w_173_2448, w_173_2452, w_173_2455, w_173_2458, w_173_2466, w_173_2472, w_173_2481, w_173_2484, w_173_2489, w_173_2497, w_173_2499, w_173_2501, w_173_2502, w_173_2507, w_173_2511, w_173_2527, w_173_2529, w_173_2543, w_173_2544, w_173_2553, w_173_2556, w_173_2565, w_173_2577, w_173_2580, w_173_2581, w_173_2584, w_173_2610, w_173_2628, w_173_2631, w_173_2634, w_173_2637, w_173_2644, w_173_2650, w_173_2660, w_173_2663, w_173_2670, w_173_2672, w_173_2678, w_173_2686, w_173_2688, w_173_2704, w_173_2711, w_173_2713, w_173_2717, w_173_2721, w_173_2722, w_173_2728, w_173_2730, w_173_2736, w_173_2745, w_173_2746, w_173_2750, w_173_2754, w_173_2760, w_173_2762, w_173_2773, w_173_2792, w_173_2794, w_173_2799, w_173_2805, w_173_2817, w_173_2830, w_173_2831, w_173_2835, w_173_2836, w_173_2838, w_173_2843, w_173_2846, w_173_2855, w_173_2856, w_173_2857, w_173_2859, w_173_2870, w_173_2882, w_173_2897, w_173_2911, w_173_2922, w_173_2923, w_173_2926, w_173_2931, w_173_2933, w_173_2934, w_173_2937, w_173_2952, w_173_2953, w_173_2965, w_173_2980, w_173_2981, w_173_2986, w_173_2988, w_173_2989, w_173_2991, w_173_3040, w_173_3047, w_173_3050, w_173_3058, w_173_3071, w_173_3072, w_173_3082, w_173_3102, w_173_3105, w_173_3113, w_173_3126, w_173_3127, w_173_3137, w_173_3138, w_173_3149, w_173_3154, w_173_3159, w_173_3160, w_173_3168, w_173_3176, w_173_3178, w_173_3188, w_173_3192, w_173_3198, w_173_3202, w_173_3210, w_173_3213, w_173_3217, w_173_3222, w_173_3229, w_173_3243, w_173_3248, w_173_3251, w_173_3252, w_173_3254, w_173_3260, w_173_3264, w_173_3265, w_173_3280, w_173_3287, w_173_3289, w_173_3290, w_173_3298, w_173_3310, w_173_3312, w_173_3318, w_173_3323, w_173_3326, w_173_3332, w_173_3333, w_173_3343, w_173_3344, w_173_3345, w_173_3351, w_173_3358, w_173_3360, w_173_3391, w_173_3400, w_173_3401, w_173_3402, w_173_3403, w_173_3404, w_173_3405, w_173_3406, w_173_3408, w_173_3410, w_173_3411, w_173_3412, w_173_3413, w_173_3414, w_173_3415, w_173_3416, w_173_3418;
  wire w_174_003, w_174_004, w_174_006, w_174_007, w_174_011, w_174_016, w_174_019, w_174_020, w_174_021, w_174_027, w_174_030, w_174_031, w_174_035, w_174_036, w_174_048, w_174_069, w_174_073, w_174_079, w_174_081, w_174_089, w_174_094, w_174_099, w_174_101, w_174_103, w_174_106, w_174_116, w_174_123, w_174_128, w_174_132, w_174_152, w_174_153, w_174_159, w_174_161, w_174_162, w_174_164, w_174_165, w_174_170, w_174_172, w_174_173, w_174_176, w_174_184, w_174_185, w_174_190, w_174_192, w_174_196, w_174_197, w_174_204, w_174_205, w_174_207, w_174_210, w_174_215, w_174_220, w_174_222, w_174_225, w_174_227, w_174_230, w_174_231, w_174_239, w_174_241, w_174_242, w_174_247, w_174_259, w_174_264, w_174_267, w_174_270, w_174_281, w_174_284, w_174_293, w_174_296, w_174_299, w_174_300, w_174_301, w_174_304, w_174_316, w_174_318, w_174_319, w_174_320, w_174_325, w_174_329, w_174_331, w_174_338, w_174_343, w_174_344, w_174_346, w_174_348, w_174_359, w_174_361, w_174_362, w_174_366, w_174_370, w_174_373, w_174_375, w_174_381, w_174_383, w_174_386, w_174_393, w_174_396, w_174_397, w_174_398, w_174_403, w_174_406, w_174_408, w_174_411, w_174_415, w_174_419, w_174_427, w_174_434, w_174_435, w_174_440, w_174_442, w_174_455, w_174_458, w_174_461, w_174_469, w_174_482, w_174_484, w_174_492, w_174_493, w_174_495, w_174_498, w_174_500, w_174_510, w_174_536, w_174_539, w_174_541, w_174_542, w_174_546, w_174_549, w_174_550, w_174_551, w_174_552, w_174_553, w_174_559, w_174_566, w_174_568, w_174_570, w_174_581, w_174_583, w_174_584, w_174_591, w_174_593, w_174_598, w_174_604, w_174_606, w_174_609, w_174_611, w_174_612, w_174_615, w_174_621, w_174_624, w_174_626, w_174_642, w_174_651, w_174_652, w_174_653, w_174_655, w_174_658, w_174_659, w_174_661, w_174_670, w_174_674, w_174_681, w_174_683, w_174_685, w_174_687, w_174_692, w_174_699, w_174_701, w_174_703, w_174_713, w_174_716, w_174_717, w_174_725, w_174_727, w_174_730, w_174_731, w_174_733, w_174_736, w_174_737, w_174_739, w_174_741, w_174_742, w_174_746, w_174_753, w_174_756, w_174_757, w_174_759, w_174_761, w_174_762, w_174_764, w_174_768, w_174_778, w_174_785, w_174_786, w_174_790, w_174_791, w_174_792, w_174_800, w_174_803, w_174_805, w_174_809, w_174_811, w_174_823, w_174_826, w_174_836, w_174_840, w_174_842, w_174_854, w_174_861, w_174_866, w_174_869, w_174_873, w_174_878, w_174_883, w_174_884, w_174_885, w_174_886, w_174_890, w_174_891, w_174_896, w_174_897, w_174_904, w_174_906, w_174_911, w_174_912, w_174_913, w_174_917, w_174_919, w_174_923, w_174_925, w_174_928, w_174_934, w_174_939, w_174_941, w_174_948, w_174_954, w_174_968, w_174_972, w_174_976, w_174_983, w_174_987, w_174_993, w_174_997, w_174_999, w_174_1002, w_174_1008, w_174_1017, w_174_1019, w_174_1024, w_174_1028, w_174_1030, w_174_1031, w_174_1034, w_174_1040, w_174_1056, w_174_1069, w_174_1070, w_174_1071, w_174_1072, w_174_1073, w_174_1075, w_174_1084, w_174_1086, w_174_1088, w_174_1090, w_174_1092, w_174_1096, w_174_1097, w_174_1098, w_174_1111, w_174_1113, w_174_1115, w_174_1119, w_174_1120, w_174_1121, w_174_1129, w_174_1131, w_174_1137, w_174_1142, w_174_1149, w_174_1150, w_174_1154, w_174_1155, w_174_1163, w_174_1165, w_174_1171, w_174_1179, w_174_1180, w_174_1181, w_174_1190, w_174_1192, w_174_1193, w_174_1201, w_174_1202, w_174_1204, w_174_1205, w_174_1218, w_174_1221, w_174_1223, w_174_1225, w_174_1227, w_174_1228, w_174_1229, w_174_1239, w_174_1245, w_174_1248, w_174_1249, w_174_1250, w_174_1255, w_174_1256, w_174_1260, w_174_1261, w_174_1263, w_174_1264, w_174_1272, w_174_1283, w_174_1284, w_174_1297, w_174_1299, w_174_1300, w_174_1302, w_174_1304, w_174_1305, w_174_1318, w_174_1319, w_174_1326, w_174_1327, w_174_1328, w_174_1330, w_174_1334, w_174_1342, w_174_1345, w_174_1347, w_174_1352, w_174_1357, w_174_1361, w_174_1364, w_174_1366, w_174_1367, w_174_1368, w_174_1369, w_174_1376, w_174_1382, w_174_1388, w_174_1401, w_174_1402, w_174_1403, w_174_1404, w_174_1405, w_174_1406, w_174_1415, w_174_1419, w_174_1427, w_174_1428, w_174_1429, w_174_1439, w_174_1446, w_174_1448, w_174_1453, w_174_1458, w_174_1464, w_174_1465, w_174_1466, w_174_1467, w_174_1472, w_174_1477, w_174_1478, w_174_1481, w_174_1482, w_174_1483, w_174_1484, w_174_1487, w_174_1489, w_174_1491, w_174_1492, w_174_1493, w_174_1497, w_174_1503, w_174_1506, w_174_1507, w_174_1515, w_174_1516, w_174_1518, w_174_1525, w_174_1528, w_174_1530, w_174_1531, w_174_1532, w_174_1535, w_174_1541, w_174_1551, w_174_1553, w_174_1555, w_174_1557, w_174_1560, w_174_1564, w_174_1565, w_174_1569, w_174_1579, w_174_1586, w_174_1596, w_174_1602, w_174_1604, w_174_1608, w_174_1610, w_174_1620, w_174_1629, w_174_1640, w_174_1647, w_174_1654, w_174_1664, w_174_1670, w_174_1674, w_174_1676, w_174_1682, w_174_1699, w_174_1700, w_174_1705, w_174_1709, w_174_1712, w_174_1721, w_174_1729, w_174_1742, w_174_1752, w_174_1758, w_174_1760, w_174_1771, w_174_1778, w_174_1781, w_174_1790, w_174_1794, w_174_1810, w_174_1811, w_174_1812, w_174_1824, w_174_1837, w_174_1838, w_174_1842, w_174_1844, w_174_1853, w_174_1858, w_174_1870, w_174_1885, w_174_1896, w_174_1908, w_174_1909, w_174_1910, w_174_1913, w_174_1920, w_174_1921, w_174_1928, w_174_1937, w_174_1941, w_174_1946, w_174_1965, w_174_1969, w_174_1974, w_174_1979, w_174_1980, w_174_1990, w_174_1991, w_174_1994, w_174_1997, w_174_1999, w_174_2004, w_174_2005, w_174_2007, w_174_2015, w_174_2030, w_174_2043, w_174_2050, w_174_2055, w_174_2059, w_174_2060, w_174_2069, w_174_2076, w_174_2079, w_174_2084, w_174_2089, w_174_2090, w_174_2094, w_174_2099, w_174_2115, w_174_2131, w_174_2144, w_174_2150, w_174_2151, w_174_2159, w_174_2160, w_174_2162, w_174_2166, w_174_2169, w_174_2173, w_174_2178, w_174_2179, w_174_2185, w_174_2193, w_174_2199, w_174_2200, w_174_2218, w_174_2219, w_174_2247, w_174_2250, w_174_2251, w_174_2252, w_174_2256, w_174_2278, w_174_2292, w_174_2294, w_174_2299, w_174_2330, w_174_2333, w_174_2334, w_174_2336, w_174_2342, w_174_2357, w_174_2359, w_174_2361, w_174_2365, w_174_2372, w_174_2385, w_174_2387, w_174_2392, w_174_2393, w_174_2396, w_174_2398, w_174_2406, w_174_2409, w_174_2417, w_174_2419, w_174_2422, w_174_2426, w_174_2432, w_174_2434, w_174_2435, w_174_2437, w_174_2448, w_174_2451, w_174_2453, w_174_2454, w_174_2455, w_174_2471, w_174_2475, w_174_2486, w_174_2488, w_174_2493, w_174_2498, w_174_2499, w_174_2506, w_174_2509, w_174_2511, w_174_2519, w_174_2522, w_174_2527, w_174_2544, w_174_2547, w_174_2555, w_174_2566, w_174_2576, w_174_2584, w_174_2587, w_174_2588, w_174_2589, w_174_2591, w_174_2592, w_174_2612, w_174_2613, w_174_2625, w_174_2626, w_174_2634, w_174_2655, w_174_2657, w_174_2663, w_174_2676, w_174_2691, w_174_2695, w_174_2696, w_174_2701, w_174_2703, w_174_2706, w_174_2711, w_174_2718, w_174_2719, w_174_2725, w_174_2728, w_174_2740, w_174_2745, w_174_2746, w_174_2748, w_174_2750, w_174_2753, w_174_2754, w_174_2760, w_174_2767, w_174_2784, w_174_2788, w_174_2798, w_174_2799, w_174_2808, w_174_2814, w_174_2818, w_174_2824, w_174_2826, w_174_2827, w_174_2831, w_174_2837, w_174_2842, w_174_2844, w_174_2851, w_174_2855, w_174_2860, w_174_2862, w_174_2864, w_174_2866, w_174_2868, w_174_2876, w_174_2909, w_174_2946, w_174_2947, w_174_2949, w_174_2953, w_174_2962, w_174_2968, w_174_2971, w_174_2980, w_174_2982, w_174_2988, w_174_2991, w_174_2992, w_174_2994, w_174_3000, w_174_3008, w_174_3032, w_174_3054, w_174_3057, w_174_3071, w_174_3072, w_174_3073, w_174_3074, w_174_3093, w_174_3109, w_174_3115, w_174_3128, w_174_3139, w_174_3155, w_174_3157, w_174_3166, w_174_3176, w_174_3177, w_174_3178, w_174_3189, w_174_3194, w_174_3214, w_174_3225, w_174_3228, w_174_3233, w_174_3241, w_174_3253, w_174_3255, w_174_3291, w_174_3294, w_174_3301, w_174_3304, w_174_3313, w_174_3314, w_174_3318, w_174_3321, w_174_3324, w_174_3327, w_174_3328, w_174_3329, w_174_3332, w_174_3338, w_174_3340, w_174_3343, w_174_3345, w_174_3351, w_174_3354, w_174_3359, w_174_3360, w_174_3366, w_174_3369, w_174_3393, w_174_3395, w_174_3399, w_174_3400, w_174_3405, w_174_3408, w_174_3418, w_174_3419, w_174_3433, w_174_3434, w_174_3440;
  wire w_175_000, w_175_003, w_175_005, w_175_006, w_175_007, w_175_012, w_175_013, w_175_016, w_175_018, w_175_019, w_175_020, w_175_021, w_175_022, w_175_025, w_175_026, w_175_028, w_175_029, w_175_030, w_175_032, w_175_033, w_175_034, w_175_036, w_175_037, w_175_038, w_175_042, w_175_048, w_175_049, w_175_050, w_175_051, w_175_052, w_175_053, w_175_054, w_175_055, w_175_056, w_175_057, w_175_058, w_175_060, w_175_061, w_175_063, w_175_064, w_175_065, w_175_066, w_175_067, w_175_068, w_175_071, w_175_072, w_175_074, w_175_075, w_175_079, w_175_081, w_175_084, w_175_085, w_175_087, w_175_088, w_175_089, w_175_091, w_175_092, w_175_093, w_175_094, w_175_098, w_175_100, w_175_101, w_175_102, w_175_103, w_175_104, w_175_106, w_175_107, w_175_108, w_175_109, w_175_110, w_175_111, w_175_113, w_175_115, w_175_116, w_175_121, w_175_124, w_175_125, w_175_126, w_175_127, w_175_128, w_175_130, w_175_131, w_175_133, w_175_136, w_175_137, w_175_140, w_175_141, w_175_142, w_175_144, w_175_145, w_175_148, w_175_149, w_175_152, w_175_154, w_175_155, w_175_156, w_175_158, w_175_161, w_175_162, w_175_163, w_175_165, w_175_166, w_175_168, w_175_169, w_175_170, w_175_172, w_175_173, w_175_177, w_175_180, w_175_184, w_175_193, w_175_195, w_175_196, w_175_197, w_175_198, w_175_203, w_175_206, w_175_209, w_175_210, w_175_211, w_175_212, w_175_213, w_175_214, w_175_215, w_175_218, w_175_219, w_175_220, w_175_222, w_175_223, w_175_225, w_175_228, w_175_229, w_175_230, w_175_231, w_175_232, w_175_233, w_175_234, w_175_237, w_175_239, w_175_240, w_175_241, w_175_242, w_175_243, w_175_244, w_175_245, w_175_246, w_175_248, w_175_250, w_175_251, w_175_253, w_175_256, w_175_262, w_175_264, w_175_266, w_175_268, w_175_271, w_175_272, w_175_275, w_175_276, w_175_277, w_175_279, w_175_281, w_175_282, w_175_284, w_175_286, w_175_287, w_175_288, w_175_292, w_175_295, w_175_296, w_175_299, w_175_300, w_175_303, w_175_304, w_175_307, w_175_308, w_175_309, w_175_310, w_175_311, w_175_312, w_175_315, w_175_316, w_175_318, w_175_320, w_175_322, w_175_324, w_175_327, w_175_328, w_175_329, w_175_333, w_175_334, w_175_335, w_175_336, w_175_337, w_175_338, w_175_339, w_175_341, w_175_342, w_175_344, w_175_345, w_175_346, w_175_349, w_175_350, w_175_351, w_175_352, w_175_353, w_175_354, w_175_355, w_175_357, w_175_360, w_175_361, w_175_362, w_175_363, w_175_366, w_175_368, w_175_369, w_175_371, w_175_373, w_175_377, w_175_379, w_175_383, w_175_384, w_175_386, w_175_387, w_175_388, w_175_389, w_175_392, w_175_394, w_175_395, w_175_396, w_175_397, w_175_400, w_175_401, w_175_402, w_175_406, w_175_407, w_175_408, w_175_409, w_175_415, w_175_416, w_175_419, w_175_421, w_175_426, w_175_427, w_175_429, w_175_430, w_175_431, w_175_432, w_175_435, w_175_436, w_175_439, w_175_440, w_175_444, w_175_445, w_175_446, w_175_449, w_175_450, w_175_451, w_175_452, w_175_455, w_175_457, w_175_458, w_175_464, w_175_465, w_175_466, w_175_467, w_175_469, w_175_470, w_175_471, w_175_474, w_175_475, w_175_476, w_175_478, w_175_479, w_175_482, w_175_485, w_175_489, w_175_492, w_175_495, w_175_496, w_175_498, w_175_500, w_175_501, w_175_502, w_175_503, w_175_505, w_175_507, w_175_508, w_175_510, w_175_512, w_175_514, w_175_516, w_175_517, w_175_519, w_175_520, w_175_523, w_175_524, w_175_525, w_175_526, w_175_530, w_175_533, w_175_534, w_175_535, w_175_538, w_175_543, w_175_544, w_175_546, w_175_547, w_175_548, w_175_550, w_175_554, w_175_556, w_175_557, w_175_558, w_175_560, w_175_562, w_175_565, w_175_566, w_175_567, w_175_569, w_175_572, w_175_573, w_175_576, w_175_578, w_175_579, w_175_581, w_175_584, w_175_585, w_175_587, w_175_588, w_175_589, w_175_590, w_175_592, w_175_594, w_175_595, w_175_597, w_175_598, w_175_599, w_175_603, w_175_604, w_175_605, w_175_608, w_175_610, w_175_612, w_175_614, w_175_615, w_175_617, w_175_619, w_175_620, w_175_621, w_175_622, w_175_623, w_175_624, w_175_626, w_175_628, w_175_631, w_175_632, w_175_633, w_175_634, w_175_635, w_175_638, w_175_639, w_175_640, w_175_642, w_175_644, w_175_646, w_175_648, w_175_650, w_175_652, w_175_653, w_175_654, w_175_657, w_175_658, w_175_660, w_175_665, w_175_666, w_175_670, w_175_673, w_175_675, w_175_679, w_175_680, w_175_682, w_175_684, w_175_686, w_175_690, w_175_691, w_175_692, w_175_694, w_175_695, w_175_697, w_175_699, w_175_700, w_175_704, w_175_706, w_175_709, w_175_718, w_175_719, w_175_720, w_175_721, w_175_722, w_175_723, w_175_726, w_175_727, w_175_728, w_175_729, w_175_730, w_175_733, w_175_734, w_175_735, w_175_737, w_175_739, w_175_744, w_175_747, w_175_748, w_175_749, w_175_750, w_175_751, w_175_755, w_175_757, w_175_758, w_175_760, w_175_763, w_175_765, w_175_767, w_175_770, w_175_771, w_175_773, w_175_774, w_175_777, w_175_778, w_175_779, w_175_781, w_175_784, w_175_785, w_175_787, w_175_789, w_175_791, w_175_792, w_175_793, w_175_796, w_175_799, w_175_800, w_175_802, w_175_803, w_175_804, w_175_806, w_175_807, w_175_809, w_175_811, w_175_812, w_175_813, w_175_814, w_175_815, w_175_816, w_175_817, w_175_819, w_175_820, w_175_822, w_175_824, w_175_825, w_175_827, w_175_828, w_175_833, w_175_834, w_175_838, w_175_839, w_175_840, w_175_842, w_175_845, w_175_848, w_175_849, w_175_851, w_175_852, w_175_854, w_175_857, w_175_861, w_175_863, w_175_864, w_175_866, w_175_867, w_175_870, w_175_873, w_175_874, w_175_876, w_175_879, w_175_880, w_175_881, w_175_882, w_175_883, w_175_884, w_175_886, w_175_887, w_175_889, w_175_893, w_175_894, w_175_895, w_175_896, w_175_898, w_175_899, w_175_900, w_175_903, w_175_904, w_175_908, w_175_909, w_175_910, w_175_913, w_175_914, w_175_916, w_175_917, w_175_919, w_175_920, w_175_921, w_175_923, w_175_925, w_175_926, w_175_927, w_175_929, w_175_930, w_175_931, w_175_932, w_175_933, w_175_934, w_175_935, w_175_936, w_175_938, w_175_941, w_175_942, w_175_943, w_175_944, w_175_945, w_175_946, w_175_947, w_175_948, w_175_949, w_175_950, w_175_952, w_175_953, w_175_955, w_175_956, w_175_957, w_175_959, w_175_960, w_175_961, w_175_962, w_175_964, w_175_965, w_175_966, w_175_967, w_175_973;
  wire w_176_000, w_176_001, w_176_002, w_176_003, w_176_004, w_176_005, w_176_006, w_176_007, w_176_008, w_176_009, w_176_010, w_176_011, w_176_012, w_176_013, w_176_014, w_176_015, w_176_016, w_176_017, w_176_018, w_176_019, w_176_020, w_176_021, w_176_022, w_176_023, w_176_024, w_176_025, w_176_026, w_176_027, w_176_028, w_176_029, w_176_030, w_176_031, w_176_032, w_176_033, w_176_034, w_176_035, w_176_036, w_176_037, w_176_038, w_176_039, w_176_040, w_176_041, w_176_042, w_176_043, w_176_044, w_176_045, w_176_046, w_176_047, w_176_048, w_176_049, w_176_050, w_176_051, w_176_052, w_176_053, w_176_054, w_176_055, w_176_056, w_176_057, w_176_058, w_176_059, w_176_060, w_176_061, w_176_062, w_176_063, w_176_064, w_176_065, w_176_066, w_176_067, w_176_068, w_176_069, w_176_070, w_176_072, w_176_073, w_176_074, w_176_075, w_176_076, w_176_077, w_176_078, w_176_079, w_176_080;
  wire w_177_012, w_177_021, w_177_024, w_177_032, w_177_033, w_177_035, w_177_037, w_177_039, w_177_040, w_177_044, w_177_045, w_177_046, w_177_048, w_177_056, w_177_060, w_177_061, w_177_071, w_177_078, w_177_080, w_177_081, w_177_083, w_177_085, w_177_087, w_177_088, w_177_090, w_177_095, w_177_100, w_177_101, w_177_102, w_177_109, w_177_110, w_177_115, w_177_120, w_177_121, w_177_122, w_177_138, w_177_143, w_177_144, w_177_147, w_177_149, w_177_150, w_177_157, w_177_158, w_177_163, w_177_165, w_177_167, w_177_168, w_177_169, w_177_174, w_177_176, w_177_180, w_177_181, w_177_183, w_177_186, w_177_189, w_177_196, w_177_197, w_177_198, w_177_205, w_177_208, w_177_213, w_177_221, w_177_222, w_177_223, w_177_225, w_177_233, w_177_234, w_177_237, w_177_240, w_177_241, w_177_242, w_177_243, w_177_247, w_177_248, w_177_249, w_177_250, w_177_253, w_177_256, w_177_261, w_177_266, w_177_268, w_177_270, w_177_280, w_177_288, w_177_290, w_177_291, w_177_300, w_177_301, w_177_307, w_177_309, w_177_315, w_177_331, w_177_334, w_177_337, w_177_340, w_177_341, w_177_344, w_177_351, w_177_355, w_177_357, w_177_362, w_177_364, w_177_368, w_177_369, w_177_374, w_177_375, w_177_377, w_177_384, w_177_391, w_177_394, w_177_400, w_177_401, w_177_405, w_177_407, w_177_415, w_177_423, w_177_427, w_177_433, w_177_434, w_177_437, w_177_438, w_177_444, w_177_446, w_177_447, w_177_448, w_177_451, w_177_453, w_177_457, w_177_460, w_177_462, w_177_463, w_177_466, w_177_468, w_177_469, w_177_472, w_177_477, w_177_479, w_177_482, w_177_483, w_177_487, w_177_496, w_177_498, w_177_499, w_177_500, w_177_503, w_177_508, w_177_510, w_177_511, w_177_516, w_177_517, w_177_518, w_177_520, w_177_521, w_177_527, w_177_531, w_177_533, w_177_539, w_177_552, w_177_553, w_177_555, w_177_559, w_177_561, w_177_564, w_177_565, w_177_581, w_177_582, w_177_586, w_177_587, w_177_589, w_177_605, w_177_608, w_177_613, w_177_616, w_177_619, w_177_622, w_177_623, w_177_629, w_177_633, w_177_635, w_177_641, w_177_645, w_177_646, w_177_650, w_177_651, w_177_652, w_177_653, w_177_664, w_177_669, w_177_674, w_177_681, w_177_690, w_177_700, w_177_703, w_177_705, w_177_706, w_177_707, w_177_711, w_177_721, w_177_725, w_177_727, w_177_728, w_177_734, w_177_736, w_177_744, w_177_745, w_177_746, w_177_747, w_177_748, w_177_752, w_177_758, w_177_765, w_177_769, w_177_777, w_177_779, w_177_780, w_177_781, w_177_783, w_177_784, w_177_787, w_177_790, w_177_797, w_177_800, w_177_809, w_177_810, w_177_814, w_177_828, w_177_840, w_177_843, w_177_853, w_177_862, w_177_865, w_177_874, w_177_875, w_177_887, w_177_889, w_177_891, w_177_894, w_177_895, w_177_897, w_177_899, w_177_900, w_177_912, w_177_918, w_177_919, w_177_923, w_177_924, w_177_941, w_177_947, w_177_957, w_177_959, w_177_962, w_177_963, w_177_975, w_177_981, w_177_987, w_177_988, w_177_991, w_177_992, w_177_1001, w_177_1007, w_177_1013, w_177_1014, w_177_1019, w_177_1020, w_177_1024, w_177_1027, w_177_1033, w_177_1034, w_177_1035, w_177_1039, w_177_1043, w_177_1048, w_177_1051, w_177_1052, w_177_1054, w_177_1055, w_177_1057, w_177_1060, w_177_1062, w_177_1063, w_177_1064, w_177_1066, w_177_1078, w_177_1083, w_177_1086, w_177_1089, w_177_1090, w_177_1093, w_177_1094, w_177_1097, w_177_1102, w_177_1111, w_177_1118, w_177_1120, w_177_1121, w_177_1125, w_177_1127, w_177_1128, w_177_1133, w_177_1144, w_177_1146, w_177_1147, w_177_1154, w_177_1157, w_177_1158, w_177_1159, w_177_1164, w_177_1168, w_177_1172, w_177_1174, w_177_1179, w_177_1183, w_177_1187, w_177_1188, w_177_1191, w_177_1195, w_177_1202, w_177_1203, w_177_1204, w_177_1205, w_177_1210, w_177_1212, w_177_1216, w_177_1217, w_177_1221, w_177_1231, w_177_1233, w_177_1238, w_177_1241, w_177_1242, w_177_1244, w_177_1245, w_177_1247, w_177_1251, w_177_1254, w_177_1255, w_177_1256, w_177_1258, w_177_1260, w_177_1262, w_177_1263, w_177_1272, w_177_1276, w_177_1278, w_177_1280, w_177_1281, w_177_1283, w_177_1285, w_177_1302, w_177_1306, w_177_1313, w_177_1321, w_177_1323, w_177_1324, w_177_1327, w_177_1329, w_177_1337, w_177_1344, w_177_1345, w_177_1347, w_177_1348, w_177_1350, w_177_1354, w_177_1357, w_177_1363, w_177_1368, w_177_1371, w_177_1372, w_177_1375, w_177_1378, w_177_1379, w_177_1380, w_177_1385, w_177_1391, w_177_1404, w_177_1407, w_177_1408, w_177_1413, w_177_1416, w_177_1423, w_177_1427, w_177_1430, w_177_1433, w_177_1434, w_177_1436, w_177_1437, w_177_1442, w_177_1445, w_177_1452, w_177_1454, w_177_1455, w_177_1467, w_177_1470, w_177_1474, w_177_1477, w_177_1478, w_177_1479, w_177_1483, w_177_1485, w_177_1486, w_177_1490, w_177_1491, w_177_1505, w_177_1507, w_177_1520, w_177_1527, w_177_1531, w_177_1532, w_177_1536, w_177_1541, w_177_1543, w_177_1546, w_177_1547, w_177_1549, w_177_1550, w_177_1554, w_177_1555, w_177_1560, w_177_1562, w_177_1563, w_177_1575, w_177_1580, w_177_1587, w_177_1589, w_177_1590, w_177_1591, w_177_1592, w_177_1602, w_177_1603, w_177_1609, w_177_1614, w_177_1617, w_177_1619, w_177_1621, w_177_1631, w_177_1634, w_177_1637, w_177_1638, w_177_1640, w_177_1643, w_177_1645, w_177_1648, w_177_1649, w_177_1660, w_177_1664, w_177_1667, w_177_1672, w_177_1676, w_177_1685, w_177_1686, w_177_1689, w_177_1690, w_177_1692, w_177_1694, w_177_1698, w_177_1700, w_177_1708, w_177_1709, w_177_1712, w_177_1713, w_177_1716, w_177_1718, w_177_1721, w_177_1724, w_177_1725, w_177_1735, w_177_1736, w_177_1740, w_177_1743, w_177_1749, w_177_1750, w_177_1752, w_177_1753, w_177_1759, w_177_1762, w_177_1764, w_177_1768, w_177_1770, w_177_1773, w_177_1776, w_177_1780, w_177_1781, w_177_1785, w_177_1788, w_177_1802, w_177_1804, w_177_1807, w_177_1808, w_177_1811, w_177_1812, w_177_1815, w_177_1817, w_177_1821, w_177_1824, w_177_1825, w_177_1827, w_177_1836, w_177_1841, w_177_1849, w_177_1851, w_177_1856, w_177_1859, w_177_1860, w_177_1865, w_177_1868, w_177_1870, w_177_1873, w_177_1876, w_177_1894, w_177_1895, w_177_1897, w_177_1898, w_177_1900, w_177_1901, w_177_1918, w_177_1920, w_177_1925, w_177_1935, w_177_1941, w_177_1949, w_177_1957, w_177_1963, w_177_1970, w_177_1972, w_177_1978, w_177_1982, w_177_1985, w_177_1987, w_177_1989, w_177_1993, w_177_2009, w_177_2017, w_177_2018, w_177_2020, w_177_2027, w_177_2035, w_177_2038, w_177_2047, w_177_2054, w_177_2059, w_177_2060, w_177_2065, w_177_2074, w_177_2081, w_177_2098, w_177_2100, w_177_2101, w_177_2104, w_177_2108, w_177_2114, w_177_2122, w_177_2124, w_177_2125, w_177_2126, w_177_2134, w_177_2161, w_177_2177, w_177_2184, w_177_2187, w_177_2188, w_177_2193, w_177_2198, w_177_2202, w_177_2203, w_177_2220, w_177_2224, w_177_2226, w_177_2230, w_177_2233, w_177_2244, w_177_2247, w_177_2251, w_177_2254, w_177_2269, w_177_2277, w_177_2280, w_177_2283, w_177_2290, w_177_2291, w_177_2296, w_177_2297, w_177_2309, w_177_2317, w_177_2319, w_177_2325, w_177_2332, w_177_2345, w_177_2363, w_177_2383, w_177_2396, w_177_2404, w_177_2408, w_177_2416, w_177_2417, w_177_2431, w_177_2442, w_177_2447, w_177_2456, w_177_2457, w_177_2459, w_177_2463, w_177_2464, w_177_2474, w_177_2478, w_177_2484, w_177_2499, w_177_2503, w_177_2518, w_177_2522, w_177_2525, w_177_2544, w_177_2552, w_177_2555, w_177_2557, w_177_2567, w_177_2582, w_177_2583, w_177_2585, w_177_2589, w_177_2598, w_177_2602, w_177_2614, w_177_2628, w_177_2645, w_177_2648, w_177_2649, w_177_2657, w_177_2661, w_177_2675, w_177_2685, w_177_2687, w_177_2689, w_177_2701, w_177_2702, w_177_2708, w_177_2709, w_177_2716, w_177_2733, w_177_2743, w_177_2748, w_177_2750, w_177_2752, w_177_2753, w_177_2765, w_177_2773, w_177_2776, w_177_2785, w_177_2798, w_177_2802, w_177_2806, w_177_2811, w_177_2814, w_177_2815, w_177_2817, w_177_2829, w_177_2831, w_177_2833, w_177_2839, w_177_2863, w_177_2904, w_177_2911, w_177_2914, w_177_2928, w_177_2929, w_177_2934, w_177_2941, w_177_2946, w_177_2954, w_177_2958, w_177_2976, w_177_2978, w_177_2982, w_177_3003, w_177_3008, w_177_3011, w_177_3013, w_177_3015, w_177_3017, w_177_3021, w_177_3025, w_177_3036, w_177_3039, w_177_3042, w_177_3044, w_177_3047, w_177_3053, w_177_3058, w_177_3067, w_177_3068, w_177_3084, w_177_3086, w_177_3087, w_177_3093;
  wire w_178_004, w_178_006, w_178_008, w_178_010, w_178_012, w_178_013, w_178_015, w_178_016, w_178_017, w_178_020, w_178_021, w_178_024, w_178_025, w_178_027, w_178_033, w_178_034, w_178_035, w_178_036, w_178_042, w_178_044, w_178_046, w_178_047, w_178_048, w_178_049, w_178_050, w_178_052, w_178_053, w_178_054, w_178_055, w_178_056, w_178_063, w_178_064, w_178_067, w_178_068, w_178_072, w_178_075, w_178_076, w_178_078, w_178_079, w_178_080, w_178_083, w_178_086, w_178_087, w_178_088, w_178_089, w_178_090, w_178_093, w_178_094, w_178_095, w_178_098, w_178_100, w_178_103, w_178_107, w_178_108, w_178_110, w_178_112, w_178_117, w_178_118, w_178_120, w_178_122, w_178_123, w_178_124, w_178_128, w_178_129, w_178_130, w_178_132, w_178_134, w_178_139, w_178_140, w_178_142, w_178_144, w_178_145, w_178_146, w_178_147, w_178_148, w_178_150, w_178_151, w_178_152, w_178_153, w_178_155, w_178_156, w_178_159, w_178_160, w_178_161, w_178_162, w_178_163, w_178_165, w_178_167, w_178_168, w_178_169, w_178_170, w_178_172, w_178_174, w_178_177, w_178_178, w_178_179, w_178_180, w_178_181, w_178_183, w_178_187, w_178_188, w_178_189, w_178_191, w_178_192, w_178_193, w_178_195, w_178_197, w_178_198, w_178_199, w_178_200, w_178_204, w_178_205, w_178_206, w_178_213, w_178_215, w_178_216, w_178_217, w_178_218, w_178_219, w_178_222, w_178_223, w_178_224, w_178_226, w_178_230, w_178_233, w_178_241, w_178_242, w_178_246, w_178_247, w_178_248, w_178_251, w_178_252, w_178_257, w_178_259, w_178_262, w_178_263, w_178_264, w_178_267, w_178_268, w_178_273, w_178_276, w_178_279, w_178_280, w_178_286, w_178_287, w_178_288, w_178_289, w_178_290, w_178_294, w_178_296, w_178_299, w_178_300, w_178_303, w_178_307, w_178_309, w_178_310, w_178_314, w_178_315, w_178_317, w_178_318, w_178_319, w_178_320, w_178_324, w_178_325, w_178_326, w_178_327, w_178_330, w_178_331, w_178_332, w_178_336, w_178_337, w_178_340, w_178_341, w_178_343, w_178_345, w_178_349, w_178_350, w_178_356, w_178_357, w_178_358, w_178_360, w_178_361, w_178_363, w_178_364, w_178_365, w_178_366, w_178_370, w_178_372, w_178_373, w_178_374, w_178_392, w_178_395, w_178_400, w_178_402, w_178_406, w_178_415, w_178_422, w_178_423, w_178_428, w_178_432, w_178_434, w_178_438, w_178_439, w_178_442, w_178_443, w_178_444, w_178_446, w_178_448, w_178_451, w_178_452, w_178_453, w_178_460, w_178_461, w_178_464, w_178_466, w_178_468, w_178_469, w_178_471, w_178_473, w_178_476, w_178_478, w_178_479, w_178_480, w_178_484, w_178_485, w_178_488, w_178_490, w_178_496, w_178_501, w_178_502, w_178_507, w_178_513, w_178_514, w_178_518, w_178_519, w_178_523, w_178_527, w_178_532, w_178_534, w_178_544, w_178_550, w_178_551, w_178_552, w_178_553, w_178_559, w_178_562, w_178_563, w_178_564, w_178_565, w_178_567, w_178_568, w_178_569, w_178_570, w_178_571, w_178_574, w_178_582, w_178_583, w_178_584, w_178_589, w_178_593, w_178_597, w_178_603, w_178_605, w_178_606, w_178_610, w_178_611, w_178_616, w_178_617, w_178_618, w_178_623, w_178_624, w_178_631, w_178_632, w_178_637, w_178_638, w_178_639, w_178_641, w_178_643, w_178_644, w_178_645, w_178_646, w_178_647, w_178_648, w_178_649, w_178_650, w_178_653, w_178_654, w_178_655, w_178_658, w_178_660, w_178_662, w_178_667, w_178_668, w_178_669, w_178_670, w_178_671, w_178_673, w_178_674, w_178_675, w_178_678, w_178_679, w_178_680, w_178_686, w_178_688, w_178_693, w_178_694, w_178_696, w_178_700, w_178_701, w_178_703, w_178_705, w_178_709, w_178_715, w_178_719, w_178_724, w_178_725, w_178_726, w_178_730, w_178_733, w_178_734, w_178_736, w_178_737, w_178_742, w_178_744, w_178_749, w_178_750, w_178_756, w_178_758, w_178_760, w_178_763, w_178_765, w_178_768, w_178_769, w_178_770, w_178_771, w_178_775, w_178_778, w_178_784, w_178_786, w_178_787, w_178_788, w_178_790, w_178_792, w_178_793, w_178_801, w_178_807, w_178_808, w_178_810, w_178_817, w_178_820, w_178_821, w_178_822, w_178_830, w_178_832, w_178_836, w_178_839, w_178_840, w_178_841, w_178_846, w_178_849, w_178_850, w_178_851, w_178_852, w_178_855, w_178_857, w_178_858, w_178_859, w_178_861, w_178_866, w_178_868, w_178_869, w_178_870, w_178_873, w_178_875, w_178_877, w_178_887, w_178_888, w_178_889, w_178_895, w_178_898, w_178_903, w_178_904, w_178_905, w_178_906, w_178_909, w_178_915, w_178_921, w_178_923, w_178_929, w_178_930, w_178_932, w_178_934, w_178_936, w_178_942, w_178_943, w_178_944, w_178_948, w_178_950, w_178_953, w_178_954, w_178_955, w_178_957, w_178_959, w_178_963, w_178_965, w_178_968, w_178_969, w_178_971, w_178_972, w_178_973, w_178_977, w_178_978, w_178_982, w_178_985, w_178_986, w_178_987, w_178_988, w_178_989, w_178_993, w_178_994, w_178_995, w_178_997, w_178_999, w_178_1002, w_178_1004, w_178_1009, w_178_1011, w_178_1013, w_178_1015, w_178_1016, w_178_1018, w_178_1019, w_178_1020, w_178_1023, w_178_1024, w_178_1028, w_178_1029, w_178_1030, w_178_1032, w_178_1035, w_178_1036, w_178_1038, w_178_1039, w_178_1040, w_178_1044, w_178_1048, w_178_1051, w_178_1053, w_178_1056, w_178_1060, w_178_1062, w_178_1065, w_178_1067, w_178_1068, w_178_1073, w_178_1077, w_178_1078, w_178_1080, w_178_1082, w_178_1083, w_178_1087, w_178_1089, w_178_1094, w_178_1097, w_178_1098, w_178_1101, w_178_1103, w_178_1105, w_178_1106, w_178_1110, w_178_1112, w_178_1113, w_178_1116, w_178_1117, w_178_1118, w_178_1124, w_178_1127, w_178_1128, w_178_1129, w_178_1132, w_178_1136, w_178_1137, w_178_1144, w_178_1150, w_178_1151, w_178_1155, w_178_1158, w_178_1160, w_178_1161, w_178_1165, w_178_1167, w_178_1168, w_178_1171, w_178_1173, w_178_1174, w_178_1181, w_178_1186, w_178_1187, w_178_1191, w_178_1194, w_178_1195, w_178_1200, w_178_1201, w_178_1205, w_178_1208, w_178_1213, w_178_1214, w_178_1215, w_178_1216, w_178_1217, w_178_1219, w_178_1221, w_178_1222, w_178_1225, w_178_1227, w_178_1228, w_178_1229, w_178_1231, w_178_1234, w_178_1235, w_178_1236, w_178_1237, w_178_1238, w_178_1243, w_178_1244, w_178_1245, w_178_1246, w_178_1254, w_178_1257, w_178_1262, w_178_1264, w_178_1266, w_178_1272, w_178_1274, w_178_1278, w_178_1279, w_178_1281, w_178_1282, w_178_1283, w_178_1288, w_178_1294, w_178_1295, w_178_1296, w_178_1297, w_178_1299, w_178_1304, w_178_1306, w_178_1307, w_178_1309, w_178_1311, w_178_1313, w_178_1317, w_178_1320, w_178_1322, w_178_1329, w_178_1332, w_178_1334, w_178_1335, w_178_1343, w_178_1344, w_178_1345, w_178_1347, w_178_1355, w_178_1357, w_178_1362, w_178_1363, w_178_1364, w_178_1367, w_178_1369, w_178_1370, w_178_1371, w_178_1372, w_178_1379, w_178_1380, w_178_1381, w_178_1384, w_178_1387, w_178_1390, w_178_1391, w_178_1394, w_178_1395, w_178_1397, w_178_1402, w_178_1403, w_178_1404, w_178_1406, w_178_1408, w_178_1409, w_178_1412, w_178_1419, w_178_1420, w_178_1422, w_178_1432, w_178_1435, w_178_1436, w_178_1439, w_178_1442, w_178_1444, w_178_1446, w_178_1447, w_178_1449, w_178_1453, w_178_1456, w_178_1457, w_178_1459, w_178_1460, w_178_1461, w_178_1462, w_178_1463, w_178_1464, w_178_1465, w_178_1470, w_178_1471, w_178_1473, w_178_1476, w_178_1477, w_178_1478, w_178_1479, w_178_1481, w_178_1486, w_178_1487, w_178_1489, w_178_1491, w_178_1499, w_178_1503, w_178_1504, w_178_1505, w_178_1506, w_178_1508, w_178_1510, w_178_1513, w_178_1517, w_178_1518, w_178_1519, w_178_1520, w_178_1523, w_178_1524, w_178_1528, w_178_1532, w_178_1533, w_178_1534, w_178_1535, w_178_1536, w_178_1539, w_178_1541, w_178_1542, w_178_1543, w_178_1545;
  wire w_179_000, w_179_001, w_179_002, w_179_004, w_179_006, w_179_007, w_179_010, w_179_011, w_179_015, w_179_017, w_179_020, w_179_021, w_179_023, w_179_024, w_179_028, w_179_033, w_179_034, w_179_036, w_179_037, w_179_041, w_179_043, w_179_047, w_179_050, w_179_051, w_179_053, w_179_054, w_179_055, w_179_056, w_179_057, w_179_058, w_179_061, w_179_062, w_179_063, w_179_065, w_179_067, w_179_071, w_179_074, w_179_076, w_179_077, w_179_078, w_179_080, w_179_082, w_179_088, w_179_089, w_179_094, w_179_095, w_179_096, w_179_099, w_179_102, w_179_105, w_179_111, w_179_112, w_179_117, w_179_120, w_179_121, w_179_124, w_179_134, w_179_137, w_179_139, w_179_144, w_179_145, w_179_146, w_179_147, w_179_153, w_179_155, w_179_156, w_179_157, w_179_160, w_179_162, w_179_169, w_179_171, w_179_172, w_179_173, w_179_179, w_179_181, w_179_183, w_179_186, w_179_188, w_179_189, w_179_194, w_179_195, w_179_198, w_179_199, w_179_200, w_179_202, w_179_203, w_179_204, w_179_205, w_179_207, w_179_210, w_179_211, w_179_212, w_179_217, w_179_224, w_179_225, w_179_226, w_179_228, w_179_230, w_179_235, w_179_236, w_179_239, w_179_240, w_179_241, w_179_242, w_179_248, w_179_249, w_179_250, w_179_253, w_179_256, w_179_262, w_179_263, w_179_264, w_179_268, w_179_270, w_179_273, w_179_276, w_179_278, w_179_280, w_179_282, w_179_283, w_179_291, w_179_292, w_179_293, w_179_296, w_179_298, w_179_299, w_179_307, w_179_310, w_179_311, w_179_313, w_179_314, w_179_315, w_179_319, w_179_324, w_179_326, w_179_327, w_179_330, w_179_332, w_179_333, w_179_334, w_179_336, w_179_339, w_179_340, w_179_342, w_179_343, w_179_345, w_179_349, w_179_350, w_179_351, w_179_356, w_179_357, w_179_360, w_179_362, w_179_367, w_179_372, w_179_374, w_179_376, w_179_377, w_179_378, w_179_380, w_179_383, w_179_386, w_179_387, w_179_390, w_179_396, w_179_398, w_179_400, w_179_401, w_179_403, w_179_404, w_179_406, w_179_407, w_179_408, w_179_412, w_179_421, w_179_427, w_179_428, w_179_431, w_179_433, w_179_435, w_179_437, w_179_439, w_179_441, w_179_447, w_179_449, w_179_451, w_179_452, w_179_453, w_179_454, w_179_458, w_179_461, w_179_463, w_179_466, w_179_469, w_179_470, w_179_471, w_179_473, w_179_481, w_179_482, w_179_484, w_179_489, w_179_493, w_179_495, w_179_496, w_179_497, w_179_500, w_179_501, w_179_502, w_179_507, w_179_509, w_179_517, w_179_523, w_179_524, w_179_525, w_179_527, w_179_528, w_179_529, w_179_531, w_179_534, w_179_539, w_179_546, w_179_549, w_179_556, w_179_558, w_179_559, w_179_560, w_179_561, w_179_563, w_179_564, w_179_567, w_179_568, w_179_570, w_179_576, w_179_578, w_179_581, w_179_582, w_179_585, w_179_587, w_179_588, w_179_592, w_179_594, w_179_595, w_179_597, w_179_598, w_179_600, w_179_603, w_179_604, w_179_609, w_179_615, w_179_616, w_179_617, w_179_619, w_179_620, w_179_621, w_179_622, w_179_633, w_179_635, w_179_637, w_179_638, w_179_640, w_179_641, w_179_646, w_179_648, w_179_649, w_179_653, w_179_654, w_179_655, w_179_656, w_179_658, w_179_660, w_179_661, w_179_664, w_179_666, w_179_677, w_179_678, w_179_679, w_179_684, w_179_686, w_179_689, w_179_691, w_179_693, w_179_694, w_179_696, w_179_697, w_179_701, w_179_705, w_179_712, w_179_718, w_179_720, w_179_723, w_179_726, w_179_728, w_179_729, w_179_735, w_179_736, w_179_737, w_179_740, w_179_741, w_179_742, w_179_743, w_179_745, w_179_746, w_179_749, w_179_752, w_179_754, w_179_756, w_179_757, w_179_759, w_179_762, w_179_763, w_179_766, w_179_771, w_179_772, w_179_776, w_179_782, w_179_783, w_179_784, w_179_788, w_179_789, w_179_791, w_179_792, w_179_794, w_179_796, w_179_802, w_179_803, w_179_806, w_179_808, w_179_809, w_179_811, w_179_813, w_179_814, w_179_817, w_179_818, w_179_820, w_179_822, w_179_826, w_179_828, w_179_829, w_179_833, w_179_836, w_179_837, w_179_838, w_179_841, w_179_842, w_179_844, w_179_847, w_179_852, w_179_854, w_179_855, w_179_856, w_179_857, w_179_858, w_179_859, w_179_862, w_179_868, w_179_874, w_179_879, w_179_883, w_179_885, w_179_887, w_179_888, w_179_891, w_179_897, w_179_898, w_179_900, w_179_901, w_179_903, w_179_904, w_179_905, w_179_908, w_179_909, w_179_920, w_179_921, w_179_923, w_179_925, w_179_928, w_179_929, w_179_938, w_179_939, w_179_942, w_179_943, w_179_947, w_179_948, w_179_949, w_179_953, w_179_962, w_179_966, w_179_970, w_179_973, w_179_977, w_179_980, w_179_981, w_179_982, w_179_985, w_179_988, w_179_989, w_179_990, w_179_992, w_179_998, w_179_1000, w_179_1001, w_179_1008, w_179_1012, w_179_1013, w_179_1014, w_179_1016, w_179_1023, w_179_1027, w_179_1028, w_179_1029, w_179_1030, w_179_1033, w_179_1035, w_179_1038, w_179_1039, w_179_1043, w_179_1046, w_179_1048, w_179_1050, w_179_1053, w_179_1056, w_179_1057, w_179_1059, w_179_1063, w_179_1066, w_179_1068, w_179_1072, w_179_1073, w_179_1074, w_179_1081, w_179_1084, w_179_1085, w_179_1089, w_179_1091, w_179_1092, w_179_1097, w_179_1098, w_179_1099, w_179_1106, w_179_1107, w_179_1110, w_179_1132, w_179_1141, w_179_1144, w_179_1148, w_179_1149, w_179_1151, w_179_1160, w_179_1162, w_179_1165, w_179_1167, w_179_1177, w_179_1187, w_179_1188, w_179_1189, w_179_1192, w_179_1197, w_179_1212, w_179_1224, w_179_1228, w_179_1229, w_179_1230, w_179_1234, w_179_1239, w_179_1243, w_179_1247, w_179_1253, w_179_1256, w_179_1259, w_179_1262, w_179_1265, w_179_1266, w_179_1268, w_179_1269, w_179_1270, w_179_1274, w_179_1275, w_179_1281, w_179_1286, w_179_1289, w_179_1295, w_179_1296, w_179_1302, w_179_1303, w_179_1304, w_179_1320, w_179_1323, w_179_1325, w_179_1332, w_179_1334, w_179_1340, w_179_1343, w_179_1346, w_179_1347, w_179_1355, w_179_1357, w_179_1362, w_179_1366, w_179_1367, w_179_1368, w_179_1370, w_179_1373, w_179_1375, w_179_1376, w_179_1379, w_179_1380, w_179_1381, w_179_1388, w_179_1389, w_179_1390, w_179_1401, w_179_1404, w_179_1409, w_179_1422, w_179_1423, w_179_1424, w_179_1431, w_179_1434, w_179_1440, w_179_1449, w_179_1452, w_179_1455, w_179_1460, w_179_1465, w_179_1472, w_179_1473, w_179_1483, w_179_1496, w_179_1502, w_179_1509, w_179_1513, w_179_1522, w_179_1525, w_179_1526, w_179_1528, w_179_1530, w_179_1533, w_179_1534, w_179_1536, w_179_1537, w_179_1543, w_179_1545, w_179_1546, w_179_1547, w_179_1549, w_179_1553, w_179_1554, w_179_1557, w_179_1559, w_179_1562, w_179_1564, w_179_1565, w_179_1569, w_179_1583, w_179_1585, w_179_1588, w_179_1590, w_179_1591, w_179_1594, w_179_1596, w_179_1597, w_179_1598, w_179_1599, w_179_1600, w_179_1607, w_179_1614, w_179_1615, w_179_1617, w_179_1618, w_179_1619, w_179_1625, w_179_1627, w_179_1629, w_179_1632, w_179_1638, w_179_1641, w_179_1645, w_179_1647, w_179_1649, w_179_1654, w_179_1656, w_179_1658, w_179_1667, w_179_1670, w_179_1675, w_179_1681, w_179_1688, w_179_1689, w_179_1692, w_179_1695, w_179_1697, w_179_1698, w_179_1701, w_179_1702, w_179_1705, w_179_1711, w_179_1715, w_179_1718, w_179_1719, w_179_1726, w_179_1729, w_179_1730, w_179_1732, w_179_1738, w_179_1743, w_179_1746, w_179_1747, w_179_1748, w_179_1749, w_179_1752, w_179_1753, w_179_1760, w_179_1763, w_179_1769, w_179_1773, w_179_1774, w_179_1778, w_179_1788, w_179_1789, w_179_1791, w_179_1796, w_179_1799, w_179_1801, w_179_1804, w_179_1807, w_179_1808, w_179_1810, w_179_1812, w_179_1816, w_179_1817, w_179_1818, w_179_1819, w_179_1821, w_179_1826, w_179_1829, w_179_1834, w_179_1836, w_179_1838, w_179_1839, w_179_1846, w_179_1848, w_179_1850, w_179_1851, w_179_1852, w_179_1858, w_179_1864, w_179_1865, w_179_1866, w_179_1870, w_179_1872, w_179_1873, w_179_1881, w_179_1886, w_179_1888, w_179_1889, w_179_1892, w_179_1893, w_179_1894, w_179_1895, w_179_1896, w_179_1899, w_179_1900, w_179_1907, w_179_1908, w_179_1909, w_179_1910, w_179_1916, w_179_1925, w_179_1927, w_179_1933, w_179_1940, w_179_1943, w_179_1945, w_179_1947, w_179_1948, w_179_1949, w_179_1950, w_179_1951, w_179_1952, w_179_1954;
  wire w_180_002, w_180_003, w_180_004, w_180_006, w_180_008, w_180_009, w_180_010, w_180_011, w_180_012, w_180_013, w_180_014, w_180_015, w_180_016, w_180_018, w_180_021, w_180_024, w_180_026, w_180_028, w_180_030, w_180_036, w_180_037, w_180_041, w_180_043, w_180_052, w_180_054, w_180_055, w_180_058, w_180_059, w_180_060, w_180_061, w_180_063, w_180_067, w_180_068, w_180_070, w_180_072, w_180_073, w_180_074, w_180_075, w_180_079, w_180_080, w_180_082, w_180_083, w_180_086, w_180_087, w_180_089, w_180_090, w_180_094, w_180_095, w_180_096, w_180_097, w_180_098, w_180_100, w_180_103, w_180_104, w_180_105, w_180_106, w_180_107, w_180_109, w_180_112, w_180_113, w_180_115, w_180_118, w_180_121, w_180_124, w_180_125, w_180_126, w_180_128, w_180_131, w_180_132, w_180_133, w_180_134, w_180_135, w_180_136, w_180_137, w_180_138, w_180_139, w_180_140, w_180_141, w_180_147, w_180_148, w_180_151, w_180_152, w_180_153, w_180_155, w_180_157, w_180_158, w_180_159, w_180_160, w_180_163, w_180_164, w_180_168, w_180_170, w_180_171, w_180_173, w_180_176, w_180_180, w_180_181, w_180_182, w_180_185, w_180_186, w_180_191, w_180_195, w_180_196, w_180_198, w_180_199, w_180_200, w_180_201, w_180_205, w_180_207, w_180_208, w_180_213, w_180_215, w_180_217, w_180_218, w_180_222, w_180_224, w_180_225, w_180_229, w_180_230, w_180_231, w_180_232, w_180_233, w_180_234, w_180_235, w_180_236, w_180_237, w_180_238, w_180_239, w_180_240, w_180_241, w_180_242, w_180_244, w_180_245, w_180_246, w_180_248, w_180_251, w_180_252, w_180_254, w_180_255, w_180_257, w_180_258, w_180_263, w_180_264, w_180_265, w_180_267, w_180_271, w_180_273, w_180_275, w_180_276, w_180_278, w_180_279, w_180_282, w_180_287, w_180_289, w_180_291, w_180_293, w_180_294, w_180_295, w_180_297, w_180_299, w_180_301, w_180_302, w_180_304, w_180_305, w_180_306, w_180_307, w_180_309, w_180_310, w_180_314, w_180_319, w_180_321, w_180_322, w_180_324, w_180_326, w_180_331, w_180_332, w_180_333, w_180_334, w_180_335, w_180_337, w_180_340, w_180_342, w_180_343, w_180_352, w_180_354, w_180_355, w_180_356, w_180_357, w_180_358, w_180_360, w_180_361, w_180_362, w_180_367, w_180_369, w_180_371, w_180_374, w_180_378, w_180_381, w_180_382, w_180_383, w_180_385, w_180_388, w_180_391, w_180_392, w_180_395, w_180_397, w_180_400, w_180_401, w_180_402, w_180_403, w_180_404, w_180_406, w_180_407, w_180_408, w_180_413, w_180_414, w_180_417, w_180_420, w_180_421, w_180_422, w_180_423, w_180_430, w_180_431, w_180_433, w_180_440, w_180_442, w_180_443, w_180_446, w_180_450, w_180_452, w_180_455, w_180_456, w_180_458, w_180_459, w_180_461, w_180_466, w_180_469, w_180_471, w_180_474, w_180_475, w_180_478, w_180_479, w_180_481, w_180_482, w_180_485, w_180_486, w_180_487, w_180_488, w_180_491, w_180_493, w_180_495, w_180_496, w_180_497, w_180_499, w_180_500, w_180_502, w_180_503, w_180_505, w_180_506, w_180_507, w_180_508, w_180_510, w_180_513, w_180_515, w_180_520, w_180_524, w_180_525, w_180_526, w_180_527, w_180_533, w_180_534, w_180_537, w_180_538, w_180_539, w_180_540, w_180_541, w_180_543, w_180_550, w_180_560, w_180_561, w_180_564, w_180_565, w_180_566, w_180_567, w_180_569, w_180_572, w_180_573, w_180_575, w_180_576, w_180_579, w_180_584, w_180_588, w_180_593, w_180_594, w_180_595, w_180_598, w_180_604, w_180_606, w_180_607, w_180_608, w_180_609, w_180_610, w_180_613, w_180_619, w_180_625, w_180_627, w_180_630, w_180_631, w_180_633, w_180_635, w_180_642, w_180_644, w_180_646, w_180_647, w_180_651, w_180_655, w_180_657, w_180_658, w_180_660, w_180_662, w_180_667, w_180_669, w_180_672, w_180_673, w_180_677, w_180_679, w_180_683, w_180_684, w_180_685, w_180_687, w_180_688, w_180_689, w_180_690, w_180_691, w_180_693, w_180_694, w_180_695, w_180_697, w_180_698, w_180_699, w_180_700, w_180_703, w_180_705, w_180_707, w_180_709, w_180_712, w_180_713, w_180_715, w_180_717, w_180_719, w_180_721, w_180_722, w_180_723, w_180_725, w_180_727, w_180_728, w_180_731, w_180_735, w_180_736, w_180_737, w_180_742, w_180_743, w_180_744, w_180_745, w_180_747, w_180_748, w_180_749, w_180_750, w_180_751, w_180_752, w_180_753, w_180_754, w_180_755, w_180_760, w_180_761, w_180_762, w_180_766, w_180_767, w_180_769, w_180_770, w_180_775, w_180_776, w_180_780, w_180_783, w_180_784, w_180_789, w_180_796, w_180_800, w_180_802, w_180_808, w_180_811, w_180_813, w_180_814, w_180_815, w_180_816, w_180_819, w_180_820, w_180_821, w_180_822, w_180_823, w_180_826, w_180_828, w_180_834, w_180_835, w_180_838, w_180_839, w_180_844, w_180_845, w_180_846, w_180_849, w_180_850, w_180_853, w_180_854, w_180_857, w_180_859, w_180_863, w_180_867, w_180_868, w_180_873, w_180_877, w_180_880, w_180_882, w_180_884, w_180_885, w_180_889, w_180_890, w_180_893, w_180_894, w_180_895, w_180_898, w_180_899, w_180_902, w_180_904, w_180_905, w_180_909, w_180_912, w_180_913, w_180_916, w_180_917, w_180_920, w_180_922, w_180_923, w_180_925, w_180_928, w_180_930, w_180_943, w_180_946, w_180_947, w_180_950, w_180_952, w_180_954, w_180_963, w_180_965, w_180_968, w_180_973, w_180_974, w_180_976, w_180_979, w_180_981, w_180_983, w_180_985, w_180_986, w_180_989, w_180_991, w_180_997, w_180_1002, w_180_1004, w_180_1006, w_180_1008, w_180_1011, w_180_1013, w_180_1014, w_180_1015, w_180_1018, w_180_1019, w_180_1021, w_180_1022, w_180_1029, w_180_1034, w_180_1035, w_180_1038, w_180_1042, w_180_1046, w_180_1048, w_180_1052, w_180_1056, w_180_1062, w_180_1064, w_180_1068, w_180_1072, w_180_1075, w_180_1076, w_180_1080, w_180_1082, w_180_1083, w_180_1084, w_180_1088, w_180_1090, w_180_1092, w_180_1095, w_180_1098, w_180_1106, w_180_1108, w_180_1109, w_180_1113, w_180_1114, w_180_1115, w_180_1117, w_180_1122, w_180_1126, w_180_1130, w_180_1132, w_180_1135, w_180_1140, w_180_1141, w_180_1142, w_180_1147, w_180_1149, w_180_1159, w_180_1163, w_180_1170, w_180_1172, w_180_1174, w_180_1176, w_180_1178, w_180_1187, w_180_1192, w_180_1194, w_180_1196, w_180_1197, w_180_1201, w_180_1204, w_180_1205, w_180_1206, w_180_1208, w_180_1210, w_180_1215, w_180_1224, w_180_1231, w_180_1232, w_180_1242, w_180_1248, w_180_1252, w_180_1257, w_180_1259, w_180_1262, w_180_1273, w_180_1274, w_180_1277, w_180_1282, w_180_1283, w_180_1286, w_180_1289, w_180_1291, w_180_1296, w_180_1299, w_180_1302, w_180_1307, w_180_1308, w_180_1310, w_180_1315, w_180_1317, w_180_1323, w_180_1324, w_180_1325, w_180_1326, w_180_1327, w_180_1336, w_180_1341, w_180_1346, w_180_1350, w_180_1352, w_180_1353, w_180_1356, w_180_1360, w_180_1364, w_180_1365, w_180_1368, w_180_1369, w_180_1371, w_180_1372, w_180_1373, w_180_1374, w_180_1375, w_180_1376, w_180_1377, w_180_1378, w_180_1379, w_180_1383, w_180_1384, w_180_1385, w_180_1386, w_180_1387, w_180_1388, w_180_1389, w_180_1390, w_180_1391, w_180_1392, w_180_1393, w_180_1395;
  wire w_181_000, w_181_002, w_181_004, w_181_005, w_181_006, w_181_007, w_181_009, w_181_011, w_181_012, w_181_013, w_181_015, w_181_016, w_181_018, w_181_019, w_181_022, w_181_023, w_181_024, w_181_027, w_181_030, w_181_031, w_181_032, w_181_034, w_181_036, w_181_038, w_181_040, w_181_043, w_181_047, w_181_048, w_181_052, w_181_055, w_181_057, w_181_058, w_181_060, w_181_061, w_181_062, w_181_063, w_181_066, w_181_067, w_181_069, w_181_074, w_181_077, w_181_078, w_181_079, w_181_080, w_181_084, w_181_087, w_181_089, w_181_091, w_181_094, w_181_096, w_181_099, w_181_103, w_181_107, w_181_109, w_181_110, w_181_112, w_181_117, w_181_118, w_181_121, w_181_124, w_181_125, w_181_126, w_181_127, w_181_129, w_181_133, w_181_135, w_181_136, w_181_137, w_181_139, w_181_140, w_181_141, w_181_144, w_181_147, w_181_148, w_181_150, w_181_151, w_181_153, w_181_157, w_181_160, w_181_162, w_181_164, w_181_166, w_181_167, w_181_172, w_181_173, w_181_174, w_181_176, w_181_177, w_181_178, w_181_180, w_181_182, w_181_183, w_181_184, w_181_185, w_181_187, w_181_190, w_181_191, w_181_192, w_181_196, w_181_197, w_181_199, w_181_202, w_181_204, w_181_213, w_181_214, w_181_217, w_181_221, w_181_223, w_181_224, w_181_226, w_181_227, w_181_228, w_181_229, w_181_230, w_181_234, w_181_235, w_181_236, w_181_237, w_181_244, w_181_245, w_181_250, w_181_253, w_181_254, w_181_256, w_181_257, w_181_258, w_181_262, w_181_263, w_181_264, w_181_265, w_181_266, w_181_267, w_181_269, w_181_271, w_181_273, w_181_277, w_181_278, w_181_279, w_181_280, w_181_281, w_181_283, w_181_287, w_181_288, w_181_290, w_181_291, w_181_294, w_181_295, w_181_299, w_181_300, w_181_301, w_181_302, w_181_305, w_181_306, w_181_314, w_181_322, w_181_325, w_181_327, w_181_329, w_181_330, w_181_335, w_181_336, w_181_341, w_181_346, w_181_347, w_181_348, w_181_349, w_181_350, w_181_351, w_181_353, w_181_354, w_181_357, w_181_360, w_181_362, w_181_364, w_181_365, w_181_369, w_181_371, w_181_373, w_181_374, w_181_375, w_181_376, w_181_377, w_181_380, w_181_382, w_181_383, w_181_384, w_181_385, w_181_386, w_181_387, w_181_389, w_181_391, w_181_392, w_181_393, w_181_394, w_181_397, w_181_403, w_181_404, w_181_406, w_181_409, w_181_410, w_181_413, w_181_417, w_181_418, w_181_419, w_181_420, w_181_429, w_181_433, w_181_437, w_181_438, w_181_439, w_181_441, w_181_443, w_181_444, w_181_447, w_181_448, w_181_449, w_181_456, w_181_457, w_181_459, w_181_460, w_181_462, w_181_466, w_181_468, w_181_469, w_181_471, w_181_476, w_181_477, w_181_478, w_181_479, w_181_482, w_181_483, w_181_486, w_181_487, w_181_491, w_181_494, w_181_496, w_181_497, w_181_500, w_181_501, w_181_502, w_181_505, w_181_508, w_181_519, w_181_520, w_181_521, w_181_522, w_181_525, w_181_527, w_181_528, w_181_529, w_181_530, w_181_531, w_181_542, w_181_543, w_181_544, w_181_546, w_181_549, w_181_551, w_181_554, w_181_556, w_181_563, w_181_565, w_181_566, w_181_567, w_181_569, w_181_570, w_181_571, w_181_576, w_181_578, w_181_579, w_181_588, w_181_589, w_181_590, w_181_591, w_181_592, w_181_593, w_181_594, w_181_595, w_181_597, w_181_598, w_181_599, w_181_600, w_181_602, w_181_604, w_181_607, w_181_608, w_181_610, w_181_611, w_181_615, w_181_616, w_181_617, w_181_621, w_181_623, w_181_625, w_181_626, w_181_629, w_181_631, w_181_632, w_181_633, w_181_635, w_181_636, w_181_638, w_181_645, w_181_647, w_181_648, w_181_649, w_181_650, w_181_652, w_181_660, w_181_668, w_181_669, w_181_670, w_181_671, w_181_672, w_181_673, w_181_674, w_181_675, w_181_677, w_181_678, w_181_681, w_181_683, w_181_685, w_181_686, w_181_690, w_181_693, w_181_698, w_181_704, w_181_707, w_181_708, w_181_710, w_181_713, w_181_714, w_181_718, w_181_719, w_181_720, w_181_722, w_181_723, w_181_727, w_181_730, w_181_731, w_181_734, w_181_736, w_181_737, w_181_740, w_181_741, w_181_743, w_181_745, w_181_746, w_181_755, w_181_756, w_181_758, w_181_759, w_181_760, w_181_761, w_181_762, w_181_763, w_181_764, w_181_766, w_181_767, w_181_774, w_181_775, w_181_776, w_181_778, w_181_779, w_181_780, w_181_782, w_181_784, w_181_791, w_181_794, w_181_796, w_181_798, w_181_800, w_181_803, w_181_813, w_181_817, w_181_818, w_181_819, w_181_820, w_181_821, w_181_823, w_181_824, w_181_825, w_181_826, w_181_828, w_181_831, w_181_832, w_181_833, w_181_834, w_181_835, w_181_836, w_181_837, w_181_838, w_181_839, w_181_840, w_181_841, w_181_842, w_181_843, w_181_844, w_181_845, w_181_846, w_181_847, w_181_848, w_181_849, w_181_852, w_181_853, w_181_856, w_181_863, w_181_864, w_181_866, w_181_868, w_181_869, w_181_871, w_181_872, w_181_873, w_181_877, w_181_878, w_181_879, w_181_881, w_181_882, w_181_883, w_181_884, w_181_886, w_181_887, w_181_889, w_181_891, w_181_892, w_181_893, w_181_898, w_181_900, w_181_905, w_181_906, w_181_910, w_181_911, w_181_912, w_181_913, w_181_917, w_181_920, w_181_921, w_181_924, w_181_927, w_181_929, w_181_930, w_181_931, w_181_936, w_181_937, w_181_938, w_181_940, w_181_942, w_181_943, w_181_944, w_181_945, w_181_946, w_181_947, w_181_948, w_181_949, w_181_950, w_181_951, w_181_955, w_181_956, w_181_957, w_181_958, w_181_960, w_181_963, w_181_964, w_181_965, w_181_966, w_181_967, w_181_968, w_181_971, w_181_972, w_181_973, w_181_977, w_181_978, w_181_980, w_181_981, w_181_982, w_181_983, w_181_985, w_181_986, w_181_989, w_181_990, w_181_992, w_181_993, w_181_994, w_181_1000, w_181_1002, w_181_1006, w_181_1007, w_181_1008, w_181_1012, w_181_1014, w_181_1016, w_181_1019, w_181_1020, w_181_1021, w_181_1022, w_181_1025, w_181_1026, w_181_1027, w_181_1029, w_181_1030, w_181_1032, w_181_1033, w_181_1034, w_181_1035, w_181_1037, w_181_1038, w_181_1041, w_181_1047, w_181_1057, w_181_1061, w_181_1062, w_181_1066, w_181_1067, w_181_1068, w_181_1070, w_181_1071, w_181_1079, w_181_1083, w_181_1084, w_181_1087, w_181_1090, w_181_1091, w_181_1097, w_181_1101, w_181_1103, w_181_1106, w_181_1108, w_181_1109, w_181_1110, w_181_1111, w_181_1112, w_181_1113, w_181_1114, w_181_1118, w_181_1119, w_181_1121, w_181_1125, w_181_1127, w_181_1128, w_181_1135, w_181_1136, w_181_1137, w_181_1139, w_181_1141, w_181_1146, w_181_1152, w_181_1154, w_181_1156, w_181_1159, w_181_1168, w_181_1169, w_181_1171, w_181_1174, w_181_1175, w_181_1177, w_181_1181, w_181_1182, w_181_1187, w_181_1194, w_181_1196, w_181_1197, w_181_1198;
  wire w_182_000, w_182_003, w_182_005, w_182_008, w_182_010, w_182_011, w_182_013, w_182_018, w_182_021, w_182_024, w_182_025, w_182_026, w_182_028, w_182_030, w_182_031, w_182_033, w_182_035, w_182_039, w_182_040, w_182_043, w_182_045, w_182_047, w_182_048, w_182_050, w_182_051, w_182_055, w_182_059, w_182_061, w_182_063, w_182_064, w_182_066, w_182_068, w_182_071, w_182_072, w_182_077, w_182_078, w_182_087, w_182_088, w_182_090, w_182_098, w_182_099, w_182_105, w_182_106, w_182_110, w_182_112, w_182_113, w_182_114, w_182_117, w_182_124, w_182_126, w_182_129, w_182_130, w_182_134, w_182_135, w_182_136, w_182_141, w_182_147, w_182_149, w_182_150, w_182_153, w_182_155, w_182_156, w_182_159, w_182_161, w_182_162, w_182_163, w_182_164, w_182_166, w_182_167, w_182_170, w_182_175, w_182_176, w_182_179, w_182_182, w_182_184, w_182_187, w_182_191, w_182_196, w_182_198, w_182_199, w_182_202, w_182_205, w_182_206, w_182_209, w_182_211, w_182_212, w_182_213, w_182_216, w_182_218, w_182_219, w_182_222, w_182_224, w_182_226, w_182_227, w_182_230, w_182_242, w_182_244, w_182_245, w_182_248, w_182_251, w_182_256, w_182_258, w_182_263, w_182_266, w_182_267, w_182_268, w_182_275, w_182_278, w_182_285, w_182_286, w_182_287, w_182_288, w_182_289, w_182_290, w_182_295, w_182_296, w_182_297, w_182_299, w_182_301, w_182_307, w_182_313, w_182_320, w_182_323, w_182_326, w_182_334, w_182_337, w_182_340, w_182_346, w_182_348, w_182_350, w_182_353, w_182_356, w_182_361, w_182_367, w_182_369, w_182_371, w_182_374, w_182_375, w_182_377, w_182_380, w_182_382, w_182_383, w_182_386, w_182_387, w_182_389, w_182_397, w_182_398, w_182_406, w_182_409, w_182_414, w_182_416, w_182_418, w_182_421, w_182_422, w_182_423, w_182_424, w_182_426, w_182_428, w_182_434, w_182_436, w_182_438, w_182_439, w_182_442, w_182_443, w_182_445, w_182_446, w_182_458, w_182_460, w_182_464, w_182_465, w_182_468, w_182_469, w_182_471, w_182_474, w_182_476, w_182_478, w_182_482, w_182_484, w_182_489, w_182_490, w_182_491, w_182_492, w_182_494, w_182_500, w_182_501, w_182_503, w_182_506, w_182_509, w_182_510, w_182_514, w_182_516, w_182_517, w_182_518, w_182_520, w_182_521, w_182_525, w_182_533, w_182_541, w_182_543, w_182_545, w_182_548, w_182_550, w_182_554, w_182_555, w_182_556, w_182_557, w_182_558, w_182_566, w_182_567, w_182_568, w_182_571, w_182_574, w_182_575, w_182_576, w_182_578, w_182_581, w_182_582, w_182_585, w_182_587, w_182_588, w_182_594, w_182_599, w_182_600, w_182_602, w_182_605, w_182_606, w_182_607, w_182_611, w_182_613, w_182_616, w_182_629, w_182_630, w_182_634, w_182_635, w_182_638, w_182_640, w_182_642, w_182_644, w_182_646, w_182_649, w_182_653, w_182_656, w_182_657, w_182_658, w_182_664, w_182_667, w_182_670, w_182_671, w_182_675, w_182_678, w_182_679, w_182_680, w_182_682, w_182_691, w_182_693, w_182_696, w_182_697, w_182_700, w_182_703, w_182_706, w_182_709, w_182_712, w_182_716, w_182_718, w_182_721, w_182_727, w_182_732, w_182_735, w_182_738, w_182_740, w_182_741, w_182_743, w_182_746, w_182_748, w_182_749, w_182_750, w_182_754, w_182_755, w_182_757, w_182_763, w_182_767, w_182_768, w_182_769, w_182_772, w_182_773, w_182_776, w_182_778, w_182_782, w_182_783, w_182_786, w_182_787, w_182_789, w_182_792, w_182_793, w_182_797, w_182_799, w_182_801, w_182_803, w_182_806, w_182_808, w_182_810, w_182_811, w_182_814, w_182_815, w_182_817, w_182_820, w_182_822, w_182_823, w_182_827, w_182_831, w_182_833, w_182_837, w_182_840, w_182_843, w_182_845, w_182_846, w_182_847, w_182_848, w_182_850, w_182_853, w_182_855, w_182_858, w_182_859, w_182_860, w_182_865, w_182_866, w_182_869, w_182_870, w_182_872, w_182_875, w_182_877, w_182_879, w_182_886, w_182_891, w_182_894, w_182_897, w_182_898, w_182_900, w_182_901, w_182_902, w_182_903, w_182_913, w_182_914, w_182_916, w_182_918, w_182_919, w_182_920, w_182_921, w_182_922, w_182_930, w_182_934, w_182_935, w_182_938, w_182_939, w_182_940, w_182_941, w_182_943, w_182_944, w_182_946, w_182_954, w_182_955, w_182_956, w_182_958, w_182_960, w_182_962, w_182_963, w_182_969, w_182_970, w_182_972, w_182_973, w_182_974, w_182_976, w_182_977, w_182_980, w_182_981, w_182_986, w_182_989, w_182_993, w_182_995, w_182_997, w_182_998, w_182_999, w_182_1000, w_182_1004, w_182_1006, w_182_1009, w_182_1012, w_182_1014, w_182_1018, w_182_1021, w_182_1023, w_182_1024, w_182_1025, w_182_1026, w_182_1028, w_182_1031, w_182_1033, w_182_1034, w_182_1037, w_182_1038, w_182_1039, w_182_1040, w_182_1043, w_182_1046, w_182_1051, w_182_1052, w_182_1055, w_182_1056, w_182_1058, w_182_1060, w_182_1061, w_182_1062, w_182_1068, w_182_1070, w_182_1071, w_182_1073, w_182_1075, w_182_1076, w_182_1077, w_182_1082, w_182_1088, w_182_1090, w_182_1091, w_182_1096, w_182_1097, w_182_1101, w_182_1105, w_182_1106, w_182_1107, w_182_1108, w_182_1109, w_182_1112, w_182_1114, w_182_1116, w_182_1119, w_182_1120, w_182_1129, w_182_1136, w_182_1137, w_182_1141, w_182_1142, w_182_1144, w_182_1145, w_182_1148, w_182_1149, w_182_1150, w_182_1152, w_182_1154, w_182_1161, w_182_1162, w_182_1164, w_182_1165, w_182_1166, w_182_1180, w_182_1182, w_182_1184, w_182_1185, w_182_1186, w_182_1189, w_182_1197, w_182_1203, w_182_1206, w_182_1207, w_182_1208, w_182_1209, w_182_1210, w_182_1213, w_182_1214, w_182_1220, w_182_1226, w_182_1235, w_182_1236, w_182_1247, w_182_1250, w_182_1251, w_182_1253, w_182_1260, w_182_1261, w_182_1264, w_182_1270, w_182_1275, w_182_1276, w_182_1281, w_182_1282, w_182_1285, w_182_1291, w_182_1295, w_182_1297, w_182_1300, w_182_1301, w_182_1302, w_182_1303, w_182_1304, w_182_1305, w_182_1306, w_182_1309, w_182_1312, w_182_1316, w_182_1319, w_182_1323, w_182_1328, w_182_1333, w_182_1335, w_182_1336, w_182_1338, w_182_1339, w_182_1340, w_182_1341, w_182_1344, w_182_1347, w_182_1349, w_182_1353, w_182_1354, w_182_1362, w_182_1363, w_182_1369, w_182_1372, w_182_1373, w_182_1376, w_182_1379, w_182_1382, w_182_1384, w_182_1387, w_182_1390, w_182_1391, w_182_1397, w_182_1398, w_182_1400, w_182_1402, w_182_1406, w_182_1407, w_182_1410, w_182_1415, w_182_1416, w_182_1418, w_182_1428, w_182_1431, w_182_1432, w_182_1438, w_182_1440, w_182_1456, w_182_1459, w_182_1463, w_182_1464, w_182_1466, w_182_1470, w_182_1473, w_182_1478, w_182_1480, w_182_1482, w_182_1483, w_182_1486, w_182_1488, w_182_1492, w_182_1493, w_182_1494, w_182_1495, w_182_1496, w_182_1497, w_182_1498, w_182_1500, w_182_1503, w_182_1505, w_182_1506, w_182_1507, w_182_1508, w_182_1511, w_182_1515, w_182_1518, w_182_1521, w_182_1522, w_182_1524, w_182_1526, w_182_1528, w_182_1533, w_182_1534, w_182_1536, w_182_1537, w_182_1539, w_182_1540, w_182_1542, w_182_1545, w_182_1547, w_182_1548, w_182_1549, w_182_1550, w_182_1556, w_182_1558, w_182_1561, w_182_1568, w_182_1571, w_182_1576, w_182_1577, w_182_1578, w_182_1579, w_182_1583, w_182_1590, w_182_1593, w_182_1594, w_182_1599, w_182_1603, w_182_1604, w_182_1607, w_182_1610, w_182_1611, w_182_1618, w_182_1619, w_182_1620, w_182_1621, w_182_1622, w_182_1623, w_182_1624, w_182_1625, w_182_1626, w_182_1628;
  wire w_183_000, w_183_003, w_183_005, w_183_008, w_183_009, w_183_013, w_183_019, w_183_021, w_183_022, w_183_026, w_183_027, w_183_029, w_183_031, w_183_032, w_183_036, w_183_037, w_183_042, w_183_043, w_183_045, w_183_049, w_183_050, w_183_052, w_183_053, w_183_054, w_183_055, w_183_064, w_183_067, w_183_069, w_183_070, w_183_071, w_183_072, w_183_079, w_183_081, w_183_085, w_183_090, w_183_093, w_183_095, w_183_096, w_183_097, w_183_101, w_183_102, w_183_104, w_183_107, w_183_117, w_183_119, w_183_121, w_183_122, w_183_126, w_183_127, w_183_129, w_183_130, w_183_141, w_183_142, w_183_146, w_183_156, w_183_158, w_183_159, w_183_165, w_183_169, w_183_173, w_183_180, w_183_183, w_183_184, w_183_187, w_183_189, w_183_190, w_183_193, w_183_197, w_183_198, w_183_200, w_183_206, w_183_207, w_183_210, w_183_215, w_183_218, w_183_220, w_183_225, w_183_226, w_183_231, w_183_232, w_183_236, w_183_241, w_183_242, w_183_243, w_183_245, w_183_249, w_183_251, w_183_252, w_183_255, w_183_256, w_183_260, w_183_262, w_183_263, w_183_264, w_183_266, w_183_269, w_183_272, w_183_274, w_183_276, w_183_277, w_183_278, w_183_283, w_183_289, w_183_290, w_183_292, w_183_299, w_183_300, w_183_314, w_183_328, w_183_329, w_183_330, w_183_331, w_183_334, w_183_335, w_183_338, w_183_341, w_183_345, w_183_348, w_183_349, w_183_353, w_183_355, w_183_357, w_183_358, w_183_362, w_183_363, w_183_367, w_183_369, w_183_371, w_183_373, w_183_374, w_183_376, w_183_384, w_183_390, w_183_391, w_183_393, w_183_394, w_183_395, w_183_396, w_183_401, w_183_402, w_183_403, w_183_407, w_183_408, w_183_409, w_183_410, w_183_411, w_183_412, w_183_414, w_183_417, w_183_418, w_183_419, w_183_421, w_183_422, w_183_424, w_183_425, w_183_426, w_183_427, w_183_428, w_183_429, w_183_430, w_183_431, w_183_436, w_183_437, w_183_442, w_183_443, w_183_444, w_183_445, w_183_446, w_183_447, w_183_448, w_183_453, w_183_456, w_183_458, w_183_461, w_183_462, w_183_463, w_183_464, w_183_468, w_183_470, w_183_471, w_183_473, w_183_476, w_183_479, w_183_480, w_183_483, w_183_485, w_183_486, w_183_488, w_183_490, w_183_495, w_183_496, w_183_505, w_183_508, w_183_511, w_183_512, w_183_521, w_183_526, w_183_533, w_183_535, w_183_537, w_183_540, w_183_546, w_183_548, w_183_550, w_183_557, w_183_560, w_183_565, w_183_575, w_183_579, w_183_580, w_183_585, w_183_590, w_183_591, w_183_593, w_183_595, w_183_597, w_183_604, w_183_605, w_183_608, w_183_609, w_183_619, w_183_620, w_183_621, w_183_623, w_183_626, w_183_628, w_183_629, w_183_637, w_183_640, w_183_646, w_183_651, w_183_652, w_183_656, w_183_658, w_183_660, w_183_662, w_183_665, w_183_666, w_183_667, w_183_671, w_183_674, w_183_675, w_183_678, w_183_680, w_183_681, w_183_684, w_183_685, w_183_690, w_183_691, w_183_693, w_183_694, w_183_696, w_183_697, w_183_698, w_183_699, w_183_701, w_183_702, w_183_710, w_183_712, w_183_713, w_183_714, w_183_716, w_183_717, w_183_720, w_183_721, w_183_727, w_183_729, w_183_731, w_183_733, w_183_748, w_183_752, w_183_759, w_183_763, w_183_764, w_183_771, w_183_776, w_183_777, w_183_778, w_183_782, w_183_788, w_183_799, w_183_811, w_183_818, w_183_822, w_183_825, w_183_828, w_183_830, w_183_837, w_183_838, w_183_839, w_183_840, w_183_846, w_183_847, w_183_848, w_183_850, w_183_854, w_183_855, w_183_856, w_183_857, w_183_858, w_183_860, w_183_862, w_183_863, w_183_866, w_183_869, w_183_870, w_183_873, w_183_877, w_183_879, w_183_883, w_183_886, w_183_889, w_183_891, w_183_896, w_183_901, w_183_902, w_183_921, w_183_925, w_183_928, w_183_930, w_183_931, w_183_936, w_183_937, w_183_939, w_183_941, w_183_947, w_183_948, w_183_960, w_183_963, w_183_965, w_183_966, w_183_967, w_183_969, w_183_974, w_183_975, w_183_979, w_183_984, w_183_986, w_183_992, w_183_993, w_183_996, w_183_997, w_183_998, w_183_1004, w_183_1006, w_183_1011, w_183_1016, w_183_1022, w_183_1033, w_183_1038, w_183_1045, w_183_1046, w_183_1053, w_183_1055, w_183_1056, w_183_1058, w_183_1059, w_183_1061, w_183_1065, w_183_1067, w_183_1068, w_183_1071, w_183_1072, w_183_1078, w_183_1079, w_183_1084, w_183_1089, w_183_1098, w_183_1099, w_183_1103, w_183_1104, w_183_1110, w_183_1114, w_183_1119, w_183_1120, w_183_1123, w_183_1125, w_183_1133, w_183_1138, w_183_1139, w_183_1140, w_183_1141, w_183_1146, w_183_1149, w_183_1154, w_183_1155, w_183_1159, w_183_1165, w_183_1173, w_183_1176, w_183_1181, w_183_1188, w_183_1189, w_183_1191, w_183_1195, w_183_1202, w_183_1205, w_183_1206, w_183_1216, w_183_1221, w_183_1230, w_183_1233, w_183_1237, w_183_1239, w_183_1240, w_183_1241, w_183_1250, w_183_1252, w_183_1253, w_183_1254, w_183_1258, w_183_1265, w_183_1268, w_183_1269, w_183_1281, w_183_1284, w_183_1285, w_183_1288, w_183_1289, w_183_1291, w_183_1298, w_183_1301, w_183_1303, w_183_1305, w_183_1309, w_183_1311, w_183_1312, w_183_1315, w_183_1317, w_183_1323, w_183_1325, w_183_1330, w_183_1331, w_183_1333, w_183_1337, w_183_1341, w_183_1342, w_183_1354, w_183_1358, w_183_1359, w_183_1372, w_183_1378, w_183_1381, w_183_1382, w_183_1396, w_183_1401, w_183_1403, w_183_1408, w_183_1410, w_183_1411, w_183_1412, w_183_1413, w_183_1420, w_183_1422, w_183_1424, w_183_1425, w_183_1431, w_183_1433, w_183_1438, w_183_1441, w_183_1444, w_183_1447, w_183_1448, w_183_1450, w_183_1452, w_183_1455, w_183_1459, w_183_1461, w_183_1462, w_183_1464, w_183_1466, w_183_1472, w_183_1478, w_183_1482, w_183_1486, w_183_1492, w_183_1494, w_183_1496, w_183_1497, w_183_1506, w_183_1509, w_183_1511, w_183_1517, w_183_1521, w_183_1522, w_183_1524, w_183_1525, w_183_1528, w_183_1529, w_183_1531, w_183_1535, w_183_1536, w_183_1537, w_183_1538, w_183_1547, w_183_1552, w_183_1554, w_183_1560, w_183_1561, w_183_1568, w_183_1574, w_183_1577, w_183_1580, w_183_1582, w_183_1583, w_183_1584, w_183_1585, w_183_1589, w_183_1593, w_183_1595, w_183_1605, w_183_1607, w_183_1609, w_183_1611, w_183_1619, w_183_1626, w_183_1627, w_183_1630, w_183_1632, w_183_1636, w_183_1640, w_183_1644, w_183_1655, w_183_1657, w_183_1658, w_183_1665, w_183_1667, w_183_1668, w_183_1669, w_183_1673, w_183_1683, w_183_1688, w_183_1690, w_183_1691, w_183_1696, w_183_1699, w_183_1703, w_183_1711, w_183_1723, w_183_1724, w_183_1726, w_183_1728, w_183_1730, w_183_1736, w_183_1738, w_183_1740, w_183_1743, w_183_1745, w_183_1748, w_183_1749, w_183_1750, w_183_1751, w_183_1753, w_183_1759, w_183_1761, w_183_1765, w_183_1771, w_183_1772, w_183_1775, w_183_1777, w_183_1782, w_183_1783, w_183_1786, w_183_1787, w_183_1789, w_183_1795, w_183_1796, w_183_1803, w_183_1810, w_183_1811, w_183_1813, w_183_1814, w_183_1817, w_183_1826, w_183_1833, w_183_1842, w_183_1851, w_183_1852, w_183_1853, w_183_1856, w_183_1858, w_183_1863, w_183_1869, w_183_1870, w_183_1877, w_183_1881, w_183_1889, w_183_1893, w_183_1903, w_183_1906, w_183_1911, w_183_1913, w_183_1917, w_183_1919, w_183_1920, w_183_1922, w_183_1924, w_183_1927, w_183_1931, w_183_1932, w_183_1936, w_183_1938, w_183_1946, w_183_1947, w_183_1950, w_183_1951, w_183_1963, w_183_1966, w_183_1973, w_183_1974, w_183_1975, w_183_1976, w_183_1982, w_183_1984, w_183_1986, w_183_1988, w_183_1994, w_183_1998, w_183_2000, w_183_2001, w_183_2002, w_183_2004, w_183_2005, w_183_2009, w_183_2012, w_183_2024, w_183_2028, w_183_2034, w_183_2039, w_183_2040, w_183_2041, w_183_2045, w_183_2047, w_183_2049, w_183_2054, w_183_2055, w_183_2057, w_183_2059, w_183_2064, w_183_2072, w_183_2078, w_183_2086, w_183_2089, w_183_2090, w_183_2097, w_183_2102, w_183_2114, w_183_2117;
  wire w_184_000, w_184_001, w_184_006, w_184_007, w_184_009, w_184_011, w_184_019, w_184_021, w_184_024, w_184_030, w_184_036, w_184_041, w_184_042, w_184_045, w_184_051, w_184_052, w_184_053, w_184_056, w_184_057, w_184_060, w_184_063, w_184_068, w_184_073, w_184_077, w_184_078, w_184_079, w_184_080, w_184_082, w_184_084, w_184_085, w_184_090, w_184_091, w_184_098, w_184_110, w_184_111, w_184_119, w_184_120, w_184_125, w_184_136, w_184_137, w_184_138, w_184_142, w_184_143, w_184_146, w_184_147, w_184_151, w_184_159, w_184_162, w_184_166, w_184_173, w_184_176, w_184_178, w_184_179, w_184_180, w_184_181, w_184_182, w_184_194, w_184_197, w_184_200, w_184_202, w_184_203, w_184_204, w_184_208, w_184_211, w_184_212, w_184_213, w_184_222, w_184_228, w_184_232, w_184_237, w_184_248, w_184_249, w_184_250, w_184_253, w_184_256, w_184_263, w_184_270, w_184_272, w_184_273, w_184_278, w_184_279, w_184_281, w_184_284, w_184_289, w_184_292, w_184_294, w_184_297, w_184_304, w_184_305, w_184_308, w_184_312, w_184_314, w_184_332, w_184_347, w_184_349, w_184_350, w_184_360, w_184_365, w_184_373, w_184_382, w_184_385, w_184_388, w_184_394, w_184_398, w_184_400, w_184_402, w_184_406, w_184_408, w_184_409, w_184_411, w_184_421, w_184_434, w_184_437, w_184_448, w_184_462, w_184_464, w_184_469, w_184_471, w_184_478, w_184_486, w_184_490, w_184_497, w_184_499, w_184_503, w_184_504, w_184_508, w_184_510, w_184_511, w_184_521, w_184_522, w_184_526, w_184_528, w_184_529, w_184_538, w_184_541, w_184_555, w_184_579, w_184_581, w_184_586, w_184_587, w_184_588, w_184_592, w_184_597, w_184_599, w_184_602, w_184_604, w_184_605, w_184_609, w_184_616, w_184_619, w_184_623, w_184_626, w_184_628, w_184_629, w_184_636, w_184_637, w_184_639, w_184_646, w_184_652, w_184_653, w_184_659, w_184_660, w_184_663, w_184_666, w_184_671, w_184_673, w_184_674, w_184_675, w_184_677, w_184_684, w_184_686, w_184_687, w_184_690, w_184_701, w_184_705, w_184_709, w_184_710, w_184_714, w_184_715, w_184_717, w_184_720, w_184_725, w_184_728, w_184_733, w_184_737, w_184_740, w_184_741, w_184_742, w_184_746, w_184_749, w_184_751, w_184_753, w_184_754, w_184_757, w_184_758, w_184_767, w_184_774, w_184_776, w_184_778, w_184_782, w_184_784, w_184_791, w_184_794, w_184_799, w_184_800, w_184_804, w_184_808, w_184_811, w_184_815, w_184_816, w_184_819, w_184_829, w_184_830, w_184_831, w_184_834, w_184_835, w_184_837, w_184_840, w_184_842, w_184_844, w_184_845, w_184_848, w_184_850, w_184_853, w_184_855, w_184_856, w_184_862, w_184_871, w_184_876, w_184_878, w_184_879, w_184_885, w_184_901, w_184_904, w_184_910, w_184_913, w_184_915, w_184_920, w_184_921, w_184_924, w_184_928, w_184_931, w_184_933, w_184_935, w_184_939, w_184_942, w_184_947, w_184_950, w_184_953, w_184_957, w_184_958, w_184_959, w_184_963, w_184_964, w_184_966, w_184_967, w_184_969, w_184_971, w_184_972, w_184_975, w_184_980, w_184_986, w_184_990, w_184_993, w_184_1002, w_184_1006, w_184_1010, w_184_1011, w_184_1013, w_184_1014, w_184_1017, w_184_1024, w_184_1028, w_184_1029, w_184_1033, w_184_1038, w_184_1042, w_184_1048, w_184_1055, w_184_1058, w_184_1063, w_184_1066, w_184_1069, w_184_1071, w_184_1072, w_184_1073, w_184_1082, w_184_1083, w_184_1086, w_184_1090, w_184_1094, w_184_1101, w_184_1105, w_184_1108, w_184_1113, w_184_1115, w_184_1117, w_184_1123, w_184_1126, w_184_1130, w_184_1135, w_184_1137, w_184_1138, w_184_1141, w_184_1148, w_184_1149, w_184_1162, w_184_1163, w_184_1166, w_184_1167, w_184_1169, w_184_1178, w_184_1190, w_184_1192, w_184_1195, w_184_1196, w_184_1200, w_184_1202, w_184_1204, w_184_1206, w_184_1208, w_184_1213, w_184_1219, w_184_1223, w_184_1225, w_184_1226, w_184_1228, w_184_1242, w_184_1245, w_184_1251, w_184_1253, w_184_1254, w_184_1258, w_184_1262, w_184_1273, w_184_1274, w_184_1277, w_184_1281, w_184_1285, w_184_1294, w_184_1295, w_184_1297, w_184_1304, w_184_1308, w_184_1309, w_184_1312, w_184_1315, w_184_1317, w_184_1318, w_184_1320, w_184_1322, w_184_1323, w_184_1324, w_184_1332, w_184_1333, w_184_1340, w_184_1341, w_184_1343, w_184_1349, w_184_1350, w_184_1357, w_184_1364, w_184_1366, w_184_1373, w_184_1380, w_184_1382, w_184_1385, w_184_1387, w_184_1392, w_184_1397, w_184_1407, w_184_1409, w_184_1414, w_184_1416, w_184_1420, w_184_1426, w_184_1427, w_184_1431, w_184_1433, w_184_1434, w_184_1444, w_184_1450, w_184_1452, w_184_1459, w_184_1462, w_184_1463, w_184_1466, w_184_1469, w_184_1475, w_184_1481, w_184_1482, w_184_1484, w_184_1486, w_184_1488, w_184_1492, w_184_1493, w_184_1496, w_184_1500, w_184_1505, w_184_1507, w_184_1512, w_184_1514, w_184_1530, w_184_1534, w_184_1539, w_184_1542, w_184_1543, w_184_1547, w_184_1550, w_184_1551, w_184_1552, w_184_1554, w_184_1558, w_184_1559, w_184_1560, w_184_1563, w_184_1564, w_184_1565, w_184_1567, w_184_1569, w_184_1574, w_184_1577, w_184_1578, w_184_1582, w_184_1586, w_184_1587, w_184_1595, w_184_1598, w_184_1604, w_184_1608, w_184_1612, w_184_1617, w_184_1618, w_184_1625, w_184_1634, w_184_1635, w_184_1636, w_184_1640, w_184_1644, w_184_1655, w_184_1656, w_184_1657, w_184_1661, w_184_1665, w_184_1667, w_184_1668, w_184_1669, w_184_1680, w_184_1682, w_184_1687, w_184_1689, w_184_1690, w_184_1691, w_184_1693, w_184_1699, w_184_1703, w_184_1708, w_184_1713, w_184_1714, w_184_1716, w_184_1719, w_184_1720, w_184_1722, w_184_1725, w_184_1741, w_184_1746, w_184_1750, w_184_1752, w_184_1760, w_184_1765, w_184_1767, w_184_1770, w_184_1773, w_184_1774, w_184_1777, w_184_1780, w_184_1784, w_184_1793, w_184_1801, w_184_1803, w_184_1804, w_184_1805, w_184_1807, w_184_1808, w_184_1813, w_184_1822, w_184_1823, w_184_1831, w_184_1835, w_184_1843, w_184_1847, w_184_1848, w_184_1853, w_184_1860, w_184_1863, w_184_1865, w_184_1867, w_184_1868, w_184_1873, w_184_1875, w_184_1876, w_184_1877, w_184_1882, w_184_1889, w_184_1892, w_184_1899, w_184_1904, w_184_1907, w_184_1912, w_184_1915, w_184_1917, w_184_1918, w_184_1920, w_184_1922, w_184_1930, w_184_1932, w_184_1938, w_184_1941, w_184_1946, w_184_1947, w_184_1949, w_184_1952, w_184_1953, w_184_1957, w_184_1961, w_184_1965, w_184_1970, w_184_1977, w_184_1980, w_184_1981, w_184_1983, w_184_1986, w_184_1987, w_184_1995, w_184_1996, w_184_1997, w_184_2001, w_184_2002, w_184_2008, w_184_2015, w_184_2016, w_184_2017, w_184_2019, w_184_2020, w_184_2021, w_184_2023, w_184_2032, w_184_2035, w_184_2036, w_184_2039, w_184_2045, w_184_2050, w_184_2055, w_184_2058, w_184_2069, w_184_2070, w_184_2071, w_184_2074, w_184_2076, w_184_2079, w_184_2080, w_184_2083, w_184_2093, w_184_2098, w_184_2099, w_184_2101, w_184_2103, w_184_2104, w_184_2123, w_184_2126, w_184_2139, w_184_2157, w_184_2158, w_184_2172, w_184_2180, w_184_2192, w_184_2194, w_184_2209, w_184_2211, w_184_2222, w_184_2224, w_184_2228, w_184_2235, w_184_2241, w_184_2246, w_184_2253, w_184_2267, w_184_2273, w_184_2282, w_184_2287, w_184_2290, w_184_2302, w_184_2369, w_184_2375, w_184_2384, w_184_2389, w_184_2403, w_184_2404, w_184_2407, w_184_2423, w_184_2428, w_184_2437, w_184_2442, w_184_2444, w_184_2446, w_184_2449, w_184_2452, w_184_2456, w_184_2472, w_184_2474, w_184_2475, w_184_2476, w_184_2479, w_184_2481, w_184_2499, w_184_2507, w_184_2523, w_184_2524, w_184_2525, w_184_2538, w_184_2543, w_184_2548, w_184_2560, w_184_2562, w_184_2563, w_184_2581, w_184_2593, w_184_2596, w_184_2602, w_184_2613, w_184_2616, w_184_2621, w_184_2625, w_184_2640, w_184_2645, w_184_2648, w_184_2670, w_184_2671, w_184_2679, w_184_2685, w_184_2694, w_184_2702, w_184_2707, w_184_2711, w_184_2716, w_184_2718, w_184_2721, w_184_2724, w_184_2725, w_184_2734, w_184_2736, w_184_2748, w_184_2754, w_184_2757, w_184_2761, w_184_2781, w_184_2793, w_184_2794, w_184_2795, w_184_2807, w_184_2817, w_184_2820, w_184_2821, w_184_2826, w_184_2829, w_184_2831, w_184_2834, w_184_2838, w_184_2847, w_184_2848, w_184_2853, w_184_2857, w_184_2862, w_184_2874, w_184_2882, w_184_2883;
  wire w_185_005, w_185_006, w_185_007, w_185_009, w_185_011, w_185_012, w_185_016, w_185_018, w_185_019, w_185_022, w_185_025, w_185_029, w_185_033, w_185_035, w_185_036, w_185_037, w_185_038, w_185_044, w_185_045, w_185_047, w_185_048, w_185_049, w_185_050, w_185_052, w_185_058, w_185_062, w_185_064, w_185_065, w_185_066, w_185_074, w_185_076, w_185_079, w_185_081, w_185_084, w_185_085, w_185_094, w_185_096, w_185_102, w_185_105, w_185_107, w_185_112, w_185_121, w_185_122, w_185_123, w_185_125, w_185_130, w_185_133, w_185_134, w_185_140, w_185_146, w_185_147, w_185_148, w_185_149, w_185_152, w_185_154, w_185_156, w_185_160, w_185_163, w_185_164, w_185_175, w_185_177, w_185_178, w_185_179, w_185_180, w_185_195, w_185_200, w_185_202, w_185_203, w_185_205, w_185_206, w_185_208, w_185_209, w_185_213, w_185_225, w_185_229, w_185_245, w_185_246, w_185_249, w_185_251, w_185_252, w_185_256, w_185_259, w_185_266, w_185_268, w_185_269, w_185_275, w_185_276, w_185_279, w_185_283, w_185_286, w_185_287, w_185_288, w_185_294, w_185_295, w_185_299, w_185_304, w_185_305, w_185_306, w_185_311, w_185_312, w_185_314, w_185_315, w_185_316, w_185_318, w_185_320, w_185_324, w_185_325, w_185_326, w_185_330, w_185_334, w_185_335, w_185_340, w_185_351, w_185_362, w_185_363, w_185_364, w_185_371, w_185_377, w_185_381, w_185_390, w_185_395, w_185_396, w_185_398, w_185_399, w_185_403, w_185_405, w_185_406, w_185_415, w_185_416, w_185_417, w_185_418, w_185_420, w_185_422, w_185_423, w_185_425, w_185_427, w_185_428, w_185_431, w_185_434, w_185_438, w_185_443, w_185_447, w_185_449, w_185_451, w_185_452, w_185_456, w_185_462, w_185_464, w_185_469, w_185_472, w_185_474, w_185_475, w_185_482, w_185_485, w_185_491, w_185_497, w_185_502, w_185_503, w_185_505, w_185_508, w_185_509, w_185_521, w_185_536, w_185_541, w_185_546, w_185_547, w_185_552, w_185_557, w_185_562, w_185_563, w_185_564, w_185_572, w_185_578, w_185_579, w_185_581, w_185_582, w_185_583, w_185_587, w_185_588, w_185_597, w_185_598, w_185_604, w_185_609, w_185_610, w_185_611, w_185_615, w_185_620, w_185_621, w_185_622, w_185_631, w_185_633, w_185_635, w_185_636, w_185_640, w_185_641, w_185_643, w_185_645, w_185_649, w_185_653, w_185_655, w_185_656, w_185_657, w_185_659, w_185_675, w_185_676, w_185_677, w_185_683, w_185_694, w_185_699, w_185_700, w_185_702, w_185_703, w_185_704, w_185_707, w_185_719, w_185_722, w_185_727, w_185_728, w_185_729, w_185_731, w_185_732, w_185_742, w_185_745, w_185_749, w_185_751, w_185_753, w_185_754, w_185_755, w_185_759, w_185_764, w_185_765, w_185_767, w_185_769, w_185_771, w_185_773, w_185_774, w_185_775, w_185_776, w_185_780, w_185_781, w_185_783, w_185_784, w_185_787, w_185_789, w_185_790, w_185_796, w_185_800, w_185_803, w_185_807, w_185_808, w_185_819, w_185_822, w_185_830, w_185_835, w_185_837, w_185_841, w_185_842, w_185_844, w_185_845, w_185_847, w_185_850, w_185_853, w_185_859, w_185_874, w_185_878, w_185_882, w_185_891, w_185_895, w_185_900, w_185_903, w_185_905, w_185_907, w_185_908, w_185_911, w_185_912, w_185_914, w_185_925, w_185_928, w_185_929, w_185_933, w_185_935, w_185_936, w_185_937, w_185_938, w_185_939, w_185_950, w_185_952, w_185_955, w_185_962, w_185_969, w_185_977, w_185_978, w_185_983, w_185_987, w_185_993, w_185_1005, w_185_1011, w_185_1012, w_185_1016, w_185_1022, w_185_1024, w_185_1025, w_185_1037, w_185_1039, w_185_1042, w_185_1043, w_185_1053, w_185_1055, w_185_1056, w_185_1070, w_185_1072, w_185_1082, w_185_1092, w_185_1098, w_185_1100, w_185_1106, w_185_1117, w_185_1119, w_185_1121, w_185_1125, w_185_1129, w_185_1131, w_185_1136, w_185_1138, w_185_1139, w_185_1140, w_185_1147, w_185_1149, w_185_1152, w_185_1155, w_185_1159, w_185_1161, w_185_1165, w_185_1168, w_185_1172, w_185_1175, w_185_1180, w_185_1185, w_185_1187, w_185_1188, w_185_1191, w_185_1193, w_185_1194, w_185_1201, w_185_1205, w_185_1210, w_185_1212, w_185_1216, w_185_1217, w_185_1221, w_185_1222, w_185_1223, w_185_1230, w_185_1233, w_185_1235, w_185_1246, w_185_1250, w_185_1252, w_185_1260, w_185_1264, w_185_1266, w_185_1268, w_185_1269, w_185_1272, w_185_1273, w_185_1274, w_185_1275, w_185_1281, w_185_1284, w_185_1285, w_185_1287, w_185_1292, w_185_1293, w_185_1297, w_185_1302, w_185_1310, w_185_1317, w_185_1318, w_185_1320, w_185_1321, w_185_1323, w_185_1325, w_185_1332, w_185_1341, w_185_1346, w_185_1347, w_185_1348, w_185_1355, w_185_1357, w_185_1362, w_185_1366, w_185_1369, w_185_1371, w_185_1372, w_185_1374, w_185_1376, w_185_1377, w_185_1378, w_185_1380, w_185_1385, w_185_1386, w_185_1387, w_185_1393, w_185_1396, w_185_1402, w_185_1404, w_185_1405, w_185_1409, w_185_1410, w_185_1413, w_185_1415, w_185_1420, w_185_1422, w_185_1430, w_185_1433, w_185_1435, w_185_1436, w_185_1437, w_185_1440, w_185_1443, w_185_1444, w_185_1445, w_185_1446, w_185_1449, w_185_1452, w_185_1454, w_185_1455, w_185_1460, w_185_1461, w_185_1472, w_185_1474, w_185_1477, w_185_1478, w_185_1481, w_185_1482, w_185_1489, w_185_1491, w_185_1495, w_185_1499, w_185_1501, w_185_1509, w_185_1513, w_185_1521, w_185_1531, w_185_1539, w_185_1544, w_185_1550, w_185_1559, w_185_1560, w_185_1562, w_185_1564, w_185_1566, w_185_1567, w_185_1569, w_185_1570, w_185_1572, w_185_1573, w_185_1580, w_185_1588, w_185_1590, w_185_1592, w_185_1593, w_185_1596, w_185_1597, w_185_1599, w_185_1601, w_185_1602, w_185_1606, w_185_1612, w_185_1622, w_185_1626, w_185_1632, w_185_1635, w_185_1636, w_185_1638, w_185_1645, w_185_1646, w_185_1648, w_185_1651, w_185_1653, w_185_1656, w_185_1661, w_185_1664, w_185_1665, w_185_1667, w_185_1670, w_185_1672, w_185_1674, w_185_1680, w_185_1682, w_185_1683, w_185_1686, w_185_1689, w_185_1703, w_185_1704, w_185_1709, w_185_1722, w_185_1723, w_185_1727, w_185_1729, w_185_1735, w_185_1742, w_185_1748, w_185_1752, w_185_1760, w_185_1783, w_185_1792, w_185_1793, w_185_1794, w_185_1795, w_185_1801, w_185_1802, w_185_1803, w_185_1806, w_185_1810, w_185_1812, w_185_1813, w_185_1827, w_185_1831, w_185_1832, w_185_1833, w_185_1836, w_185_1840, w_185_1849, w_185_1854, w_185_1855, w_185_1859, w_185_1860, w_185_1861, w_185_1863, w_185_1868, w_185_1872, w_185_1873, w_185_1876, w_185_1878, w_185_1880, w_185_1882, w_185_1883, w_185_1888, w_185_1893, w_185_1897, w_185_1903, w_185_1907, w_185_1913, w_185_1917, w_185_1918, w_185_1919, w_185_1921, w_185_1927, w_185_1930, w_185_1931, w_185_1933, w_185_1944, w_185_1946, w_185_1947, w_185_1952, w_185_1956, w_185_1962, w_185_1965, w_185_1969, w_185_1979, w_185_1980, w_185_1984, w_185_1986, w_185_1989, w_185_1992, w_185_1997, w_185_2000, w_185_2009, w_185_2015, w_185_2017, w_185_2028, w_185_2032, w_185_2035, w_185_2036, w_185_2038, w_185_2039, w_185_2041, w_185_2045, w_185_2049, w_185_2050, w_185_2052, w_185_2053, w_185_2054, w_185_2065, w_185_2066, w_185_2074, w_185_2077, w_185_2078, w_185_2081, w_185_2085, w_185_2089, w_185_2096, w_185_2101, w_185_2102, w_185_2109, w_185_2110, w_185_2111, w_185_2118, w_185_2123, w_185_2127, w_185_2133, w_185_2134, w_185_2166, w_185_2172, w_185_2177, w_185_2178, w_185_2202, w_185_2207, w_185_2211, w_185_2221, w_185_2224, w_185_2225, w_185_2229, w_185_2235, w_185_2248, w_185_2250, w_185_2253, w_185_2256, w_185_2262, w_185_2268, w_185_2279, w_185_2295, w_185_2296, w_185_2299, w_185_2306, w_185_2308, w_185_2309, w_185_2311, w_185_2312, w_185_2316, w_185_2322, w_185_2324, w_185_2326, w_185_2332, w_185_2341, w_185_2355, w_185_2365, w_185_2380, w_185_2384, w_185_2388, w_185_2390, w_185_2398, w_185_2402, w_185_2405, w_185_2414, w_185_2419, w_185_2421, w_185_2436, w_185_2439, w_185_2441, w_185_2455, w_185_2461, w_185_2465, w_185_2468, w_185_2471, w_185_2501, w_185_2503, w_185_2508, w_185_2527, w_185_2542, w_185_2549, w_185_2560, w_185_2562, w_185_2565, w_185_2571, w_185_2576, w_185_2581, w_185_2583, w_185_2584, w_185_2587, w_185_2589, w_185_2607, w_185_2617, w_185_2621, w_185_2635, w_185_2636, w_185_2658, w_185_2671, w_185_2679, w_185_2691, w_185_2692, w_185_2702, w_185_2703, w_185_2717, w_185_2720, w_185_2723, w_185_2726, w_185_2729, w_185_2730, w_185_2731, w_185_2734, w_185_2738, w_185_2745, w_185_2756, w_185_2766, w_185_2769, w_185_2784, w_185_2785, w_185_2813, w_185_2818, w_185_2820, w_185_2828, w_185_2830, w_185_2856;
  wire w_186_000, w_186_001, w_186_003, w_186_004, w_186_005, w_186_009, w_186_014, w_186_015, w_186_017, w_186_027, w_186_028, w_186_033, w_186_034, w_186_039, w_186_041, w_186_042, w_186_044, w_186_047, w_186_048, w_186_053, w_186_056, w_186_063, w_186_064, w_186_066, w_186_068, w_186_083, w_186_085, w_186_087, w_186_091, w_186_092, w_186_097, w_186_104, w_186_105, w_186_107, w_186_109, w_186_111, w_186_113, w_186_117, w_186_118, w_186_121, w_186_124, w_186_129, w_186_132, w_186_135, w_186_137, w_186_140, w_186_141, w_186_145, w_186_146, w_186_147, w_186_153, w_186_154, w_186_161, w_186_163, w_186_166, w_186_167, w_186_174, w_186_175, w_186_181, w_186_182, w_186_183, w_186_184, w_186_185, w_186_186, w_186_188, w_186_193, w_186_199, w_186_201, w_186_206, w_186_207, w_186_211, w_186_212, w_186_213, w_186_223, w_186_225, w_186_226, w_186_232, w_186_235, w_186_245, w_186_249, w_186_250, w_186_251, w_186_252, w_186_255, w_186_258, w_186_267, w_186_273, w_186_280, w_186_285, w_186_288, w_186_289, w_186_291, w_186_292, w_186_293, w_186_296, w_186_297, w_186_302, w_186_304, w_186_309, w_186_310, w_186_311, w_186_312, w_186_313, w_186_314, w_186_315, w_186_316, w_186_319, w_186_326, w_186_327, w_186_330, w_186_331, w_186_338, w_186_339, w_186_343, w_186_346, w_186_349, w_186_353, w_186_355, w_186_358, w_186_359, w_186_360, w_186_362, w_186_363, w_186_364, w_186_368, w_186_369, w_186_371, w_186_373, w_186_374, w_186_377, w_186_382, w_186_389, w_186_396, w_186_399, w_186_403, w_186_409, w_186_412, w_186_420, w_186_423, w_186_425, w_186_428, w_186_429, w_186_430, w_186_432, w_186_436, w_186_437, w_186_439, w_186_440, w_186_447, w_186_448, w_186_449, w_186_452, w_186_453, w_186_454, w_186_456, w_186_457, w_186_464, w_186_465, w_186_469, w_186_470, w_186_472, w_186_475, w_186_477, w_186_481, w_186_484, w_186_488, w_186_489, w_186_491, w_186_495, w_186_498, w_186_503, w_186_504, w_186_506, w_186_507, w_186_510, w_186_514, w_186_515, w_186_516, w_186_520, w_186_521, w_186_527, w_186_530, w_186_532, w_186_533, w_186_538, w_186_543, w_186_544, w_186_546, w_186_548, w_186_551, w_186_552, w_186_558, w_186_563, w_186_564, w_186_566, w_186_568, w_186_572, w_186_575, w_186_579, w_186_583, w_186_585, w_186_586, w_186_591, w_186_596, w_186_598, w_186_602, w_186_603, w_186_604, w_186_605, w_186_606, w_186_615, w_186_616, w_186_619, w_186_622, w_186_623, w_186_624, w_186_625, w_186_626, w_186_629, w_186_630, w_186_632, w_186_636, w_186_642, w_186_644, w_186_650, w_186_653, w_186_654, w_186_656, w_186_657, w_186_658, w_186_662, w_186_663, w_186_665, w_186_676, w_186_679, w_186_680, w_186_681, w_186_685, w_186_687, w_186_689, w_186_690, w_186_691, w_186_692, w_186_693, w_186_694, w_186_697, w_186_698, w_186_704, w_186_708, w_186_711, w_186_712, w_186_717, w_186_718, w_186_720, w_186_725, w_186_727, w_186_732, w_186_736, w_186_739, w_186_741, w_186_747, w_186_754, w_186_755, w_186_757, w_186_764, w_186_766, w_186_770, w_186_774, w_186_776, w_186_779, w_186_780, w_186_783, w_186_784, w_186_790, w_186_793, w_186_797, w_186_799, w_186_802, w_186_804, w_186_806, w_186_812, w_186_813, w_186_814, w_186_817, w_186_818, w_186_820, w_186_821, w_186_824, w_186_825, w_186_826, w_186_831, w_186_833, w_186_835, w_186_842, w_186_852, w_186_857, w_186_860, w_186_868, w_186_875, w_186_878, w_186_881, w_186_884, w_186_898, w_186_901, w_186_904, w_186_909, w_186_910, w_186_912, w_186_916, w_186_921, w_186_922, w_186_924, w_186_928, w_186_931, w_186_936, w_186_938, w_186_939, w_186_940, w_186_941, w_186_943, w_186_944, w_186_948, w_186_949, w_186_951, w_186_952, w_186_953, w_186_954, w_186_956, w_186_961, w_186_964, w_186_966, w_186_967, w_186_968, w_186_969, w_186_973, w_186_975, w_186_976, w_186_984, w_186_985, w_186_986, w_186_987, w_186_990, w_186_991, w_186_993, w_186_994, w_186_995, w_186_996, w_186_1009, w_186_1011, w_186_1012, w_186_1015, w_186_1016, w_186_1020, w_186_1021, w_186_1023, w_186_1024, w_186_1028, w_186_1029, w_186_1030, w_186_1032, w_186_1033, w_186_1034, w_186_1037, w_186_1038, w_186_1039, w_186_1041, w_186_1043, w_186_1049, w_186_1050, w_186_1052, w_186_1053, w_186_1058, w_186_1059, w_186_1060, w_186_1062, w_186_1073, w_186_1074, w_186_1077, w_186_1079, w_186_1080, w_186_1084, w_186_1085, w_186_1092, w_186_1101, w_186_1102, w_186_1104, w_186_1105, w_186_1109, w_186_1114, w_186_1119, w_186_1125, w_186_1127, w_186_1130, w_186_1132, w_186_1139, w_186_1142, w_186_1144, w_186_1152, w_186_1153, w_186_1156, w_186_1157, w_186_1158, w_186_1159, w_186_1160, w_186_1165, w_186_1167, w_186_1168, w_186_1172, w_186_1173, w_186_1174, w_186_1175, w_186_1179, w_186_1180, w_186_1182, w_186_1183, w_186_1187, w_186_1189, w_186_1190, w_186_1192, w_186_1193, w_186_1196, w_186_1199, w_186_1201, w_186_1205, w_186_1206, w_186_1207, w_186_1213, w_186_1217, w_186_1218, w_186_1221, w_186_1222, w_186_1224, w_186_1225, w_186_1227, w_186_1232, w_186_1236, w_186_1249, w_186_1251, w_186_1254, w_186_1255, w_186_1256, w_186_1259, w_186_1267, w_186_1277, w_186_1279, w_186_1284, w_186_1287, w_186_1290, w_186_1292, w_186_1297, w_186_1298, w_186_1299, w_186_1300, w_186_1303, w_186_1308, w_186_1309, w_186_1313, w_186_1314, w_186_1316, w_186_1319, w_186_1324, w_186_1325, w_186_1326, w_186_1330, w_186_1333, w_186_1334, w_186_1335, w_186_1336, w_186_1337, w_186_1339, w_186_1341, w_186_1347, w_186_1349, w_186_1352, w_186_1353, w_186_1354, w_186_1355, w_186_1358, w_186_1362, w_186_1363, w_186_1364, w_186_1365, w_186_1371, w_186_1372, w_186_1373, w_186_1374, w_186_1376, w_186_1378, w_186_1383, w_186_1385, w_186_1386, w_186_1387, w_186_1388, w_186_1389, w_186_1393, w_186_1395, w_186_1396, w_186_1397, w_186_1402, w_186_1405, w_186_1407, w_186_1408, w_186_1412, w_186_1414, w_186_1418, w_186_1420, w_186_1423, w_186_1427, w_186_1430, w_186_1434, w_186_1438, w_186_1446, w_186_1453, w_186_1459, w_186_1464, w_186_1466, w_186_1469, w_186_1470, w_186_1473, w_186_1477, w_186_1480, w_186_1482, w_186_1483, w_186_1486, w_186_1488, w_186_1491, w_186_1493, w_186_1494, w_186_1495, w_186_1496, w_186_1497, w_186_1501, w_186_1502, w_186_1505, w_186_1507, w_186_1510, w_186_1515, w_186_1517, w_186_1518, w_186_1521, w_186_1524, w_186_1525, w_186_1527, w_186_1531, w_186_1532, w_186_1538, w_186_1544, w_186_1546, w_186_1550, w_186_1551, w_186_1552, w_186_1553, w_186_1555, w_186_1558, w_186_1559, w_186_1565, w_186_1567, w_186_1570, w_186_1571, w_186_1577, w_186_1578, w_186_1579, w_186_1582, w_186_1584, w_186_1585, w_186_1589, w_186_1592, w_186_1596, w_186_1598, w_186_1602, w_186_1603, w_186_1604, w_186_1607, w_186_1609, w_186_1611, w_186_1612, w_186_1613, w_186_1621, w_186_1628, w_186_1631, w_186_1633, w_186_1637, w_186_1642, w_186_1643, w_186_1644, w_186_1647, w_186_1654, w_186_1657, w_186_1661, w_186_1662, w_186_1663, w_186_1664, w_186_1665, w_186_1666;
  wire w_187_000, w_187_006, w_187_008, w_187_012, w_187_024, w_187_025, w_187_031, w_187_037, w_187_040, w_187_041, w_187_048, w_187_052, w_187_056, w_187_063, w_187_064, w_187_067, w_187_070, w_187_073, w_187_075, w_187_076, w_187_077, w_187_078, w_187_079, w_187_082, w_187_083, w_187_088, w_187_090, w_187_095, w_187_105, w_187_106, w_187_110, w_187_115, w_187_118, w_187_121, w_187_125, w_187_136, w_187_139, w_187_142, w_187_147, w_187_164, w_187_166, w_187_170, w_187_172, w_187_173, w_187_176, w_187_179, w_187_185, w_187_188, w_187_194, w_187_195, w_187_198, w_187_200, w_187_202, w_187_214, w_187_218, w_187_219, w_187_221, w_187_232, w_187_244, w_187_245, w_187_253, w_187_255, w_187_262, w_187_265, w_187_268, w_187_272, w_187_274, w_187_276, w_187_278, w_187_279, w_187_284, w_187_289, w_187_292, w_187_298, w_187_299, w_187_308, w_187_312, w_187_313, w_187_314, w_187_316, w_187_320, w_187_323, w_187_326, w_187_329, w_187_330, w_187_331, w_187_333, w_187_336, w_187_339, w_187_343, w_187_346, w_187_352, w_187_355, w_187_360, w_187_370, w_187_372, w_187_373, w_187_380, w_187_381, w_187_384, w_187_391, w_187_392, w_187_398, w_187_400, w_187_404, w_187_411, w_187_412, w_187_413, w_187_416, w_187_418, w_187_420, w_187_421, w_187_422, w_187_426, w_187_432, w_187_433, w_187_434, w_187_436, w_187_439, w_187_442, w_187_462, w_187_465, w_187_472, w_187_477, w_187_479, w_187_483, w_187_488, w_187_489, w_187_490, w_187_491, w_187_493, w_187_494, w_187_495, w_187_498, w_187_503, w_187_510, w_187_512, w_187_514, w_187_519, w_187_521, w_187_522, w_187_524, w_187_527, w_187_530, w_187_533, w_187_534, w_187_535, w_187_538, w_187_539, w_187_549, w_187_551, w_187_552, w_187_557, w_187_564, w_187_567, w_187_569, w_187_580, w_187_582, w_187_583, w_187_591, w_187_596, w_187_601, w_187_602, w_187_604, w_187_605, w_187_607, w_187_608, w_187_611, w_187_613, w_187_615, w_187_616, w_187_617, w_187_624, w_187_627, w_187_631, w_187_639, w_187_641, w_187_646, w_187_647, w_187_648, w_187_654, w_187_655, w_187_667, w_187_684, w_187_686, w_187_689, w_187_695, w_187_696, w_187_697, w_187_698, w_187_702, w_187_703, w_187_704, w_187_709, w_187_710, w_187_719, w_187_727, w_187_729, w_187_731, w_187_737, w_187_744, w_187_745, w_187_756, w_187_757, w_187_764, w_187_766, w_187_767, w_187_771, w_187_776, w_187_782, w_187_784, w_187_785, w_187_788, w_187_790, w_187_793, w_187_795, w_187_796, w_187_798, w_187_800, w_187_812, w_187_815, w_187_816, w_187_819, w_187_838, w_187_842, w_187_847, w_187_848, w_187_853, w_187_856, w_187_857, w_187_858, w_187_859, w_187_862, w_187_863, w_187_866, w_187_868, w_187_869, w_187_877, w_187_880, w_187_882, w_187_886, w_187_887, w_187_890, w_187_892, w_187_895, w_187_899, w_187_902, w_187_905, w_187_906, w_187_907, w_187_913, w_187_915, w_187_916, w_187_917, w_187_919, w_187_923, w_187_925, w_187_927, w_187_932, w_187_935, w_187_937, w_187_938, w_187_940, w_187_942, w_187_951, w_187_958, w_187_959, w_187_961, w_187_962, w_187_965, w_187_966, w_187_968, w_187_980, w_187_982, w_187_983, w_187_987, w_187_988, w_187_991, w_187_997, w_187_998, w_187_1002, w_187_1003, w_187_1004, w_187_1005, w_187_1006, w_187_1009, w_187_1010, w_187_1012, w_187_1015, w_187_1018, w_187_1024, w_187_1026, w_187_1034, w_187_1036, w_187_1037, w_187_1044, w_187_1046, w_187_1053, w_187_1055, w_187_1056, w_187_1062, w_187_1063, w_187_1069, w_187_1072, w_187_1074, w_187_1083, w_187_1088, w_187_1095, w_187_1101, w_187_1113, w_187_1116, w_187_1121, w_187_1130, w_187_1134, w_187_1136, w_187_1137, w_187_1140, w_187_1143, w_187_1147, w_187_1148, w_187_1151, w_187_1153, w_187_1165, w_187_1167, w_187_1170, w_187_1171, w_187_1179, w_187_1182, w_187_1187, w_187_1188, w_187_1198, w_187_1203, w_187_1210, w_187_1212, w_187_1215, w_187_1219, w_187_1221, w_187_1226, w_187_1229, w_187_1233, w_187_1234, w_187_1235, w_187_1240, w_187_1242, w_187_1243, w_187_1246, w_187_1247, w_187_1248, w_187_1254, w_187_1255, w_187_1264, w_187_1265, w_187_1270, w_187_1271, w_187_1277, w_187_1286, w_187_1288, w_187_1291, w_187_1292, w_187_1294, w_187_1307, w_187_1309, w_187_1316, w_187_1318, w_187_1322, w_187_1325, w_187_1326, w_187_1333, w_187_1335, w_187_1339, w_187_1340, w_187_1342, w_187_1344, w_187_1346, w_187_1347, w_187_1349, w_187_1351, w_187_1352, w_187_1353, w_187_1354, w_187_1359, w_187_1360, w_187_1366, w_187_1370, w_187_1373, w_187_1374, w_187_1377, w_187_1380, w_187_1385, w_187_1386, w_187_1388, w_187_1389, w_187_1390, w_187_1393, w_187_1398, w_187_1400, w_187_1405, w_187_1407, w_187_1410, w_187_1411, w_187_1412, w_187_1418, w_187_1421, w_187_1428, w_187_1431, w_187_1433, w_187_1434, w_187_1443, w_187_1445, w_187_1447, w_187_1449, w_187_1450, w_187_1454, w_187_1462, w_187_1466, w_187_1467, w_187_1469, w_187_1470, w_187_1472, w_187_1476, w_187_1477, w_187_1478, w_187_1481, w_187_1485, w_187_1488, w_187_1492, w_187_1498, w_187_1540, w_187_1546, w_187_1548, w_187_1563, w_187_1565, w_187_1572, w_187_1574, w_187_1579, w_187_1595, w_187_1598, w_187_1617, w_187_1638, w_187_1641, w_187_1643, w_187_1648, w_187_1657, w_187_1663, w_187_1664, w_187_1674, w_187_1675, w_187_1688, w_187_1689, w_187_1691, w_187_1694, w_187_1726, w_187_1728, w_187_1732, w_187_1742, w_187_1744, w_187_1750, w_187_1752, w_187_1757, w_187_1767, w_187_1773, w_187_1782, w_187_1803, w_187_1808, w_187_1812, w_187_1813, w_187_1825, w_187_1847, w_187_1851, w_187_1854, w_187_1855, w_187_1858, w_187_1862, w_187_1866, w_187_1872, w_187_1875, w_187_1885, w_187_1888, w_187_1894, w_187_1901, w_187_1904, w_187_1905, w_187_1908, w_187_1926, w_187_1927, w_187_1929, w_187_1930, w_187_1931, w_187_1943, w_187_1960, w_187_1976, w_187_1981, w_187_1985, w_187_1999, w_187_2012, w_187_2013, w_187_2017, w_187_2030, w_187_2037, w_187_2053, w_187_2070, w_187_2073, w_187_2078, w_187_2082, w_187_2093, w_187_2094, w_187_2104, w_187_2111, w_187_2113, w_187_2125, w_187_2127, w_187_2128, w_187_2154, w_187_2155, w_187_2160, w_187_2161, w_187_2163, w_187_2167, w_187_2171, w_187_2174, w_187_2180, w_187_2181, w_187_2188, w_187_2195, w_187_2201, w_187_2205, w_187_2214, w_187_2219, w_187_2221, w_187_2224, w_187_2230, w_187_2233, w_187_2234, w_187_2241, w_187_2250, w_187_2271, w_187_2297, w_187_2299, w_187_2302, w_187_2303, w_187_2307, w_187_2323, w_187_2332, w_187_2353, w_187_2355, w_187_2363, w_187_2366, w_187_2367, w_187_2377, w_187_2392, w_187_2395, w_187_2399, w_187_2433, w_187_2435, w_187_2437, w_187_2440, w_187_2442, w_187_2457, w_187_2464, w_187_2470, w_187_2472, w_187_2485, w_187_2490, w_187_2504, w_187_2509, w_187_2528, w_187_2530, w_187_2532, w_187_2536, w_187_2538, w_187_2542, w_187_2546, w_187_2548, w_187_2554, w_187_2571, w_187_2577, w_187_2579, w_187_2590, w_187_2592, w_187_2593, w_187_2595, w_187_2611, w_187_2621, w_187_2631, w_187_2635, w_187_2639, w_187_2653, w_187_2654, w_187_2658, w_187_2662, w_187_2687, w_187_2696, w_187_2713, w_187_2726, w_187_2729, w_187_2732, w_187_2752, w_187_2755, w_187_2757, w_187_2758, w_187_2759, w_187_2760, w_187_2762, w_187_2772, w_187_2776, w_187_2798, w_187_2807, w_187_2811, w_187_2830, w_187_2837, w_187_2838, w_187_2841, w_187_2843, w_187_2848, w_187_2856, w_187_2858, w_187_2867, w_187_2874, w_187_2876, w_187_2881, w_187_2890, w_187_2893, w_187_2899, w_187_2901, w_187_2908, w_187_2912, w_187_2916, w_187_2918, w_187_2920, w_187_2924, w_187_2938, w_187_2940, w_187_2952, w_187_2959, w_187_2960, w_187_2963, w_187_2968, w_187_2973, w_187_2975, w_187_3003, w_187_3005, w_187_3015, w_187_3022, w_187_3023, w_187_3038, w_187_3039, w_187_3046, w_187_3057, w_187_3068, w_187_3076, w_187_3092, w_187_3104, w_187_3110, w_187_3121, w_187_3123, w_187_3142, w_187_3148, w_187_3156, w_187_3159, w_187_3174, w_187_3188, w_187_3191, w_187_3192, w_187_3194, w_187_3202, w_187_3205, w_187_3214, w_187_3215, w_187_3242, w_187_3250, w_187_3257, w_187_3263, w_187_3265, w_187_3267, w_187_3275, w_187_3285, w_187_3291, w_187_3293, w_187_3299, w_187_3311, w_187_3312, w_187_3314, w_187_3315, w_187_3319, w_187_3339, w_187_3359, w_187_3371, w_187_3377, w_187_3381, w_187_3388, w_187_3389, w_187_3395, w_187_3410, w_187_3415, w_187_3424, w_187_3438, w_187_3443, w_187_3444, w_187_3448, w_187_3453, w_187_3474;
  wire w_188_001, w_188_003, w_188_004, w_188_007, w_188_010, w_188_013, w_188_017, w_188_019, w_188_020, w_188_021, w_188_022, w_188_024, w_188_025, w_188_028, w_188_030, w_188_031, w_188_033, w_188_035, w_188_036, w_188_042, w_188_049, w_188_054, w_188_057, w_188_060, w_188_061, w_188_062, w_188_064, w_188_065, w_188_068, w_188_070, w_188_072, w_188_075, w_188_076, w_188_078, w_188_079, w_188_081, w_188_083, w_188_086, w_188_087, w_188_089, w_188_091, w_188_092, w_188_094, w_188_097, w_188_099, w_188_103, w_188_104, w_188_105, w_188_108, w_188_110, w_188_112, w_188_114, w_188_117, w_188_118, w_188_122, w_188_124, w_188_131, w_188_133, w_188_135, w_188_136, w_188_141, w_188_142, w_188_144, w_188_145, w_188_147, w_188_148, w_188_150, w_188_158, w_188_159, w_188_161, w_188_162, w_188_164, w_188_167, w_188_168, w_188_169, w_188_171, w_188_172, w_188_174, w_188_179, w_188_181, w_188_185, w_188_188, w_188_189, w_188_190, w_188_192, w_188_195, w_188_199, w_188_200, w_188_201, w_188_205, w_188_210, w_188_211, w_188_213, w_188_215, w_188_218, w_188_219, w_188_220, w_188_221, w_188_223, w_188_225, w_188_226, w_188_227, w_188_233, w_188_236, w_188_239, w_188_240, w_188_241, w_188_245, w_188_247, w_188_248, w_188_254, w_188_256, w_188_257, w_188_259, w_188_260, w_188_262, w_188_263, w_188_267, w_188_268, w_188_273, w_188_274, w_188_276, w_188_280, w_188_282, w_188_283, w_188_285, w_188_290, w_188_295, w_188_296, w_188_297, w_188_298, w_188_300, w_188_302, w_188_303, w_188_304, w_188_305, w_188_310, w_188_311, w_188_314, w_188_315, w_188_316, w_188_318, w_188_319, w_188_320, w_188_325, w_188_326, w_188_330, w_188_331, w_188_332, w_188_333, w_188_334, w_188_336, w_188_337, w_188_338, w_188_339, w_188_341, w_188_344, w_188_347, w_188_349, w_188_354, w_188_356, w_188_358, w_188_359, w_188_361, w_188_362, w_188_363, w_188_364, w_188_365, w_188_369, w_188_370, w_188_372, w_188_375, w_188_376, w_188_377, w_188_378, w_188_379, w_188_381, w_188_382, w_188_383, w_188_384, w_188_385, w_188_387, w_188_390, w_188_392, w_188_393, w_188_396, w_188_397, w_188_399, w_188_403, w_188_406, w_188_409, w_188_410, w_188_413, w_188_415, w_188_417, w_188_418, w_188_420, w_188_423, w_188_424, w_188_426, w_188_428, w_188_429, w_188_430, w_188_431, w_188_434, w_188_437, w_188_439, w_188_440, w_188_441, w_188_442, w_188_445, w_188_446, w_188_447, w_188_448, w_188_452, w_188_453, w_188_454, w_188_457, w_188_458, w_188_459, w_188_461, w_188_462, w_188_466, w_188_468, w_188_472, w_188_475, w_188_477, w_188_481, w_188_484, w_188_485, w_188_488, w_188_489, w_188_490, w_188_493, w_188_494, w_188_496, w_188_499, w_188_500, w_188_501, w_188_502, w_188_503, w_188_504, w_188_505, w_188_507, w_188_509, w_188_518, w_188_521, w_188_524, w_188_525, w_188_527, w_188_530, w_188_531, w_188_532, w_188_533, w_188_538, w_188_542, w_188_543, w_188_545, w_188_547, w_188_553, w_188_559, w_188_560, w_188_564, w_188_566, w_188_572, w_188_575, w_188_577, w_188_578, w_188_581, w_188_589, w_188_590, w_188_591, w_188_593, w_188_595, w_188_603, w_188_604, w_188_609, w_188_610, w_188_613, w_188_615, w_188_618, w_188_619, w_188_621, w_188_623, w_188_625, w_188_627, w_188_628, w_188_629, w_188_632, w_188_634, w_188_635, w_188_637, w_188_638, w_188_646, w_188_649, w_188_651, w_188_652, w_188_653, w_188_656, w_188_661, w_188_662, w_188_669, w_188_672, w_188_673, w_188_674, w_188_675, w_188_680, w_188_681, w_188_683, w_188_686, w_188_687, w_188_691, w_188_692, w_188_693, w_188_703, w_188_706, w_188_710, w_188_712, w_188_715, w_188_717, w_188_719, w_188_720, w_188_721, w_188_723, w_188_724, w_188_726, w_188_728, w_188_732, w_188_733, w_188_735, w_188_737, w_188_739, w_188_745, w_188_746, w_188_749, w_188_755, w_188_759, w_188_762, w_188_763, w_188_765, w_188_772, w_188_774, w_188_776, w_188_778, w_188_779, w_188_781, w_188_784, w_188_785, w_188_786, w_188_791, w_188_792, w_188_793, w_188_794, w_188_795, w_188_796, w_188_798, w_188_799, w_188_805, w_188_811, w_188_814, w_188_816, w_188_817, w_188_820, w_188_821, w_188_824, w_188_825, w_188_826, w_188_828, w_188_830, w_188_831, w_188_832, w_188_833, w_188_836, w_188_839, w_188_840, w_188_842, w_188_843, w_188_845, w_188_846, w_188_849, w_188_850, w_188_851, w_188_852, w_188_853, w_188_854, w_188_859, w_188_861, w_188_862, w_188_865, w_188_866, w_188_867, w_188_868, w_188_870, w_188_871, w_188_872, w_188_876, w_188_877, w_188_878, w_188_879, w_188_880, w_188_881, w_188_884, w_188_886, w_188_889, w_188_890, w_188_892, w_188_893, w_188_897, w_188_899, w_188_903, w_188_905, w_188_906, w_188_910, w_188_912, w_188_913, w_188_914, w_188_921, w_188_924, w_188_925, w_188_927, w_188_928, w_188_930, w_188_933, w_188_936, w_188_938, w_188_939, w_188_943, w_188_946, w_188_948, w_188_960, w_188_961, w_188_962, w_188_963, w_188_964, w_188_967, w_188_970, w_188_971, w_188_973, w_188_974, w_188_978, w_188_982, w_188_987, w_188_990, w_188_994, w_188_995, w_188_1004, w_188_1006, w_188_1008, w_188_1010, w_188_1011, w_188_1012, w_188_1017, w_188_1018, w_188_1024, w_188_1031, w_188_1032, w_188_1034, w_188_1035, w_188_1040, w_188_1044, w_188_1045, w_188_1046, w_188_1053, w_188_1057, w_188_1062, w_188_1063, w_188_1066, w_188_1067, w_188_1068, w_188_1069, w_188_1071, w_188_1073, w_188_1076, w_188_1077, w_188_1078, w_188_1080, w_188_1083, w_188_1086, w_188_1092, w_188_1099, w_188_1101, w_188_1105, w_188_1106, w_188_1110, w_188_1113, w_188_1115, w_188_1119, w_188_1120, w_188_1122, w_188_1126, w_188_1127, w_188_1130, w_188_1132, w_188_1135, w_188_1136, w_188_1137, w_188_1138, w_188_1142, w_188_1143, w_188_1146, w_188_1147, w_188_1150, w_188_1152, w_188_1158, w_188_1161, w_188_1163, w_188_1164, w_188_1166, w_188_1167, w_188_1169, w_188_1176, w_188_1178, w_188_1179, w_188_1180, w_188_1182, w_188_1184, w_188_1186, w_188_1191, w_188_1195, w_188_1197, w_188_1202, w_188_1208, w_188_1211, w_188_1212, w_188_1218, w_188_1219, w_188_1222, w_188_1227, w_188_1230, w_188_1232, w_188_1235, w_188_1238, w_188_1239, w_188_1240, w_188_1245, w_188_1248, w_188_1252, w_188_1255, w_188_1259, w_188_1262, w_188_1263, w_188_1270, w_188_1272, w_188_1274, w_188_1275, w_188_1279, w_188_1280, w_188_1285, w_188_1289, w_188_1291, w_188_1292, w_188_1294, w_188_1295, w_188_1302, w_188_1305, w_188_1311, w_188_1312, w_188_1313, w_188_1314, w_188_1315, w_188_1319, w_188_1320, w_188_1323, w_188_1330, w_188_1332, w_188_1336, w_188_1337;
  wire w_189_001, w_189_005, w_189_006, w_189_008, w_189_011, w_189_014, w_189_015, w_189_016, w_189_017, w_189_019, w_189_021, w_189_022, w_189_026, w_189_027, w_189_029, w_189_031, w_189_032, w_189_033, w_189_034, w_189_035, w_189_036, w_189_037, w_189_039, w_189_040, w_189_044, w_189_045, w_189_046, w_189_047, w_189_048, w_189_051, w_189_052, w_189_053, w_189_057, w_189_058, w_189_059, w_189_061, w_189_062, w_189_065, w_189_066, w_189_067, w_189_068, w_189_069, w_189_070, w_189_071, w_189_073, w_189_074, w_189_075, w_189_076, w_189_079, w_189_080, w_189_081, w_189_083, w_189_084, w_189_085, w_189_086, w_189_087, w_189_088, w_189_090, w_189_091, w_189_092, w_189_096, w_189_098, w_189_099, w_189_100, w_189_102, w_189_103, w_189_104, w_189_105, w_189_106, w_189_108, w_189_109, w_189_110, w_189_111, w_189_112, w_189_113, w_189_115, w_189_116, w_189_118, w_189_119, w_189_120, w_189_121, w_189_122, w_189_125, w_189_126, w_189_127, w_189_129, w_189_131, w_189_132, w_189_135, w_189_137, w_189_140, w_189_141, w_189_142, w_189_143, w_189_146, w_189_147, w_189_148, w_189_151, w_189_152, w_189_155, w_189_156, w_189_157, w_189_160, w_189_162, w_189_164, w_189_165, w_189_167, w_189_168, w_189_171, w_189_173, w_189_174, w_189_175, w_189_177, w_189_178, w_189_179, w_189_182, w_189_183, w_189_184, w_189_185, w_189_189, w_189_190, w_189_192, w_189_193, w_189_195, w_189_196, w_189_197, w_189_199, w_189_200, w_189_201, w_189_202, w_189_204, w_189_207, w_189_209, w_189_211, w_189_213, w_189_215, w_189_220, w_189_221, w_189_223, w_189_224, w_189_226, w_189_227, w_189_228, w_189_229, w_189_230, w_189_232, w_189_234, w_189_235, w_189_236, w_189_239, w_189_243, w_189_244, w_189_245, w_189_247, w_189_249, w_189_250, w_189_251, w_189_252, w_189_254, w_189_255, w_189_257, w_189_259, w_189_260, w_189_262, w_189_263, w_189_269, w_189_270, w_189_271, w_189_274, w_189_276, w_189_278, w_189_281, w_189_282, w_189_284, w_189_285, w_189_289, w_189_290, w_189_291, w_189_293, w_189_294, w_189_295, w_189_298, w_189_300, w_189_301, w_189_302, w_189_304, w_189_305, w_189_307, w_189_310, w_189_311, w_189_313, w_189_315, w_189_316, w_189_317, w_189_318, w_189_320, w_189_323, w_189_324, w_189_325, w_189_326, w_189_328, w_189_329, w_189_330, w_189_331, w_189_332, w_189_333, w_189_336, w_189_338, w_189_339, w_189_341, w_189_343, w_189_345, w_189_346, w_189_347, w_189_348, w_189_349, w_189_350, w_189_351, w_189_352, w_189_353, w_189_354, w_189_355, w_189_356, w_189_357, w_189_358, w_189_359, w_189_360, w_189_362, w_189_363, w_189_365, w_189_366, w_189_367, w_189_368, w_189_373, w_189_375, w_189_377, w_189_378, w_189_380, w_189_382, w_189_383, w_189_386, w_189_389, w_189_392, w_189_402, w_189_404, w_189_406, w_189_407, w_189_408, w_189_409, w_189_414, w_189_417, w_189_418, w_189_420, w_189_421, w_189_423, w_189_424, w_189_425, w_189_428, w_189_430, w_189_431, w_189_432, w_189_435, w_189_436, w_189_437, w_189_438, w_189_440, w_189_441, w_189_442, w_189_443, w_189_444, w_189_445, w_189_447, w_189_449, w_189_450, w_189_451, w_189_452, w_189_453, w_189_455, w_189_456, w_189_458, w_189_459, w_189_461, w_189_462, w_189_464, w_189_465, w_189_466, w_189_467, w_189_468, w_189_469, w_189_471, w_189_475, w_189_476, w_189_477, w_189_478, w_189_479, w_189_480, w_189_485, w_189_486, w_189_488, w_189_489, w_189_490, w_189_491, w_189_492, w_189_493, w_189_494, w_189_496, w_189_501, w_189_504, w_189_505, w_189_507, w_189_509, w_189_510, w_189_511, w_189_512, w_189_513, w_189_514, w_189_516, w_189_517, w_189_518, w_189_520, w_189_521, w_189_523, w_189_524, w_189_525, w_189_528, w_189_529, w_189_530, w_189_533, w_189_536, w_189_539, w_189_540, w_189_541, w_189_542, w_189_543, w_189_544, w_189_545, w_189_547, w_189_548, w_189_550, w_189_551, w_189_554, w_189_555, w_189_556, w_189_557, w_189_559, w_189_560, w_189_562, w_189_563, w_189_565, w_189_567, w_189_570, w_189_571, w_189_572, w_189_574, w_189_575, w_189_576, w_189_577, w_189_579, w_189_582, w_189_583, w_189_584, w_189_586, w_189_589, w_189_590, w_189_591, w_189_592, w_189_593, w_189_595, w_189_597, w_189_598, w_189_599, w_189_602, w_189_603, w_189_605, w_189_609, w_189_610, w_189_613, w_189_614, w_189_615, w_189_617, w_189_618, w_189_621, w_189_622, w_189_623, w_189_624, w_189_625, w_189_626, w_189_628, w_189_629, w_189_631, w_189_632, w_189_633, w_189_634, w_189_635, w_189_636, w_189_641, w_189_642, w_189_644, w_189_649, w_189_650, w_189_651, w_189_652, w_189_653, w_189_655, w_189_656, w_189_658, w_189_660, w_189_661, w_189_663, w_189_664, w_189_665, w_189_667, w_189_668, w_189_672, w_189_675, w_189_676, w_189_678, w_189_680, w_189_682, w_189_683, w_189_686, w_189_689, w_189_692, w_189_697, w_189_699, w_189_702, w_189_706, w_189_707, w_189_708, w_189_709, w_189_711, w_189_712, w_189_714, w_189_716, w_189_718, w_189_719, w_189_721, w_189_722, w_189_723, w_189_724, w_189_725, w_189_726, w_189_727, w_189_728, w_189_729, w_189_730;
  wire w_190_004, w_190_013, w_190_014, w_190_015, w_190_016, w_190_019, w_190_028, w_190_030, w_190_036, w_190_037, w_190_062, w_190_081, w_190_084, w_190_095, w_190_099, w_190_103, w_190_107, w_190_113, w_190_118, w_190_119, w_190_124, w_190_131, w_190_152, w_190_154, w_190_161, w_190_165, w_190_167, w_190_173, w_190_176, w_190_181, w_190_182, w_190_192, w_190_193, w_190_206, w_190_207, w_190_210, w_190_212, w_190_213, w_190_216, w_190_217, w_190_224, w_190_230, w_190_233, w_190_234, w_190_250, w_190_254, w_190_255, w_190_257, w_190_264, w_190_266, w_190_268, w_190_274, w_190_277, w_190_279, w_190_280, w_190_284, w_190_287, w_190_303, w_190_304, w_190_305, w_190_308, w_190_311, w_190_312, w_190_327, w_190_334, w_190_336, w_190_341, w_190_346, w_190_350, w_190_354, w_190_355, w_190_358, w_190_369, w_190_374, w_190_381, w_190_385, w_190_388, w_190_389, w_190_397, w_190_400, w_190_402, w_190_405, w_190_406, w_190_411, w_190_415, w_190_416, w_190_417, w_190_423, w_190_425, w_190_426, w_190_432, w_190_433, w_190_435, w_190_436, w_190_441, w_190_442, w_190_449, w_190_450, w_190_453, w_190_454, w_190_459, w_190_464, w_190_466, w_190_468, w_190_472, w_190_474, w_190_478, w_190_479, w_190_488, w_190_497, w_190_501, w_190_505, w_190_506, w_190_508, w_190_510, w_190_511, w_190_512, w_190_513, w_190_519, w_190_522, w_190_528, w_190_539, w_190_543, w_190_545, w_190_547, w_190_548, w_190_550, w_190_555, w_190_562, w_190_564, w_190_565, w_190_569, w_190_571, w_190_574, w_190_575, w_190_576, w_190_577, w_190_580, w_190_582, w_190_592, w_190_593, w_190_597, w_190_603, w_190_608, w_190_612, w_190_613, w_190_621, w_190_628, w_190_629, w_190_632, w_190_634, w_190_642, w_190_647, w_190_652, w_190_658, w_190_660, w_190_662, w_190_663, w_190_664, w_190_668, w_190_671, w_190_672, w_190_674, w_190_676, w_190_678, w_190_682, w_190_685, w_190_687, w_190_691, w_190_692, w_190_700, w_190_701, w_190_704, w_190_705, w_190_709, w_190_711, w_190_713, w_190_717, w_190_718, w_190_720, w_190_725, w_190_732, w_190_734, w_190_735, w_190_744, w_190_753, w_190_762, w_190_764, w_190_773, w_190_776, w_190_791, w_190_808, w_190_809, w_190_812, w_190_815, w_190_820, w_190_821, w_190_822, w_190_825, w_190_827, w_190_837, w_190_840, w_190_844, w_190_851, w_190_854, w_190_855, w_190_859, w_190_862, w_190_866, w_190_878, w_190_881, w_190_891, w_190_896, w_190_899, w_190_903, w_190_918, w_190_922, w_190_925, w_190_926, w_190_943, w_190_951, w_190_953, w_190_955, w_190_956, w_190_960, w_190_963, w_190_964, w_190_972, w_190_977, w_190_978, w_190_984, w_190_988, w_190_991, w_190_998, w_190_1001, w_190_1006, w_190_1009, w_190_1011, w_190_1012, w_190_1023, w_190_1024, w_190_1027, w_190_1029, w_190_1031, w_190_1035, w_190_1036, w_190_1038, w_190_1039, w_190_1042, w_190_1046, w_190_1064, w_190_1066, w_190_1068, w_190_1076, w_190_1081, w_190_1085, w_190_1101, w_190_1105, w_190_1117, w_190_1118, w_190_1128, w_190_1131, w_190_1132, w_190_1140, w_190_1141, w_190_1146, w_190_1168, w_190_1170, w_190_1171, w_190_1186, w_190_1187, w_190_1189, w_190_1191, w_190_1194, w_190_1202, w_190_1205, w_190_1209, w_190_1211, w_190_1213, w_190_1222, w_190_1224, w_190_1235, w_190_1238, w_190_1242, w_190_1245, w_190_1248, w_190_1249, w_190_1250, w_190_1252, w_190_1254, w_190_1257, w_190_1261, w_190_1278, w_190_1281, w_190_1282, w_190_1283, w_190_1292, w_190_1298, w_190_1301, w_190_1303, w_190_1304, w_190_1306, w_190_1308, w_190_1310, w_190_1317, w_190_1327, w_190_1328, w_190_1332, w_190_1336, w_190_1339, w_190_1342, w_190_1345, w_190_1346, w_190_1347, w_190_1355, w_190_1368, w_190_1370, w_190_1372, w_190_1379, w_190_1383, w_190_1388, w_190_1392, w_190_1397, w_190_1400, w_190_1407, w_190_1417, w_190_1420, w_190_1423, w_190_1428, w_190_1439, w_190_1440, w_190_1445, w_190_1451, w_190_1460, w_190_1468, w_190_1472, w_190_1476, w_190_1483, w_190_1488, w_190_1495, w_190_1501, w_190_1507, w_190_1511, w_190_1512, w_190_1520, w_190_1524, w_190_1525, w_190_1542, w_190_1544, w_190_1547, w_190_1548, w_190_1549, w_190_1551, w_190_1552, w_190_1558, w_190_1559, w_190_1563, w_190_1570, w_190_1576, w_190_1577, w_190_1579, w_190_1583, w_190_1584, w_190_1592, w_190_1593, w_190_1598, w_190_1601, w_190_1604, w_190_1608, w_190_1612, w_190_1615, w_190_1616, w_190_1618, w_190_1625, w_190_1630, w_190_1634, w_190_1637, w_190_1639, w_190_1649, w_190_1653, w_190_1662, w_190_1675, w_190_1682, w_190_1683, w_190_1688, w_190_1692, w_190_1699, w_190_1702, w_190_1703, w_190_1704, w_190_1708, w_190_1709, w_190_1712, w_190_1729, w_190_1738, w_190_1739, w_190_1742, w_190_1743, w_190_1746, w_190_1748, w_190_1755, w_190_1758, w_190_1759, w_190_1769, w_190_1770, w_190_1778, w_190_1782, w_190_1793, w_190_1794, w_190_1795, w_190_1797, w_190_1798, w_190_1803, w_190_1807, w_190_1810, w_190_1816, w_190_1819, w_190_1820, w_190_1822, w_190_1823, w_190_1827, w_190_1829, w_190_1831, w_190_1835, w_190_1836, w_190_1842, w_190_1854, w_190_1855, w_190_1864, w_190_1865, w_190_1876, w_190_1877, w_190_1883, w_190_1892, w_190_1894, w_190_1905, w_190_1907, w_190_1908, w_190_1911, w_190_1913, w_190_1917, w_190_1919, w_190_1925, w_190_1926, w_190_1927, w_190_1928, w_190_1929, w_190_1930, w_190_1948, w_190_1954, w_190_1955, w_190_1960, w_190_1964, w_190_1973, w_190_1980, w_190_1983, w_190_1984, w_190_1986, w_190_1987, w_190_1989, w_190_1990, w_190_1992, w_190_1999, w_190_2000, w_190_2007, w_190_2009, w_190_2013, w_190_2017, w_190_2026, w_190_2027, w_190_2032, w_190_2033, w_190_2034, w_190_2036, w_190_2038, w_190_2039, w_190_2044, w_190_2046, w_190_2053, w_190_2055, w_190_2061, w_190_2064, w_190_2068, w_190_2069, w_190_2072, w_190_2080, w_190_2087, w_190_2095, w_190_2101, w_190_2104, w_190_2105, w_190_2109, w_190_2113, w_190_2117, w_190_2120, w_190_2122, w_190_2124, w_190_2125, w_190_2129, w_190_2137, w_190_2139, w_190_2159, w_190_2171, w_190_2176, w_190_2190, w_190_2201, w_190_2209, w_190_2212, w_190_2229, w_190_2232, w_190_2235, w_190_2241, w_190_2242, w_190_2244, w_190_2259, w_190_2297, w_190_2310, w_190_2311, w_190_2325, w_190_2349, w_190_2350, w_190_2360, w_190_2368, w_190_2380, w_190_2383, w_190_2397, w_190_2401, w_190_2409, w_190_2414, w_190_2419, w_190_2430, w_190_2438, w_190_2445, w_190_2448, w_190_2454, w_190_2486, w_190_2487, w_190_2491, w_190_2493, w_190_2497, w_190_2519, w_190_2520, w_190_2523, w_190_2534, w_190_2538, w_190_2539, w_190_2541, w_190_2583, w_190_2591, w_190_2600, w_190_2611, w_190_2616, w_190_2621, w_190_2638, w_190_2639, w_190_2642, w_190_2659, w_190_2667, w_190_2669, w_190_2673, w_190_2698, w_190_2705, w_190_2711, w_190_2715, w_190_2719, w_190_2732, w_190_2741, w_190_2746, w_190_2771, w_190_2773, w_190_2776, w_190_2793, w_190_2805, w_190_2806, w_190_2809, w_190_2815, w_190_2819, w_190_2824, w_190_2825, w_190_2826, w_190_2827, w_190_2828, w_190_2829, w_190_2830, w_190_2831, w_190_2832, w_190_2833, w_190_2835, w_190_2837, w_190_2838, w_190_2839, w_190_2840, w_190_2841, w_190_2842, w_190_2843, w_190_2845;
  wire w_191_003, w_191_005, w_191_007, w_191_009, w_191_011, w_191_012, w_191_016, w_191_019, w_191_024, w_191_025, w_191_029, w_191_030, w_191_032, w_191_034, w_191_037, w_191_040, w_191_047, w_191_049, w_191_050, w_191_051, w_191_057, w_191_058, w_191_061, w_191_066, w_191_071, w_191_072, w_191_074, w_191_075, w_191_082, w_191_088, w_191_091, w_191_094, w_191_095, w_191_099, w_191_103, w_191_104, w_191_110, w_191_113, w_191_121, w_191_122, w_191_123, w_191_129, w_191_131, w_191_133, w_191_134, w_191_136, w_191_138, w_191_139, w_191_142, w_191_147, w_191_150, w_191_154, w_191_172, w_191_178, w_191_180, w_191_191, w_191_195, w_191_199, w_191_204, w_191_205, w_191_207, w_191_217, w_191_223, w_191_226, w_191_229, w_191_237, w_191_243, w_191_250, w_191_253, w_191_257, w_191_260, w_191_266, w_191_270, w_191_271, w_191_278, w_191_283, w_191_285, w_191_289, w_191_293, w_191_297, w_191_301, w_191_304, w_191_306, w_191_311, w_191_317, w_191_329, w_191_333, w_191_336, w_191_338, w_191_340, w_191_341, w_191_344, w_191_345, w_191_346, w_191_349, w_191_352, w_191_356, w_191_359, w_191_366, w_191_374, w_191_377, w_191_384, w_191_395, w_191_398, w_191_400, w_191_404, w_191_405, w_191_409, w_191_412, w_191_413, w_191_415, w_191_423, w_191_427, w_191_431, w_191_433, w_191_435, w_191_436, w_191_438, w_191_445, w_191_446, w_191_447, w_191_450, w_191_454, w_191_461, w_191_464, w_191_467, w_191_468, w_191_472, w_191_474, w_191_477, w_191_479, w_191_483, w_191_487, w_191_488, w_191_496, w_191_509, w_191_513, w_191_515, w_191_534, w_191_541, w_191_544, w_191_545, w_191_546, w_191_551, w_191_552, w_191_594, w_191_600, w_191_605, w_191_608, w_191_617, w_191_631, w_191_638, w_191_640, w_191_647, w_191_660, w_191_663, w_191_687, w_191_699, w_191_723, w_191_725, w_191_729, w_191_733, w_191_738, w_191_755, w_191_757, w_191_759, w_191_767, w_191_771, w_191_800, w_191_801, w_191_828, w_191_832, w_191_833, w_191_874, w_191_880, w_191_890, w_191_904, w_191_912, w_191_916, w_191_919, w_191_922, w_191_937, w_191_949, w_191_969, w_191_970, w_191_976, w_191_979, w_191_981, w_191_986, w_191_991, w_191_996, w_191_1002, w_191_1006, w_191_1011, w_191_1013, w_191_1014, w_191_1030, w_191_1048, w_191_1054, w_191_1061, w_191_1066, w_191_1074, w_191_1079, w_191_1084, w_191_1088, w_191_1094, w_191_1101, w_191_1112, w_191_1116, w_191_1122, w_191_1123, w_191_1126, w_191_1132, w_191_1133, w_191_1143, w_191_1155, w_191_1157, w_191_1158, w_191_1162, w_191_1169, w_191_1171, w_191_1174, w_191_1184, w_191_1186, w_191_1188, w_191_1190, w_191_1204, w_191_1211, w_191_1221, w_191_1229, w_191_1234, w_191_1245, w_191_1247, w_191_1252, w_191_1253, w_191_1279, w_191_1296, w_191_1303, w_191_1325, w_191_1337, w_191_1349, w_191_1353, w_191_1357, w_191_1360, w_191_1367, w_191_1370, w_191_1373, w_191_1375, w_191_1380, w_191_1382, w_191_1385, w_191_1408, w_191_1413, w_191_1420, w_191_1429, w_191_1431, w_191_1445, w_191_1462, w_191_1463, w_191_1464, w_191_1474, w_191_1475, w_191_1481, w_191_1488, w_191_1492, w_191_1500, w_191_1508, w_191_1515, w_191_1522, w_191_1529, w_191_1531, w_191_1563, w_191_1570, w_191_1579, w_191_1591, w_191_1593, w_191_1643, w_191_1655, w_191_1656, w_191_1658, w_191_1668, w_191_1672, w_191_1678, w_191_1679, w_191_1696, w_191_1702, w_191_1708, w_191_1710, w_191_1712, w_191_1724, w_191_1755, w_191_1758, w_191_1780, w_191_1793, w_191_1801, w_191_1813, w_191_1815, w_191_1825, w_191_1828, w_191_1832, w_191_1838, w_191_1849, w_191_1856, w_191_1870, w_191_1878, w_191_1883, w_191_1887, w_191_1890, w_191_1892, w_191_1898, w_191_1917, w_191_1919, w_191_1923, w_191_1934, w_191_1936, w_191_1941, w_191_1945, w_191_1972, w_191_1975, w_191_1984, w_191_1988, w_191_1993, w_191_1995, w_191_1997, w_191_1998, w_191_2008, w_191_2012, w_191_2019, w_191_2025, w_191_2029, w_191_2031, w_191_2032, w_191_2033, w_191_2039, w_191_2042, w_191_2047, w_191_2051, w_191_2058, w_191_2059, w_191_2071, w_191_2079, w_191_2100, w_191_2102, w_191_2123, w_191_2127, w_191_2131, w_191_2146, w_191_2147, w_191_2158, w_191_2165, w_191_2180, w_191_2182, w_191_2199, w_191_2200, w_191_2209, w_191_2217, w_191_2218, w_191_2222, w_191_2232, w_191_2235, w_191_2237, w_191_2244, w_191_2260, w_191_2261, w_191_2269, w_191_2270, w_191_2271, w_191_2287, w_191_2297, w_191_2302, w_191_2304, w_191_2311, w_191_2314, w_191_2317, w_191_2324, w_191_2326, w_191_2348, w_191_2351, w_191_2358, w_191_2366, w_191_2370, w_191_2387, w_191_2391, w_191_2397, w_191_2404, w_191_2417, w_191_2425, w_191_2427, w_191_2429, w_191_2436, w_191_2449, w_191_2463, w_191_2468, w_191_2472, w_191_2478, w_191_2481, w_191_2489, w_191_2492, w_191_2508, w_191_2534, w_191_2536, w_191_2538, w_191_2543, w_191_2548, w_191_2551, w_191_2554, w_191_2567, w_191_2568, w_191_2571, w_191_2572, w_191_2573, w_191_2584, w_191_2599, w_191_2612, w_191_2619, w_191_2624, w_191_2647, w_191_2651, w_191_2666, w_191_2688, w_191_2696, w_191_2705, w_191_2722, w_191_2729, w_191_2733, w_191_2734, w_191_2755, w_191_2761, w_191_2774, w_191_2791, w_191_2792, w_191_2798, w_191_2892, w_191_2906, w_191_2925, w_191_2927, w_191_2939, w_191_2940, w_191_2952, w_191_2956, w_191_2965, w_191_2975, w_191_2977, w_191_2989, w_191_2999, w_191_3004, w_191_3007, w_191_3018, w_191_3024, w_191_3030, w_191_3040, w_191_3055, w_191_3056, w_191_3063, w_191_3068, w_191_3082, w_191_3083, w_191_3093, w_191_3096, w_191_3099, w_191_3106, w_191_3117, w_191_3124, w_191_3134, w_191_3135, w_191_3136, w_191_3139, w_191_3142, w_191_3146, w_191_3150, w_191_3173, w_191_3179, w_191_3183, w_191_3205, w_191_3208, w_191_3216, w_191_3248, w_191_3253, w_191_3254, w_191_3256, w_191_3260, w_191_3263, w_191_3266, w_191_3285, w_191_3287, w_191_3289, w_191_3293, w_191_3295, w_191_3307, w_191_3309, w_191_3315, w_191_3317, w_191_3320, w_191_3330, w_191_3334, w_191_3346, w_191_3347, w_191_3349, w_191_3351, w_191_3364, w_191_3371, w_191_3376, w_191_3379, w_191_3389, w_191_3391, w_191_3412, w_191_3420, w_191_3426, w_191_3434, w_191_3435, w_191_3440, w_191_3442, w_191_3448, w_191_3457, w_191_3469, w_191_3471, w_191_3473, w_191_3489, w_191_3493, w_191_3498, w_191_3499, w_191_3502, w_191_3503, w_191_3507, w_191_3510, w_191_3511, w_191_3512, w_191_3534, w_191_3545, w_191_3551, w_191_3553, w_191_3560, w_191_3568, w_191_3571, w_191_3573, w_191_3574, w_191_3575, w_191_3579, w_191_3591, w_191_3598, w_191_3610, w_191_3611, w_191_3616, w_191_3622, w_191_3632, w_191_3640, w_191_3644, w_191_3659, w_191_3673, w_191_3681, w_191_3684, w_191_3700, w_191_3726, w_191_3728, w_191_3729, w_191_3739, w_191_3748, w_191_3749, w_191_3752, w_191_3757, w_191_3761, w_191_3762, w_191_3767, w_191_3775, w_191_3784, w_191_3785, w_191_3788, w_191_3792, w_191_3794, w_191_3795, w_191_3796, w_191_3800, w_191_3805, w_191_3829, w_191_3832, w_191_3839, w_191_3840, w_191_3846, w_191_3862, w_191_3863, w_191_3879, w_191_3904, w_191_3909, w_191_3922, w_191_3985, w_191_3997, w_191_4002, w_191_4018, w_191_4022, w_191_4028, w_191_4029, w_191_4038, w_191_4041, w_191_4045, w_191_4071, w_191_4081, w_191_4091, w_191_4099, w_191_4101, w_191_4111, w_191_4127, w_191_4131, w_191_4143, w_191_4150, w_191_4154, w_191_4155, w_191_4160, w_191_4161, w_191_4176, w_191_4181, w_191_4198, w_191_4199, w_191_4206, w_191_4220, w_191_4226, w_191_4250, w_191_4257, w_191_4260, w_191_4264, w_191_4266, w_191_4273, w_191_4284, w_191_4292, w_191_4293, w_191_4298, w_191_4300, w_191_4310, w_191_4316, w_191_4327, w_191_4330, w_191_4337, w_191_4339, w_191_4342, w_191_4344, w_191_4345, w_191_4353, w_191_4356, w_191_4357, w_191_4361, w_191_4367, w_191_4368, w_191_4378, w_191_4387, w_191_4389, w_191_4393, w_191_4399, w_191_4404, w_191_4405, w_191_4406, w_191_4410, w_191_4423, w_191_4427, w_191_4429, w_191_4430, w_191_4435;
  wire w_192_001, w_192_009, w_192_015, w_192_019, w_192_025, w_192_031, w_192_037, w_192_049, w_192_051, w_192_060, w_192_061, w_192_084, w_192_105, w_192_108, w_192_118, w_192_121, w_192_123, w_192_131, w_192_134, w_192_143, w_192_150, w_192_152, w_192_157, w_192_160, w_192_167, w_192_180, w_192_191, w_192_198, w_192_202, w_192_205, w_192_210, w_192_217, w_192_218, w_192_227, w_192_239, w_192_270, w_192_273, w_192_297, w_192_299, w_192_301, w_192_308, w_192_313, w_192_326, w_192_328, w_192_329, w_192_336, w_192_345, w_192_346, w_192_361, w_192_368, w_192_374, w_192_376, w_192_413, w_192_415, w_192_416, w_192_418, w_192_421, w_192_429, w_192_431, w_192_446, w_192_449, w_192_453, w_192_457, w_192_466, w_192_471, w_192_495, w_192_496, w_192_500, w_192_505, w_192_510, w_192_516, w_192_532, w_192_545, w_192_549, w_192_555, w_192_559, w_192_560, w_192_565, w_192_575, w_192_579, w_192_585, w_192_592, w_192_594, w_192_602, w_192_605, w_192_606, w_192_614, w_192_633, w_192_643, w_192_644, w_192_650, w_192_669, w_192_671, w_192_672, w_192_690, w_192_699, w_192_701, w_192_706, w_192_711, w_192_717, w_192_735, w_192_748, w_192_772, w_192_779, w_192_780, w_192_783, w_192_786, w_192_794, w_192_799, w_192_801, w_192_805, w_192_814, w_192_815, w_192_821, w_192_823, w_192_834, w_192_840, w_192_846, w_192_852, w_192_855, w_192_858, w_192_860, w_192_878, w_192_885, w_192_893, w_192_896, w_192_900, w_192_902, w_192_907, w_192_908, w_192_909, w_192_921, w_192_922, w_192_932, w_192_933, w_192_946, w_192_948, w_192_950, w_192_953, w_192_958, w_192_959, w_192_973, w_192_974, w_192_980, w_192_989, w_192_990, w_192_994, w_192_996, w_192_1006, w_192_1011, w_192_1012, w_192_1023, w_192_1030, w_192_1031, w_192_1035, w_192_1036, w_192_1038, w_192_1042, w_192_1053, w_192_1056, w_192_1057, w_192_1059, w_192_1060, w_192_1065, w_192_1085, w_192_1103, w_192_1108, w_192_1111, w_192_1121, w_192_1164, w_192_1168, w_192_1175, w_192_1192, w_192_1199, w_192_1224, w_192_1230, w_192_1239, w_192_1253, w_192_1257, w_192_1270, w_192_1272, w_192_1276, w_192_1277, w_192_1279, w_192_1280, w_192_1285, w_192_1286, w_192_1296, w_192_1307, w_192_1312, w_192_1318, w_192_1319, w_192_1330, w_192_1333, w_192_1344, w_192_1346, w_192_1356, w_192_1371, w_192_1376, w_192_1404, w_192_1405, w_192_1437, w_192_1450, w_192_1459, w_192_1482, w_192_1501, w_192_1506, w_192_1508, w_192_1517, w_192_1546, w_192_1547, w_192_1548, w_192_1563, w_192_1585, w_192_1588, w_192_1604, w_192_1607, w_192_1608, w_192_1612, w_192_1616, w_192_1617, w_192_1625, w_192_1661, w_192_1668, w_192_1674, w_192_1682, w_192_1696, w_192_1699, w_192_1703, w_192_1704, w_192_1706, w_192_1710, w_192_1711, w_192_1732, w_192_1741, w_192_1744, w_192_1748, w_192_1754, w_192_1757, w_192_1760, w_192_1766, w_192_1774, w_192_1776, w_192_1778, w_192_1804, w_192_1821, w_192_1826, w_192_1854, w_192_1918, w_192_1925, w_192_1936, w_192_1942, w_192_1948, w_192_1965, w_192_1969, w_192_1970, w_192_1973, w_192_1983, w_192_1995, w_192_2022, w_192_2025, w_192_2027, w_192_2036, w_192_2044, w_192_2045, w_192_2049, w_192_2055, w_192_2068, w_192_2069, w_192_2074, w_192_2075, w_192_2078, w_192_2087, w_192_2098, w_192_2105, w_192_2106, w_192_2116, w_192_2125, w_192_2130, w_192_2131, w_192_2135, w_192_2139, w_192_2142, w_192_2145, w_192_2162, w_192_2164, w_192_2170, w_192_2173, w_192_2182, w_192_2196, w_192_2206, w_192_2214, w_192_2218, w_192_2221, w_192_2244, w_192_2245, w_192_2259, w_192_2260, w_192_2261, w_192_2264, w_192_2286, w_192_2288, w_192_2297, w_192_2300, w_192_2312, w_192_2313, w_192_2315, w_192_2316, w_192_2318, w_192_2333, w_192_2362, w_192_2366, w_192_2369, w_192_2377, w_192_2389, w_192_2399, w_192_2402, w_192_2412, w_192_2414, w_192_2429, w_192_2442, w_192_2452, w_192_2456, w_192_2463, w_192_2464, w_192_2478, w_192_2487, w_192_2494, w_192_2500, w_192_2502, w_192_2514, w_192_2522, w_192_2523, w_192_2525, w_192_2526, w_192_2529, w_192_2545, w_192_2554, w_192_2567, w_192_2589, w_192_2596, w_192_2608, w_192_2610, w_192_2613, w_192_2616, w_192_2617, w_192_2647, w_192_2648, w_192_2651, w_192_2652, w_192_2656, w_192_2657, w_192_2659, w_192_2665, w_192_2685, w_192_2694, w_192_2695, w_192_2703, w_192_2709, w_192_2714, w_192_2732, w_192_2743, w_192_2762, w_192_2767, w_192_2770, w_192_2771, w_192_2774, w_192_2778, w_192_2788, w_192_2789, w_192_2791, w_192_2796, w_192_2803, w_192_2805, w_192_2807, w_192_2813, w_192_2815, w_192_2826, w_192_2845, w_192_2846, w_192_2851, w_192_2865, w_192_2882, w_192_2887, w_192_2893, w_192_2897, w_192_2899, w_192_2907, w_192_2925, w_192_2930, w_192_2933, w_192_2938, w_192_2947, w_192_2948, w_192_2956, w_192_2959, w_192_2961, w_192_2970, w_192_2987, w_192_2990, w_192_2991, w_192_2992, w_192_3003, w_192_3014, w_192_3016, w_192_3017, w_192_3021, w_192_3024, w_192_3025, w_192_3038, w_192_3044, w_192_3045, w_192_3046, w_192_3057, w_192_3060, w_192_3068, w_192_3069, w_192_3083, w_192_3104, w_192_3117, w_192_3129, w_192_3132, w_192_3146, w_192_3155, w_192_3160, w_192_3163, w_192_3167, w_192_3169, w_192_3172, w_192_3176, w_192_3183, w_192_3188, w_192_3189, w_192_3197, w_192_3202, w_192_3219, w_192_3222, w_192_3227, w_192_3228, w_192_3233, w_192_3235, w_192_3238, w_192_3244, w_192_3247, w_192_3249, w_192_3267, w_192_3269, w_192_3274, w_192_3279, w_192_3287, w_192_3317, w_192_3328, w_192_3331, w_192_3347, w_192_3348, w_192_3350, w_192_3354, w_192_3363, w_192_3364, w_192_3367, w_192_3374, w_192_3381, w_192_3382, w_192_3392, w_192_3403, w_192_3410, w_192_3421, w_192_3449, w_192_3459, w_192_3460, w_192_3461, w_192_3468, w_192_3476, w_192_3483, w_192_3491, w_192_3501, w_192_3513, w_192_3514, w_192_3518, w_192_3529, w_192_3530, w_192_3544, w_192_3552, w_192_3576, w_192_3584, w_192_3585, w_192_3588, w_192_3591, w_192_3595, w_192_3603, w_192_3613, w_192_3624, w_192_3633, w_192_3636, w_192_3645, w_192_3648, w_192_3658, w_192_3665, w_192_3671, w_192_3674, w_192_3701, w_192_3713, w_192_3714, w_192_3720, w_192_3725, w_192_3734, w_192_3738, w_192_3748, w_192_3755, w_192_3763, w_192_3767, w_192_3771, w_192_3774, w_192_3781, w_192_3791, w_192_3795, w_192_3803, w_192_3817, w_192_3820, w_192_3823, w_192_3829, w_192_3851, w_192_3857, w_192_3865, w_192_3873, w_192_3877, w_192_3887, w_192_3892, w_192_3904, w_192_3932, w_192_3933, w_192_3952, w_192_3957, w_192_3964, w_192_4019, w_192_4022, w_192_4025, w_192_4027, w_192_4040, w_192_4041, w_192_4053, w_192_4055, w_192_4062, w_192_4079, w_192_4093, w_192_4100, w_192_4109, w_192_4112, w_192_4115, w_192_4121, w_192_4125, w_192_4147, w_192_4161, w_192_4174, w_192_4183, w_192_4244, w_192_4251, w_192_4256, w_192_4264, w_192_4269, w_192_4274, w_192_4284, w_192_4289, w_192_4292, w_192_4307, w_192_4318, w_192_4323, w_192_4339, w_192_4343, w_192_4352, w_192_4365, w_192_4370, w_192_4374, w_192_4394, w_192_4396, w_192_4409, w_192_4411, w_192_4420, w_192_4424, w_192_4440, w_192_4444, w_192_4451, w_192_4457, w_192_4461, w_192_4471, w_192_4481, w_192_4487, w_192_4488, w_192_4492, w_192_4496, w_192_4498, w_192_4510, w_192_4511, w_192_4528, w_192_4531, w_192_4532, w_192_4539, w_192_4549, w_192_4551, w_192_4562, w_192_4574, w_192_4582, w_192_4586, w_192_4596, w_192_4601, w_192_4604, w_192_4611, w_192_4621, w_192_4622, w_192_4629, w_192_4638, w_192_4641, w_192_4644, w_192_4658, w_192_4667, w_192_4674, w_192_4675, w_192_4681, w_192_4695, w_192_4702, w_192_4715, w_192_4717, w_192_4724, w_192_4726, w_192_4731, w_192_4732, w_192_4742, w_192_4759, w_192_4797, w_192_4831, w_192_4835, w_192_4836, w_192_4837, w_192_4839, w_192_4840, w_192_4848, w_192_4859, w_192_4863, w_192_4865, w_192_4869, w_192_4870, w_192_4871, w_192_4885, w_192_4886, w_192_4888, w_192_4891, w_192_4897, w_192_4902, w_192_4905, w_192_4914, w_192_4915, w_192_4916, w_192_4927, w_192_4939, w_192_4948, w_192_4954, w_192_4960, w_192_4961, w_192_4962, w_192_4963, w_192_4964, w_192_4965, w_192_4969, w_192_4970, w_192_4971, w_192_4972, w_192_4973, w_192_4974, w_192_4975, w_192_4976, w_192_4977, w_192_4978, w_192_4979, w_192_4980, w_192_4982;
  wire w_193_001, w_193_002, w_193_004, w_193_005, w_193_006, w_193_011, w_193_013, w_193_015, w_193_020, w_193_022, w_193_025, w_193_030, w_193_032, w_193_043, w_193_046, w_193_058, w_193_060, w_193_061, w_193_063, w_193_066, w_193_070, w_193_074, w_193_077, w_193_083, w_193_084, w_193_085, w_193_087, w_193_091, w_193_092, w_193_094, w_193_097, w_193_099, w_193_101, w_193_116, w_193_117, w_193_121, w_193_127, w_193_128, w_193_129, w_193_130, w_193_131, w_193_133, w_193_136, w_193_138, w_193_141, w_193_142, w_193_144, w_193_148, w_193_149, w_193_159, w_193_160, w_193_162, w_193_163, w_193_165, w_193_173, w_193_176, w_193_178, w_193_181, w_193_184, w_193_186, w_193_190, w_193_196, w_193_199, w_193_200, w_193_203, w_193_205, w_193_207, w_193_210, w_193_212, w_193_214, w_193_217, w_193_223, w_193_226, w_193_228, w_193_236, w_193_238, w_193_239, w_193_241, w_193_250, w_193_255, w_193_256, w_193_262, w_193_270, w_193_273, w_193_275, w_193_284, w_193_293, w_193_294, w_193_295, w_193_300, w_193_302, w_193_306, w_193_308, w_193_320, w_193_334, w_193_341, w_193_342, w_193_344, w_193_352, w_193_354, w_193_358, w_193_360, w_193_365, w_193_369, w_193_375, w_193_377, w_193_381, w_193_384, w_193_386, w_193_391, w_193_398, w_193_401, w_193_402, w_193_416, w_193_419, w_193_424, w_193_425, w_193_434, w_193_436, w_193_440, w_193_441, w_193_446, w_193_449, w_193_451, w_193_457, w_193_467, w_193_469, w_193_470, w_193_472, w_193_475, w_193_477, w_193_480, w_193_484, w_193_487, w_193_488, w_193_489, w_193_491, w_193_492, w_193_497, w_193_500, w_193_504, w_193_505, w_193_508, w_193_514, w_193_517, w_193_520, w_193_525, w_193_528, w_193_533, w_193_534, w_193_541, w_193_547, w_193_550, w_193_551, w_193_554, w_193_560, w_193_564, w_193_567, w_193_574, w_193_576, w_193_578, w_193_579, w_193_580, w_193_582, w_193_586, w_193_597, w_193_598, w_193_609, w_193_610, w_193_615, w_193_620, w_193_623, w_193_624, w_193_630, w_193_634, w_193_637, w_193_639, w_193_644, w_193_654, w_193_655, w_193_660, w_193_666, w_193_669, w_193_673, w_193_679, w_193_686, w_193_687, w_193_688, w_193_689, w_193_692, w_193_694, w_193_696, w_193_698, w_193_708, w_193_713, w_193_717, w_193_722, w_193_724, w_193_725, w_193_730, w_193_733, w_193_735, w_193_738, w_193_739, w_193_743, w_193_747, w_193_749, w_193_752, w_193_753, w_193_754, w_193_762, w_193_764, w_193_776, w_193_781, w_193_785, w_193_786, w_193_787, w_193_794, w_193_800, w_193_807, w_193_808, w_193_814, w_193_820, w_193_821, w_193_822, w_193_824, w_193_827, w_193_840, w_193_847, w_193_848, w_193_850, w_193_853, w_193_855, w_193_858, w_193_859, w_193_863, w_193_865, w_193_870, w_193_875, w_193_876, w_193_879, w_193_880, w_193_887, w_193_888, w_193_890, w_193_891, w_193_893, w_193_902, w_193_913, w_193_914, w_193_917, w_193_918, w_193_919, w_193_921, w_193_923, w_193_928, w_193_932, w_193_937, w_193_942, w_193_956, w_193_957, w_193_958, w_193_961, w_193_963, w_193_966, w_193_967, w_193_975, w_193_977, w_193_979, w_193_985, w_193_986, w_193_989, w_193_992, w_193_1001, w_193_1004, w_193_1008, w_193_1024, w_193_1028, w_193_1031, w_193_1034, w_193_1038, w_193_1043, w_193_1048, w_193_1051, w_193_1052, w_193_1056, w_193_1057, w_193_1061, w_193_1065, w_193_1068, w_193_1072, w_193_1073, w_193_1081, w_193_1085, w_193_1088, w_193_1090, w_193_1093, w_193_1094, w_193_1101, w_193_1104, w_193_1106, w_193_1112, w_193_1114, w_193_1117, w_193_1121, w_193_1133, w_193_1142, w_193_1146, w_193_1147, w_193_1154, w_193_1158, w_193_1164, w_193_1175, w_193_1176, w_193_1177, w_193_1179, w_193_1183, w_193_1188, w_193_1199, w_193_1200, w_193_1201, w_193_1202, w_193_1210, w_193_1212, w_193_1230, w_193_1234, w_193_1243, w_193_1244, w_193_1257, w_193_1258, w_193_1259, w_193_1260, w_193_1261, w_193_1263, w_193_1264, w_193_1266, w_193_1272, w_193_1274, w_193_1277, w_193_1281, w_193_1282, w_193_1288, w_193_1289, w_193_1291, w_193_1292, w_193_1296, w_193_1297, w_193_1311, w_193_1317, w_193_1320, w_193_1327, w_193_1328, w_193_1330, w_193_1333, w_193_1334, w_193_1346, w_193_1349, w_193_1354, w_193_1356, w_193_1357, w_193_1365, w_193_1368, w_193_1370, w_193_1377, w_193_1384, w_193_1386, w_193_1387, w_193_1388, w_193_1397, w_193_1400, w_193_1414, w_193_1416, w_193_1418, w_193_1419, w_193_1421, w_193_1428, w_193_1433, w_193_1435, w_193_1439, w_193_1441, w_193_1444, w_193_1446, w_193_1447, w_193_1463, w_193_1470, w_193_1474, w_193_1475, w_193_1477, w_193_1478, w_193_1479, w_193_1485, w_193_1487, w_193_1490, w_193_1495, w_193_1507, w_193_1510, w_193_1512, w_193_1516, w_193_1517, w_193_1523, w_193_1530, w_193_1531, w_193_1533, w_193_1534, w_193_1537, w_193_1543, w_193_1544, w_193_1548, w_193_1549, w_193_1553, w_193_1554, w_193_1557, w_193_1560, w_193_1564, w_193_1573, w_193_1587, w_193_1590, w_193_1592, w_193_1603, w_193_1604, w_193_1609, w_193_1615, w_193_1616, w_193_1618, w_193_1625, w_193_1626, w_193_1634, w_193_1635, w_193_1644, w_193_1646, w_193_1648, w_193_1651, w_193_1656, w_193_1660, w_193_1662, w_193_1667, w_193_1668, w_193_1677, w_193_1686, w_193_1689, w_193_1692, w_193_1700, w_193_1706, w_193_1712, w_193_1714, w_193_1715, w_193_1721, w_193_1738, w_193_1743, w_193_1747, w_193_1760, w_193_1761, w_193_1765, w_193_1766, w_193_1767, w_193_1768, w_193_1769, w_193_1777, w_193_1796, w_193_1798, w_193_1818, w_193_1822, w_193_1830, w_193_1831, w_193_1838, w_193_1843, w_193_1846, w_193_1894, w_193_1897, w_193_1898, w_193_1900, w_193_1926, w_193_1936, w_193_1940, w_193_1942, w_193_1958, w_193_1961, w_193_1968, w_193_1975, w_193_1985, w_193_1986, w_193_1988, w_193_2001, w_193_2022, w_193_2023, w_193_2029, w_193_2043, w_193_2045, w_193_2058, w_193_2066, w_193_2075, w_193_2077, w_193_2100, w_193_2101, w_193_2120, w_193_2122, w_193_2125, w_193_2126, w_193_2128, w_193_2143, w_193_2154, w_193_2163, w_193_2173, w_193_2180, w_193_2187, w_193_2214, w_193_2216, w_193_2229, w_193_2238, w_193_2241, w_193_2242, w_193_2243, w_193_2245, w_193_2276, w_193_2284, w_193_2289, w_193_2299, w_193_2303, w_193_2309, w_193_2317, w_193_2327, w_193_2328, w_193_2345, w_193_2347, w_193_2377, w_193_2383, w_193_2386, w_193_2390, w_193_2404, w_193_2408, w_193_2409, w_193_2410, w_193_2416, w_193_2424, w_193_2425, w_193_2450, w_193_2452, w_193_2455, w_193_2471, w_193_2487, w_193_2509, w_193_2517, w_193_2519, w_193_2524, w_193_2525, w_193_2531, w_193_2533, w_193_2537, w_193_2541, w_193_2565, w_193_2571, w_193_2580, w_193_2581, w_193_2595, w_193_2602, w_193_2611, w_193_2612, w_193_2622, w_193_2629, w_193_2639, w_193_2641, w_193_2648, w_193_2662, w_193_2665, w_193_2683, w_193_2702, w_193_2712, w_193_2719, w_193_2731, w_193_2737, w_193_2747, w_193_2749, w_193_2760, w_193_2778, w_193_2779, w_193_2789, w_193_2809, w_193_2810, w_193_2839, w_193_2848, w_193_2852, w_193_2853, w_193_2861, w_193_2874, w_193_2876, w_193_2880, w_193_2887, w_193_2893, w_193_2909, w_193_2910, w_193_2914, w_193_2915, w_193_2919, w_193_2925, w_193_2930, w_193_2939, w_193_2952, w_193_2963, w_193_2964, w_193_2983, w_193_2986, w_193_2987, w_193_2996, w_193_3002, w_193_3008, w_193_3020, w_193_3023, w_193_3029, w_193_3030, w_193_3033, w_193_3049, w_193_3076, w_193_3118, w_193_3122, w_193_3124, w_193_3136, w_193_3138, w_193_3140, w_193_3149, w_193_3152, w_193_3153, w_193_3161, w_193_3175, w_193_3177, w_193_3181, w_193_3203, w_193_3205, w_193_3207, w_193_3211, w_193_3214, w_193_3216, w_193_3221, w_193_3228, w_193_3238, w_193_3249, w_193_3254, w_193_3255;
  wire w_194_005, w_194_011, w_194_018, w_194_021, w_194_022, w_194_023, w_194_027, w_194_029, w_194_030, w_194_031, w_194_034, w_194_035, w_194_038, w_194_039, w_194_040, w_194_042, w_194_048, w_194_053, w_194_060, w_194_068, w_194_075, w_194_076, w_194_081, w_194_082, w_194_084, w_194_091, w_194_095, w_194_099, w_194_102, w_194_103, w_194_109, w_194_110, w_194_112, w_194_118, w_194_122, w_194_128, w_194_133, w_194_136, w_194_138, w_194_146, w_194_148, w_194_153, w_194_158, w_194_161, w_194_165, w_194_167, w_194_168, w_194_171, w_194_185, w_194_188, w_194_189, w_194_199, w_194_203, w_194_209, w_194_210, w_194_221, w_194_227, w_194_233, w_194_234, w_194_243, w_194_244, w_194_246, w_194_251, w_194_252, w_194_269, w_194_273, w_194_274, w_194_278, w_194_281, w_194_283, w_194_285, w_194_289, w_194_294, w_194_297, w_194_298, w_194_299, w_194_305, w_194_309, w_194_313, w_194_314, w_194_317, w_194_318, w_194_321, w_194_323, w_194_326, w_194_329, w_194_330, w_194_339, w_194_347, w_194_352, w_194_355, w_194_362, w_194_363, w_194_364, w_194_376, w_194_381, w_194_383, w_194_387, w_194_397, w_194_400, w_194_402, w_194_405, w_194_406, w_194_410, w_194_413, w_194_419, w_194_425, w_194_426, w_194_429, w_194_430, w_194_439, w_194_441, w_194_448, w_194_451, w_194_459, w_194_463, w_194_466, w_194_470, w_194_478, w_194_479, w_194_480, w_194_481, w_194_482, w_194_483, w_194_486, w_194_487, w_194_489, w_194_495, w_194_497, w_194_500, w_194_504, w_194_508, w_194_510, w_194_514, w_194_515, w_194_523, w_194_528, w_194_531, w_194_539, w_194_543, w_194_544, w_194_550, w_194_551, w_194_552, w_194_554, w_194_557, w_194_561, w_194_570, w_194_575, w_194_578, w_194_584, w_194_585, w_194_589, w_194_590, w_194_595, w_194_597, w_194_602, w_194_605, w_194_606, w_194_607, w_194_609, w_194_611, w_194_612, w_194_616, w_194_621, w_194_624, w_194_626, w_194_634, w_194_638, w_194_640, w_194_645, w_194_646, w_194_649, w_194_653, w_194_654, w_194_657, w_194_660, w_194_661, w_194_665, w_194_674, w_194_676, w_194_682, w_194_688, w_194_691, w_194_695, w_194_700, w_194_701, w_194_703, w_194_707, w_194_709, w_194_710, w_194_717, w_194_720, w_194_729, w_194_735, w_194_749, w_194_751, w_194_753, w_194_754, w_194_755, w_194_761, w_194_771, w_194_773, w_194_775, w_194_776, w_194_777, w_194_782, w_194_788, w_194_790, w_194_793, w_194_796, w_194_810, w_194_813, w_194_817, w_194_818, w_194_819, w_194_820, w_194_821, w_194_823, w_194_824, w_194_825, w_194_827, w_194_837, w_194_838, w_194_839, w_194_841, w_194_843, w_194_847, w_194_851, w_194_857, w_194_862, w_194_865, w_194_867, w_194_868, w_194_871, w_194_875, w_194_876, w_194_877, w_194_878, w_194_886, w_194_887, w_194_891, w_194_895, w_194_896, w_194_902, w_194_903, w_194_907, w_194_909, w_194_917, w_194_928, w_194_930, w_194_931, w_194_935, w_194_942, w_194_945, w_194_947, w_194_949, w_194_952, w_194_973, w_194_977, w_194_978, w_194_986, w_194_990, w_194_993, w_194_994, w_194_1000, w_194_1010, w_194_1011, w_194_1012, w_194_1013, w_194_1023, w_194_1029, w_194_1030, w_194_1033, w_194_1048, w_194_1049, w_194_1052, w_194_1066, w_194_1067, w_194_1078, w_194_1080, w_194_1108, w_194_1114, w_194_1117, w_194_1122, w_194_1123, w_194_1128, w_194_1159, w_194_1160, w_194_1165, w_194_1170, w_194_1190, w_194_1207, w_194_1208, w_194_1214, w_194_1225, w_194_1229, w_194_1233, w_194_1237, w_194_1254, w_194_1275, w_194_1278, w_194_1293, w_194_1319, w_194_1323, w_194_1326, w_194_1332, w_194_1339, w_194_1346, w_194_1348, w_194_1349, w_194_1354, w_194_1379, w_194_1385, w_194_1397, w_194_1399, w_194_1405, w_194_1409, w_194_1417, w_194_1422, w_194_1434, w_194_1451, w_194_1452, w_194_1459, w_194_1460, w_194_1466, w_194_1475, w_194_1481, w_194_1485, w_194_1492, w_194_1493, w_194_1496, w_194_1500, w_194_1508, w_194_1509, w_194_1515, w_194_1536, w_194_1545, w_194_1568, w_194_1577, w_194_1591, w_194_1593, w_194_1598, w_194_1609, w_194_1612, w_194_1622, w_194_1638, w_194_1640, w_194_1641, w_194_1642, w_194_1654, w_194_1669, w_194_1672, w_194_1679, w_194_1682, w_194_1716, w_194_1722, w_194_1726, w_194_1751, w_194_1758, w_194_1764, w_194_1776, w_194_1778, w_194_1793, w_194_1811, w_194_1814, w_194_1817, w_194_1823, w_194_1831, w_194_1841, w_194_1861, w_194_1866, w_194_1868, w_194_1883, w_194_1891, w_194_1892, w_194_1906, w_194_1914, w_194_1919, w_194_1924, w_194_1931, w_194_1933, w_194_1949, w_194_1962, w_194_1964, w_194_1965, w_194_1966, w_194_1973, w_194_1985, w_194_1986, w_194_1995, w_194_1998, w_194_1999, w_194_2006, w_194_2016, w_194_2023, w_194_2030, w_194_2032, w_194_2036, w_194_2051, w_194_2061, w_194_2063, w_194_2113, w_194_2118, w_194_2127, w_194_2130, w_194_2132, w_194_2136, w_194_2140, w_194_2150, w_194_2151, w_194_2155, w_194_2156, w_194_2171, w_194_2179, w_194_2190, w_194_2191, w_194_2193, w_194_2195, w_194_2202, w_194_2203, w_194_2209, w_194_2211, w_194_2213, w_194_2215, w_194_2220, w_194_2229, w_194_2237, w_194_2249, w_194_2259, w_194_2261, w_194_2264, w_194_2269, w_194_2283, w_194_2297, w_194_2301, w_194_2311, w_194_2320, w_194_2325, w_194_2326, w_194_2344, w_194_2352, w_194_2358, w_194_2367, w_194_2368, w_194_2373, w_194_2375, w_194_2382, w_194_2414, w_194_2452, w_194_2456, w_194_2458, w_194_2465, w_194_2474, w_194_2485, w_194_2492, w_194_2507, w_194_2515, w_194_2520, w_194_2521, w_194_2533, w_194_2535, w_194_2536, w_194_2540, w_194_2545, w_194_2546, w_194_2550, w_194_2554, w_194_2556, w_194_2559, w_194_2562, w_194_2577, w_194_2578, w_194_2579, w_194_2584, w_194_2585, w_194_2592, w_194_2598, w_194_2602, w_194_2603, w_194_2607, w_194_2609, w_194_2610, w_194_2624, w_194_2643, w_194_2648, w_194_2669, w_194_2678, w_194_2680, w_194_2683, w_194_2685, w_194_2686, w_194_2691, w_194_2703, w_194_2709, w_194_2714, w_194_2717, w_194_2731, w_194_2740, w_194_2741, w_194_2743, w_194_2746, w_194_2756, w_194_2764, w_194_2768, w_194_2772, w_194_2779, w_194_2786, w_194_2795, w_194_2796, w_194_2798, w_194_2804, w_194_2808, w_194_2810, w_194_2825, w_194_2849, w_194_2855, w_194_2857, w_194_2868, w_194_2874, w_194_2879, w_194_2883, w_194_2886, w_194_2889, w_194_2890, w_194_2902, w_194_2905, w_194_2908, w_194_2929, w_194_2936, w_194_2941, w_194_2948, w_194_2951, w_194_2965, w_194_2981, w_194_2987, w_194_2997, w_194_3012, w_194_3024, w_194_3035, w_194_3042, w_194_3043, w_194_3049, w_194_3054, w_194_3060, w_194_3069, w_194_3071, w_194_3086, w_194_3088, w_194_3089, w_194_3090, w_194_3094, w_194_3099, w_194_3108, w_194_3111, w_194_3117, w_194_3118, w_194_3119, w_194_3120, w_194_3122, w_194_3123, w_194_3133, w_194_3136, w_194_3142, w_194_3150, w_194_3153, w_194_3157, w_194_3165, w_194_3166, w_194_3169, w_194_3176, w_194_3187, w_194_3215, w_194_3220, w_194_3224, w_194_3225, w_194_3241, w_194_3243, w_194_3253, w_194_3262, w_194_3277, w_194_3288, w_194_3297, w_194_3303, w_194_3305, w_194_3306, w_194_3322, w_194_3325, w_194_3329, w_194_3340, w_194_3347, w_194_3351, w_194_3356, w_194_3358, w_194_3368, w_194_3370, w_194_3372, w_194_3380, w_194_3387, w_194_3395, w_194_3397, w_194_3420, w_194_3426, w_194_3432, w_194_3440, w_194_3443, w_194_3453, w_194_3457, w_194_3484, w_194_3486, w_194_3518, w_194_3520, w_194_3521, w_194_3529, w_194_3534, w_194_3569, w_194_3574, w_194_3575, w_194_3576, w_194_3588, w_194_3592, w_194_3605, w_194_3606, w_194_3607, w_194_3608, w_194_3609, w_194_3614, w_194_3645, w_194_3669, w_194_3670, w_194_3672, w_194_3673, w_194_3682, w_194_3683, w_194_3697, w_194_3700, w_194_3717, w_194_3722, w_194_3727, w_194_3743, w_194_3746, w_194_3753, w_194_3757, w_194_3759, w_194_3776, w_194_3788, w_194_3799, w_194_3800, w_194_3801, w_194_3821, w_194_3822, w_194_3832, w_194_3834, w_194_3838, w_194_3844, w_194_3846, w_194_3858, w_194_3865, w_194_3866, w_194_3874, w_194_3875, w_194_3884, w_194_3891, w_194_3900, w_194_3915, w_194_3918, w_194_3922, w_194_3950, w_194_3955, w_194_3964, w_194_3966, w_194_3976, w_194_3985, w_194_3992, w_194_4000, w_194_4002, w_194_4003, w_194_4010, w_194_4012, w_194_4033, w_194_4060, w_194_4064, w_194_4070;
  wire w_195_000, w_195_001, w_195_002, w_195_003, w_195_004, w_195_005, w_195_006, w_195_007, w_195_008, w_195_009, w_195_010, w_195_011, w_195_012, w_195_013, w_195_014, w_195_015, w_195_016, w_195_017, w_195_018, w_195_019, w_195_020, w_195_021, w_195_022, w_195_023, w_195_024, w_195_025, w_195_026, w_195_027, w_195_028, w_195_029, w_195_030, w_195_031, w_195_032, w_195_033, w_195_034, w_195_035, w_195_036, w_195_037, w_195_038, w_195_039, w_195_040, w_195_041, w_195_042, w_195_043, w_195_044, w_195_045, w_195_046, w_195_047, w_195_048, w_195_049, w_195_050, w_195_051, w_195_052, w_195_053, w_195_054, w_195_055, w_195_056, w_195_057, w_195_058, w_195_059, w_195_060, w_195_061, w_195_062, w_195_063, w_195_064, w_195_065, w_195_066, w_195_067, w_195_068, w_195_069, w_195_070, w_195_071, w_195_072, w_195_073, w_195_074, w_195_075, w_195_076, w_195_077, w_195_078, w_195_079, w_195_080, w_195_081, w_195_082, w_195_083, w_195_084, w_195_085, w_195_086, w_195_087, w_195_088, w_195_089, w_195_090, w_195_091, w_195_092, w_195_093, w_195_094, w_195_095, w_195_097, w_195_098, w_195_099, w_195_100, w_195_101, w_195_102, w_195_103, w_195_104, w_195_105, w_195_106, w_195_107, w_195_108, w_195_109, w_195_110, w_195_111, w_195_112, w_195_113, w_195_114, w_195_115, w_195_116, w_195_117, w_195_118, w_195_119, w_195_120, w_195_121, w_195_122, w_195_123, w_195_124, w_195_125, w_195_126, w_195_127, w_195_128, w_195_129, w_195_130, w_195_131, w_195_132, w_195_133, w_195_134, w_195_135, w_195_136, w_195_137, w_195_138, w_195_139, w_195_140, w_195_141;
  wire w_196_000, w_196_001, w_196_002, w_196_003, w_196_004, w_196_005, w_196_006, w_196_007, w_196_008, w_196_009, w_196_010, w_196_011, w_196_012, w_196_013, w_196_014, w_196_015, w_196_016, w_196_017, w_196_018, w_196_019, w_196_020, w_196_021, w_196_022, w_196_023, w_196_024, w_196_025, w_196_026, w_196_027, w_196_028, w_196_029, w_196_030, w_196_031, w_196_032, w_196_033, w_196_034, w_196_035, w_196_036, w_196_037, w_196_038, w_196_039, w_196_040, w_196_041, w_196_042, w_196_043, w_196_044, w_196_045, w_196_046, w_196_047, w_196_048, w_196_049, w_196_050, w_196_051, w_196_052, w_196_053, w_196_054, w_196_055, w_196_056, w_196_057, w_196_058, w_196_059, w_196_060, w_196_061, w_196_062, w_196_063, w_196_064, w_196_065, w_196_066, w_196_067, w_196_068, w_196_069, w_196_070, w_196_071, w_196_072, w_196_073, w_196_074, w_196_075, w_196_076, w_196_077, w_196_078, w_196_079, w_196_080, w_196_081, w_196_082, w_196_083, w_196_084, w_196_085, w_196_086, w_196_087, w_196_088, w_196_089, w_196_090, w_196_091, w_196_092, w_196_093, w_196_094, w_196_095, w_196_096, w_196_097, w_196_098, w_196_099, w_196_100, w_196_101, w_196_102, w_196_103, w_196_104, w_196_105, w_196_106, w_196_107, w_196_108, w_196_109, w_196_110, w_196_112, w_196_113, w_196_114, w_196_115, w_196_116, w_196_117, w_196_118, w_196_119, w_196_120, w_196_121, w_196_122, w_196_126, w_196_127, w_196_128, w_196_129, w_196_131;
  wire w_197_008, w_197_009, w_197_011, w_197_017, w_197_018, w_197_022, w_197_025, w_197_027, w_197_029, w_197_031, w_197_038, w_197_039, w_197_042, w_197_044, w_197_046, w_197_047, w_197_052, w_197_054, w_197_057, w_197_060, w_197_072, w_197_073, w_197_076, w_197_081, w_197_084, w_197_085, w_197_089, w_197_092, w_197_094, w_197_095, w_197_097, w_197_098, w_197_100, w_197_101, w_197_104, w_197_111, w_197_113, w_197_114, w_197_116, w_197_117, w_197_119, w_197_121, w_197_122, w_197_123, w_197_124, w_197_125, w_197_126, w_197_130, w_197_131, w_197_134, w_197_136, w_197_140, w_197_142, w_197_144, w_197_149, w_197_151, w_197_152, w_197_153, w_197_154, w_197_159, w_197_163, w_197_172, w_197_182, w_197_186, w_197_189, w_197_190, w_197_193, w_197_199, w_197_200, w_197_201, w_197_203, w_197_204, w_197_208, w_197_210, w_197_211, w_197_213, w_197_218, w_197_219, w_197_222, w_197_225, w_197_229, w_197_231, w_197_236, w_197_238, w_197_239, w_197_243, w_197_244, w_197_246, w_197_247, w_197_253, w_197_255, w_197_265, w_197_273, w_197_275, w_197_277, w_197_278, w_197_279, w_197_282, w_197_287, w_197_291, w_197_292, w_197_294, w_197_301, w_197_303, w_197_308, w_197_316, w_197_320, w_197_321, w_197_323, w_197_325, w_197_331, w_197_332, w_197_338, w_197_339, w_197_342, w_197_344, w_197_345, w_197_353, w_197_354, w_197_355, w_197_357, w_197_359, w_197_360, w_197_361, w_197_367, w_197_371, w_197_372, w_197_380, w_197_381, w_197_384, w_197_388, w_197_395, w_197_397, w_197_401, w_197_403, w_197_405, w_197_416, w_197_418, w_197_421, w_197_423, w_197_429, w_197_433, w_197_436, w_197_438, w_197_439, w_197_445, w_197_447, w_197_450, w_197_451, w_197_462, w_197_468, w_197_469, w_197_471, w_197_475, w_197_482, w_197_483, w_197_485, w_197_487, w_197_489, w_197_490, w_197_491, w_197_496, w_197_498, w_197_500, w_197_501, w_197_504, w_197_512, w_197_516, w_197_517, w_197_519, w_197_523, w_197_526, w_197_527, w_197_533, w_197_534, w_197_535, w_197_538, w_197_539, w_197_541, w_197_543, w_197_548, w_197_549, w_197_550, w_197_560, w_197_563, w_197_570, w_197_573, w_197_574, w_197_575, w_197_577, w_197_580, w_197_584, w_197_585, w_197_588, w_197_595, w_197_600, w_197_605, w_197_608, w_197_611, w_197_614, w_197_615, w_197_621, w_197_622, w_197_628, w_197_631, w_197_633, w_197_649, w_197_653, w_197_655, w_197_661, w_197_663, w_197_665, w_197_677, w_197_685, w_197_687, w_197_694, w_197_696, w_197_707, w_197_711, w_197_714, w_197_716, w_197_720, w_197_737, w_197_738, w_197_739, w_197_744, w_197_745, w_197_746, w_197_750, w_197_757, w_197_759, w_197_762, w_197_763, w_197_765, w_197_767, w_197_769, w_197_773, w_197_774, w_197_775, w_197_776, w_197_778, w_197_782, w_197_785, w_197_788, w_197_792, w_197_797, w_197_803, w_197_805, w_197_806, w_197_807, w_197_808, w_197_812, w_197_815, w_197_816, w_197_823, w_197_824, w_197_827, w_197_830, w_197_831, w_197_834, w_197_847, w_197_849, w_197_861, w_197_863, w_197_866, w_197_867, w_197_871, w_197_885, w_197_887, w_197_893, w_197_896, w_197_906, w_197_907, w_197_909, w_197_914, w_197_919, w_197_924, w_197_926, w_197_927, w_197_928, w_197_929, w_197_931, w_197_940, w_197_942, w_197_943, w_197_947, w_197_949, w_197_958, w_197_974, w_197_976, w_197_979, w_197_980, w_197_983, w_197_986, w_197_989, w_197_992, w_197_994, w_197_995, w_197_999, w_197_1012, w_197_1013, w_197_1014, w_197_1018, w_197_1019, w_197_1027, w_197_1030, w_197_1032, w_197_1033, w_197_1035, w_197_1045, w_197_1053, w_197_1056, w_197_1059, w_197_1065, w_197_1066, w_197_1068, w_197_1074, w_197_1087, w_197_1090, w_197_1097, w_197_1100, w_197_1101, w_197_1107, w_197_1112, w_197_1115, w_197_1125, w_197_1129, w_197_1132, w_197_1134, w_197_1136, w_197_1137, w_197_1146, w_197_1154, w_197_1157, w_197_1163, w_197_1175, w_197_1177, w_197_1186, w_197_1191, w_197_1204, w_197_1205, w_197_1206, w_197_1214, w_197_1221, w_197_1222, w_197_1228, w_197_1229, w_197_1233, w_197_1235, w_197_1237, w_197_1238, w_197_1243, w_197_1244, w_197_1255, w_197_1256, w_197_1257, w_197_1261, w_197_1264, w_197_1265, w_197_1266, w_197_1267, w_197_1269, w_197_1275, w_197_1278, w_197_1281, w_197_1283, w_197_1284, w_197_1289, w_197_1291, w_197_1295, w_197_1301, w_197_1304, w_197_1305, w_197_1315, w_197_1317, w_197_1326, w_197_1327, w_197_1329, w_197_1336, w_197_1337, w_197_1338, w_197_1340, w_197_1348, w_197_1350, w_197_1356, w_197_1365, w_197_1366, w_197_1367, w_197_1368, w_197_1370, w_197_1371, w_197_1373, w_197_1382, w_197_1384, w_197_1385, w_197_1386, w_197_1390, w_197_1391, w_197_1394, w_197_1395, w_197_1397, w_197_1407, w_197_1408, w_197_1413, w_197_1419, w_197_1422, w_197_1427, w_197_1431, w_197_1437, w_197_1438, w_197_1440, w_197_1442, w_197_1445, w_197_1447, w_197_1450, w_197_1452, w_197_1457, w_197_1458, w_197_1462, w_197_1469, w_197_1474, w_197_1487, w_197_1488, w_197_1491, w_197_1492, w_197_1495, w_197_1498, w_197_1501, w_197_1505, w_197_1506, w_197_1513, w_197_1515, w_197_1516, w_197_1522, w_197_1523, w_197_1526, w_197_1530, w_197_1537, w_197_1538, w_197_1539, w_197_1540, w_197_1541, w_197_1543, w_197_1546, w_197_1547, w_197_1552, w_197_1554, w_197_1565, w_197_1568, w_197_1570, w_197_1580, w_197_1584, w_197_1585, w_197_1588, w_197_1589, w_197_1593, w_197_1594, w_197_1595, w_197_1597, w_197_1603, w_197_1607, w_197_1609, w_197_1616, w_197_1618, w_197_1622, w_197_1623, w_197_1625, w_197_1627, w_197_1629, w_197_1637, w_197_1641, w_197_1644, w_197_1645, w_197_1647, w_197_1649, w_197_1650, w_197_1655, w_197_1667, w_197_1668, w_197_1689, w_197_1691, w_197_1694, w_197_1695, w_197_1697, w_197_1700, w_197_1708, w_197_1710, w_197_1716, w_197_1719, w_197_1727, w_197_1728, w_197_1730, w_197_1733, w_197_1735, w_197_1749, w_197_1758, w_197_1760, w_197_1764, w_197_1766, w_197_1769, w_197_1772, w_197_1779, w_197_1781, w_197_1785, w_197_1788, w_197_1791, w_197_1793, w_197_1798, w_197_1801, w_197_1805, w_197_1808, w_197_1810, w_197_1811, w_197_1813, w_197_1814, w_197_1817, w_197_1832, w_197_1833, w_197_1843, w_197_1845, w_197_1852, w_197_1856, w_197_1859, w_197_1861, w_197_1862, w_197_1865, w_197_1866, w_197_1868, w_197_1869, w_197_1872, w_197_1879, w_197_1882, w_197_1884, w_197_1886, w_197_1890, w_197_1906, w_197_1910, w_197_1912, w_197_1916, w_197_1931, w_197_1932, w_197_1933, w_197_1934, w_197_1935, w_197_1943, w_197_1952, w_197_1954, w_197_1958, w_197_1961, w_197_1966, w_197_1967, w_197_1968, w_197_1969, w_197_1979, w_197_1980, w_197_1983, w_197_1990, w_197_1993, w_197_1999, w_197_2010, w_197_2011, w_197_2012, w_197_2014, w_197_2021, w_197_2024, w_197_2027, w_197_2034, w_197_2036, w_197_2038, w_197_2039, w_197_2040, w_197_2044, w_197_2048, w_197_2049, w_197_2053, w_197_2056, w_197_2057, w_197_2058, w_197_2059, w_197_2064, w_197_2065, w_197_2081, w_197_2084, w_197_2100, w_197_2102, w_197_2105, w_197_2108, w_197_2109, w_197_2112, w_197_2115, w_197_2117, w_197_2126, w_197_2129, w_197_2131, w_197_2140, w_197_2142, w_197_2143, w_197_2147, w_197_2151, w_197_2158, w_197_2160, w_197_2161, w_197_2162, w_197_2163, w_197_2165, w_197_2167, w_197_2170, w_197_2171, w_197_2175, w_197_2176, w_197_2177;
  wire w_198_002, w_198_004, w_198_007, w_198_009, w_198_010, w_198_011, w_198_014, w_198_018, w_198_019, w_198_026, w_198_027, w_198_034, w_198_041, w_198_042, w_198_048, w_198_051, w_198_052, w_198_057, w_198_060, w_198_061, w_198_062, w_198_068, w_198_070, w_198_071, w_198_076, w_198_077, w_198_079, w_198_083, w_198_084, w_198_086, w_198_088, w_198_092, w_198_094, w_198_099, w_198_102, w_198_105, w_198_106, w_198_107, w_198_109, w_198_110, w_198_113, w_198_115, w_198_118, w_198_121, w_198_128, w_198_137, w_198_138, w_198_139, w_198_140, w_198_144, w_198_145, w_198_146, w_198_150, w_198_151, w_198_153, w_198_156, w_198_161, w_198_162, w_198_169, w_198_175, w_198_176, w_198_178, w_198_181, w_198_184, w_198_187, w_198_188, w_198_191, w_198_195, w_198_199, w_198_200, w_198_202, w_198_205, w_198_206, w_198_207, w_198_208, w_198_210, w_198_218, w_198_220, w_198_221, w_198_226, w_198_228, w_198_233, w_198_237, w_198_238, w_198_241, w_198_245, w_198_248, w_198_251, w_198_256, w_198_258, w_198_262, w_198_264, w_198_265, w_198_267, w_198_269, w_198_270, w_198_272, w_198_274, w_198_277, w_198_279, w_198_286, w_198_287, w_198_288, w_198_293, w_198_294, w_198_295, w_198_297, w_198_299, w_198_304, w_198_307, w_198_309, w_198_310, w_198_312, w_198_316, w_198_318, w_198_320, w_198_324, w_198_325, w_198_329, w_198_330, w_198_331, w_198_333, w_198_334, w_198_335, w_198_337, w_198_338, w_198_340, w_198_342, w_198_344, w_198_346, w_198_347, w_198_350, w_198_353, w_198_356, w_198_358, w_198_360, w_198_361, w_198_369, w_198_371, w_198_374, w_198_378, w_198_380, w_198_387, w_198_389, w_198_391, w_198_394, w_198_400, w_198_410, w_198_415, w_198_418, w_198_419, w_198_421, w_198_423, w_198_425, w_198_428, w_198_429, w_198_437, w_198_438, w_198_442, w_198_444, w_198_451, w_198_456, w_198_458, w_198_463, w_198_468, w_198_473, w_198_474, w_198_476, w_198_477, w_198_482, w_198_487, w_198_489, w_198_492, w_198_496, w_198_497, w_198_498, w_198_499, w_198_500, w_198_503, w_198_504, w_198_505, w_198_506, w_198_508, w_198_514, w_198_517, w_198_522, w_198_527, w_198_535, w_198_538, w_198_543, w_198_547, w_198_550, w_198_552, w_198_554, w_198_559, w_198_562, w_198_571, w_198_578, w_198_583, w_198_589, w_198_590, w_198_596, w_198_599, w_198_608, w_198_609, w_198_610, w_198_611, w_198_612, w_198_617, w_198_618, w_198_631, w_198_644, w_198_648, w_198_653, w_198_654, w_198_658, w_198_659, w_198_661, w_198_675, w_198_676, w_198_679, w_198_685, w_198_688, w_198_691, w_198_696, w_198_703, w_198_707, w_198_718, w_198_719, w_198_720, w_198_726, w_198_728, w_198_732, w_198_733, w_198_735, w_198_737, w_198_738, w_198_740, w_198_745, w_198_746, w_198_748, w_198_753, w_198_761, w_198_765, w_198_767, w_198_770, w_198_778, w_198_782, w_198_783, w_198_792, w_198_794, w_198_795, w_198_797, w_198_800, w_198_801, w_198_803, w_198_806, w_198_810, w_198_817, w_198_819, w_198_823, w_198_825, w_198_832, w_198_835, w_198_836, w_198_843, w_198_844, w_198_849, w_198_852, w_198_854, w_198_860, w_198_865, w_198_866, w_198_869, w_198_872, w_198_874, w_198_879, w_198_882, w_198_883, w_198_884, w_198_887, w_198_900, w_198_904, w_198_905, w_198_906, w_198_908, w_198_909, w_198_911, w_198_913, w_198_915, w_198_919, w_198_922, w_198_929, w_198_930, w_198_931, w_198_932, w_198_934, w_198_936, w_198_938, w_198_942, w_198_944, w_198_946, w_198_949, w_198_953, w_198_962, w_198_964, w_198_965, w_198_972, w_198_982, w_198_985, w_198_986, w_198_994, w_198_1001, w_198_1004, w_198_1006, w_198_1009, w_198_1024, w_198_1042, w_198_1047, w_198_1052, w_198_1056, w_198_1059, w_198_1077, w_198_1079, w_198_1083, w_198_1085, w_198_1092, w_198_1093, w_198_1096, w_198_1097, w_198_1098, w_198_1100, w_198_1102, w_198_1106, w_198_1107, w_198_1109, w_198_1121, w_198_1123, w_198_1125, w_198_1126, w_198_1130, w_198_1131, w_198_1141, w_198_1145, w_198_1148, w_198_1155, w_198_1156, w_198_1162, w_198_1163, w_198_1164, w_198_1171, w_198_1178, w_198_1179, w_198_1186, w_198_1196, w_198_1202, w_198_1205, w_198_1215, w_198_1219, w_198_1220, w_198_1222, w_198_1226, w_198_1227, w_198_1229, w_198_1230, w_198_1237, w_198_1248, w_198_1256, w_198_1257, w_198_1261, w_198_1272, w_198_1275, w_198_1284, w_198_1289, w_198_1292, w_198_1293, w_198_1297, w_198_1303, w_198_1314, w_198_1316, w_198_1318, w_198_1320, w_198_1326, w_198_1343, w_198_1345, w_198_1352, w_198_1354, w_198_1362, w_198_1366, w_198_1368, w_198_1370, w_198_1384, w_198_1385, w_198_1387, w_198_1388, w_198_1390, w_198_1392, w_198_1393, w_198_1395, w_198_1396, w_198_1399, w_198_1401, w_198_1404, w_198_1407, w_198_1408, w_198_1410, w_198_1414, w_198_1416, w_198_1424, w_198_1430, w_198_1431, w_198_1439, w_198_1442, w_198_1445, w_198_1467, w_198_1471, w_198_1476, w_198_1478, w_198_1479, w_198_1484, w_198_1486, w_198_1490, w_198_1496, w_198_1497, w_198_1498, w_198_1506, w_198_1515, w_198_1519, w_198_1533, w_198_1534, w_198_1540, w_198_1542, w_198_1543, w_198_1546, w_198_1549, w_198_1555, w_198_1558, w_198_1559, w_198_1561, w_198_1572, w_198_1583, w_198_1584, w_198_1590, w_198_1592, w_198_1593, w_198_1595, w_198_1598, w_198_1601, w_198_1602, w_198_1605, w_198_1606, w_198_1629, w_198_1630, w_198_1635, w_198_1642, w_198_1643, w_198_1648, w_198_1656, w_198_1658, w_198_1661, w_198_1670, w_198_1672, w_198_1685, w_198_1687, w_198_1693, w_198_1694, w_198_1697, w_198_1700, w_198_1710, w_198_1711, w_198_1718, w_198_1719, w_198_1726, w_198_1737, w_198_1738, w_198_1741, w_198_1747, w_198_1749, w_198_1750, w_198_1751, w_198_1758, w_198_1761, w_198_1765, w_198_1766, w_198_1769, w_198_1775, w_198_1778, w_198_1787, w_198_1804, w_198_1812, w_198_1815, w_198_1822, w_198_1824, w_198_1825, w_198_1826, w_198_1828, w_198_1829, w_198_1833, w_198_1837, w_198_1843, w_198_1847, w_198_1853, w_198_1857, w_198_1861, w_198_1882, w_198_1892, w_198_1893, w_198_1894, w_198_1900, w_198_1905, w_198_1907, w_198_1919, w_198_1920, w_198_1923, w_198_1925, w_198_1926, w_198_1931, w_198_1932, w_198_1934, w_198_1937, w_198_1943, w_198_1946, w_198_1947, w_198_1949, w_198_1959, w_198_1964, w_198_1966, w_198_1973, w_198_1983, w_198_1986, w_198_1989, w_198_1992, w_198_1997, w_198_2000, w_198_2004, w_198_2010, w_198_2012, w_198_2020, w_198_2025, w_198_2030, w_198_2033, w_198_2036, w_198_2037, w_198_2039, w_198_2043, w_198_2049, w_198_2057, w_198_2062, w_198_2079, w_198_2083, w_198_2089, w_198_2090, w_198_2092, w_198_2094, w_198_2106, w_198_2113, w_198_2116, w_198_2118, w_198_2120, w_198_2122, w_198_2123, w_198_2130, w_198_2131, w_198_2132, w_198_2134, w_198_2135, w_198_2142, w_198_2148, w_198_2150, w_198_2155, w_198_2159, w_198_2165, w_198_2166, w_198_2170, w_198_2171, w_198_2174, w_198_2183, w_198_2187, w_198_2189, w_198_2190, w_198_2191, w_198_2203, w_198_2209, w_198_2211, w_198_2223, w_198_2226, w_198_2233, w_198_2235, w_198_2240, w_198_2242, w_198_2243, w_198_2247, w_198_2248, w_198_2250, w_198_2252, w_198_2255, w_198_2256, w_198_2258, w_198_2260, w_198_2270, w_198_2276, w_198_2277;
  wire w_199_003, w_199_004, w_199_006, w_199_009, w_199_013, w_199_015, w_199_019, w_199_025, w_199_029, w_199_033, w_199_035, w_199_036, w_199_037, w_199_040, w_199_041, w_199_042, w_199_044, w_199_046, w_199_048, w_199_050, w_199_051, w_199_057, w_199_059, w_199_064, w_199_065, w_199_067, w_199_068, w_199_069, w_199_071, w_199_072, w_199_075, w_199_080, w_199_081, w_199_083, w_199_084, w_199_088, w_199_090, w_199_092, w_199_094, w_199_098, w_199_100, w_199_102, w_199_104, w_199_105, w_199_107, w_199_108, w_199_112, w_199_113, w_199_115, w_199_120, w_199_125, w_199_127, w_199_129, w_199_131, w_199_132, w_199_133, w_199_138, w_199_141, w_199_143, w_199_144, w_199_146, w_199_150, w_199_167, w_199_170, w_199_172, w_199_174, w_199_175, w_199_176, w_199_177, w_199_183, w_199_184, w_199_185, w_199_188, w_199_193, w_199_196, w_199_202, w_199_209, w_199_210, w_199_213, w_199_216, w_199_218, w_199_222, w_199_224, w_199_227, w_199_228, w_199_237, w_199_242, w_199_244, w_199_245, w_199_247, w_199_248, w_199_252, w_199_261, w_199_263, w_199_272, w_199_276, w_199_277, w_199_279, w_199_282, w_199_287, w_199_288, w_199_299, w_199_300, w_199_301, w_199_303, w_199_305, w_199_311, w_199_318, w_199_319, w_199_324, w_199_326, w_199_330, w_199_334, w_199_335, w_199_336, w_199_338, w_199_340, w_199_342, w_199_347, w_199_348, w_199_352, w_199_354, w_199_360, w_199_361, w_199_363, w_199_364, w_199_365, w_199_369, w_199_370, w_199_375, w_199_381, w_199_387, w_199_390, w_199_393, w_199_396, w_199_397, w_199_398, w_199_401, w_199_405, w_199_410, w_199_414, w_199_415, w_199_416, w_199_417, w_199_421, w_199_422, w_199_423, w_199_425, w_199_428, w_199_431, w_199_432, w_199_433, w_199_435, w_199_438, w_199_442, w_199_448, w_199_450, w_199_456, w_199_461, w_199_465, w_199_470, w_199_476, w_199_479, w_199_480, w_199_481, w_199_484, w_199_485, w_199_488, w_199_490, w_199_494, w_199_496, w_199_497, w_199_499, w_199_502, w_199_505, w_199_506, w_199_508, w_199_509, w_199_510, w_199_511, w_199_514, w_199_515, w_199_517, w_199_519, w_199_521, w_199_525, w_199_526, w_199_529, w_199_531, w_199_532, w_199_533, w_199_535, w_199_537, w_199_539, w_199_540, w_199_544, w_199_550, w_199_551, w_199_555, w_199_557, w_199_559, w_199_560, w_199_561, w_199_563, w_199_564, w_199_570, w_199_571, w_199_574, w_199_579, w_199_583, w_199_586, w_199_590, w_199_593, w_199_594, w_199_600, w_199_602, w_199_606, w_199_613, w_199_621, w_199_624, w_199_630, w_199_631, w_199_632, w_199_635, w_199_636, w_199_638, w_199_641, w_199_642, w_199_647, w_199_658, w_199_659, w_199_660, w_199_661, w_199_668, w_199_670, w_199_681, w_199_682, w_199_686, w_199_687, w_199_689, w_199_690, w_199_691, w_199_693, w_199_694, w_199_697, w_199_698, w_199_704, w_199_705, w_199_707, w_199_708, w_199_713, w_199_714, w_199_715, w_199_719, w_199_721, w_199_728, w_199_729, w_199_730, w_199_732, w_199_733, w_199_737, w_199_741, w_199_750, w_199_754, w_199_760, w_199_764, w_199_770, w_199_771, w_199_775, w_199_777, w_199_778, w_199_781, w_199_782, w_199_783, w_199_786, w_199_789, w_199_790, w_199_792, w_199_793, w_199_797, w_199_798, w_199_799, w_199_800, w_199_802, w_199_803, w_199_811, w_199_812, w_199_813, w_199_815, w_199_817, w_199_818, w_199_821, w_199_822, w_199_823, w_199_831, w_199_834, w_199_839, w_199_841, w_199_846, w_199_849, w_199_850, w_199_853, w_199_857, w_199_867, w_199_872, w_199_873, w_199_874, w_199_875, w_199_878, w_199_880, w_199_885, w_199_888, w_199_889, w_199_892, w_199_893, w_199_898, w_199_899, w_199_900, w_199_902, w_199_905, w_199_908, w_199_909, w_199_912, w_199_914, w_199_918, w_199_919, w_199_921, w_199_927, w_199_929, w_199_930, w_199_935, w_199_936, w_199_940, w_199_942, w_199_943, w_199_951, w_199_954, w_199_955, w_199_956, w_199_959, w_199_963, w_199_965, w_199_975, w_199_976, w_199_983, w_199_985, w_199_988, w_199_990, w_199_992, w_199_997, w_199_999, w_199_1001, w_199_1002, w_199_1005, w_199_1009, w_199_1011, w_199_1012, w_199_1013, w_199_1014, w_199_1018, w_199_1019, w_199_1020, w_199_1022, w_199_1028, w_199_1029, w_199_1030, w_199_1031, w_199_1033, w_199_1035, w_199_1037, w_199_1038, w_199_1042, w_199_1043, w_199_1046, w_199_1049, w_199_1051, w_199_1053, w_199_1054, w_199_1057, w_199_1060, w_199_1067, w_199_1070, w_199_1072, w_199_1076, w_199_1080, w_199_1081, w_199_1083, w_199_1085, w_199_1090, w_199_1097, w_199_1098, w_199_1099, w_199_1103, w_199_1108, w_199_1112, w_199_1116, w_199_1117, w_199_1119, w_199_1123, w_199_1124, w_199_1136, w_199_1138, w_199_1141, w_199_1142, w_199_1143, w_199_1145, w_199_1146, w_199_1147, w_199_1148, w_199_1156, w_199_1158, w_199_1166, w_199_1167, w_199_1168, w_199_1175, w_199_1176, w_199_1177, w_199_1178, w_199_1180, w_199_1185, w_199_1186, w_199_1187, w_199_1190, w_199_1193, w_199_1194, w_199_1208, w_199_1213, w_199_1215, w_199_1217, w_199_1221, w_199_1223, w_199_1224, w_199_1227, w_199_1228, w_199_1230, w_199_1236, w_199_1237, w_199_1239, w_199_1242, w_199_1244, w_199_1246, w_199_1253, w_199_1254, w_199_1255, w_199_1258, w_199_1259, w_199_1260, w_199_1268, w_199_1272, w_199_1277, w_199_1282, w_199_1286, w_199_1293, w_199_1297, w_199_1299, w_199_1303, w_199_1308, w_199_1315, w_199_1320, w_199_1321, w_199_1324, w_199_1325, w_199_1328, w_199_1332, w_199_1334, w_199_1335, w_199_1337, w_199_1344, w_199_1349, w_199_1350, w_199_1351, w_199_1356, w_199_1357, w_199_1360, w_199_1361, w_199_1362, w_199_1369, w_199_1375, w_199_1376, w_199_1378, w_199_1379, w_199_1380, w_199_1382, w_199_1388, w_199_1391, w_199_1392, w_199_1394, w_199_1403, w_199_1406, w_199_1407, w_199_1408, w_199_1409, w_199_1410, w_199_1412, w_199_1417, w_199_1418, w_199_1423, w_199_1425, w_199_1427, w_199_1428, w_199_1433, w_199_1435, w_199_1436, w_199_1438, w_199_1441, w_199_1442, w_199_1443, w_199_1444, w_199_1448, w_199_1449, w_199_1451, w_199_1453, w_199_1454, w_199_1456, w_199_1459, w_199_1460, w_199_1461, w_199_1464, w_199_1465, w_199_1466, w_199_1471, w_199_1472, w_199_1476, w_199_1477, w_199_1480, w_199_1485, w_199_1488, w_199_1490, w_199_1492, w_199_1493, w_199_1495, w_199_1497, w_199_1499, w_199_1500, w_199_1508, w_199_1511, w_199_1512, w_199_1514, w_199_1521, w_199_1529, w_199_1537, w_199_1541, w_199_1544, w_199_1547, w_199_1548, w_199_1551, w_199_1558, w_199_1561, w_199_1570, w_199_1571, w_199_1572, w_199_1579, w_199_1580, w_199_1585, w_199_1586, w_199_1589, w_199_1593, w_199_1594, w_199_1595, w_199_1599, w_199_1601, w_199_1606, w_199_1609, w_199_1610, w_199_1612, w_199_1614, w_199_1621, w_199_1623, w_199_1627, w_199_1629, w_199_1630;
  wire w_200_005, w_200_010, w_200_012, w_200_025, w_200_026, w_200_027, w_200_028, w_200_031, w_200_032, w_200_040, w_200_042, w_200_043, w_200_045, w_200_047, w_200_052, w_200_061, w_200_065, w_200_067, w_200_068, w_200_070, w_200_072, w_200_077, w_200_078, w_200_079, w_200_080, w_200_082, w_200_090, w_200_095, w_200_098, w_200_101, w_200_103, w_200_104, w_200_113, w_200_114, w_200_122, w_200_134, w_200_135, w_200_142, w_200_145, w_200_147, w_200_153, w_200_164, w_200_169, w_200_170, w_200_171, w_200_173, w_200_178, w_200_181, w_200_182, w_200_185, w_200_187, w_200_189, w_200_191, w_200_204, w_200_210, w_200_212, w_200_214, w_200_219, w_200_222, w_200_224, w_200_225, w_200_231, w_200_233, w_200_238, w_200_246, w_200_256, w_200_262, w_200_267, w_200_272, w_200_274, w_200_277, w_200_281, w_200_287, w_200_289, w_200_294, w_200_295, w_200_296, w_200_299, w_200_303, w_200_306, w_200_307, w_200_314, w_200_317, w_200_322, w_200_323, w_200_324, w_200_331, w_200_334, w_200_344, w_200_348, w_200_349, w_200_358, w_200_362, w_200_365, w_200_371, w_200_376, w_200_387, w_200_388, w_200_390, w_200_396, w_200_397, w_200_398, w_200_401, w_200_403, w_200_407, w_200_414, w_200_419, w_200_439, w_200_443, w_200_449, w_200_462, w_200_469, w_200_471, w_200_480, w_200_486, w_200_490, w_200_498, w_200_499, w_200_502, w_200_504, w_200_505, w_200_506, w_200_507, w_200_510, w_200_511, w_200_515, w_200_521, w_200_527, w_200_529, w_200_530, w_200_533, w_200_534, w_200_538, w_200_541, w_200_542, w_200_556, w_200_562, w_200_565, w_200_571, w_200_575, w_200_593, w_200_602, w_200_605, w_200_608, w_200_612, w_200_615, w_200_623, w_200_625, w_200_626, w_200_632, w_200_635, w_200_641, w_200_644, w_200_646, w_200_647, w_200_648, w_200_649, w_200_655, w_200_656, w_200_661, w_200_665, w_200_668, w_200_673, w_200_681, w_200_685, w_200_686, w_200_688, w_200_689, w_200_692, w_200_696, w_200_697, w_200_700, w_200_705, w_200_707, w_200_710, w_200_712, w_200_716, w_200_720, w_200_725, w_200_729, w_200_737, w_200_746, w_200_747, w_200_752, w_200_755, w_200_756, w_200_758, w_200_769, w_200_771, w_200_775, w_200_776, w_200_780, w_200_784, w_200_800, w_200_802, w_200_808, w_200_813, w_200_821, w_200_823, w_200_826, w_200_831, w_200_835, w_200_836, w_200_837, w_200_840, w_200_843, w_200_847, w_200_848, w_200_858, w_200_862, w_200_866, w_200_870, w_200_871, w_200_872, w_200_873, w_200_876, w_200_878, w_200_879, w_200_887, w_200_888, w_200_891, w_200_898, w_200_901, w_200_905, w_200_912, w_200_918, w_200_920, w_200_922, w_200_925, w_200_926, w_200_930, w_200_934, w_200_936, w_200_938, w_200_941, w_200_943, w_200_948, w_200_950, w_200_951, w_200_955, w_200_963, w_200_972, w_200_980, w_200_984, w_200_987, w_200_992, w_200_993, w_200_1007, w_200_1011, w_200_1017, w_200_1019, w_200_1020, w_200_1022, w_200_1025, w_200_1027, w_200_1028, w_200_1031, w_200_1033, w_200_1040, w_200_1043, w_200_1045, w_200_1054, w_200_1055, w_200_1057, w_200_1064, w_200_1069, w_200_1071, w_200_1077, w_200_1078, w_200_1080, w_200_1087, w_200_1092, w_200_1096, w_200_1101, w_200_1103, w_200_1105, w_200_1108, w_200_1110, w_200_1120, w_200_1122, w_200_1128, w_200_1133, w_200_1135, w_200_1136, w_200_1137, w_200_1138, w_200_1141, w_200_1143, w_200_1150, w_200_1152, w_200_1153, w_200_1154, w_200_1155, w_200_1158, w_200_1159, w_200_1165, w_200_1176, w_200_1177, w_200_1181, w_200_1189, w_200_1193, w_200_1200, w_200_1206, w_200_1208, w_200_1212, w_200_1213, w_200_1217, w_200_1219, w_200_1223, w_200_1225, w_200_1228, w_200_1231, w_200_1235, w_200_1242, w_200_1244, w_200_1246, w_200_1253, w_200_1255, w_200_1260, w_200_1270, w_200_1274, w_200_1282, w_200_1285, w_200_1290, w_200_1292, w_200_1294, w_200_1295, w_200_1302, w_200_1304, w_200_1308, w_200_1309, w_200_1319, w_200_1325, w_200_1327, w_200_1333, w_200_1347, w_200_1354, w_200_1361, w_200_1366, w_200_1369, w_200_1381, w_200_1383, w_200_1389, w_200_1390, w_200_1392, w_200_1393, w_200_1394, w_200_1402, w_200_1413, w_200_1420, w_200_1422, w_200_1424, w_200_1427, w_200_1428, w_200_1429, w_200_1430, w_200_1431, w_200_1441, w_200_1442, w_200_1451, w_200_1452, w_200_1454, w_200_1458, w_200_1459, w_200_1462, w_200_1466, w_200_1467, w_200_1472, w_200_1480, w_200_1493, w_200_1506, w_200_1510, w_200_1517, w_200_1522, w_200_1523, w_200_1524, w_200_1531, w_200_1533, w_200_1535, w_200_1536, w_200_1539, w_200_1541, w_200_1543, w_200_1545, w_200_1549, w_200_1563, w_200_1567, w_200_1569, w_200_1573, w_200_1574, w_200_1578, w_200_1583, w_200_1588, w_200_1589, w_200_1597, w_200_1604, w_200_1607, w_200_1611, w_200_1613, w_200_1615, w_200_1620, w_200_1625, w_200_1631, w_200_1635, w_200_1636, w_200_1643, w_200_1650, w_200_1658, w_200_1659, w_200_1663, w_200_1668, w_200_1677, w_200_1680, w_200_1682, w_200_1688, w_200_1701, w_200_1703, w_200_1704, w_200_1712, w_200_1716, w_200_1720, w_200_1730, w_200_1732, w_200_1734, w_200_1735, w_200_1737, w_200_1748, w_200_1753, w_200_1756, w_200_1760, w_200_1761, w_200_1763, w_200_1767, w_200_1768, w_200_1771, w_200_1772, w_200_1781, w_200_1785, w_200_1788, w_200_1790, w_200_1791, w_200_1793, w_200_1802, w_200_1804, w_200_1805, w_200_1808, w_200_1812, w_200_1815, w_200_1817, w_200_1818, w_200_1819, w_200_1824, w_200_1826, w_200_1843, w_200_1846, w_200_1853, w_200_1854, w_200_1855, w_200_1856, w_200_1863, w_200_1869, w_200_1870, w_200_1873, w_200_1875, w_200_1888, w_200_1890, w_200_1893, w_200_1894, w_200_1897, w_200_1907, w_200_1908, w_200_1916, w_200_1917, w_200_1926, w_200_1929, w_200_1930, w_200_1934, w_200_1937, w_200_1939, w_200_1940, w_200_1941, w_200_1945, w_200_1946, w_200_1950, w_200_1953, w_200_1958, w_200_1973, w_200_1979, w_200_1980, w_200_1981, w_200_1986, w_200_1988, w_200_1990, w_200_1992, w_200_1993, w_200_1997, w_200_2001, w_200_2002, w_200_2003, w_200_2004, w_200_2009, w_200_2013, w_200_2017, w_200_2022, w_200_2023, w_200_2032, w_200_2035, w_200_2037, w_200_2038, w_200_2047, w_200_2051, w_200_2054, w_200_2064, w_200_2080, w_200_2084, w_200_2105, w_200_2106, w_200_2113, w_200_2116, w_200_2118, w_200_2120, w_200_2136, w_200_2144, w_200_2146, w_200_2154, w_200_2157, w_200_2167, w_200_2188, w_200_2194, w_200_2211, w_200_2214, w_200_2223, w_200_2228, w_200_2235, w_200_2240, w_200_2245, w_200_2256, w_200_2261, w_200_2269, w_200_2276, w_200_2280, w_200_2287, w_200_2288, w_200_2308, w_200_2310, w_200_2341, w_200_2347, w_200_2348, w_200_2356, w_200_2361, w_200_2363, w_200_2366, w_200_2375, w_200_2396, w_200_2402, w_200_2408, w_200_2416, w_200_2422, w_200_2452, w_200_2453, w_200_2454, w_200_2463, w_200_2487, w_200_2488, w_200_2494, w_200_2499, w_200_2503, w_200_2511, w_200_2515, w_200_2531, w_200_2542, w_200_2544, w_200_2550, w_200_2568, w_200_2576, w_200_2586, w_200_2591, w_200_2594, w_200_2599, w_200_2601, w_200_2606, w_200_2621, w_200_2624, w_200_2629, w_200_2641, w_200_2650, w_200_2652, w_200_2657, w_200_2664, w_200_2672, w_200_2675, w_200_2680, w_200_2687, w_200_2693, w_200_2703, w_200_2709, w_200_2711, w_200_2720, w_200_2726, w_200_2736, w_200_2738, w_200_2745, w_200_2769, w_200_2773, w_200_2779, w_200_2783, w_200_2787, w_200_2793, w_200_2799, w_200_2802, w_200_2807, w_200_2812, w_200_2815, w_200_2821, w_200_2832, w_200_2837, w_200_2850, w_200_2869, w_200_2871, w_200_2877, w_200_2885, w_200_2888, w_200_2890, w_200_2893, w_200_2902, w_200_2907, w_200_2912, w_200_2915;
  wire w_201_006, w_201_008, w_201_009, w_201_023, w_201_024, w_201_025, w_201_030, w_201_031, w_201_038, w_201_045, w_201_051, w_201_052, w_201_061, w_201_065, w_201_066, w_201_067, w_201_072, w_201_075, w_201_089, w_201_100, w_201_110, w_201_115, w_201_117, w_201_121, w_201_127, w_201_128, w_201_130, w_201_139, w_201_144, w_201_146, w_201_149, w_201_152, w_201_161, w_201_165, w_201_166, w_201_168, w_201_170, w_201_173, w_201_175, w_201_185, w_201_189, w_201_190, w_201_193, w_201_194, w_201_196, w_201_200, w_201_202, w_201_203, w_201_205, w_201_207, w_201_208, w_201_209, w_201_211, w_201_222, w_201_225, w_201_228, w_201_230, w_201_233, w_201_234, w_201_238, w_201_240, w_201_243, w_201_251, w_201_263, w_201_267, w_201_278, w_201_279, w_201_281, w_201_285, w_201_289, w_201_291, w_201_301, w_201_303, w_201_310, w_201_312, w_201_318, w_201_329, w_201_334, w_201_335, w_201_341, w_201_348, w_201_350, w_201_351, w_201_356, w_201_382, w_201_391, w_201_406, w_201_407, w_201_408, w_201_413, w_201_422, w_201_424, w_201_427, w_201_428, w_201_430, w_201_431, w_201_433, w_201_439, w_201_440, w_201_441, w_201_448, w_201_454, w_201_459, w_201_464, w_201_468, w_201_471, w_201_477, w_201_478, w_201_479, w_201_484, w_201_488, w_201_489, w_201_490, w_201_494, w_201_495, w_201_496, w_201_497, w_201_501, w_201_509, w_201_523, w_201_529, w_201_539, w_201_540, w_201_546, w_201_547, w_201_550, w_201_554, w_201_565, w_201_568, w_201_569, w_201_575, w_201_584, w_201_587, w_201_588, w_201_593, w_201_602, w_201_607, w_201_612, w_201_613, w_201_615, w_201_622, w_201_633, w_201_640, w_201_643, w_201_645, w_201_649, w_201_651, w_201_659, w_201_662, w_201_664, w_201_668, w_201_675, w_201_681, w_201_685, w_201_689, w_201_699, w_201_705, w_201_715, w_201_717, w_201_718, w_201_722, w_201_726, w_201_732, w_201_734, w_201_736, w_201_739, w_201_752, w_201_758, w_201_759, w_201_764, w_201_765, w_201_766, w_201_767, w_201_780, w_201_783, w_201_784, w_201_786, w_201_788, w_201_794, w_201_795, w_201_800, w_201_803, w_201_807, w_201_808, w_201_810, w_201_811, w_201_815, w_201_820, w_201_823, w_201_824, w_201_828, w_201_831, w_201_835, w_201_838, w_201_840, w_201_843, w_201_854, w_201_855, w_201_859, w_201_862, w_201_864, w_201_865, w_201_869, w_201_870, w_201_871, w_201_875, w_201_878, w_201_884, w_201_886, w_201_887, w_201_888, w_201_891, w_201_899, w_201_901, w_201_906, w_201_908, w_201_917, w_201_919, w_201_920, w_201_923, w_201_927, w_201_932, w_201_937, w_201_938, w_201_949, w_201_953, w_201_965, w_201_967, w_201_986, w_201_991, w_201_996, w_201_997, w_201_1000, w_201_1004, w_201_1015, w_201_1021, w_201_1022, w_201_1024, w_201_1030, w_201_1032, w_201_1036, w_201_1037, w_201_1038, w_201_1044, w_201_1047, w_201_1051, w_201_1060, w_201_1062, w_201_1068, w_201_1081, w_201_1082, w_201_1083, w_201_1091, w_201_1106, w_201_1107, w_201_1110, w_201_1118, w_201_1124, w_201_1126, w_201_1132, w_201_1134, w_201_1138, w_201_1141, w_201_1147, w_201_1158, w_201_1163, w_201_1164, w_201_1165, w_201_1167, w_201_1169, w_201_1170, w_201_1177, w_201_1180, w_201_1184, w_201_1191, w_201_1193, w_201_1196, w_201_1198, w_201_1200, w_201_1211, w_201_1214, w_201_1217, w_201_1222, w_201_1223, w_201_1224, w_201_1227, w_201_1232, w_201_1233, w_201_1234, w_201_1239, w_201_1240, w_201_1247, w_201_1248, w_201_1264, w_201_1265, w_201_1267, w_201_1275, w_201_1276, w_201_1280, w_201_1285, w_201_1289, w_201_1290, w_201_1299, w_201_1303, w_201_1305, w_201_1309, w_201_1316, w_201_1320, w_201_1327, w_201_1333, w_201_1335, w_201_1336, w_201_1344, w_201_1345, w_201_1347, w_201_1348, w_201_1349, w_201_1351, w_201_1355, w_201_1360, w_201_1364, w_201_1365, w_201_1368, w_201_1370, w_201_1371, w_201_1372, w_201_1377, w_201_1378, w_201_1388, w_201_1389, w_201_1391, w_201_1393, w_201_1399, w_201_1401, w_201_1404, w_201_1406, w_201_1408, w_201_1413, w_201_1422, w_201_1430, w_201_1431, w_201_1433, w_201_1435, w_201_1442, w_201_1444, w_201_1448, w_201_1453, w_201_1456, w_201_1458, w_201_1459, w_201_1464, w_201_1466, w_201_1470, w_201_1471, w_201_1480, w_201_1488, w_201_1491, w_201_1494, w_201_1497, w_201_1499, w_201_1505, w_201_1508, w_201_1517, w_201_1522, w_201_1524, w_201_1529, w_201_1530, w_201_1531, w_201_1533, w_201_1535, w_201_1545, w_201_1548, w_201_1550, w_201_1552, w_201_1553, w_201_1554, w_201_1564, w_201_1566, w_201_1569, w_201_1572, w_201_1574, w_201_1577, w_201_1586, w_201_1587, w_201_1590, w_201_1602, w_201_1604, w_201_1607, w_201_1612, w_201_1613, w_201_1614, w_201_1616, w_201_1618, w_201_1626, w_201_1628, w_201_1630, w_201_1633, w_201_1640, w_201_1642, w_201_1643, w_201_1645, w_201_1654, w_201_1658, w_201_1659, w_201_1665, w_201_1671, w_201_1674, w_201_1680, w_201_1685, w_201_1694, w_201_1695, w_201_1698, w_201_1702, w_201_1707, w_201_1708, w_201_1709, w_201_1711, w_201_1714, w_201_1724, w_201_1725, w_201_1728, w_201_1730, w_201_1731, w_201_1734, w_201_1742, w_201_1745, w_201_1746, w_201_1747, w_201_1752, w_201_1753, w_201_1756, w_201_1759, w_201_1763, w_201_1764, w_201_1766, w_201_1767, w_201_1771, w_201_1772, w_201_1776, w_201_1784, w_201_1789, w_201_1790, w_201_1791, w_201_1795, w_201_1796, w_201_1797, w_201_1803, w_201_1805, w_201_1807, w_201_1810, w_201_1813, w_201_1819, w_201_1821, w_201_1822, w_201_1831, w_201_1833, w_201_1838, w_201_1846, w_201_1853, w_201_1855, w_201_1860, w_201_1861, w_201_1870, w_201_1877, w_201_1878, w_201_1886, w_201_1889, w_201_1895, w_201_1896, w_201_1898, w_201_1901, w_201_1915, w_201_1926, w_201_1936, w_201_1939, w_201_1948, w_201_1950, w_201_1963, w_201_1968, w_201_1973, w_201_1977, w_201_1981, w_201_1985, w_201_1990, w_201_1999, w_201_2003, w_201_2006, w_201_2018, w_201_2019, w_201_2021, w_201_2026, w_201_2030, w_201_2034, w_201_2035, w_201_2041, w_201_2044, w_201_2045, w_201_2047, w_201_2050, w_201_2059, w_201_2061, w_201_2065, w_201_2066, w_201_2068, w_201_2070, w_201_2073, w_201_2075, w_201_2085, w_201_2087, w_201_2092, w_201_2094, w_201_2095, w_201_2098, w_201_2100, w_201_2102, w_201_2105, w_201_2125, w_201_2126, w_201_2131, w_201_2135, w_201_2137, w_201_2149, w_201_2151, w_201_2152, w_201_2160, w_201_2161, w_201_2166, w_201_2169, w_201_2177, w_201_2182, w_201_2188, w_201_2190, w_201_2195, w_201_2204, w_201_2205, w_201_2217, w_201_2228, w_201_2229, w_201_2231, w_201_2241, w_201_2253, w_201_2254, w_201_2259, w_201_2262, w_201_2269, w_201_2275, w_201_2276, w_201_2279, w_201_2281, w_201_2287, w_201_2296, w_201_2298, w_201_2336, w_201_2355, w_201_2372, w_201_2375, w_201_2382, w_201_2388, w_201_2392, w_201_2421, w_201_2425, w_201_2437, w_201_2439, w_201_2443, w_201_2445, w_201_2449, w_201_2454, w_201_2460, w_201_2463, w_201_2466, w_201_2481, w_201_2493, w_201_2494, w_201_2498, w_201_2505, w_201_2507, w_201_2511, w_201_2526, w_201_2528, w_201_2539, w_201_2542, w_201_2543, w_201_2547, w_201_2561, w_201_2572, w_201_2591, w_201_2596, w_201_2608, w_201_2615, w_201_2616, w_201_2617, w_201_2622, w_201_2628, w_201_2640, w_201_2654, w_201_2660, w_201_2667, w_201_2668, w_201_2670, w_201_2674, w_201_2675, w_201_2678, w_201_2681, w_201_2683, w_201_2688;
  wire w_202_000, w_202_001, w_202_002, w_202_003, w_202_004, w_202_006, w_202_007, w_202_008, w_202_009, w_202_010, w_202_012, w_202_013, w_202_014, w_202_015, w_202_016, w_202_017, w_202_020, w_202_022, w_202_023, w_202_024, w_202_025, w_202_026, w_202_027, w_202_029, w_202_030, w_202_031, w_202_032, w_202_033, w_202_034, w_202_035, w_202_036, w_202_037, w_202_039, w_202_040, w_202_043, w_202_045, w_202_046, w_202_048, w_202_049, w_202_051, w_202_056, w_202_057, w_202_059, w_202_060, w_202_061, w_202_062, w_202_063, w_202_065, w_202_066, w_202_067, w_202_068, w_202_069, w_202_070, w_202_072, w_202_073, w_202_074, w_202_075, w_202_077, w_202_078, w_202_079, w_202_081, w_202_084, w_202_085, w_202_087, w_202_088, w_202_089, w_202_091, w_202_092, w_202_094, w_202_096, w_202_097, w_202_098, w_202_099, w_202_100, w_202_101, w_202_102, w_202_104, w_202_105, w_202_106, w_202_110, w_202_111, w_202_112, w_202_114, w_202_115, w_202_116, w_202_117, w_202_119, w_202_121, w_202_122, w_202_124, w_202_125, w_202_126, w_202_130, w_202_132, w_202_133, w_202_136, w_202_137, w_202_138, w_202_139, w_202_141, w_202_142, w_202_144, w_202_146, w_202_147, w_202_148, w_202_150, w_202_152, w_202_154, w_202_155, w_202_156, w_202_157, w_202_158, w_202_160, w_202_162, w_202_165, w_202_166, w_202_167, w_202_168, w_202_169, w_202_170, w_202_173, w_202_174, w_202_175, w_202_177, w_202_180, w_202_181, w_202_182, w_202_183, w_202_184, w_202_185, w_202_188, w_202_189, w_202_191, w_202_192, w_202_194, w_202_195, w_202_196, w_202_198, w_202_199, w_202_200, w_202_201, w_202_202, w_202_205, w_202_208, w_202_209, w_202_210, w_202_211, w_202_212, w_202_214, w_202_216, w_202_217, w_202_218, w_202_219, w_202_221, w_202_222, w_202_224, w_202_227, w_202_230, w_202_233, w_202_234, w_202_236, w_202_237, w_202_239, w_202_240, w_202_242, w_202_243, w_202_245, w_202_246, w_202_250, w_202_251, w_202_252, w_202_253, w_202_254, w_202_258, w_202_259, w_202_263, w_202_264, w_202_265, w_202_266, w_202_267, w_202_268, w_202_269, w_202_270, w_202_271, w_202_273, w_202_274, w_202_275, w_202_276, w_202_278, w_202_279, w_202_281, w_202_282, w_202_285, w_202_287, w_202_288, w_202_290, w_202_291, w_202_293, w_202_294, w_202_298, w_202_299, w_202_300, w_202_304, w_202_306, w_202_307, w_202_308, w_202_309, w_202_311, w_202_313, w_202_314, w_202_316, w_202_317, w_202_318, w_202_319, w_202_322, w_202_325, w_202_326, w_202_327, w_202_328, w_202_333, w_202_335, w_202_336, w_202_339, w_202_340, w_202_341, w_202_342, w_202_344, w_202_347, w_202_348, w_202_349, w_202_351, w_202_352, w_202_353, w_202_356, w_202_358, w_202_360, w_202_361, w_202_362, w_202_366, w_202_368, w_202_369, w_202_371, w_202_374, w_202_375, w_202_376, w_202_377, w_202_378, w_202_379, w_202_380, w_202_382, w_202_383, w_202_387, w_202_389, w_202_393, w_202_395, w_202_396, w_202_398, w_202_399, w_202_400, w_202_401, w_202_402, w_202_403, w_202_404, w_202_406, w_202_407, w_202_408, w_202_409, w_202_411, w_202_412, w_202_413, w_202_415, w_202_418, w_202_420, w_202_421, w_202_422, w_202_424, w_202_425, w_202_426, w_202_428, w_202_429, w_202_435, w_202_437, w_202_438, w_202_439, w_202_441, w_202_442, w_202_444, w_202_445, w_202_446, w_202_447, w_202_448, w_202_450, w_202_453, w_202_454, w_202_456, w_202_457, w_202_458, w_202_459, w_202_460, w_202_461, w_202_465, w_202_466, w_202_467, w_202_468, w_202_469, w_202_470, w_202_471, w_202_478, w_202_479, w_202_480, w_202_481, w_202_484, w_202_485, w_202_486, w_202_487, w_202_489, w_202_490, w_202_493, w_202_494, w_202_495, w_202_497, w_202_498, w_202_499, w_202_500, w_202_501, w_202_502, w_202_504, w_202_505, w_202_506, w_202_508, w_202_509, w_202_510, w_202_514, w_202_515, w_202_516, w_202_518, w_202_521, w_202_522, w_202_524, w_202_525, w_202_526, w_202_527, w_202_529, w_202_531, w_202_535, w_202_539, w_202_540, w_202_541, w_202_542, w_202_544, w_202_545, w_202_546, w_202_547, w_202_549, w_202_551, w_202_552, w_202_553, w_202_554, w_202_558, w_202_560, w_202_562, w_202_563, w_202_565, w_202_567, w_202_569, w_202_570, w_202_571, w_202_572, w_202_573, w_202_575, w_202_576, w_202_577, w_202_578, w_202_580, w_202_582, w_202_585, w_202_586, w_202_590, w_202_591, w_202_592, w_202_594, w_202_595, w_202_596, w_202_597, w_202_598, w_202_599, w_202_601, w_202_604, w_202_606, w_202_607, w_202_608, w_202_609, w_202_611, w_202_613, w_202_614, w_202_615, w_202_618, w_202_619, w_202_621, w_202_622, w_202_624, w_202_626, w_202_627, w_202_632, w_202_633, w_202_634, w_202_635, w_202_638, w_202_639, w_202_640, w_202_642, w_202_643, w_202_644, w_202_646, w_202_648, w_202_649, w_202_652, w_202_653, w_202_656, w_202_661, w_202_663, w_202_664, w_202_665;
  wire w_203_000, w_203_006, w_203_012, w_203_017, w_203_021, w_203_025, w_203_039, w_203_043, w_203_044, w_203_047, w_203_050, w_203_057, w_203_065, w_203_066, w_203_080, w_203_086, w_203_091, w_203_098, w_203_101, w_203_103, w_203_109, w_203_125, w_203_132, w_203_136, w_203_142, w_203_153, w_203_155, w_203_159, w_203_160, w_203_162, w_203_164, w_203_166, w_203_173, w_203_175, w_203_176, w_203_179, w_203_186, w_203_190, w_203_191, w_203_192, w_203_199, w_203_200, w_203_201, w_203_204, w_203_210, w_203_216, w_203_217, w_203_220, w_203_223, w_203_229, w_203_232, w_203_240, w_203_241, w_203_242, w_203_243, w_203_244, w_203_247, w_203_250, w_203_254, w_203_255, w_203_261, w_203_263, w_203_267, w_203_269, w_203_270, w_203_272, w_203_274, w_203_282, w_203_292, w_203_294, w_203_295, w_203_307, w_203_311, w_203_313, w_203_315, w_203_319, w_203_321, w_203_322, w_203_324, w_203_325, w_203_326, w_203_327, w_203_336, w_203_340, w_203_344, w_203_368, w_203_376, w_203_377, w_203_379, w_203_385, w_203_388, w_203_391, w_203_398, w_203_400, w_203_405, w_203_407, w_203_411, w_203_422, w_203_426, w_203_429, w_203_430, w_203_433, w_203_436, w_203_441, w_203_442, w_203_444, w_203_451, w_203_452, w_203_459, w_203_466, w_203_467, w_203_478, w_203_481, w_203_482, w_203_497, w_203_498, w_203_499, w_203_505, w_203_508, w_203_517, w_203_536, w_203_550, w_203_553, w_203_558, w_203_561, w_203_564, w_203_583, w_203_592, w_203_594, w_203_600, w_203_601, w_203_603, w_203_604, w_203_612, w_203_619, w_203_620, w_203_626, w_203_640, w_203_641, w_203_656, w_203_659, w_203_665, w_203_666, w_203_673, w_203_674, w_203_677, w_203_685, w_203_695, w_203_704, w_203_705, w_203_707, w_203_708, w_203_711, w_203_720, w_203_726, w_203_731, w_203_736, w_203_739, w_203_740, w_203_741, w_203_743, w_203_749, w_203_752, w_203_753, w_203_754, w_203_758, w_203_771, w_203_774, w_203_775, w_203_777, w_203_781, w_203_783, w_203_785, w_203_801, w_203_806, w_203_809, w_203_810, w_203_814, w_203_821, w_203_830, w_203_838, w_203_843, w_203_845, w_203_850, w_203_856, w_203_858, w_203_859, w_203_861, w_203_867, w_203_868, w_203_869, w_203_874, w_203_878, w_203_881, w_203_882, w_203_884, w_203_893, w_203_894, w_203_902, w_203_907, w_203_909, w_203_910, w_203_912, w_203_915, w_203_916, w_203_917, w_203_922, w_203_928, w_203_930, w_203_937, w_203_946, w_203_947, w_203_948, w_203_953, w_203_954, w_203_956, w_203_962, w_203_970, w_203_980, w_203_983, w_203_987, w_203_993, w_203_995, w_203_999, w_203_1007, w_203_1015, w_203_1027, w_203_1029, w_203_1035, w_203_1036, w_203_1037, w_203_1040, w_203_1042, w_203_1047, w_203_1048, w_203_1049, w_203_1052, w_203_1054, w_203_1064, w_203_1067, w_203_1069, w_203_1076, w_203_1081, w_203_1082, w_203_1087, w_203_1090, w_203_1092, w_203_1094, w_203_1099, w_203_1108, w_203_1111, w_203_1129, w_203_1131, w_203_1143, w_203_1150, w_203_1152, w_203_1153, w_203_1155, w_203_1160, w_203_1161, w_203_1162, w_203_1164, w_203_1169, w_203_1170, w_203_1172, w_203_1174, w_203_1175, w_203_1177, w_203_1179, w_203_1182, w_203_1185, w_203_1187, w_203_1189, w_203_1194, w_203_1198, w_203_1200, w_203_1203, w_203_1204, w_203_1208, w_203_1212, w_203_1215, w_203_1216, w_203_1217, w_203_1221, w_203_1222, w_203_1227, w_203_1237, w_203_1259, w_203_1270, w_203_1272, w_203_1275, w_203_1276, w_203_1279, w_203_1282, w_203_1289, w_203_1296, w_203_1299, w_203_1300, w_203_1301, w_203_1306, w_203_1316, w_203_1320, w_203_1323, w_203_1333, w_203_1334, w_203_1341, w_203_1349, w_203_1356, w_203_1357, w_203_1359, w_203_1365, w_203_1366, w_203_1368, w_203_1369, w_203_1370, w_203_1372, w_203_1375, w_203_1376, w_203_1380, w_203_1384, w_203_1388, w_203_1390, w_203_1394, w_203_1396, w_203_1398, w_203_1403, w_203_1407, w_203_1408, w_203_1409, w_203_1414, w_203_1417, w_203_1427, w_203_1428, w_203_1434, w_203_1439, w_203_1455, w_203_1457, w_203_1458, w_203_1466, w_203_1470, w_203_1510, w_203_1513, w_203_1517, w_203_1522, w_203_1523, w_203_1540, w_203_1544, w_203_1549, w_203_1554, w_203_1559, w_203_1570, w_203_1583, w_203_1584, w_203_1585, w_203_1589, w_203_1622, w_203_1632, w_203_1636, w_203_1638, w_203_1647, w_203_1662, w_203_1664, w_203_1665, w_203_1672, w_203_1673, w_203_1675, w_203_1677, w_203_1681, w_203_1687, w_203_1694, w_203_1695, w_203_1707, w_203_1712, w_203_1719, w_203_1728, w_203_1731, w_203_1741, w_203_1752, w_203_1753, w_203_1754, w_203_1756, w_203_1781, w_203_1799, w_203_1801, w_203_1802, w_203_1808, w_203_1811, w_203_1818, w_203_1828, w_203_1829, w_203_1840, w_203_1845, w_203_1852, w_203_1856, w_203_1860, w_203_1868, w_203_1869, w_203_1884, w_203_1886, w_203_1906, w_203_1908, w_203_1936, w_203_1939, w_203_1956, w_203_1960, w_203_1966, w_203_1977, w_203_1988, w_203_1992, w_203_1999, w_203_2002, w_203_2023, w_203_2033, w_203_2043, w_203_2045, w_203_2058, w_203_2064, w_203_2067, w_203_2075, w_203_2090, w_203_2096, w_203_2097, w_203_2098, w_203_2108, w_203_2109, w_203_2115, w_203_2139, w_203_2153, w_203_2160, w_203_2166, w_203_2175, w_203_2176, w_203_2178, w_203_2179, w_203_2181, w_203_2186, w_203_2200, w_203_2203, w_203_2207, w_203_2217, w_203_2219, w_203_2221, w_203_2228, w_203_2238, w_203_2243, w_203_2257, w_203_2270, w_203_2275, w_203_2282, w_203_2284, w_203_2298, w_203_2320, w_203_2330, w_203_2339, w_203_2342, w_203_2349, w_203_2353, w_203_2355, w_203_2358, w_203_2360, w_203_2373, w_203_2378, w_203_2379, w_203_2381, w_203_2395, w_203_2410, w_203_2416, w_203_2424, w_203_2442, w_203_2444, w_203_2458, w_203_2473, w_203_2518, w_203_2520, w_203_2531, w_203_2536, w_203_2539, w_203_2549, w_203_2551, w_203_2559, w_203_2565, w_203_2577, w_203_2585, w_203_2588, w_203_2598, w_203_2602, w_203_2605, w_203_2606, w_203_2610, w_203_2612, w_203_2619, w_203_2621, w_203_2623, w_203_2635, w_203_2637, w_203_2639, w_203_2673, w_203_2674, w_203_2678, w_203_2692, w_203_2714, w_203_2717, w_203_2722, w_203_2730, w_203_2731, w_203_2750, w_203_2761, w_203_2773, w_203_2781, w_203_2787, w_203_2802, w_203_2822, w_203_2840, w_203_2845, w_203_2849, w_203_2856, w_203_2859, w_203_2861, w_203_2872, w_203_2879, w_203_2880, w_203_2882, w_203_2887, w_203_2889, w_203_2892, w_203_2894, w_203_2901, w_203_2907, w_203_2909, w_203_2915, w_203_2942, w_203_2945, w_203_2947, w_203_2950, w_203_2951, w_203_2962, w_203_2964, w_203_2978, w_203_2979, w_203_2987, w_203_2989, w_203_3004, w_203_3007, w_203_3021, w_203_3041, w_203_3043, w_203_3044, w_203_3059, w_203_3073, w_203_3076, w_203_3079, w_203_3111, w_203_3112, w_203_3121, w_203_3128, w_203_3154, w_203_3159, w_203_3164, w_203_3178, w_203_3183, w_203_3207, w_203_3208, w_203_3224, w_203_3234, w_203_3265, w_203_3267, w_203_3271, w_203_3280, w_203_3284, w_203_3285, w_203_3289, w_203_3299, w_203_3308, w_203_3341, w_203_3350, w_203_3351, w_203_3359, w_203_3363, w_203_3365, w_203_3393, w_203_3405, w_203_3412, w_203_3416, w_203_3436, w_203_3437, w_203_3438, w_203_3455, w_203_3456, w_203_3466, w_203_3473, w_203_3481, w_203_3486, w_203_3493, w_203_3497, w_203_3498, w_203_3532, w_203_3533, w_203_3537, w_203_3555, w_203_3559, w_203_3563, w_203_3569;
  wire w_204_003, w_204_004, w_204_005, w_204_009, w_204_017, w_204_018, w_204_027, w_204_029, w_204_031, w_204_032, w_204_036, w_204_040, w_204_041, w_204_046, w_204_048, w_204_054, w_204_063, w_204_064, w_204_066, w_204_067, w_204_068, w_204_069, w_204_070, w_204_073, w_204_075, w_204_079, w_204_080, w_204_085, w_204_086, w_204_089, w_204_096, w_204_098, w_204_099, w_204_100, w_204_101, w_204_102, w_204_106, w_204_108, w_204_110, w_204_111, w_204_113, w_204_116, w_204_120, w_204_121, w_204_122, w_204_123, w_204_124, w_204_127, w_204_131, w_204_134, w_204_137, w_204_138, w_204_144, w_204_145, w_204_150, w_204_151, w_204_152, w_204_155, w_204_156, w_204_157, w_204_159, w_204_160, w_204_165, w_204_167, w_204_168, w_204_169, w_204_174, w_204_176, w_204_177, w_204_179, w_204_181, w_204_185, w_204_186, w_204_187, w_204_189, w_204_190, w_204_192, w_204_196, w_204_202, w_204_207, w_204_208, w_204_209, w_204_211, w_204_212, w_204_213, w_204_217, w_204_220, w_204_221, w_204_222, w_204_227, w_204_234, w_204_236, w_204_243, w_204_246, w_204_247, w_204_248, w_204_250, w_204_252, w_204_253, w_204_255, w_204_256, w_204_269, w_204_270, w_204_273, w_204_275, w_204_277, w_204_278, w_204_282, w_204_283, w_204_285, w_204_288, w_204_289, w_204_291, w_204_294, w_204_295, w_204_296, w_204_299, w_204_300, w_204_302, w_204_308, w_204_309, w_204_310, w_204_313, w_204_314, w_204_315, w_204_319, w_204_320, w_204_322, w_204_325, w_204_329, w_204_335, w_204_339, w_204_340, w_204_347, w_204_349, w_204_352, w_204_353, w_204_356, w_204_359, w_204_362, w_204_363, w_204_364, w_204_368, w_204_369, w_204_370, w_204_371, w_204_372, w_204_376, w_204_377, w_204_378, w_204_392, w_204_393, w_204_394, w_204_399, w_204_400, w_204_403, w_204_405, w_204_409, w_204_419, w_204_421, w_204_426, w_204_428, w_204_430, w_204_433, w_204_441, w_204_443, w_204_445, w_204_446, w_204_450, w_204_452, w_204_461, w_204_464, w_204_467, w_204_469, w_204_472, w_204_473, w_204_477, w_204_478, w_204_479, w_204_482, w_204_483, w_204_488, w_204_492, w_204_493, w_204_495, w_204_496, w_204_502, w_204_507, w_204_509, w_204_511, w_204_512, w_204_514, w_204_521, w_204_522, w_204_532, w_204_541, w_204_542, w_204_544, w_204_549, w_204_560, w_204_563, w_204_565, w_204_567, w_204_571, w_204_575, w_204_576, w_204_577, w_204_582, w_204_583, w_204_588, w_204_590, w_204_592, w_204_593, w_204_594, w_204_596, w_204_598, w_204_604, w_204_605, w_204_607, w_204_610, w_204_611, w_204_614, w_204_616, w_204_619, w_204_620, w_204_623, w_204_624, w_204_625, w_204_629, w_204_631, w_204_641, w_204_642, w_204_646, w_204_650, w_204_653, w_204_656, w_204_662, w_204_663, w_204_664, w_204_668, w_204_669, w_204_675, w_204_678, w_204_682, w_204_684, w_204_685, w_204_691, w_204_698, w_204_700, w_204_701, w_204_704, w_204_706, w_204_712, w_204_715, w_204_717, w_204_719, w_204_722, w_204_723, w_204_724, w_204_730, w_204_731, w_204_732, w_204_734, w_204_738, w_204_739, w_204_741, w_204_742, w_204_743, w_204_744, w_204_747, w_204_751, w_204_752, w_204_754, w_204_767, w_204_770, w_204_772, w_204_773, w_204_781, w_204_785, w_204_786, w_204_795, w_204_803, w_204_804, w_204_807, w_204_817, w_204_820, w_204_822, w_204_834, w_204_836, w_204_838, w_204_839, w_204_842, w_204_851, w_204_852, w_204_855, w_204_858, w_204_859, w_204_868, w_204_869, w_204_871, w_204_872, w_204_875, w_204_878, w_204_881, w_204_884, w_204_887, w_204_888, w_204_891, w_204_892, w_204_893, w_204_895, w_204_896, w_204_898, w_204_904, w_204_905, w_204_912, w_204_916, w_204_918, w_204_921, w_204_926, w_204_927, w_204_928, w_204_930, w_204_934, w_204_937, w_204_938, w_204_944, w_204_946, w_204_947, w_204_953, w_204_954, w_204_955, w_204_957, w_204_958, w_204_962, w_204_963, w_204_966, w_204_967, w_204_970, w_204_977, w_204_987, w_204_988, w_204_990, w_204_991, w_204_992, w_204_994, w_204_998, w_204_1000, w_204_1004, w_204_1007, w_204_1008, w_204_1009, w_204_1012, w_204_1013, w_204_1016, w_204_1020, w_204_1021, w_204_1024, w_204_1029, w_204_1030, w_204_1032, w_204_1036, w_204_1039, w_204_1042, w_204_1043, w_204_1047, w_204_1051, w_204_1052, w_204_1053, w_204_1060, w_204_1062, w_204_1066, w_204_1067, w_204_1070, w_204_1073, w_204_1074, w_204_1075, w_204_1081, w_204_1083, w_204_1088, w_204_1089, w_204_1090, w_204_1095, w_204_1096, w_204_1098, w_204_1099, w_204_1101, w_204_1105, w_204_1109, w_204_1113, w_204_1114, w_204_1119, w_204_1124, w_204_1127, w_204_1129, w_204_1130, w_204_1131, w_204_1137, w_204_1139, w_204_1140, w_204_1141, w_204_1142, w_204_1143, w_204_1144, w_204_1146, w_204_1147, w_204_1148, w_204_1153, w_204_1155, w_204_1157, w_204_1158, w_204_1177, w_204_1180, w_204_1182, w_204_1191, w_204_1197, w_204_1201, w_204_1207, w_204_1213, w_204_1215, w_204_1238, w_204_1239, w_204_1242, w_204_1251, w_204_1253, w_204_1255, w_204_1259, w_204_1261, w_204_1265, w_204_1268, w_204_1273, w_204_1275, w_204_1277, w_204_1280, w_204_1283, w_204_1285, w_204_1286, w_204_1287, w_204_1288, w_204_1289, w_204_1292, w_204_1293, w_204_1299, w_204_1301, w_204_1303, w_204_1304, w_204_1306, w_204_1309, w_204_1311, w_204_1315, w_204_1319, w_204_1320, w_204_1321, w_204_1324, w_204_1331, w_204_1333, w_204_1338, w_204_1342, w_204_1349, w_204_1355, w_204_1356, w_204_1365, w_204_1368, w_204_1373, w_204_1374, w_204_1378, w_204_1379, w_204_1386, w_204_1388, w_204_1393, w_204_1400, w_204_1411, w_204_1412, w_204_1415, w_204_1416, w_204_1424, w_204_1431, w_204_1432, w_204_1437, w_204_1438, w_204_1441, w_204_1444, w_204_1446, w_204_1456, w_204_1457, w_204_1467, w_204_1471, w_204_1472, w_204_1473, w_204_1477, w_204_1478, w_204_1481, w_204_1482, w_204_1483, w_204_1497, w_204_1505, w_204_1508, w_204_1513, w_204_1516, w_204_1518, w_204_1519, w_204_1527, w_204_1530, w_204_1533, w_204_1534, w_204_1536, w_204_1542, w_204_1544, w_204_1552, w_204_1553, w_204_1556, w_204_1563, w_204_1567, w_204_1568, w_204_1570, w_204_1571, w_204_1574, w_204_1575, w_204_1576;
  wire w_205_001, w_205_002, w_205_003, w_205_005, w_205_011, w_205_012, w_205_013, w_205_014, w_205_016, w_205_017, w_205_018, w_205_019, w_205_022, w_205_023, w_205_024, w_205_026, w_205_027, w_205_030, w_205_031, w_205_032, w_205_033, w_205_034, w_205_035, w_205_036, w_205_038, w_205_039, w_205_040, w_205_042, w_205_043, w_205_045, w_205_046, w_205_049, w_205_050, w_205_052, w_205_053, w_205_054, w_205_055, w_205_056, w_205_057, w_205_058, w_205_059, w_205_060, w_205_061, w_205_063, w_205_064, w_205_065, w_205_066, w_205_067, w_205_068, w_205_070, w_205_071, w_205_075, w_205_080, w_205_082, w_205_083, w_205_084, w_205_085, w_205_089, w_205_095, w_205_096, w_205_097, w_205_099, w_205_102, w_205_104, w_205_106, w_205_109, w_205_111, w_205_115, w_205_116, w_205_117, w_205_118, w_205_120, w_205_121, w_205_126, w_205_128, w_205_132, w_205_134, w_205_135, w_205_136, w_205_138, w_205_139, w_205_142, w_205_143, w_205_144, w_205_145, w_205_146, w_205_149, w_205_150, w_205_151, w_205_153, w_205_154, w_205_156, w_205_157, w_205_158, w_205_159, w_205_161, w_205_162, w_205_163, w_205_166, w_205_167, w_205_169, w_205_170, w_205_172, w_205_173, w_205_175, w_205_180, w_205_182, w_205_183, w_205_184, w_205_190, w_205_191, w_205_192, w_205_193, w_205_194, w_205_195, w_205_196, w_205_197, w_205_198, w_205_200, w_205_201, w_205_202, w_205_204, w_205_205, w_205_206, w_205_210, w_205_211, w_205_212, w_205_213, w_205_214, w_205_217, w_205_218, w_205_219, w_205_221, w_205_223, w_205_224, w_205_225, w_205_226, w_205_228, w_205_230, w_205_231, w_205_233, w_205_234, w_205_235, w_205_238, w_205_239, w_205_241, w_205_242, w_205_245, w_205_246, w_205_247, w_205_248, w_205_249, w_205_251, w_205_254, w_205_255, w_205_259, w_205_264, w_205_265, w_205_268, w_205_271, w_205_274, w_205_277, w_205_280, w_205_282, w_205_283, w_205_290, w_205_291, w_205_292, w_205_293, w_205_294, w_205_295, w_205_297, w_205_298, w_205_302, w_205_303, w_205_305, w_205_308, w_205_309, w_205_311, w_205_314, w_205_315, w_205_316, w_205_317, w_205_320, w_205_322, w_205_323, w_205_324, w_205_328, w_205_329, w_205_330, w_205_331, w_205_332, w_205_334, w_205_335, w_205_338, w_205_340, w_205_341, w_205_344, w_205_345, w_205_347, w_205_348, w_205_349, w_205_352, w_205_357, w_205_359, w_205_360, w_205_362, w_205_363, w_205_368, w_205_370, w_205_371, w_205_372, w_205_375, w_205_376, w_205_377, w_205_378, w_205_379, w_205_381, w_205_383, w_205_385, w_205_386, w_205_387, w_205_392, w_205_395, w_205_399, w_205_400, w_205_402, w_205_403, w_205_406, w_205_409, w_205_413, w_205_415, w_205_416, w_205_417, w_205_418, w_205_419, w_205_421, w_205_424, w_205_425, w_205_430, w_205_436, w_205_437, w_205_438, w_205_440, w_205_442, w_205_444, w_205_445, w_205_446, w_205_447, w_205_449, w_205_451, w_205_452, w_205_453, w_205_455, w_205_457, w_205_459, w_205_461, w_205_462, w_205_467, w_205_468, w_205_471, w_205_472, w_205_473, w_205_475, w_205_477, w_205_479, w_205_481, w_205_482, w_205_485, w_205_487, w_205_489, w_205_490, w_205_491, w_205_494, w_205_496, w_205_498, w_205_501, w_205_502, w_205_504, w_205_506, w_205_511, w_205_514, w_205_518, w_205_520, w_205_521, w_205_524, w_205_528, w_205_529, w_205_530, w_205_534, w_205_535, w_205_537, w_205_540, w_205_542, w_205_543, w_205_544, w_205_546, w_205_547, w_205_551, w_205_552, w_205_553, w_205_554, w_205_557, w_205_559, w_205_561, w_205_565, w_205_566, w_205_567, w_205_569, w_205_570, w_205_579, w_205_581, w_205_583, w_205_585, w_205_586, w_205_587, w_205_589, w_205_591, w_205_592, w_205_593, w_205_596, w_205_598, w_205_600, w_205_601, w_205_604, w_205_606, w_205_607, w_205_608, w_205_613, w_205_615, w_205_616, w_205_618, w_205_620, w_205_623, w_205_626, w_205_627, w_205_628, w_205_634, w_205_635, w_205_636, w_205_638, w_205_643, w_205_645, w_205_646, w_205_647, w_205_649, w_205_650, w_205_652, w_205_653, w_205_654, w_205_655, w_205_656, w_205_659, w_205_660, w_205_661, w_205_662, w_205_663, w_205_665, w_205_666, w_205_669, w_205_670, w_205_672, w_205_673, w_205_674, w_205_680, w_205_681, w_205_682, w_205_684, w_205_685, w_205_689, w_205_691, w_205_692, w_205_694, w_205_695, w_205_697, w_205_699, w_205_700, w_205_701, w_205_702, w_205_704, w_205_705, w_205_708, w_205_709, w_205_710, w_205_714, w_205_716, w_205_717, w_205_718, w_205_721, w_205_724, w_205_725, w_205_727, w_205_730, w_205_734, w_205_737, w_205_739, w_205_741, w_205_744, w_205_745, w_205_746, w_205_748, w_205_753, w_205_755, w_205_758, w_205_765, w_205_766, w_205_771, w_205_774, w_205_775, w_205_779, w_205_781, w_205_785, w_205_789, w_205_791, w_205_792, w_205_793, w_205_795, w_205_796, w_205_797, w_205_798, w_205_800, w_205_801, w_205_802, w_205_804, w_205_805, w_205_806, w_205_810, w_205_813, w_205_816, w_205_817, w_205_818, w_205_819, w_205_822, w_205_824, w_205_826, w_205_827, w_205_828, w_205_829, w_205_832, w_205_834, w_205_835, w_205_836, w_205_837, w_205_841, w_205_842, w_205_843, w_205_847, w_205_848, w_205_849, w_205_850, w_205_853, w_205_854, w_205_856, w_205_857, w_205_858, w_205_861, w_205_863, w_205_864, w_205_866, w_205_867, w_205_868, w_205_869, w_205_872, w_205_875, w_205_876, w_205_877, w_205_878, w_205_879, w_205_880, w_205_889, w_205_890, w_205_891, w_205_892, w_205_893, w_205_895, w_205_898, w_205_899, w_205_901, w_205_903, w_205_904, w_205_907, w_205_909, w_205_910, w_205_911, w_205_913, w_205_914, w_205_915, w_205_918, w_205_921, w_205_922, w_205_924, w_205_925, w_205_926, w_205_927, w_205_928, w_205_929, w_205_930;
  wire w_206_000, w_206_002, w_206_003, w_206_004, w_206_005, w_206_007, w_206_008, w_206_009, w_206_010, w_206_013, w_206_014, w_206_016, w_206_018, w_206_019, w_206_021, w_206_029, w_206_031, w_206_034, w_206_036, w_206_039, w_206_040, w_206_041, w_206_042, w_206_046, w_206_050, w_206_051, w_206_052, w_206_054, w_206_055, w_206_056, w_206_061, w_206_062, w_206_064, w_206_066, w_206_067, w_206_068, w_206_069, w_206_070, w_206_071, w_206_075, w_206_077, w_206_079, w_206_080, w_206_083, w_206_087, w_206_088, w_206_091, w_206_092, w_206_095, w_206_096, w_206_098, w_206_099, w_206_100, w_206_101, w_206_103, w_206_104, w_206_108, w_206_110, w_206_112, w_206_114, w_206_115, w_206_118, w_206_119, w_206_120, w_206_121, w_206_122, w_206_123, w_206_124, w_206_131, w_206_134, w_206_135, w_206_136, w_206_137, w_206_138, w_206_139, w_206_143, w_206_144, w_206_145, w_206_146, w_206_149, w_206_151, w_206_152, w_206_159, w_206_162, w_206_164, w_206_165, w_206_167, w_206_168, w_206_169, w_206_170, w_206_171, w_206_172, w_206_178, w_206_181, w_206_182, w_206_183, w_206_184, w_206_186, w_206_188, w_206_189, w_206_192, w_206_193, w_206_197, w_206_198, w_206_199, w_206_200, w_206_202, w_206_203, w_206_204, w_206_205, w_206_207, w_206_208, w_206_209, w_206_211, w_206_212, w_206_213, w_206_214, w_206_218, w_206_220, w_206_222, w_206_223, w_206_224, w_206_225, w_206_228, w_206_230, w_206_231, w_206_232, w_206_235, w_206_238, w_206_239, w_206_242, w_206_243, w_206_244, w_206_246, w_206_247, w_206_248, w_206_250, w_206_252, w_206_253, w_206_255, w_206_256, w_206_257, w_206_260, w_206_261, w_206_265, w_206_267, w_206_268, w_206_269, w_206_271, w_206_273, w_206_278, w_206_280, w_206_281, w_206_283, w_206_286, w_206_288, w_206_290, w_206_291, w_206_294, w_206_297, w_206_298, w_206_300, w_206_301, w_206_302, w_206_306, w_206_308, w_206_312, w_206_314, w_206_315, w_206_319, w_206_320, w_206_321, w_206_322, w_206_324, w_206_325, w_206_326, w_206_328, w_206_329, w_206_331, w_206_332, w_206_334, w_206_335, w_206_336, w_206_339, w_206_342, w_206_343, w_206_345, w_206_346, w_206_347, w_206_348, w_206_353, w_206_354, w_206_356, w_206_357, w_206_358, w_206_359, w_206_363, w_206_364, w_206_365, w_206_366, w_206_367, w_206_369, w_206_375, w_206_376, w_206_379, w_206_380, w_206_382, w_206_385, w_206_386, w_206_387, w_206_389, w_206_392, w_206_398, w_206_403, w_206_404, w_206_405, w_206_406, w_206_408, w_206_410, w_206_412, w_206_414, w_206_417, w_206_418, w_206_421, w_206_422, w_206_423, w_206_425, w_206_428, w_206_430, w_206_432, w_206_433, w_206_435, w_206_438, w_206_441, w_206_444, w_206_445, w_206_448, w_206_451, w_206_457, w_206_458, w_206_459, w_206_460, w_206_462, w_206_467, w_206_472, w_206_473, w_206_476, w_206_479, w_206_483, w_206_486, w_206_487, w_206_488, w_206_493, w_206_494, w_206_496, w_206_498, w_206_501, w_206_510, w_206_513, w_206_514, w_206_518, w_206_519, w_206_522, w_206_530, w_206_532, w_206_533, w_206_535, w_206_537, w_206_538, w_206_539, w_206_548, w_206_549, w_206_550, w_206_551, w_206_553, w_206_554, w_206_558, w_206_559, w_206_563, w_206_564, w_206_566, w_206_567, w_206_568, w_206_571, w_206_576, w_206_578, w_206_579, w_206_580, w_206_581, w_206_582, w_206_584, w_206_585, w_206_586, w_206_588, w_206_589, w_206_591, w_206_592, w_206_594, w_206_597, w_206_600, w_206_601, w_206_603, w_206_605, w_206_606, w_206_607, w_206_608, w_206_611, w_206_612, w_206_613, w_206_617, w_206_622, w_206_624, w_206_626, w_206_627, w_206_628, w_206_631, w_206_633, w_206_635, w_206_636, w_206_637, w_206_639, w_206_640, w_206_642, w_206_643, w_206_646, w_206_650, w_206_651, w_206_654, w_206_656, w_206_658, w_206_659, w_206_660, w_206_661, w_206_667, w_206_668, w_206_671, w_206_672, w_206_673, w_206_674, w_206_677, w_206_678, w_206_679, w_206_680, w_206_683, w_206_687, w_206_692, w_206_693, w_206_700, w_206_702, w_206_704, w_206_707, w_206_713, w_206_714, w_206_719, w_206_721, w_206_724, w_206_728, w_206_729, w_206_730, w_206_731, w_206_732, w_206_733, w_206_734, w_206_735, w_206_739, w_206_741, w_206_742, w_206_743, w_206_744, w_206_745, w_206_746, w_206_753, w_206_754, w_206_755, w_206_757, w_206_759, w_206_760, w_206_761, w_206_763, w_206_766, w_206_767, w_206_769, w_206_770, w_206_772, w_206_774, w_206_777, w_206_778, w_206_783, w_206_785, w_206_788, w_206_790, w_206_794, w_206_795, w_206_801, w_206_802, w_206_803, w_206_804, w_206_806, w_206_808, w_206_809, w_206_810, w_206_811, w_206_813, w_206_815, w_206_821, w_206_822, w_206_823, w_206_829, w_206_830, w_206_831, w_206_832, w_206_833, w_206_836, w_206_837, w_206_838, w_206_840, w_206_841, w_206_842, w_206_843, w_206_845, w_206_846, w_206_847, w_206_853, w_206_861, w_206_862, w_206_868, w_206_869, w_206_870, w_206_875, w_206_876, w_206_877, w_206_878, w_206_880, w_206_883, w_206_884, w_206_887, w_206_891, w_206_896, w_206_901, w_206_905, w_206_912, w_206_914, w_206_918, w_206_920;
  wire w_207_000, w_207_004, w_207_007, w_207_008, w_207_011, w_207_012, w_207_013, w_207_014, w_207_015, w_207_016, w_207_022, w_207_023, w_207_024, w_207_025, w_207_030, w_207_034, w_207_040, w_207_042, w_207_044, w_207_046, w_207_048, w_207_051, w_207_052, w_207_056, w_207_065, w_207_066, w_207_069, w_207_073, w_207_076, w_207_080, w_207_081, w_207_082, w_207_091, w_207_093, w_207_094, w_207_100, w_207_102, w_207_104, w_207_106, w_207_108, w_207_109, w_207_110, w_207_116, w_207_121, w_207_126, w_207_129, w_207_131, w_207_132, w_207_133, w_207_135, w_207_137, w_207_140, w_207_144, w_207_150, w_207_151, w_207_154, w_207_155, w_207_156, w_207_158, w_207_160, w_207_161, w_207_163, w_207_164, w_207_179, w_207_180, w_207_181, w_207_182, w_207_185, w_207_188, w_207_189, w_207_191, w_207_192, w_207_193, w_207_196, w_207_199, w_207_203, w_207_204, w_207_205, w_207_206, w_207_215, w_207_217, w_207_221, w_207_223, w_207_225, w_207_226, w_207_231, w_207_233, w_207_235, w_207_239, w_207_241, w_207_246, w_207_247, w_207_252, w_207_254, w_207_255, w_207_257, w_207_259, w_207_262, w_207_266, w_207_267, w_207_276, w_207_277, w_207_280, w_207_281, w_207_283, w_207_286, w_207_287, w_207_291, w_207_292, w_207_294, w_207_295, w_207_298, w_207_301, w_207_303, w_207_306, w_207_310, w_207_311, w_207_314, w_207_315, w_207_319, w_207_321, w_207_323, w_207_324, w_207_325, w_207_327, w_207_328, w_207_329, w_207_330, w_207_333, w_207_335, w_207_337, w_207_343, w_207_347, w_207_355, w_207_356, w_207_358, w_207_374, w_207_375, w_207_376, w_207_379, w_207_381, w_207_382, w_207_389, w_207_390, w_207_394, w_207_396, w_207_397, w_207_398, w_207_399, w_207_405, w_207_406, w_207_409, w_207_410, w_207_411, w_207_412, w_207_415, w_207_418, w_207_420, w_207_426, w_207_428, w_207_431, w_207_433, w_207_436, w_207_446, w_207_449, w_207_450, w_207_452, w_207_456, w_207_458, w_207_461, w_207_462, w_207_465, w_207_466, w_207_468, w_207_471, w_207_473, w_207_475, w_207_481, w_207_484, w_207_492, w_207_498, w_207_499, w_207_506, w_207_509, w_207_512, w_207_514, w_207_515, w_207_519, w_207_523, w_207_527, w_207_528, w_207_534, w_207_536, w_207_537, w_207_538, w_207_539, w_207_540, w_207_542, w_207_546, w_207_553, w_207_554, w_207_559, w_207_563, w_207_568, w_207_569, w_207_572, w_207_573, w_207_581, w_207_594, w_207_595, w_207_598, w_207_601, w_207_602, w_207_604, w_207_605, w_207_606, w_207_608, w_207_612, w_207_613, w_207_616, w_207_621, w_207_627, w_207_628, w_207_630, w_207_633, w_207_638, w_207_641, w_207_642, w_207_643, w_207_644, w_207_647, w_207_648, w_207_651, w_207_654, w_207_655, w_207_656, w_207_657, w_207_658, w_207_660, w_207_661, w_207_664, w_207_666, w_207_668, w_207_672, w_207_677, w_207_683, w_207_688, w_207_689, w_207_697, w_207_701, w_207_703, w_207_707, w_207_709, w_207_710, w_207_711, w_207_716, w_207_718, w_207_721, w_207_725, w_207_727, w_207_728, w_207_733, w_207_734, w_207_735, w_207_740, w_207_741, w_207_742, w_207_752, w_207_757, w_207_761, w_207_766, w_207_770, w_207_774, w_207_775, w_207_776, w_207_781, w_207_788, w_207_789, w_207_793, w_207_794, w_207_796, w_207_802, w_207_803, w_207_807, w_207_810, w_207_817, w_207_820, w_207_821, w_207_824, w_207_831, w_207_837, w_207_849, w_207_852, w_207_853, w_207_855, w_207_856, w_207_861, w_207_862, w_207_864, w_207_867, w_207_871, w_207_874, w_207_876, w_207_880, w_207_884, w_207_889, w_207_892, w_207_896, w_207_897, w_207_900, w_207_902, w_207_903, w_207_905, w_207_907, w_207_911, w_207_913, w_207_916, w_207_933, w_207_934, w_207_935, w_207_938, w_207_941, w_207_942, w_207_943, w_207_946, w_207_955, w_207_956, w_207_957, w_207_959, w_207_965, w_207_966, w_207_967, w_207_968, w_207_974, w_207_975, w_207_976, w_207_978, w_207_979, w_207_984, w_207_986, w_207_988, w_207_990, w_207_992, w_207_996, w_207_997, w_207_1010, w_207_1011, w_207_1015, w_207_1020, w_207_1021, w_207_1022, w_207_1023, w_207_1027, w_207_1031, w_207_1033, w_207_1038, w_207_1040, w_207_1049, w_207_1051, w_207_1052, w_207_1053, w_207_1056, w_207_1057, w_207_1072, w_207_1073, w_207_1075, w_207_1082, w_207_1083, w_207_1085, w_207_1086, w_207_1089, w_207_1092, w_207_1093, w_207_1097, w_207_1102, w_207_1103, w_207_1104, w_207_1109, w_207_1114, w_207_1127, w_207_1128, w_207_1135, w_207_1137, w_207_1142, w_207_1146, w_207_1153, w_207_1155, w_207_1163, w_207_1166, w_207_1169, w_207_1171, w_207_1179, w_207_1186, w_207_1190, w_207_1191, w_207_1195, w_207_1202, w_207_1207, w_207_1211, w_207_1212, w_207_1219, w_207_1220, w_207_1225, w_207_1226, w_207_1228, w_207_1234, w_207_1236, w_207_1237, w_207_1238, w_207_1241, w_207_1242, w_207_1243, w_207_1244, w_207_1246, w_207_1251, w_207_1254, w_207_1265, w_207_1271, w_207_1273, w_207_1277, w_207_1279, w_207_1280, w_207_1285, w_207_1286, w_207_1288, w_207_1296, w_207_1300, w_207_1301, w_207_1303, w_207_1304, w_207_1309, w_207_1310, w_207_1312, w_207_1314, w_207_1319, w_207_1320, w_207_1327, w_207_1331, w_207_1332, w_207_1334, w_207_1335, w_207_1340, w_207_1351, w_207_1354, w_207_1360, w_207_1362, w_207_1367, w_207_1370, w_207_1372, w_207_1376, w_207_1378, w_207_1381, w_207_1382, w_207_1385, w_207_1387, w_207_1397, w_207_1398, w_207_1403, w_207_1405, w_207_1407, w_207_1410, w_207_1414, w_207_1415, w_207_1419, w_207_1422, w_207_1425, w_207_1433, w_207_1435, w_207_1440, w_207_1444, w_207_1446, w_207_1447, w_207_1454, w_207_1456, w_207_1458, w_207_1460, w_207_1477, w_207_1479, w_207_1495, w_207_1500, w_207_1503, w_207_1504, w_207_1506, w_207_1509, w_207_1510, w_207_1511, w_207_1518, w_207_1519, w_207_1524, w_207_1527, w_207_1529, w_207_1531, w_207_1534, w_207_1536, w_207_1545, w_207_1550, w_207_1552, w_207_1554, w_207_1560, w_207_1564, w_207_1565, w_207_1568, w_207_1569, w_207_1574, w_207_1577, w_207_1578, w_207_1584, w_207_1586, w_207_1590, w_207_1591, w_207_1596, w_207_1602, w_207_1607, w_207_1608, w_207_1611, w_207_1612, w_207_1618, w_207_1620, w_207_1630, w_207_1634, w_207_1640, w_207_1643, w_207_1649, w_207_1651, w_207_1655, w_207_1658, w_207_1660, w_207_1670, w_207_1671, w_207_1672, w_207_1673, w_207_1674, w_207_1675, w_207_1676, w_207_1677, w_207_1678, w_207_1679, w_207_1682, w_207_1685, w_207_1689, w_207_1690, w_207_1691, w_207_1693, w_207_1694, w_207_1698, w_207_1700, w_207_1705, w_207_1706, w_207_1707, w_207_1709, w_207_1712, w_207_1718, w_207_1723, w_207_1730, w_207_1733, w_207_1734, w_207_1739, w_207_1740, w_207_1746, w_207_1748, w_207_1755, w_207_1758, w_207_1759, w_207_1761, w_207_1765, w_207_1775, w_207_1781, w_207_1784, w_207_1787, w_207_1789, w_207_1798, w_207_1800, w_207_1811, w_207_1816, w_207_1821, w_207_1825, w_207_1826, w_207_1827, w_207_1828, w_207_1831, w_207_1832, w_207_1833, w_207_1834, w_207_1835, w_207_1836, w_207_1837, w_207_1838, w_207_1840, w_207_1842, w_207_1843, w_207_1844, w_207_1845, w_207_1846, w_207_1848, w_207_1850, w_207_1851, w_207_1852, w_207_1853, w_207_1854, w_207_1855, w_207_1856, w_207_1857, w_207_1858, w_207_1859, w_207_1860, w_207_1864, w_207_1865, w_207_1866, w_207_1867, w_207_1868, w_207_1869, w_207_1870, w_207_1872, w_207_1874, w_207_1875, w_207_1876, w_207_1877;
  wire w_208_000, w_208_001, w_208_005, w_208_006, w_208_011, w_208_012, w_208_013, w_208_014, w_208_015, w_208_016, w_208_017, w_208_018, w_208_019, w_208_021, w_208_022, w_208_025, w_208_028, w_208_032, w_208_033, w_208_035, w_208_036, w_208_037, w_208_039, w_208_040, w_208_042, w_208_043, w_208_044, w_208_045, w_208_047, w_208_050, w_208_052, w_208_054, w_208_056, w_208_057, w_208_058, w_208_059, w_208_060, w_208_061, w_208_064, w_208_065, w_208_066, w_208_067, w_208_068, w_208_072, w_208_073, w_208_074, w_208_075, w_208_077, w_208_078, w_208_079, w_208_081, w_208_082, w_208_083, w_208_084, w_208_091, w_208_093, w_208_094, w_208_097, w_208_098, w_208_101, w_208_102, w_208_104, w_208_107, w_208_108, w_208_110, w_208_111, w_208_112, w_208_114, w_208_115, w_208_116, w_208_117, w_208_120, w_208_122, w_208_123, w_208_124, w_208_125, w_208_126, w_208_130, w_208_131, w_208_132, w_208_133, w_208_134, w_208_135, w_208_136, w_208_138, w_208_139, w_208_140, w_208_141, w_208_142, w_208_143, w_208_144, w_208_145, w_208_146, w_208_149, w_208_154, w_208_155, w_208_158, w_208_159, w_208_162, w_208_163, w_208_165, w_208_166, w_208_169, w_208_170, w_208_171, w_208_174, w_208_175, w_208_176, w_208_177, w_208_178, w_208_180, w_208_181, w_208_182, w_208_183, w_208_186, w_208_188, w_208_189, w_208_192, w_208_194, w_208_195, w_208_196, w_208_197, w_208_198, w_208_199, w_208_200, w_208_201, w_208_206, w_208_208, w_208_209, w_208_210, w_208_212, w_208_213, w_208_216, w_208_217, w_208_219, w_208_222, w_208_223, w_208_225, w_208_226, w_208_228, w_208_229, w_208_231, w_208_235, w_208_236, w_208_241, w_208_243, w_208_244, w_208_245, w_208_249, w_208_250, w_208_251, w_208_252, w_208_254, w_208_257, w_208_259, w_208_263, w_208_266, w_208_269, w_208_271, w_208_273, w_208_275, w_208_277, w_208_278, w_208_280, w_208_281, w_208_282, w_208_283, w_208_284, w_208_285, w_208_286, w_208_287, w_208_288, w_208_289, w_208_292, w_208_293, w_208_294, w_208_296, w_208_297, w_208_298, w_208_299, w_208_301, w_208_302, w_208_303, w_208_304, w_208_306, w_208_307, w_208_311, w_208_313, w_208_314, w_208_315, w_208_316, w_208_320, w_208_321, w_208_322, w_208_324, w_208_325, w_208_326, w_208_327, w_208_330, w_208_331, w_208_333, w_208_335, w_208_338, w_208_339, w_208_340, w_208_341, w_208_342, w_208_344, w_208_347, w_208_348, w_208_352, w_208_353, w_208_354, w_208_357, w_208_359, w_208_360, w_208_368, w_208_370, w_208_371, w_208_372, w_208_375, w_208_376, w_208_377, w_208_378, w_208_379, w_208_381, w_208_382, w_208_383, w_208_385, w_208_387, w_208_389, w_208_390, w_208_392, w_208_393, w_208_395, w_208_397, w_208_398, w_208_399, w_208_401, w_208_403, w_208_405, w_208_406, w_208_409, w_208_411, w_208_414, w_208_415, w_208_416, w_208_417, w_208_421, w_208_422, w_208_423, w_208_424, w_208_426, w_208_428, w_208_429, w_208_431, w_208_436, w_208_439, w_208_440, w_208_441, w_208_442, w_208_443, w_208_444, w_208_445, w_208_446, w_208_447, w_208_448, w_208_451, w_208_452, w_208_453, w_208_456, w_208_457, w_208_458, w_208_459, w_208_460, w_208_462, w_208_464, w_208_466, w_208_470, w_208_473, w_208_478, w_208_481, w_208_483, w_208_485, w_208_486, w_208_487, w_208_488, w_208_489, w_208_491, w_208_493, w_208_494, w_208_495, w_208_500, w_208_503, w_208_504, w_208_505, w_208_506, w_208_507, w_208_508, w_208_509, w_208_510, w_208_511, w_208_512, w_208_513, w_208_515, w_208_516, w_208_517, w_208_523, w_208_524, w_208_525, w_208_526, w_208_529, w_208_530, w_208_531, w_208_535, w_208_536, w_208_539, w_208_541, w_208_542, w_208_544, w_208_546, w_208_547, w_208_548, w_208_549, w_208_550, w_208_553, w_208_555, w_208_556, w_208_557, w_208_558, w_208_559, w_208_562, w_208_563, w_208_564, w_208_565, w_208_567, w_208_569, w_208_572, w_208_575, w_208_576, w_208_582, w_208_583, w_208_584, w_208_585, w_208_586, w_208_587, w_208_592, w_208_593, w_208_594, w_208_595, w_208_596, w_208_597, w_208_603, w_208_605, w_208_606, w_208_607, w_208_608, w_208_612, w_208_613, w_208_616, w_208_618, w_208_619, w_208_621, w_208_622, w_208_624, w_208_627, w_208_629, w_208_630, w_208_632, w_208_633, w_208_635, w_208_636, w_208_637, w_208_638, w_208_639, w_208_640, w_208_641, w_208_642, w_208_644, w_208_647, w_208_648, w_208_650, w_208_651, w_208_652, w_208_656, w_208_657, w_208_658, w_208_661, w_208_664, w_208_665, w_208_667, w_208_668, w_208_669, w_208_670, w_208_671, w_208_672, w_208_673, w_208_674, w_208_675, w_208_681, w_208_682, w_208_684, w_208_687, w_208_689, w_208_690, w_208_692, w_208_693, w_208_694, w_208_697, w_208_699, w_208_702, w_208_703, w_208_706, w_208_707, w_208_710, w_208_718, w_208_719, w_208_720, w_208_721, w_208_723, w_208_724, w_208_725, w_208_726, w_208_731, w_208_733, w_208_736, w_208_737, w_208_739, w_208_740, w_208_741, w_208_743, w_208_747, w_208_750, w_208_751, w_208_752, w_208_753, w_208_757, w_208_759, w_208_760, w_208_763, w_208_765, w_208_767, w_208_768, w_208_769, w_208_770, w_208_774, w_208_775, w_208_776, w_208_777, w_208_779, w_208_781, w_208_783, w_208_788, w_208_789, w_208_791, w_208_795, w_208_796;
  wire w_209_003, w_209_004, w_209_005, w_209_007, w_209_012, w_209_024, w_209_029, w_209_035, w_209_039, w_209_045, w_209_046, w_209_048, w_209_051, w_209_064, w_209_065, w_209_066, w_209_068, w_209_072, w_209_073, w_209_077, w_209_092, w_209_094, w_209_095, w_209_096, w_209_098, w_209_104, w_209_116, w_209_117, w_209_118, w_209_125, w_209_131, w_209_132, w_209_134, w_209_135, w_209_138, w_209_143, w_209_149, w_209_159, w_209_161, w_209_164, w_209_167, w_209_168, w_209_171, w_209_175, w_209_178, w_209_189, w_209_190, w_209_191, w_209_207, w_209_208, w_209_211, w_209_219, w_209_221, w_209_225, w_209_231, w_209_235, w_209_241, w_209_245, w_209_248, w_209_250, w_209_254, w_209_255, w_209_256, w_209_259, w_209_260, w_209_265, w_209_266, w_209_269, w_209_270, w_209_279, w_209_280, w_209_285, w_209_286, w_209_293, w_209_294, w_209_306, w_209_307, w_209_322, w_209_327, w_209_334, w_209_336, w_209_337, w_209_344, w_209_349, w_209_354, w_209_355, w_209_361, w_209_366, w_209_370, w_209_377, w_209_385, w_209_386, w_209_388, w_209_394, w_209_398, w_209_407, w_209_410, w_209_411, w_209_413, w_209_421, w_209_423, w_209_426, w_209_428, w_209_434, w_209_436, w_209_439, w_209_449, w_209_450, w_209_452, w_209_455, w_209_456, w_209_458, w_209_462, w_209_465, w_209_469, w_209_479, w_209_480, w_209_488, w_209_489, w_209_490, w_209_497, w_209_498, w_209_500, w_209_511, w_209_512, w_209_515, w_209_519, w_209_524, w_209_532, w_209_543, w_209_547, w_209_556, w_209_558, w_209_564, w_209_567, w_209_568, w_209_571, w_209_578, w_209_582, w_209_589, w_209_590, w_209_594, w_209_595, w_209_601, w_209_602, w_209_614, w_209_616, w_209_618, w_209_619, w_209_628, w_209_629, w_209_630, w_209_632, w_209_637, w_209_646, w_209_649, w_209_654, w_209_663, w_209_664, w_209_669, w_209_670, w_209_671, w_209_672, w_209_674, w_209_689, w_209_690, w_209_694, w_209_696, w_209_702, w_209_703, w_209_704, w_209_714, w_209_717, w_209_721, w_209_723, w_209_724, w_209_726, w_209_727, w_209_728, w_209_731, w_209_737, w_209_739, w_209_749, w_209_753, w_209_754, w_209_760, w_209_769, w_209_771, w_209_775, w_209_776, w_209_778, w_209_780, w_209_781, w_209_784, w_209_789, w_209_790, w_209_791, w_209_794, w_209_795, w_209_797, w_209_802, w_209_805, w_209_807, w_209_815, w_209_824, w_209_828, w_209_832, w_209_835, w_209_836, w_209_837, w_209_840, w_209_842, w_209_858, w_209_861, w_209_866, w_209_877, w_209_878, w_209_880, w_209_881, w_209_882, w_209_883, w_209_887, w_209_895, w_209_899, w_209_902, w_209_904, w_209_917, w_209_919, w_209_924, w_209_927, w_209_933, w_209_936, w_209_937, w_209_938, w_209_943, w_209_947, w_209_956, w_209_958, w_209_963, w_209_964, w_209_968, w_209_969, w_209_973, w_209_974, w_209_979, w_209_985, w_209_988, w_209_990, w_209_992, w_209_994, w_209_998, w_209_1000, w_209_1001, w_209_1004, w_209_1006, w_209_1007, w_209_1009, w_209_1013, w_209_1017, w_209_1018, w_209_1020, w_209_1022, w_209_1028, w_209_1036, w_209_1040, w_209_1044, w_209_1049, w_209_1056, w_209_1065, w_209_1068, w_209_1069, w_209_1072, w_209_1075, w_209_1077, w_209_1084, w_209_1087, w_209_1099, w_209_1101, w_209_1102, w_209_1103, w_209_1104, w_209_1108, w_209_1109, w_209_1113, w_209_1121, w_209_1127, w_209_1130, w_209_1140, w_209_1142, w_209_1143, w_209_1144, w_209_1145, w_209_1146, w_209_1150, w_209_1153, w_209_1158, w_209_1159, w_209_1161, w_209_1163, w_209_1165, w_209_1180, w_209_1183, w_209_1185, w_209_1186, w_209_1197, w_209_1198, w_209_1200, w_209_1204, w_209_1206, w_209_1219, w_209_1228, w_209_1229, w_209_1235, w_209_1236, w_209_1253, w_209_1260, w_209_1264, w_209_1269, w_209_1276, w_209_1286, w_209_1289, w_209_1292, w_209_1293, w_209_1303, w_209_1304, w_209_1305, w_209_1311, w_209_1314, w_209_1316, w_209_1324, w_209_1333, w_209_1339, w_209_1347, w_209_1356, w_209_1360, w_209_1366, w_209_1370, w_209_1375, w_209_1377, w_209_1381, w_209_1384, w_209_1388, w_209_1393, w_209_1394, w_209_1400, w_209_1402, w_209_1403, w_209_1409, w_209_1414, w_209_1420, w_209_1421, w_209_1434, w_209_1436, w_209_1449, w_209_1452, w_209_1454, w_209_1460, w_209_1466, w_209_1468, w_209_1477, w_209_1479, w_209_1481, w_209_1482, w_209_1483, w_209_1496, w_209_1505, w_209_1513, w_209_1521, w_209_1528, w_209_1533, w_209_1537, w_209_1539, w_209_1540, w_209_1541, w_209_1546, w_209_1547, w_209_1557, w_209_1561, w_209_1574, w_209_1587, w_209_1591, w_209_1593, w_209_1598, w_209_1600, w_209_1601, w_209_1605, w_209_1606, w_209_1607, w_209_1612, w_209_1614, w_209_1618, w_209_1623, w_209_1628, w_209_1630, w_209_1640, w_209_1641, w_209_1642, w_209_1644, w_209_1650, w_209_1653, w_209_1660, w_209_1662, w_209_1682, w_209_1689, w_209_1690, w_209_1691, w_209_1697, w_209_1711, w_209_1712, w_209_1722, w_209_1726, w_209_1751, w_209_1754, w_209_1785, w_209_1789, w_209_1790, w_209_1806, w_209_1811, w_209_1816, w_209_1817, w_209_1839, w_209_1858, w_209_1859, w_209_1861, w_209_1866, w_209_1874, w_209_1876, w_209_1878, w_209_1879, w_209_1887, w_209_1889, w_209_1896, w_209_1907, w_209_1912, w_209_1914, w_209_1920, w_209_1924, w_209_1930, w_209_1933, w_209_1938, w_209_1956, w_209_1977, w_209_1981, w_209_1991, w_209_1995, w_209_1998, w_209_1999, w_209_2007, w_209_2011, w_209_2016, w_209_2024, w_209_2032, w_209_2033, w_209_2035, w_209_2038, w_209_2040, w_209_2042, w_209_2045, w_209_2062, w_209_2074, w_209_2090, w_209_2091, w_209_2097, w_209_2103, w_209_2104, w_209_2110, w_209_2116, w_209_2120, w_209_2121, w_209_2128, w_209_2131, w_209_2136, w_209_2144, w_209_2149, w_209_2153, w_209_2156, w_209_2160, w_209_2164, w_209_2174, w_209_2178, w_209_2179, w_209_2183, w_209_2199, w_209_2204, w_209_2207, w_209_2219, w_209_2224, w_209_2230, w_209_2243, w_209_2258, w_209_2261, w_209_2265, w_209_2272, w_209_2280, w_209_2285, w_209_2296, w_209_2301, w_209_2317, w_209_2320, w_209_2323, w_209_2328, w_209_2339, w_209_2342, w_209_2345, w_209_2362, w_209_2363, w_209_2384, w_209_2417, w_209_2425, w_209_2435, w_209_2443, w_209_2468, w_209_2482, w_209_2487, w_209_2490, w_209_2500, w_209_2508, w_209_2514, w_209_2515, w_209_2518, w_209_2519, w_209_2539, w_209_2541, w_209_2547, w_209_2549, w_209_2552, w_209_2558, w_209_2562, w_209_2566, w_209_2582, w_209_2584, w_209_2587, w_209_2590, w_209_2600, w_209_2601, w_209_2607, w_209_2613, w_209_2625, w_209_2626, w_209_2633, w_209_2643, w_209_2644, w_209_2655, w_209_2666, w_209_2673, w_209_2682, w_209_2683, w_209_2685, w_209_2689, w_209_2691, w_209_2697, w_209_2699, w_209_2720, w_209_2734, w_209_2739, w_209_2748, w_209_2752, w_209_2754, w_209_2777, w_209_2784, w_209_2795, w_209_2801, w_209_2813, w_209_2823, w_209_2827, w_209_2828, w_209_2840, w_209_2851, w_209_2856, w_209_2868, w_209_2877, w_209_2886, w_209_2896, w_209_2917, w_209_2922, w_209_2923, w_209_2955, w_209_2975, w_209_2990, w_209_2995, w_209_3002, w_209_3003, w_209_3004, w_209_3007, w_209_3013, w_209_3035, w_209_3061, w_209_3066, w_209_3085, w_209_3089, w_209_3090, w_209_3092, w_209_3096, w_209_3123, w_209_3131, w_209_3133, w_209_3138, w_209_3140, w_209_3150, w_209_3157, w_209_3159, w_209_3164, w_209_3165, w_209_3176, w_209_3177, w_209_3189, w_209_3216, w_209_3248, w_209_3251, w_209_3254, w_209_3267, w_209_3272, w_209_3274, w_209_3286, w_209_3289, w_209_3312, w_209_3315;
  wire w_210_001, w_210_004, w_210_005, w_210_006, w_210_012, w_210_013, w_210_014, w_210_016, w_210_018, w_210_019, w_210_025, w_210_026, w_210_029, w_210_030, w_210_031, w_210_035, w_210_036, w_210_037, w_210_038, w_210_040, w_210_044, w_210_047, w_210_049, w_210_050, w_210_052, w_210_053, w_210_055, w_210_059, w_210_060, w_210_061, w_210_063, w_210_064, w_210_065, w_210_069, w_210_072, w_210_073, w_210_075, w_210_077, w_210_080, w_210_081, w_210_087, w_210_088, w_210_091, w_210_092, w_210_095, w_210_098, w_210_099, w_210_102, w_210_103, w_210_106, w_210_107, w_210_110, w_210_112, w_210_113, w_210_114, w_210_116, w_210_119, w_210_121, w_210_124, w_210_126, w_210_127, w_210_129, w_210_132, w_210_136, w_210_138, w_210_143, w_210_144, w_210_146, w_210_147, w_210_151, w_210_155, w_210_159, w_210_161, w_210_163, w_210_165, w_210_169, w_210_174, w_210_176, w_210_178, w_210_182, w_210_184, w_210_189, w_210_190, w_210_192, w_210_193, w_210_197, w_210_201, w_210_203, w_210_204, w_210_205, w_210_206, w_210_208, w_210_209, w_210_211, w_210_212, w_210_219, w_210_220, w_210_224, w_210_229, w_210_230, w_210_237, w_210_238, w_210_239, w_210_241, w_210_242, w_210_247, w_210_248, w_210_254, w_210_255, w_210_257, w_210_261, w_210_265, w_210_270, w_210_273, w_210_274, w_210_277, w_210_279, w_210_280, w_210_284, w_210_286, w_210_288, w_210_289, w_210_291, w_210_292, w_210_293, w_210_294, w_210_295, w_210_296, w_210_297, w_210_298, w_210_302, w_210_303, w_210_304, w_210_305, w_210_308, w_210_311, w_210_313, w_210_315, w_210_317, w_210_318, w_210_321, w_210_325, w_210_328, w_210_329, w_210_330, w_210_333, w_210_334, w_210_340, w_210_341, w_210_342, w_210_343, w_210_345, w_210_349, w_210_351, w_210_352, w_210_354, w_210_356, w_210_357, w_210_363, w_210_364, w_210_365, w_210_371, w_210_373, w_210_379, w_210_382, w_210_383, w_210_384, w_210_385, w_210_388, w_210_389, w_210_391, w_210_393, w_210_398, w_210_399, w_210_402, w_210_403, w_210_404, w_210_406, w_210_409, w_210_410, w_210_411, w_210_414, w_210_415, w_210_417, w_210_420, w_210_424, w_210_436, w_210_442, w_210_444, w_210_448, w_210_449, w_210_453, w_210_454, w_210_456, w_210_460, w_210_461, w_210_464, w_210_474, w_210_476, w_210_483, w_210_484, w_210_487, w_210_490, w_210_494, w_210_495, w_210_497, w_210_499, w_210_501, w_210_506, w_210_508, w_210_512, w_210_513, w_210_515, w_210_516, w_210_517, w_210_518, w_210_522, w_210_524, w_210_525, w_210_527, w_210_532, w_210_536, w_210_537, w_210_540, w_210_546, w_210_552, w_210_559, w_210_571, w_210_572, w_210_577, w_210_578, w_210_580, w_210_581, w_210_584, w_210_585, w_210_587, w_210_590, w_210_592, w_210_595, w_210_597, w_210_598, w_210_602, w_210_605, w_210_606, w_210_609, w_210_610, w_210_613, w_210_615, w_210_620, w_210_622, w_210_623, w_210_627, w_210_638, w_210_639, w_210_645, w_210_646, w_210_647, w_210_652, w_210_654, w_210_676, w_210_678, w_210_686, w_210_687, w_210_689, w_210_692, w_210_697, w_210_698, w_210_700, w_210_704, w_210_705, w_210_709, w_210_715, w_210_717, w_210_718, w_210_719, w_210_720, w_210_721, w_210_725, w_210_731, w_210_733, w_210_734, w_210_738, w_210_741, w_210_744, w_210_749, w_210_750, w_210_752, w_210_753, w_210_755, w_210_756, w_210_758, w_210_761, w_210_763, w_210_764, w_210_776, w_210_779, w_210_783, w_210_784, w_210_786, w_210_787, w_210_788, w_210_790, w_210_793, w_210_797, w_210_798, w_210_800, w_210_801, w_210_803, w_210_804, w_210_806, w_210_808, w_210_810, w_210_811, w_210_812, w_210_814, w_210_817, w_210_818, w_210_819, w_210_823, w_210_825, w_210_827, w_210_831, w_210_842, w_210_844, w_210_848, w_210_849, w_210_853, w_210_857, w_210_860, w_210_861, w_210_871, w_210_872, w_210_875, w_210_876, w_210_879, w_210_882, w_210_884, w_210_885, w_210_886, w_210_887, w_210_890, w_210_891, w_210_892, w_210_894, w_210_896, w_210_897, w_210_900, w_210_901, w_210_902, w_210_903, w_210_904, w_210_905, w_210_906, w_210_907, w_210_910, w_210_913, w_210_914, w_210_919, w_210_922, w_210_925, w_210_926, w_210_927, w_210_930, w_210_931, w_210_933, w_210_934, w_210_936, w_210_938, w_210_940, w_210_941, w_210_943, w_210_949, w_210_950, w_210_954, w_210_961, w_210_962, w_210_964, w_210_967, w_210_968, w_210_969, w_210_972, w_210_973, w_210_978, w_210_982, w_210_985, w_210_988, w_210_989, w_210_997, w_210_1003, w_210_1006, w_210_1008, w_210_1010, w_210_1011, w_210_1016, w_210_1017, w_210_1018, w_210_1020, w_210_1023, w_210_1025, w_210_1026, w_210_1032, w_210_1034, w_210_1036, w_210_1039, w_210_1043, w_210_1044, w_210_1048, w_210_1050, w_210_1051, w_210_1053, w_210_1055, w_210_1059, w_210_1062, w_210_1063, w_210_1064, w_210_1065, w_210_1068, w_210_1069, w_210_1072, w_210_1076, w_210_1077, w_210_1079, w_210_1085, w_210_1086, w_210_1090, w_210_1094, w_210_1100, w_210_1103, w_210_1105, w_210_1108, w_210_1112, w_210_1113, w_210_1116, w_210_1121, w_210_1122, w_210_1127, w_210_1128, w_210_1130, w_210_1131, w_210_1133, w_210_1135, w_210_1137, w_210_1138, w_210_1140, w_210_1142, w_210_1143, w_210_1145, w_210_1148, w_210_1152, w_210_1154, w_210_1156, w_210_1158, w_210_1160, w_210_1161, w_210_1162, w_210_1164, w_210_1169, w_210_1175, w_210_1176, w_210_1177, w_210_1179, w_210_1182, w_210_1192, w_210_1194, w_210_1196, w_210_1200, w_210_1201, w_210_1205, w_210_1207, w_210_1208, w_210_1209, w_210_1210, w_210_1211, w_210_1212, w_210_1219, w_210_1224, w_210_1227;
  wire w_211_011, w_211_013, w_211_025, w_211_028, w_211_031, w_211_043, w_211_044, w_211_049, w_211_051, w_211_060, w_211_074, w_211_079, w_211_080, w_211_081, w_211_083, w_211_096, w_211_099, w_211_100, w_211_106, w_211_112, w_211_130, w_211_144, w_211_145, w_211_148, w_211_156, w_211_160, w_211_163, w_211_164, w_211_168, w_211_182, w_211_201, w_211_207, w_211_208, w_211_211, w_211_217, w_211_218, w_211_231, w_211_234, w_211_238, w_211_239, w_211_246, w_211_256, w_211_259, w_211_260, w_211_265, w_211_268, w_211_270, w_211_273, w_211_278, w_211_285, w_211_288, w_211_292, w_211_294, w_211_299, w_211_302, w_211_309, w_211_324, w_211_325, w_211_340, w_211_343, w_211_344, w_211_345, w_211_347, w_211_349, w_211_369, w_211_370, w_211_373, w_211_377, w_211_381, w_211_384, w_211_386, w_211_387, w_211_388, w_211_391, w_211_397, w_211_398, w_211_404, w_211_405, w_211_409, w_211_412, w_211_429, w_211_433, w_211_435, w_211_443, w_211_444, w_211_448, w_211_449, w_211_453, w_211_464, w_211_468, w_211_478, w_211_480, w_211_483, w_211_487, w_211_492, w_211_498, w_211_502, w_211_507, w_211_517, w_211_521, w_211_524, w_211_525, w_211_526, w_211_530, w_211_532, w_211_533, w_211_536, w_211_537, w_211_539, w_211_546, w_211_551, w_211_558, w_211_561, w_211_565, w_211_567, w_211_575, w_211_578, w_211_580, w_211_584, w_211_587, w_211_588, w_211_590, w_211_593, w_211_605, w_211_614, w_211_623, w_211_625, w_211_633, w_211_637, w_211_640, w_211_643, w_211_644, w_211_647, w_211_667, w_211_676, w_211_678, w_211_684, w_211_685, w_211_687, w_211_688, w_211_694, w_211_696, w_211_698, w_211_704, w_211_714, w_211_719, w_211_722, w_211_723, w_211_726, w_211_738, w_211_757, w_211_761, w_211_764, w_211_766, w_211_769, w_211_777, w_211_778, w_211_784, w_211_794, w_211_795, w_211_804, w_211_807, w_211_813, w_211_820, w_211_821, w_211_823, w_211_826, w_211_828, w_211_837, w_211_861, w_211_864, w_211_866, w_211_875, w_211_877, w_211_880, w_211_888, w_211_889, w_211_891, w_211_896, w_211_897, w_211_900, w_211_901, w_211_906, w_211_915, w_211_917, w_211_918, w_211_947, w_211_949, w_211_951, w_211_962, w_211_966, w_211_975, w_211_980, w_211_981, w_211_985, w_211_986, w_211_987, w_211_989, w_211_994, w_211_995, w_211_1001, w_211_1005, w_211_1010, w_211_1011, w_211_1012, w_211_1020, w_211_1021, w_211_1031, w_211_1038, w_211_1040, w_211_1046, w_211_1047, w_211_1050, w_211_1056, w_211_1058, w_211_1062, w_211_1063, w_211_1073, w_211_1074, w_211_1079, w_211_1089, w_211_1092, w_211_1094, w_211_1098, w_211_1100, w_211_1101, w_211_1103, w_211_1107, w_211_1111, w_211_1112, w_211_1122, w_211_1126, w_211_1128, w_211_1137, w_211_1138, w_211_1144, w_211_1145, w_211_1150, w_211_1157, w_211_1166, w_211_1171, w_211_1177, w_211_1181, w_211_1183, w_211_1184, w_211_1185, w_211_1186, w_211_1187, w_211_1193, w_211_1199, w_211_1205, w_211_1214, w_211_1219, w_211_1221, w_211_1222, w_211_1228, w_211_1231, w_211_1233, w_211_1235, w_211_1240, w_211_1241, w_211_1245, w_211_1252, w_211_1265, w_211_1269, w_211_1274, w_211_1276, w_211_1277, w_211_1279, w_211_1281, w_211_1284, w_211_1287, w_211_1294, w_211_1296, w_211_1300, w_211_1309, w_211_1310, w_211_1316, w_211_1318, w_211_1320, w_211_1330, w_211_1355, w_211_1360, w_211_1393, w_211_1404, w_211_1410, w_211_1416, w_211_1420, w_211_1464, w_211_1467, w_211_1477, w_211_1489, w_211_1492, w_211_1493, w_211_1497, w_211_1504, w_211_1508, w_211_1533, w_211_1560, w_211_1561, w_211_1562, w_211_1567, w_211_1592, w_211_1597, w_211_1602, w_211_1623, w_211_1625, w_211_1627, w_211_1633, w_211_1647, w_211_1661, w_211_1676, w_211_1685, w_211_1713, w_211_1735, w_211_1736, w_211_1759, w_211_1774, w_211_1779, w_211_1784, w_211_1795, w_211_1806, w_211_1815, w_211_1834, w_211_1847, w_211_1858, w_211_1861, w_211_1872, w_211_1880, w_211_1881, w_211_1890, w_211_1904, w_211_1928, w_211_1929, w_211_1930, w_211_1931, w_211_1941, w_211_1943, w_211_1945, w_211_1968, w_211_1974, w_211_1983, w_211_1984, w_211_1990, w_211_2002, w_211_2014, w_211_2032, w_211_2049, w_211_2050, w_211_2055, w_211_2057, w_211_2064, w_211_2067, w_211_2071, w_211_2077, w_211_2084, w_211_2087, w_211_2088, w_211_2092, w_211_2093, w_211_2095, w_211_2115, w_211_2126, w_211_2142, w_211_2150, w_211_2155, w_211_2164, w_211_2170, w_211_2180, w_211_2190, w_211_2199, w_211_2212, w_211_2221, w_211_2222, w_211_2228, w_211_2242, w_211_2245, w_211_2249, w_211_2262, w_211_2264, w_211_2282, w_211_2284, w_211_2286, w_211_2291, w_211_2294, w_211_2298, w_211_2299, w_211_2320, w_211_2337, w_211_2339, w_211_2361, w_211_2366, w_211_2370, w_211_2381, w_211_2394, w_211_2412, w_211_2414, w_211_2416, w_211_2429, w_211_2431, w_211_2434, w_211_2435, w_211_2439, w_211_2493, w_211_2495, w_211_2497, w_211_2505, w_211_2525, w_211_2535, w_211_2536, w_211_2538, w_211_2540, w_211_2545, w_211_2553, w_211_2559, w_211_2564, w_211_2569, w_211_2574, w_211_2581, w_211_2586, w_211_2587, w_211_2606, w_211_2617, w_211_2623, w_211_2631, w_211_2644, w_211_2657, w_211_2676, w_211_2677, w_211_2681, w_211_2682, w_211_2690, w_211_2702, w_211_2703, w_211_2710, w_211_2716, w_211_2721, w_211_2731, w_211_2733, w_211_2758, w_211_2761, w_211_2779, w_211_2784, w_211_2789, w_211_2798, w_211_2802, w_211_2814, w_211_2818, w_211_2836, w_211_2841, w_211_2842, w_211_2848, w_211_2856, w_211_2885, w_211_2904, w_211_2907, w_211_2908, w_211_2909, w_211_2911, w_211_2915, w_211_2916, w_211_2917, w_211_2930, w_211_2939, w_211_2942, w_211_2950, w_211_2958, w_211_2992, w_211_3011, w_211_3027, w_211_3044, w_211_3046, w_211_3053, w_211_3066, w_211_3067, w_211_3074, w_211_3100, w_211_3108, w_211_3112, w_211_3136, w_211_3147, w_211_3154, w_211_3159, w_211_3173, w_211_3196, w_211_3202, w_211_3204, w_211_3208, w_211_3213, w_211_3221, w_211_3228, w_211_3232, w_211_3241, w_211_3249, w_211_3250, w_211_3262, w_211_3265, w_211_3271, w_211_3278, w_211_3287, w_211_3293, w_211_3296, w_211_3305, w_211_3312, w_211_3315, w_211_3317, w_211_3327, w_211_3328, w_211_3334, w_211_3344, w_211_3352, w_211_3364, w_211_3370, w_211_3371, w_211_3381, w_211_3383, w_211_3393, w_211_3401, w_211_3406, w_211_3412, w_211_3433, w_211_3441, w_211_3446, w_211_3451, w_211_3466, w_211_3469, w_211_3470, w_211_3472, w_211_3484, w_211_3493, w_211_3496, w_211_3507, w_211_3520, w_211_3528, w_211_3543, w_211_3565, w_211_3576, w_211_3581, w_211_3582, w_211_3597, w_211_3605, w_211_3606, w_211_3623, w_211_3645, w_211_3646, w_211_3653, w_211_3659, w_211_3662, w_211_3666, w_211_3667, w_211_3668, w_211_3669, w_211_3670, w_211_3671, w_211_3672, w_211_3673, w_211_3675, w_211_3677, w_211_3678, w_211_3679, w_211_3680, w_211_3681, w_211_3682, w_211_3683, w_211_3684, w_211_3685, w_211_3687;
  wire w_212_005, w_212_009, w_212_011, w_212_015, w_212_018, w_212_020, w_212_023, w_212_027, w_212_029, w_212_030, w_212_033, w_212_034, w_212_035, w_212_036, w_212_037, w_212_047, w_212_048, w_212_049, w_212_050, w_212_052, w_212_053, w_212_060, w_212_063, w_212_064, w_212_065, w_212_070, w_212_073, w_212_084, w_212_089, w_212_091, w_212_093, w_212_097, w_212_100, w_212_103, w_212_106, w_212_109, w_212_113, w_212_114, w_212_115, w_212_122, w_212_126, w_212_131, w_212_132, w_212_133, w_212_136, w_212_137, w_212_141, w_212_142, w_212_145, w_212_146, w_212_147, w_212_148, w_212_149, w_212_152, w_212_153, w_212_156, w_212_165, w_212_167, w_212_168, w_212_173, w_212_174, w_212_176, w_212_181, w_212_186, w_212_190, w_212_196, w_212_200, w_212_207, w_212_209, w_212_210, w_212_212, w_212_216, w_212_217, w_212_218, w_212_220, w_212_221, w_212_224, w_212_229, w_212_233, w_212_234, w_212_235, w_212_236, w_212_238, w_212_242, w_212_249, w_212_252, w_212_256, w_212_267, w_212_268, w_212_270, w_212_272, w_212_273, w_212_274, w_212_276, w_212_280, w_212_281, w_212_286, w_212_287, w_212_289, w_212_303, w_212_306, w_212_307, w_212_308, w_212_324, w_212_327, w_212_328, w_212_333, w_212_337, w_212_338, w_212_340, w_212_344, w_212_345, w_212_349, w_212_350, w_212_352, w_212_354, w_212_363, w_212_365, w_212_367, w_212_368, w_212_369, w_212_370, w_212_373, w_212_376, w_212_378, w_212_379, w_212_385, w_212_388, w_212_392, w_212_394, w_212_395, w_212_398, w_212_401, w_212_403, w_212_409, w_212_411, w_212_412, w_212_413, w_212_415, w_212_417, w_212_424, w_212_428, w_212_429, w_212_430, w_212_431, w_212_433, w_212_434, w_212_438, w_212_441, w_212_443, w_212_447, w_212_451, w_212_452, w_212_453, w_212_466, w_212_467, w_212_469, w_212_471, w_212_476, w_212_479, w_212_482, w_212_490, w_212_495, w_212_502, w_212_504, w_212_519, w_212_525, w_212_527, w_212_529, w_212_530, w_212_536, w_212_540, w_212_541, w_212_542, w_212_545, w_212_548, w_212_550, w_212_553, w_212_556, w_212_564, w_212_568, w_212_569, w_212_570, w_212_577, w_212_579, w_212_583, w_212_588, w_212_589, w_212_594, w_212_602, w_212_605, w_212_608, w_212_609, w_212_611, w_212_614, w_212_616, w_212_621, w_212_622, w_212_623, w_212_624, w_212_629, w_212_632, w_212_636, w_212_637, w_212_641, w_212_649, w_212_660, w_212_664, w_212_675, w_212_678, w_212_680, w_212_688, w_212_696, w_212_699, w_212_709, w_212_710, w_212_711, w_212_718, w_212_719, w_212_721, w_212_724, w_212_743, w_212_752, w_212_755, w_212_757, w_212_769, w_212_773, w_212_778, w_212_779, w_212_780, w_212_790, w_212_799, w_212_800, w_212_805, w_212_806, w_212_808, w_212_810, w_212_815, w_212_819, w_212_824, w_212_828, w_212_837, w_212_839, w_212_846, w_212_848, w_212_849, w_212_853, w_212_857, w_212_864, w_212_866, w_212_871, w_212_872, w_212_885, w_212_886, w_212_890, w_212_900, w_212_902, w_212_913, w_212_915, w_212_924, w_212_928, w_212_929, w_212_930, w_212_936, w_212_947, w_212_948, w_212_955, w_212_956, w_212_958, w_212_962, w_212_963, w_212_965, w_212_968, w_212_971, w_212_980, w_212_984, w_212_990, w_212_991, w_212_992, w_212_994, w_212_995, w_212_996, w_212_999, w_212_1000, w_212_1002, w_212_1008, w_212_1010, w_212_1026, w_212_1037, w_212_1046, w_212_1048, w_212_1057, w_212_1064, w_212_1072, w_212_1079, w_212_1080, w_212_1091, w_212_1097, w_212_1102, w_212_1108, w_212_1111, w_212_1119, w_212_1126, w_212_1131, w_212_1132, w_212_1137, w_212_1139, w_212_1143, w_212_1144, w_212_1145, w_212_1146, w_212_1147, w_212_1164, w_212_1165, w_212_1182, w_212_1184, w_212_1186, w_212_1187, w_212_1192, w_212_1198, w_212_1204, w_212_1209, w_212_1211, w_212_1212, w_212_1215, w_212_1217, w_212_1222, w_212_1223, w_212_1224, w_212_1229, w_212_1230, w_212_1245, w_212_1246, w_212_1250, w_212_1253, w_212_1254, w_212_1275, w_212_1282, w_212_1284, w_212_1288, w_212_1289, w_212_1291, w_212_1298, w_212_1303, w_212_1304, w_212_1305, w_212_1306, w_212_1307, w_212_1308, w_212_1312, w_212_1321, w_212_1323, w_212_1328, w_212_1330, w_212_1331, w_212_1343, w_212_1359, w_212_1360, w_212_1362, w_212_1368, w_212_1371, w_212_1375, w_212_1379, w_212_1381, w_212_1384, w_212_1389, w_212_1391, w_212_1393, w_212_1394, w_212_1397, w_212_1403, w_212_1406, w_212_1407, w_212_1421, w_212_1423, w_212_1438, w_212_1463, w_212_1465, w_212_1471, w_212_1479, w_212_1480, w_212_1484, w_212_1486, w_212_1490, w_212_1491, w_212_1492, w_212_1498, w_212_1508, w_212_1510, w_212_1513, w_212_1516, w_212_1519, w_212_1530, w_212_1541, w_212_1542, w_212_1544, w_212_1548, w_212_1554, w_212_1555, w_212_1561, w_212_1564, w_212_1572, w_212_1576, w_212_1579, w_212_1582, w_212_1589, w_212_1597, w_212_1598, w_212_1601, w_212_1612, w_212_1616, w_212_1618, w_212_1621, w_212_1622, w_212_1626, w_212_1631, w_212_1635, w_212_1642, w_212_1648, w_212_1652, w_212_1660, w_212_1662, w_212_1669, w_212_1672, w_212_1683, w_212_1686, w_212_1689, w_212_1690, w_212_1694, w_212_1704, w_212_1707, w_212_1711, w_212_1727, w_212_1731, w_212_1744, w_212_1748, w_212_1753, w_212_1758, w_212_1760, w_212_1762, w_212_1771, w_212_1775, w_212_1783, w_212_1790, w_212_1793, w_212_1794, w_212_1796, w_212_1807, w_212_1816, w_212_1818, w_212_1821, w_212_1822, w_212_1823, w_212_1824, w_212_1834, w_212_1835, w_212_1841, w_212_1842, w_212_1851, w_212_1855, w_212_1856, w_212_1863, w_212_1866, w_212_1868, w_212_1871, w_212_1872, w_212_1874, w_212_1881, w_212_1885, w_212_1891, w_212_1892, w_212_1895, w_212_1899, w_212_1906, w_212_1908, w_212_1918, w_212_1919, w_212_1920, w_212_1921, w_212_1924, w_212_1927, w_212_1935, w_212_1942, w_212_1945, w_212_1952, w_212_1960, w_212_1961, w_212_1964, w_212_1967, w_212_1969, w_212_1977, w_212_1978, w_212_1987, w_212_1989, w_212_1992, w_212_1997, w_212_2000, w_212_2001, w_212_2002, w_212_2004, w_212_2014, w_212_2028, w_212_2033, w_212_2034, w_212_2040, w_212_2042, w_212_2054, w_212_2057, w_212_2083, w_212_2085, w_212_2091, w_212_2092, w_212_2096, w_212_2097, w_212_2104, w_212_2112, w_212_2121, w_212_2130, w_212_2133, w_212_2134, w_212_2136, w_212_2147, w_212_2148, w_212_2149, w_212_2150, w_212_2154, w_212_2158, w_212_2160, w_212_2161, w_212_2162, w_212_2163, w_212_2164, w_212_2165, w_212_2166, w_212_2167, w_212_2168, w_212_2169, w_212_2170;
  wire w_213_005, w_213_008, w_213_009, w_213_011, w_213_014, w_213_020, w_213_026, w_213_033, w_213_034, w_213_035, w_213_037, w_213_041, w_213_042, w_213_045, w_213_048, w_213_061, w_213_063, w_213_067, w_213_070, w_213_074, w_213_077, w_213_081, w_213_084, w_213_091, w_213_097, w_213_098, w_213_101, w_213_105, w_213_107, w_213_111, w_213_117, w_213_124, w_213_126, w_213_129, w_213_133, w_213_135, w_213_137, w_213_142, w_213_147, w_213_159, w_213_161, w_213_165, w_213_175, w_213_197, w_213_198, w_213_204, w_213_206, w_213_214, w_213_225, w_213_228, w_213_230, w_213_231, w_213_237, w_213_242, w_213_244, w_213_249, w_213_257, w_213_261, w_213_262, w_213_273, w_213_283, w_213_288, w_213_289, w_213_292, w_213_301, w_213_304, w_213_305, w_213_310, w_213_312, w_213_326, w_213_343, w_213_344, w_213_345, w_213_347, w_213_363, w_213_372, w_213_378, w_213_382, w_213_383, w_213_391, w_213_400, w_213_401, w_213_402, w_213_404, w_213_410, w_213_415, w_213_418, w_213_420, w_213_424, w_213_427, w_213_433, w_213_440, w_213_442, w_213_443, w_213_445, w_213_447, w_213_454, w_213_455, w_213_461, w_213_462, w_213_467, w_213_473, w_213_476, w_213_480, w_213_490, w_213_492, w_213_493, w_213_495, w_213_501, w_213_502, w_213_508, w_213_512, w_213_514, w_213_515, w_213_517, w_213_531, w_213_532, w_213_533, w_213_534, w_213_535, w_213_537, w_213_541, w_213_549, w_213_555, w_213_559, w_213_560, w_213_563, w_213_564, w_213_565, w_213_576, w_213_581, w_213_583, w_213_585, w_213_587, w_213_589, w_213_598, w_213_608, w_213_612, w_213_620, w_213_624, w_213_629, w_213_638, w_213_642, w_213_651, w_213_661, w_213_662, w_213_667, w_213_670, w_213_673, w_213_683, w_213_684, w_213_686, w_213_696, w_213_697, w_213_701, w_213_703, w_213_707, w_213_711, w_213_714, w_213_719, w_213_720, w_213_730, w_213_738, w_213_747, w_213_750, w_213_755, w_213_756, w_213_767, w_213_770, w_213_771, w_213_774, w_213_778, w_213_788, w_213_790, w_213_794, w_213_796, w_213_798, w_213_799, w_213_806, w_213_812, w_213_815, w_213_818, w_213_819, w_213_823, w_213_825, w_213_827, w_213_832, w_213_835, w_213_839, w_213_840, w_213_841, w_213_846, w_213_849, w_213_850, w_213_854, w_213_856, w_213_857, w_213_859, w_213_860, w_213_862, w_213_871, w_213_873, w_213_876, w_213_877, w_213_881, w_213_883, w_213_884, w_213_887, w_213_902, w_213_904, w_213_905, w_213_908, w_213_913, w_213_914, w_213_919, w_213_921, w_213_924, w_213_926, w_213_936, w_213_938, w_213_945, w_213_947, w_213_949, w_213_952, w_213_953, w_213_954, w_213_955, w_213_969, w_213_977, w_213_980, w_213_986, w_213_997, w_213_1002, w_213_1004, w_213_1010, w_213_1020, w_213_1026, w_213_1031, w_213_1034, w_213_1038, w_213_1043, w_213_1046, w_213_1048, w_213_1055, w_213_1056, w_213_1058, w_213_1067, w_213_1068, w_213_1069, w_213_1083, w_213_1084, w_213_1087, w_213_1092, w_213_1095, w_213_1098, w_213_1103, w_213_1109, w_213_1115, w_213_1121, w_213_1125, w_213_1130, w_213_1135, w_213_1144, w_213_1153, w_213_1158, w_213_1160, w_213_1165, w_213_1166, w_213_1168, w_213_1172, w_213_1174, w_213_1175, w_213_1180, w_213_1186, w_213_1190, w_213_1194, w_213_1196, w_213_1197, w_213_1199, w_213_1201, w_213_1202, w_213_1204, w_213_1205, w_213_1210, w_213_1211, w_213_1212, w_213_1213, w_213_1214, w_213_1226, w_213_1228, w_213_1232, w_213_1238, w_213_1245, w_213_1248, w_213_1249, w_213_1252, w_213_1254, w_213_1259, w_213_1260, w_213_1261, w_213_1262, w_213_1265, w_213_1266, w_213_1277, w_213_1282, w_213_1285, w_213_1290, w_213_1292, w_213_1299, w_213_1302, w_213_1306, w_213_1307, w_213_1316, w_213_1320, w_213_1328, w_213_1333, w_213_1337, w_213_1338, w_213_1346, w_213_1351, w_213_1365, w_213_1374, w_213_1375, w_213_1380, w_213_1381, w_213_1385, w_213_1414, w_213_1416, w_213_1421, w_213_1423, w_213_1426, w_213_1427, w_213_1430, w_213_1433, w_213_1437, w_213_1442, w_213_1445, w_213_1446, w_213_1448, w_213_1452, w_213_1453, w_213_1464, w_213_1471, w_213_1475, w_213_1484, w_213_1486, w_213_1487, w_213_1491, w_213_1492, w_213_1495, w_213_1506, w_213_1511, w_213_1513, w_213_1516, w_213_1520, w_213_1525, w_213_1526, w_213_1529, w_213_1530, w_213_1551, w_213_1553, w_213_1558, w_213_1562, w_213_1565, w_213_1566, w_213_1576, w_213_1578, w_213_1582, w_213_1583, w_213_1586, w_213_1598, w_213_1603, w_213_1606, w_213_1608, w_213_1609, w_213_1621, w_213_1624, w_213_1625, w_213_1626, w_213_1630, w_213_1631, w_213_1633, w_213_1634, w_213_1639, w_213_1641, w_213_1643, w_213_1644, w_213_1650, w_213_1652, w_213_1666, w_213_1673, w_213_1675, w_213_1677, w_213_1678, w_213_1682, w_213_1691, w_213_1694, w_213_1698, w_213_1700, w_213_1702, w_213_1703, w_213_1711, w_213_1714, w_213_1719, w_213_1720, w_213_1735, w_213_1741, w_213_1742, w_213_1748, w_213_1751, w_213_1756, w_213_1761, w_213_1767, w_213_1768, w_213_1771, w_213_1780, w_213_1785, w_213_1788, w_213_1789, w_213_1791, w_213_1796, w_213_1805, w_213_1807, w_213_1808, w_213_1809, w_213_1810, w_213_1812, w_213_1818, w_213_1819, w_213_1828, w_213_1829, w_213_1839, w_213_1849, w_213_1852, w_213_1856, w_213_1859, w_213_1862, w_213_1863, w_213_1869, w_213_1870, w_213_1871, w_213_1874, w_213_1875, w_213_1878, w_213_1884, w_213_1887, w_213_1895, w_213_1913, w_213_1914, w_213_1917, w_213_1919, w_213_1922, w_213_1924, w_213_1927, w_213_1938, w_213_1943, w_213_1946, w_213_1951, w_213_1955, w_213_1957, w_213_1968, w_213_1973, w_213_1984, w_213_1985, w_213_1996, w_213_1997, w_213_2002, w_213_2008, w_213_2011, w_213_2023, w_213_2043, w_213_2047, w_213_2062, w_213_2066, w_213_2072, w_213_2074, w_213_2081, w_213_2087, w_213_2090, w_213_2092, w_213_2097, w_213_2099, w_213_2111, w_213_2133, w_213_2145, w_213_2149, w_213_2155, w_213_2160, w_213_2200, w_213_2221, w_213_2223, w_213_2225, w_213_2231, w_213_2236, w_213_2259, w_213_2266, w_213_2277, w_213_2284, w_213_2291, w_213_2310, w_213_2358, w_213_2361, w_213_2374, w_213_2400, w_213_2401, w_213_2408, w_213_2421, w_213_2426, w_213_2472, w_213_2473, w_213_2494, w_213_2518, w_213_2530, w_213_2540, w_213_2545, w_213_2554, w_213_2564, w_213_2571, w_213_2576, w_213_2583, w_213_2586, w_213_2598, w_213_2627, w_213_2631, w_213_2648, w_213_2656, w_213_2664, w_213_2667, w_213_2670, w_213_2676, w_213_2684, w_213_2716, w_213_2739, w_213_2744, w_213_2771, w_213_2775, w_213_2796, w_213_2805, w_213_2821, w_213_2827, w_213_2832, w_213_2847, w_213_2849, w_213_2850, w_213_2878, w_213_2896, w_213_2897, w_213_2899, w_213_2902, w_213_2916, w_213_2926, w_213_2930, w_213_2959, w_213_2962, w_213_2976, w_213_2979, w_213_2983, w_213_2990, w_213_2992;
  wire w_214_001, w_214_005, w_214_006, w_214_007, w_214_010, w_214_011, w_214_023, w_214_027, w_214_039, w_214_041, w_214_045, w_214_046, w_214_047, w_214_056, w_214_065, w_214_066, w_214_067, w_214_076, w_214_080, w_214_093, w_214_100, w_214_111, w_214_112, w_214_116, w_214_117, w_214_122, w_214_124, w_214_132, w_214_133, w_214_139, w_214_146, w_214_152, w_214_157, w_214_160, w_214_162, w_214_168, w_214_170, w_214_175, w_214_178, w_214_195, w_214_200, w_214_206, w_214_212, w_214_217, w_214_221, w_214_224, w_214_229, w_214_237, w_214_238, w_214_247, w_214_252, w_214_254, w_214_259, w_214_266, w_214_275, w_214_278, w_214_283, w_214_286, w_214_287, w_214_305, w_214_311, w_214_317, w_214_320, w_214_321, w_214_326, w_214_328, w_214_339, w_214_342, w_214_343, w_214_344, w_214_347, w_214_348, w_214_361, w_214_364, w_214_371, w_214_376, w_214_382, w_214_384, w_214_386, w_214_397, w_214_401, w_214_402, w_214_407, w_214_412, w_214_413, w_214_418, w_214_419, w_214_421, w_214_427, w_214_430, w_214_435, w_214_437, w_214_438, w_214_439, w_214_441, w_214_442, w_214_450, w_214_460, w_214_466, w_214_469, w_214_471, w_214_472, w_214_473, w_214_475, w_214_479, w_214_480, w_214_483, w_214_491, w_214_496, w_214_501, w_214_504, w_214_510, w_214_511, w_214_512, w_214_513, w_214_516, w_214_523, w_214_525, w_214_530, w_214_534, w_214_536, w_214_543, w_214_558, w_214_559, w_214_562, w_214_569, w_214_575, w_214_578, w_214_585, w_214_588, w_214_591, w_214_594, w_214_599, w_214_603, w_214_612, w_214_613, w_214_627, w_214_632, w_214_633, w_214_639, w_214_642, w_214_646, w_214_656, w_214_671, w_214_674, w_214_679, w_214_689, w_214_691, w_214_692, w_214_698, w_214_702, w_214_703, w_214_704, w_214_709, w_214_720, w_214_729, w_214_746, w_214_750, w_214_751, w_214_756, w_214_768, w_214_769, w_214_778, w_214_788, w_214_792, w_214_795, w_214_796, w_214_797, w_214_810, w_214_811, w_214_821, w_214_823, w_214_825, w_214_834, w_214_839, w_214_844, w_214_845, w_214_878, w_214_884, w_214_891, w_214_895, w_214_897, w_214_898, w_214_904, w_214_914, w_214_918, w_214_926, w_214_934, w_214_936, w_214_948, w_214_961, w_214_971, w_214_1011, w_214_1026, w_214_1027, w_214_1028, w_214_1041, w_214_1043, w_214_1048, w_214_1071, w_214_1076, w_214_1089, w_214_1093, w_214_1095, w_214_1106, w_214_1115, w_214_1124, w_214_1155, w_214_1159, w_214_1164, w_214_1167, w_214_1188, w_214_1196, w_214_1201, w_214_1227, w_214_1233, w_214_1253, w_214_1257, w_214_1264, w_214_1265, w_214_1289, w_214_1291, w_214_1294, w_214_1297, w_214_1305, w_214_1312, w_214_1318, w_214_1326, w_214_1338, w_214_1346, w_214_1365, w_214_1367, w_214_1376, w_214_1377, w_214_1380, w_214_1381, w_214_1387, w_214_1394, w_214_1395, w_214_1413, w_214_1416, w_214_1431, w_214_1441, w_214_1444, w_214_1449, w_214_1450, w_214_1453, w_214_1462, w_214_1477, w_214_1501, w_214_1504, w_214_1511, w_214_1512, w_214_1520, w_214_1525, w_214_1530, w_214_1538, w_214_1562, w_214_1564, w_214_1569, w_214_1591, w_214_1594, w_214_1600, w_214_1611, w_214_1614, w_214_1630, w_214_1631, w_214_1638, w_214_1643, w_214_1646, w_214_1665, w_214_1668, w_214_1672, w_214_1681, w_214_1683, w_214_1698, w_214_1721, w_214_1730, w_214_1735, w_214_1740, w_214_1749, w_214_1764, w_214_1773, w_214_1786, w_214_1806, w_214_1818, w_214_1820, w_214_1824, w_214_1827, w_214_1843, w_214_1853, w_214_1858, w_214_1887, w_214_1894, w_214_1898, w_214_1924, w_214_1927, w_214_1942, w_214_1948, w_214_1967, w_214_1973, w_214_1988, w_214_2009, w_214_2017, w_214_2028, w_214_2031, w_214_2043, w_214_2054, w_214_2061, w_214_2068, w_214_2104, w_214_2126, w_214_2144, w_214_2148, w_214_2172, w_214_2181, w_214_2182, w_214_2192, w_214_2197, w_214_2227, w_214_2228, w_214_2249, w_214_2251, w_214_2264, w_214_2265, w_214_2266, w_214_2268, w_214_2269, w_214_2279, w_214_2282, w_214_2284, w_214_2288, w_214_2301, w_214_2307, w_214_2312, w_214_2317, w_214_2330, w_214_2365, w_214_2368, w_214_2376, w_214_2387, w_214_2389, w_214_2392, w_214_2402, w_214_2405, w_214_2407, w_214_2411, w_214_2417, w_214_2418, w_214_2423, w_214_2438, w_214_2439, w_214_2440, w_214_2442, w_214_2468, w_214_2484, w_214_2497, w_214_2502, w_214_2510, w_214_2513, w_214_2519, w_214_2530, w_214_2533, w_214_2535, w_214_2573, w_214_2576, w_214_2585, w_214_2599, w_214_2600, w_214_2624, w_214_2625, w_214_2650, w_214_2653, w_214_2663, w_214_2666, w_214_2668, w_214_2672, w_214_2675, w_214_2678, w_214_2696, w_214_2703, w_214_2704, w_214_2707, w_214_2709, w_214_2714, w_214_2720, w_214_2723, w_214_2724, w_214_2742, w_214_2746, w_214_2760, w_214_2784, w_214_2793, w_214_2801, w_214_2806, w_214_2812, w_214_2817, w_214_2822, w_214_2834, w_214_2857, w_214_2879, w_214_2883, w_214_2891, w_214_2892, w_214_2898, w_214_2911, w_214_2923, w_214_2924, w_214_2925, w_214_2931, w_214_2933, w_214_2952, w_214_2959, w_214_2969, w_214_2970, w_214_2972, w_214_2974, w_214_2982, w_214_2998, w_214_2999, w_214_3008, w_214_3031, w_214_3033, w_214_3049, w_214_3055, w_214_3060, w_214_3062, w_214_3067, w_214_3070, w_214_3078, w_214_3090, w_214_3094, w_214_3101, w_214_3104, w_214_3117, w_214_3124, w_214_3129, w_214_3139, w_214_3163, w_214_3210, w_214_3214, w_214_3217, w_214_3221, w_214_3230, w_214_3233, w_214_3258, w_214_3261, w_214_3270, w_214_3275, w_214_3286, w_214_3295, w_214_3297, w_214_3305, w_214_3332, w_214_3346, w_214_3351, w_214_3352, w_214_3361, w_214_3366, w_214_3374, w_214_3382, w_214_3391, w_214_3395, w_214_3397, w_214_3405, w_214_3415, w_214_3417, w_214_3425, w_214_3427, w_214_3429, w_214_3430, w_214_3439, w_214_3443, w_214_3448, w_214_3452, w_214_3457, w_214_3461, w_214_3479, w_214_3488, w_214_3498, w_214_3501, w_214_3508, w_214_3536, w_214_3537, w_214_3540, w_214_3541, w_214_3550, w_214_3560, w_214_3564, w_214_3567, w_214_3570, w_214_3578, w_214_3581, w_214_3586, w_214_3588, w_214_3589, w_214_3594, w_214_3603, w_214_3606, w_214_3615, w_214_3617, w_214_3620, w_214_3629, w_214_3636, w_214_3638, w_214_3641, w_214_3658, w_214_3682, w_214_3683, w_214_3686, w_214_3692, w_214_3698, w_214_3703, w_214_3709, w_214_3738, w_214_3763, w_214_3770, w_214_3774, w_214_3777, w_214_3778, w_214_3792, w_214_3800, w_214_3807, w_214_3810, w_214_3821, w_214_3839, w_214_3849, w_214_3856, w_214_3862, w_214_3866, w_214_3882, w_214_3883, w_214_3886, w_214_3887, w_214_3889, w_214_3915, w_214_3917, w_214_3933, w_214_3940, w_214_3942, w_214_3953, w_214_3959, w_214_3972, w_214_3973, w_214_3979, w_214_3983, w_214_4006, w_214_4027, w_214_4028, w_214_4054, w_214_4059, w_214_4064, w_214_4068, w_214_4091, w_214_4094, w_214_4101, w_214_4108, w_214_4109, w_214_4120, w_214_4124, w_214_4128, w_214_4135, w_214_4149, w_214_4153, w_214_4154, w_214_4167, w_214_4177, w_214_4182, w_214_4183, w_214_4189, w_214_4197, w_214_4228, w_214_4238, w_214_4242, w_214_4288, w_214_4301, w_214_4310, w_214_4321, w_214_4329, w_214_4335, w_214_4341, w_214_4351, w_214_4356;
  wire w_215_000, w_215_001, w_215_003, w_215_005, w_215_006, w_215_007, w_215_009, w_215_010, w_215_012, w_215_013, w_215_014, w_215_015, w_215_016, w_215_017, w_215_018, w_215_019, w_215_020, w_215_021, w_215_022, w_215_023, w_215_024, w_215_025, w_215_026, w_215_027, w_215_028, w_215_029, w_215_030, w_215_031, w_215_032, w_215_033, w_215_034, w_215_035, w_215_036, w_215_037, w_215_038, w_215_039, w_215_040, w_215_041, w_215_042, w_215_043, w_215_044, w_215_045, w_215_046, w_215_047, w_215_048, w_215_049, w_215_050, w_215_051, w_215_052, w_215_053, w_215_054, w_215_055, w_215_056, w_215_057, w_215_058, w_215_059, w_215_060, w_215_061, w_215_062, w_215_063, w_215_064, w_215_065, w_215_067, w_215_068, w_215_069, w_215_070, w_215_071, w_215_072, w_215_073, w_215_074, w_215_075, w_215_076, w_215_077, w_215_078, w_215_079, w_215_080, w_215_081, w_215_082, w_215_083, w_215_084, w_215_085, w_215_086, w_215_088, w_215_089, w_215_090, w_215_091, w_215_092, w_215_093, w_215_094, w_215_095, w_215_096, w_215_097, w_215_098, w_215_099, w_215_100, w_215_101, w_215_102, w_215_103, w_215_104, w_215_105, w_215_106, w_215_107, w_215_108, w_215_109, w_215_110, w_215_111, w_215_112, w_215_113, w_215_114, w_215_116, w_215_117, w_215_118, w_215_119, w_215_120, w_215_121, w_215_122, w_215_123, w_215_124, w_215_125, w_215_126, w_215_127, w_215_128, w_215_129, w_215_130, w_215_133, w_215_134, w_215_135, w_215_136, w_215_137, w_215_139, w_215_140, w_215_141, w_215_142, w_215_144, w_215_146, w_215_147, w_215_148, w_215_149, w_215_150, w_215_152, w_215_154, w_215_155, w_215_156, w_215_157, w_215_158, w_215_159, w_215_160, w_215_162, w_215_163, w_215_164, w_215_165, w_215_166, w_215_167, w_215_168, w_215_169, w_215_170, w_215_171, w_215_172, w_215_173, w_215_174, w_215_175, w_215_176, w_215_177, w_215_178, w_215_180, w_215_181, w_215_182, w_215_184, w_215_185, w_215_186, w_215_187, w_215_188, w_215_189, w_215_191, w_215_192, w_215_193, w_215_194, w_215_195, w_215_196, w_215_197, w_215_198, w_215_199, w_215_200, w_215_201, w_215_202, w_215_203, w_215_204, w_215_205, w_215_206, w_215_207, w_215_208, w_215_210, w_215_211, w_215_212, w_215_213, w_215_214, w_215_215, w_215_216, w_215_218, w_215_219, w_215_220, w_215_221, w_215_222, w_215_223, w_215_224, w_215_225, w_215_226, w_215_227, w_215_228, w_215_229, w_215_230, w_215_231, w_215_232, w_215_233, w_215_235, w_215_236, w_215_237, w_215_238, w_215_239, w_215_240, w_215_241, w_215_242, w_215_243, w_215_244, w_215_245, w_215_246, w_215_247, w_215_249, w_215_250, w_215_251, w_215_252, w_215_253, w_215_254, w_215_255, w_215_256;
  wire w_216_001, w_216_003, w_216_012, w_216_015, w_216_018, w_216_021, w_216_026, w_216_030, w_216_037, w_216_042, w_216_043, w_216_045, w_216_051, w_216_053, w_216_055, w_216_060, w_216_067, w_216_068, w_216_081, w_216_082, w_216_094, w_216_102, w_216_106, w_216_111, w_216_112, w_216_114, w_216_115, w_216_116, w_216_120, w_216_126, w_216_133, w_216_140, w_216_143, w_216_146, w_216_149, w_216_150, w_216_151, w_216_152, w_216_153, w_216_159, w_216_167, w_216_168, w_216_171, w_216_177, w_216_178, w_216_182, w_216_195, w_216_198, w_216_207, w_216_208, w_216_209, w_216_212, w_216_215, w_216_221, w_216_227, w_216_229, w_216_242, w_216_243, w_216_257, w_216_259, w_216_262, w_216_264, w_216_272, w_216_281, w_216_282, w_216_283, w_216_289, w_216_303, w_216_304, w_216_306, w_216_309, w_216_312, w_216_313, w_216_329, w_216_330, w_216_338, w_216_342, w_216_343, w_216_351, w_216_356, w_216_359, w_216_362, w_216_367, w_216_372, w_216_373, w_216_374, w_216_379, w_216_386, w_216_394, w_216_395, w_216_397, w_216_398, w_216_404, w_216_406, w_216_409, w_216_416, w_216_434, w_216_440, w_216_453, w_216_463, w_216_476, w_216_480, w_216_486, w_216_490, w_216_492, w_216_494, w_216_495, w_216_507, w_216_512, w_216_522, w_216_523, w_216_524, w_216_525, w_216_529, w_216_531, w_216_539, w_216_541, w_216_543, w_216_544, w_216_549, w_216_556, w_216_557, w_216_566, w_216_572, w_216_577, w_216_583, w_216_587, w_216_593, w_216_603, w_216_614, w_216_623, w_216_630, w_216_636, w_216_653, w_216_662, w_216_674, w_216_676, w_216_677, w_216_686, w_216_692, w_216_696, w_216_706, w_216_709, w_216_715, w_216_729, w_216_732, w_216_737, w_216_738, w_216_739, w_216_742, w_216_754, w_216_757, w_216_761, w_216_765, w_216_766, w_216_771, w_216_780, w_216_781, w_216_782, w_216_783, w_216_785, w_216_786, w_216_790, w_216_792, w_216_798, w_216_805, w_216_813, w_216_823, w_216_831, w_216_836, w_216_841, w_216_847, w_216_848, w_216_857, w_216_862, w_216_867, w_216_869, w_216_876, w_216_882, w_216_883, w_216_884, w_216_887, w_216_888, w_216_895, w_216_897, w_216_899, w_216_901, w_216_902, w_216_905, w_216_916, w_216_923, w_216_924, w_216_926, w_216_936, w_216_937, w_216_943, w_216_944, w_216_951, w_216_958, w_216_965, w_216_979, w_216_985, w_216_1001, w_216_1004, w_216_1005, w_216_1010, w_216_1036, w_216_1040, w_216_1041, w_216_1045, w_216_1049, w_216_1052, w_216_1054, w_216_1057, w_216_1059, w_216_1062, w_216_1067, w_216_1068, w_216_1069, w_216_1072, w_216_1076, w_216_1090, w_216_1095, w_216_1103, w_216_1105, w_216_1117, w_216_1118, w_216_1119, w_216_1120, w_216_1135, w_216_1140, w_216_1145, w_216_1150, w_216_1152, w_216_1154, w_216_1158, w_216_1162, w_216_1167, w_216_1178, w_216_1181, w_216_1190, w_216_1191, w_216_1193, w_216_1196, w_216_1201, w_216_1202, w_216_1204, w_216_1212, w_216_1213, w_216_1216, w_216_1219, w_216_1227, w_216_1234, w_216_1245, w_216_1247, w_216_1248, w_216_1249, w_216_1250, w_216_1253, w_216_1254, w_216_1258, w_216_1261, w_216_1264, w_216_1267, w_216_1276, w_216_1286, w_216_1288, w_216_1290, w_216_1291, w_216_1298, w_216_1306, w_216_1310, w_216_1315, w_216_1320, w_216_1327, w_216_1338, w_216_1347, w_216_1348, w_216_1353, w_216_1356, w_216_1361, w_216_1377, w_216_1378, w_216_1384, w_216_1385, w_216_1394, w_216_1402, w_216_1403, w_216_1406, w_216_1423, w_216_1424, w_216_1426, w_216_1441, w_216_1481, w_216_1482, w_216_1503, w_216_1515, w_216_1520, w_216_1529, w_216_1550, w_216_1555, w_216_1560, w_216_1566, w_216_1574, w_216_1593, w_216_1614, w_216_1619, w_216_1627, w_216_1635, w_216_1639, w_216_1647, w_216_1651, w_216_1654, w_216_1661, w_216_1668, w_216_1672, w_216_1674, w_216_1689, w_216_1700, w_216_1706, w_216_1716, w_216_1743, w_216_1744, w_216_1764, w_216_1770, w_216_1773, w_216_1776, w_216_1783, w_216_1786, w_216_1811, w_216_1821, w_216_1823, w_216_1824, w_216_1825, w_216_1827, w_216_1828, w_216_1830, w_216_1833, w_216_1834, w_216_1836, w_216_1843, w_216_1845, w_216_1848, w_216_1849, w_216_1851, w_216_1873, w_216_1877, w_216_1887, w_216_1897, w_216_1898, w_216_1900, w_216_1902, w_216_1918, w_216_1927, w_216_1928, w_216_1939, w_216_1953, w_216_1955, w_216_1957, w_216_1960, w_216_1970, w_216_1973, w_216_1977, w_216_1985, w_216_1987, w_216_1988, w_216_1991, w_216_2003, w_216_2013, w_216_2019, w_216_2036, w_216_2048, w_216_2076, w_216_2082, w_216_2084, w_216_2094, w_216_2107, w_216_2108, w_216_2120, w_216_2141, w_216_2142, w_216_2146, w_216_2158, w_216_2167, w_216_2178, w_216_2198, w_216_2210, w_216_2213, w_216_2218, w_216_2220, w_216_2244, w_216_2252, w_216_2253, w_216_2300, w_216_2301, w_216_2314, w_216_2319, w_216_2331, w_216_2355, w_216_2357, w_216_2358, w_216_2378, w_216_2389, w_216_2393, w_216_2397, w_216_2400, w_216_2415, w_216_2451, w_216_2457, w_216_2465, w_216_2467, w_216_2472, w_216_2476, w_216_2483, w_216_2486, w_216_2488, w_216_2492, w_216_2494, w_216_2499, w_216_2510, w_216_2517, w_216_2518, w_216_2524, w_216_2544, w_216_2552, w_216_2564, w_216_2566, w_216_2576, w_216_2589, w_216_2607, w_216_2615, w_216_2626, w_216_2647, w_216_2649, w_216_2655, w_216_2670, w_216_2672, w_216_2682, w_216_2685, w_216_2703, w_216_2704, w_216_2719, w_216_2725, w_216_2733, w_216_2755, w_216_2756, w_216_2757, w_216_2768, w_216_2779, w_216_2784, w_216_2792, w_216_2810, w_216_2821, w_216_2834, w_216_2843, w_216_2846, w_216_2861, w_216_2864, w_216_2866, w_216_2868, w_216_2871, w_216_2873, w_216_2875, w_216_2876, w_216_2879, w_216_2886, w_216_2903, w_216_2940, w_216_2944, w_216_2951, w_216_2966, w_216_2967, w_216_2968, w_216_2977, w_216_2982, w_216_2986, w_216_2992, w_216_3007, w_216_3009, w_216_3010, w_216_3014, w_216_3033, w_216_3037, w_216_3039, w_216_3060, w_216_3062, w_216_3065, w_216_3078, w_216_3081, w_216_3092, w_216_3097, w_216_3105, w_216_3121, w_216_3135, w_216_3160, w_216_3162, w_216_3167, w_216_3168, w_216_3170, w_216_3172, w_216_3202, w_216_3209, w_216_3210, w_216_3214, w_216_3223, w_216_3229, w_216_3235, w_216_3238, w_216_3245, w_216_3250, w_216_3259, w_216_3263, w_216_3275, w_216_3276, w_216_3280, w_216_3289, w_216_3293, w_216_3297, w_216_3298, w_216_3309, w_216_3312, w_216_3314, w_216_3330, w_216_3344, w_216_3352, w_216_3353, w_216_3357, w_216_3359, w_216_3367, w_216_3368, w_216_3378, w_216_3380, w_216_3383, w_216_3386, w_216_3391, w_216_3396, w_216_3413, w_216_3416, w_216_3419, w_216_3424, w_216_3438, w_216_3461, w_216_3463, w_216_3467, w_216_3469, w_216_3475, w_216_3478, w_216_3503, w_216_3505, w_216_3515, w_216_3526, w_216_3541, w_216_3542, w_216_3543, w_216_3548, w_216_3570, w_216_3571, w_216_3573, w_216_3577, w_216_3583, w_216_3591, w_216_3593, w_216_3596, w_216_3632;
  wire w_217_006, w_217_010, w_217_012, w_217_013, w_217_014, w_217_020, w_217_027, w_217_028, w_217_033, w_217_035, w_217_037, w_217_038, w_217_039, w_217_051, w_217_056, w_217_062, w_217_068, w_217_069, w_217_071, w_217_073, w_217_078, w_217_082, w_217_089, w_217_100, w_217_106, w_217_120, w_217_121, w_217_135, w_217_136, w_217_142, w_217_148, w_217_150, w_217_152, w_217_154, w_217_155, w_217_160, w_217_165, w_217_168, w_217_174, w_217_185, w_217_186, w_217_201, w_217_202, w_217_203, w_217_204, w_217_209, w_217_212, w_217_219, w_217_233, w_217_243, w_217_244, w_217_249, w_217_256, w_217_259, w_217_262, w_217_266, w_217_270, w_217_275, w_217_278, w_217_286, w_217_287, w_217_288, w_217_289, w_217_300, w_217_307, w_217_308, w_217_314, w_217_322, w_217_323, w_217_326, w_217_329, w_217_338, w_217_346, w_217_351, w_217_354, w_217_355, w_217_362, w_217_363, w_217_374, w_217_375, w_217_378, w_217_379, w_217_393, w_217_395, w_217_398, w_217_404, w_217_416, w_217_418, w_217_423, w_217_425, w_217_431, w_217_432, w_217_435, w_217_444, w_217_445, w_217_458, w_217_459, w_217_464, w_217_474, w_217_482, w_217_483, w_217_484, w_217_492, w_217_494, w_217_495, w_217_499, w_217_500, w_217_501, w_217_504, w_217_509, w_217_513, w_217_516, w_217_517, w_217_520, w_217_537, w_217_541, w_217_552, w_217_554, w_217_555, w_217_562, w_217_565, w_217_577, w_217_584, w_217_587, w_217_589, w_217_593, w_217_594, w_217_598, w_217_607, w_217_620, w_217_621, w_217_623, w_217_628, w_217_634, w_217_636, w_217_638, w_217_639, w_217_643, w_217_645, w_217_646, w_217_652, w_217_655, w_217_659, w_217_672, w_217_674, w_217_676, w_217_679, w_217_683, w_217_684, w_217_688, w_217_691, w_217_697, w_217_700, w_217_702, w_217_703, w_217_714, w_217_720, w_217_727, w_217_734, w_217_742, w_217_749, w_217_750, w_217_752, w_217_753, w_217_759, w_217_762, w_217_766, w_217_767, w_217_775, w_217_777, w_217_778, w_217_780, w_217_782, w_217_783, w_217_787, w_217_789, w_217_794, w_217_795, w_217_796, w_217_804, w_217_807, w_217_810, w_217_822, w_217_823, w_217_828, w_217_841, w_217_844, w_217_851, w_217_858, w_217_861, w_217_862, w_217_863, w_217_867, w_217_873, w_217_888, w_217_889, w_217_891, w_217_895, w_217_896, w_217_911, w_217_915, w_217_921, w_217_925, w_217_928, w_217_933, w_217_936, w_217_938, w_217_939, w_217_940, w_217_943, w_217_945, w_217_952, w_217_954, w_217_956, w_217_957, w_217_959, w_217_960, w_217_962, w_217_964, w_217_979, w_217_980, w_217_984, w_217_985, w_217_990, w_217_993, w_217_994, w_217_1002, w_217_1003, w_217_1006, w_217_1009, w_217_1012, w_217_1013, w_217_1015, w_217_1023, w_217_1026, w_217_1027, w_217_1036, w_217_1037, w_217_1056, w_217_1057, w_217_1058, w_217_1059, w_217_1061, w_217_1064, w_217_1067, w_217_1069, w_217_1072, w_217_1073, w_217_1079, w_217_1081, w_217_1089, w_217_1094, w_217_1095, w_217_1099, w_217_1100, w_217_1103, w_217_1111, w_217_1113, w_217_1114, w_217_1115, w_217_1117, w_217_1119, w_217_1120, w_217_1123, w_217_1124, w_217_1133, w_217_1136, w_217_1137, w_217_1148, w_217_1149, w_217_1150, w_217_1152, w_217_1158, w_217_1159, w_217_1161, w_217_1164, w_217_1169, w_217_1180, w_217_1184, w_217_1189, w_217_1194, w_217_1196, w_217_1205, w_217_1206, w_217_1207, w_217_1208, w_217_1209, w_217_1215, w_217_1216, w_217_1221, w_217_1227, w_217_1234, w_217_1238, w_217_1241, w_217_1245, w_217_1247, w_217_1252, w_217_1256, w_217_1261, w_217_1263, w_217_1266, w_217_1267, w_217_1272, w_217_1274, w_217_1288, w_217_1289, w_217_1292, w_217_1294, w_217_1298, w_217_1299, w_217_1300, w_217_1315, w_217_1320, w_217_1323, w_217_1326, w_217_1348, w_217_1352, w_217_1353, w_217_1372, w_217_1374, w_217_1377, w_217_1396, w_217_1402, w_217_1404, w_217_1405, w_217_1409, w_217_1411, w_217_1412, w_217_1413, w_217_1418, w_217_1419, w_217_1421, w_217_1427, w_217_1436, w_217_1437, w_217_1457, w_217_1463, w_217_1468, w_217_1474, w_217_1482, w_217_1487, w_217_1492, w_217_1493, w_217_1494, w_217_1504, w_217_1505, w_217_1513, w_217_1514, w_217_1520, w_217_1522, w_217_1527, w_217_1535, w_217_1537, w_217_1538, w_217_1539, w_217_1552, w_217_1553, w_217_1559, w_217_1562, w_217_1564, w_217_1572, w_217_1575, w_217_1580, w_217_1583, w_217_1595, w_217_1604, w_217_1607, w_217_1611, w_217_1618, w_217_1620, w_217_1631, w_217_1633, w_217_1638, w_217_1640, w_217_1641, w_217_1650, w_217_1658, w_217_1665, w_217_1669, w_217_1672, w_217_1679, w_217_1684, w_217_1686, w_217_1696, w_217_1697, w_217_1701, w_217_1703, w_217_1704, w_217_1716, w_217_1717, w_217_1719, w_217_1724, w_217_1726, w_217_1730, w_217_1739, w_217_1742, w_217_1743, w_217_1749, w_217_1750, w_217_1751, w_217_1767, w_217_1775, w_217_1777, w_217_1783, w_217_1784, w_217_1785, w_217_1793, w_217_1797, w_217_1803, w_217_1805, w_217_1806, w_217_1818, w_217_1825, w_217_1829, w_217_1831, w_217_1835, w_217_1837, w_217_1852, w_217_1853, w_217_1855, w_217_1857, w_217_1860, w_217_1861, w_217_1870, w_217_1871, w_217_1888, w_217_1892, w_217_1894, w_217_1896, w_217_1913, w_217_1923, w_217_1928, w_217_1933, w_217_1938, w_217_1942, w_217_1944, w_217_1952, w_217_1959, w_217_1961, w_217_1962, w_217_1966, w_217_1967, w_217_1970, w_217_1973, w_217_1974, w_217_1978, w_217_1979, w_217_1983, w_217_1989, w_217_1992, w_217_2001, w_217_2011, w_217_2016, w_217_2018, w_217_2019, w_217_2020, w_217_2021, w_217_2033, w_217_2035, w_217_2037, w_217_2047, w_217_2056, w_217_2059, w_217_2062, w_217_2063, w_217_2064, w_217_2065, w_217_2066, w_217_2067, w_217_2069, w_217_2073, w_217_2075, w_217_2085, w_217_2094, w_217_2103, w_217_2106, w_217_2126, w_217_2135, w_217_2136, w_217_2144, w_217_2184, w_217_2194, w_217_2215, w_217_2216, w_217_2227, w_217_2235, w_217_2237, w_217_2242, w_217_2246, w_217_2247, w_217_2260, w_217_2263, w_217_2281, w_217_2290, w_217_2295, w_217_2306, w_217_2307, w_217_2308, w_217_2316, w_217_2320, w_217_2331, w_217_2333, w_217_2341, w_217_2342, w_217_2343, w_217_2345, w_217_2350, w_217_2358, w_217_2360, w_217_2373, w_217_2374, w_217_2397, w_217_2401, w_217_2404, w_217_2412, w_217_2425, w_217_2427, w_217_2440, w_217_2454, w_217_2456, w_217_2459, w_217_2463, w_217_2493, w_217_2502, w_217_2503, w_217_2504, w_217_2514, w_217_2522, w_217_2524, w_217_2542, w_217_2559, w_217_2581, w_217_2586, w_217_2594, w_217_2598, w_217_2600, w_217_2612, w_217_2613, w_217_2616, w_217_2622, w_217_2647, w_217_2657, w_217_2658, w_217_2663, w_217_2704, w_217_2708, w_217_2713, w_217_2716, w_217_2718, w_217_2729, w_217_2731, w_217_2732, w_217_2738, w_217_2745, w_217_2748, w_217_2759, w_217_2782, w_217_2784, w_217_2788, w_217_2790, w_217_2791, w_217_2800, w_217_2805, w_217_2806, w_217_2831, w_217_2833, w_217_2844, w_217_2846, w_217_2851, w_217_2856, w_217_2863, w_217_2865, w_217_2867, w_217_2883, w_217_2890;
  wire w_218_004, w_218_007, w_218_009, w_218_010, w_218_020, w_218_024, w_218_027, w_218_029, w_218_030, w_218_032, w_218_038, w_218_040, w_218_045, w_218_046, w_218_052, w_218_054, w_218_063, w_218_070, w_218_075, w_218_083, w_218_085, w_218_086, w_218_088, w_218_099, w_218_100, w_218_103, w_218_111, w_218_112, w_218_114, w_218_122, w_218_125, w_218_126, w_218_131, w_218_157, w_218_163, w_218_165, w_218_168, w_218_176, w_218_181, w_218_183, w_218_185, w_218_188, w_218_204, w_218_207, w_218_209, w_218_217, w_218_219, w_218_220, w_218_228, w_218_231, w_218_232, w_218_233, w_218_235, w_218_243, w_218_245, w_218_246, w_218_247, w_218_248, w_218_256, w_218_259, w_218_270, w_218_271, w_218_277, w_218_278, w_218_279, w_218_284, w_218_288, w_218_291, w_218_294, w_218_297, w_218_313, w_218_314, w_218_315, w_218_317, w_218_318, w_218_331, w_218_335, w_218_342, w_218_363, w_218_364, w_218_366, w_218_368, w_218_369, w_218_374, w_218_384, w_218_387, w_218_389, w_218_391, w_218_394, w_218_398, w_218_402, w_218_406, w_218_410, w_218_420, w_218_424, w_218_425, w_218_427, w_218_434, w_218_435, w_218_436, w_218_437, w_218_444, w_218_450, w_218_453, w_218_462, w_218_464, w_218_468, w_218_473, w_218_479, w_218_484, w_218_485, w_218_493, w_218_504, w_218_507, w_218_520, w_218_521, w_218_525, w_218_527, w_218_532, w_218_544, w_218_546, w_218_549, w_218_552, w_218_554, w_218_555, w_218_557, w_218_559, w_218_560, w_218_561, w_218_565, w_218_570, w_218_573, w_218_584, w_218_592, w_218_596, w_218_609, w_218_610, w_218_612, w_218_614, w_218_615, w_218_617, w_218_618, w_218_623, w_218_624, w_218_625, w_218_630, w_218_632, w_218_635, w_218_645, w_218_647, w_218_658, w_218_659, w_218_662, w_218_664, w_218_675, w_218_684, w_218_689, w_218_693, w_218_696, w_218_707, w_218_709, w_218_713, w_218_723, w_218_726, w_218_727, w_218_728, w_218_734, w_218_735, w_218_742, w_218_746, w_218_753, w_218_754, w_218_758, w_218_759, w_218_764, w_218_769, w_218_775, w_218_780, w_218_781, w_218_785, w_218_793, w_218_795, w_218_797, w_218_800, w_218_804, w_218_809, w_218_811, w_218_815, w_218_826, w_218_834, w_218_840, w_218_856, w_218_863, w_218_864, w_218_871, w_218_890, w_218_894, w_218_904, w_218_905, w_218_910, w_218_925, w_218_926, w_218_935, w_218_946, w_218_948, w_218_949, w_218_963, w_218_968, w_218_971, w_218_979, w_218_982, w_218_984, w_218_1001, w_218_1003, w_218_1006, w_218_1019, w_218_1020, w_218_1022, w_218_1023, w_218_1026, w_218_1032, w_218_1041, w_218_1042, w_218_1043, w_218_1048, w_218_1051, w_218_1052, w_218_1059, w_218_1065, w_218_1067, w_218_1069, w_218_1070, w_218_1073, w_218_1074, w_218_1075, w_218_1082, w_218_1085, w_218_1087, w_218_1088, w_218_1090, w_218_1095, w_218_1097, w_218_1100, w_218_1116, w_218_1117, w_218_1122, w_218_1123, w_218_1143, w_218_1147, w_218_1148, w_218_1151, w_218_1158, w_218_1164, w_218_1167, w_218_1168, w_218_1174, w_218_1177, w_218_1180, w_218_1191, w_218_1192, w_218_1193, w_218_1194, w_218_1204, w_218_1209, w_218_1215, w_218_1217, w_218_1218, w_218_1221, w_218_1230, w_218_1232, w_218_1234, w_218_1235, w_218_1238, w_218_1242, w_218_1245, w_218_1248, w_218_1249, w_218_1252, w_218_1253, w_218_1255, w_218_1264, w_218_1265, w_218_1267, w_218_1274, w_218_1275, w_218_1277, w_218_1279, w_218_1283, w_218_1292, w_218_1293, w_218_1295, w_218_1297, w_218_1303, w_218_1305, w_218_1308, w_218_1320, w_218_1321, w_218_1326, w_218_1327, w_218_1332, w_218_1346, w_218_1347, w_218_1349, w_218_1354, w_218_1356, w_218_1363, w_218_1367, w_218_1370, w_218_1391, w_218_1392, w_218_1399, w_218_1407, w_218_1413, w_218_1414, w_218_1418, w_218_1423, w_218_1429, w_218_1430, w_218_1434, w_218_1440, w_218_1441, w_218_1457, w_218_1459, w_218_1463, w_218_1465, w_218_1470, w_218_1478, w_218_1481, w_218_1484, w_218_1485, w_218_1492, w_218_1502, w_218_1508, w_218_1523, w_218_1524, w_218_1526, w_218_1528, w_218_1532, w_218_1534, w_218_1536, w_218_1552, w_218_1555, w_218_1560, w_218_1568, w_218_1569, w_218_1571, w_218_1574, w_218_1576, w_218_1578, w_218_1579, w_218_1582, w_218_1584, w_218_1585, w_218_1590, w_218_1593, w_218_1602, w_218_1622, w_218_1623, w_218_1626, w_218_1630, w_218_1637, w_218_1638, w_218_1643, w_218_1644, w_218_1649, w_218_1654, w_218_1660, w_218_1664, w_218_1674, w_218_1681, w_218_1684, w_218_1699, w_218_1700, w_218_1713, w_218_1717, w_218_1721, w_218_1727, w_218_1729, w_218_1737, w_218_1739, w_218_1743, w_218_1757, w_218_1765, w_218_1768, w_218_1774, w_218_1777, w_218_1780, w_218_1784, w_218_1790, w_218_1803, w_218_1804, w_218_1806, w_218_1811, w_218_1813, w_218_1814, w_218_1819, w_218_1824, w_218_1825, w_218_1841, w_218_1842, w_218_1848, w_218_1858, w_218_1861, w_218_1870, w_218_1875, w_218_1882, w_218_1886, w_218_1899, w_218_1901, w_218_1904, w_218_1909, w_218_1920, w_218_1923, w_218_1924, w_218_1927, w_218_1947, w_218_1967, w_218_1968, w_218_1985, w_218_1995, w_218_2000, w_218_2001, w_218_2006, w_218_2014, w_218_2017, w_218_2019, w_218_2027, w_218_2046, w_218_2048, w_218_2053, w_218_2056, w_218_2068, w_218_2072, w_218_2082, w_218_2103, w_218_2124, w_218_2137, w_218_2149, w_218_2158, w_218_2183, w_218_2193, w_218_2205, w_218_2212, w_218_2214, w_218_2231, w_218_2249, w_218_2254, w_218_2282, w_218_2296, w_218_2302, w_218_2307, w_218_2308, w_218_2310, w_218_2325, w_218_2330, w_218_2332, w_218_2338, w_218_2341, w_218_2356, w_218_2357, w_218_2363, w_218_2370, w_218_2386, w_218_2389, w_218_2390, w_218_2402, w_218_2411, w_218_2416, w_218_2430, w_218_2432, w_218_2445, w_218_2451, w_218_2469, w_218_2472, w_218_2482, w_218_2491, w_218_2493, w_218_2498, w_218_2510, w_218_2532, w_218_2555, w_218_2563, w_218_2569, w_218_2593, w_218_2599, w_218_2602, w_218_2622, w_218_2624, w_218_2669, w_218_2681, w_218_2686, w_218_2688, w_218_2691, w_218_2718, w_218_2721, w_218_2726, w_218_2735, w_218_2753, w_218_2764, w_218_2770, w_218_2775, w_218_2802, w_218_2807, w_218_2809, w_218_2825, w_218_2831, w_218_2844, w_218_2848, w_218_2870, w_218_2871, w_218_2885, w_218_2886, w_218_2888, w_218_2889, w_218_2903, w_218_2909, w_218_2913, w_218_2937, w_218_2944, w_218_2949, w_218_2952, w_218_2959, w_218_2968, w_218_2985, w_218_2993, w_218_2996, w_218_3003, w_218_3006, w_218_3016, w_218_3017, w_218_3022, w_218_3023, w_218_3027, w_218_3031, w_218_3037, w_218_3051, w_218_3054, w_218_3059, w_218_3062, w_218_3063, w_218_3080, w_218_3085;
  wire w_219_000, w_219_001, w_219_003, w_219_010, w_219_013, w_219_014, w_219_022, w_219_023, w_219_024, w_219_028, w_219_032, w_219_037, w_219_040, w_219_042, w_219_043, w_219_048, w_219_049, w_219_051, w_219_055, w_219_057, w_219_059, w_219_062, w_219_064, w_219_069, w_219_078, w_219_083, w_219_086, w_219_088, w_219_090, w_219_091, w_219_095, w_219_096, w_219_098, w_219_099, w_219_103, w_219_106, w_219_110, w_219_112, w_219_116, w_219_117, w_219_118, w_219_120, w_219_123, w_219_125, w_219_127, w_219_130, w_219_134, w_219_135, w_219_137, w_219_138, w_219_139, w_219_140, w_219_144, w_219_147, w_219_152, w_219_156, w_219_160, w_219_163, w_219_167, w_219_175, w_219_180, w_219_181, w_219_183, w_219_188, w_219_190, w_219_192, w_219_195, w_219_198, w_219_201, w_219_202, w_219_204, w_219_210, w_219_215, w_219_216, w_219_219, w_219_221, w_219_232, w_219_236, w_219_237, w_219_239, w_219_243, w_219_252, w_219_253, w_219_255, w_219_260, w_219_262, w_219_264, w_219_268, w_219_277, w_219_278, w_219_279, w_219_283, w_219_284, w_219_285, w_219_286, w_219_287, w_219_289, w_219_299, w_219_307, w_219_309, w_219_315, w_219_316, w_219_322, w_219_332, w_219_333, w_219_334, w_219_335, w_219_336, w_219_339, w_219_345, w_219_347, w_219_348, w_219_349, w_219_356, w_219_359, w_219_363, w_219_365, w_219_366, w_219_367, w_219_368, w_219_371, w_219_376, w_219_377, w_219_383, w_219_385, w_219_387, w_219_390, w_219_393, w_219_398, w_219_404, w_219_409, w_219_411, w_219_415, w_219_421, w_219_423, w_219_425, w_219_431, w_219_435, w_219_445, w_219_446, w_219_449, w_219_450, w_219_458, w_219_466, w_219_467, w_219_468, w_219_469, w_219_470, w_219_471, w_219_473, w_219_475, w_219_476, w_219_477, w_219_479, w_219_481, w_219_485, w_219_487, w_219_491, w_219_492, w_219_494, w_219_497, w_219_498, w_219_503, w_219_506, w_219_509, w_219_510, w_219_512, w_219_514, w_219_515, w_219_518, w_219_520, w_219_529, w_219_536, w_219_538, w_219_539, w_219_543, w_219_544, w_219_547, w_219_553, w_219_556, w_219_557, w_219_559, w_219_561, w_219_565, w_219_566, w_219_567, w_219_568, w_219_574, w_219_575, w_219_576, w_219_577, w_219_586, w_219_588, w_219_589, w_219_591, w_219_593, w_219_594, w_219_596, w_219_600, w_219_606, w_219_607, w_219_615, w_219_621, w_219_622, w_219_623, w_219_626, w_219_627, w_219_628, w_219_630, w_219_632, w_219_635, w_219_637, w_219_645, w_219_647, w_219_650, w_219_651, w_219_656, w_219_657, w_219_658, w_219_660, w_219_662, w_219_663, w_219_665, w_219_671, w_219_686, w_219_687, w_219_689, w_219_692, w_219_694, w_219_696, w_219_698, w_219_702, w_219_703, w_219_704, w_219_705, w_219_706, w_219_707, w_219_709, w_219_711, w_219_717, w_219_719, w_219_722, w_219_727, w_219_728, w_219_731, w_219_734, w_219_737, w_219_740, w_219_741, w_219_743, w_219_747, w_219_752, w_219_759, w_219_760, w_219_761, w_219_764, w_219_765, w_219_767, w_219_770, w_219_773, w_219_781, w_219_783, w_219_784, w_219_788, w_219_792, w_219_794, w_219_801, w_219_803, w_219_805, w_219_806, w_219_819, w_219_825, w_219_828, w_219_831, w_219_834, w_219_837, w_219_842, w_219_847, w_219_861, w_219_862, w_219_864, w_219_873, w_219_875, w_219_876, w_219_883, w_219_884, w_219_885, w_219_890, w_219_891, w_219_892, w_219_893, w_219_898, w_219_899, w_219_901, w_219_902, w_219_908, w_219_912, w_219_913, w_219_918, w_219_923, w_219_926, w_219_929, w_219_934, w_219_939, w_219_940, w_219_941, w_219_942, w_219_946, w_219_949, w_219_952, w_219_961, w_219_968, w_219_969, w_219_971, w_219_973, w_219_978, w_219_980, w_219_982, w_219_988, w_219_989, w_219_990, w_219_994, w_219_995, w_219_997, w_219_1008, w_219_1016, w_219_1017, w_219_1021, w_219_1022, w_219_1024, w_219_1028, w_219_1030, w_219_1032, w_219_1035, w_219_1038, w_219_1042, w_219_1046, w_219_1051, w_219_1052, w_219_1058, w_219_1059, w_219_1062, w_219_1068, w_219_1070, w_219_1076, w_219_1079, w_219_1082, w_219_1084, w_219_1087, w_219_1090, w_219_1091, w_219_1094, w_219_1096, w_219_1099, w_219_1100, w_219_1101, w_219_1103, w_219_1106, w_219_1108, w_219_1115, w_219_1121, w_219_1124, w_219_1125, w_219_1129, w_219_1130, w_219_1143, w_219_1147, w_219_1148, w_219_1151, w_219_1152, w_219_1156, w_219_1166, w_219_1170, w_219_1176, w_219_1180, w_219_1182, w_219_1195, w_219_1198, w_219_1199, w_219_1204, w_219_1210, w_219_1211, w_219_1212, w_219_1214, w_219_1216, w_219_1219, w_219_1222, w_219_1223, w_219_1227, w_219_1231, w_219_1232, w_219_1233, w_219_1236, w_219_1239, w_219_1241, w_219_1242, w_219_1244, w_219_1248, w_219_1252, w_219_1255, w_219_1260, w_219_1270, w_219_1277, w_219_1278, w_219_1280, w_219_1283, w_219_1287, w_219_1289, w_219_1294, w_219_1300, w_219_1303, w_219_1304, w_219_1308, w_219_1309, w_219_1311, w_219_1318, w_219_1319, w_219_1320, w_219_1321, w_219_1324, w_219_1338, w_219_1339, w_219_1340, w_219_1346, w_219_1349, w_219_1351, w_219_1354, w_219_1358, w_219_1361, w_219_1362, w_219_1364, w_219_1365, w_219_1367, w_219_1368, w_219_1369, w_219_1375, w_219_1378, w_219_1388, w_219_1397, w_219_1399, w_219_1400, w_219_1403, w_219_1409, w_219_1410, w_219_1411, w_219_1416, w_219_1417, w_219_1420, w_219_1422, w_219_1435, w_219_1442, w_219_1445, w_219_1449, w_219_1453, w_219_1458, w_219_1459, w_219_1460, w_219_1470, w_219_1472, w_219_1477, w_219_1479, w_219_1481, w_219_1483, w_219_1487, w_219_1489, w_219_1490, w_219_1499, w_219_1503, w_219_1504, w_219_1513, w_219_1530, w_219_1541, w_219_1543, w_219_1545, w_219_1554, w_219_1558, w_219_1564, w_219_1565, w_219_1573, w_219_1578, w_219_1583, w_219_1585, w_219_1586, w_219_1595, w_219_1602, w_219_1603, w_219_1608, w_219_1609, w_219_1610, w_219_1619, w_219_1623, w_219_1624, w_219_1629, w_219_1640, w_219_1648, w_219_1654, w_219_1657, w_219_1680, w_219_1682, w_219_1686, w_219_1697, w_219_1699, w_219_1701, w_219_1708, w_219_1709, w_219_1717, w_219_1720, w_219_1721, w_219_1729, w_219_1741, w_219_1744, w_219_1747, w_219_1751, w_219_1752, w_219_1753, w_219_1754, w_219_1755, w_219_1756, w_219_1757, w_219_1758, w_219_1762, w_219_1763, w_219_1764, w_219_1765, w_219_1766, w_219_1767, w_219_1768, w_219_1769, w_219_1771;
  wire w_220_000, w_220_004, w_220_005, w_220_006, w_220_008, w_220_009, w_220_014, w_220_018, w_220_020, w_220_030, w_220_033, w_220_036, w_220_042, w_220_043, w_220_049, w_220_054, w_220_058, w_220_060, w_220_062, w_220_064, w_220_065, w_220_067, w_220_071, w_220_079, w_220_083, w_220_092, w_220_096, w_220_099, w_220_102, w_220_108, w_220_112, w_220_124, w_220_151, w_220_159, w_220_160, w_220_164, w_220_165, w_220_179, w_220_185, w_220_186, w_220_192, w_220_199, w_220_214, w_220_215, w_220_230, w_220_231, w_220_237, w_220_238, w_220_245, w_220_250, w_220_252, w_220_256, w_220_271, w_220_274, w_220_277, w_220_279, w_220_286, w_220_293, w_220_294, w_220_304, w_220_313, w_220_321, w_220_323, w_220_326, w_220_331, w_220_345, w_220_348, w_220_355, w_220_358, w_220_364, w_220_369, w_220_386, w_220_388, w_220_395, w_220_403, w_220_405, w_220_407, w_220_410, w_220_411, w_220_413, w_220_423, w_220_430, w_220_434, w_220_440, w_220_448, w_220_454, w_220_457, w_220_461, w_220_465, w_220_467, w_220_474, w_220_476, w_220_478, w_220_482, w_220_485, w_220_486, w_220_487, w_220_490, w_220_496, w_220_499, w_220_503, w_220_514, w_220_518, w_220_526, w_220_527, w_220_538, w_220_540, w_220_542, w_220_547, w_220_548, w_220_553, w_220_555, w_220_559, w_220_560, w_220_569, w_220_574, w_220_581, w_220_582, w_220_585, w_220_586, w_220_589, w_220_592, w_220_594, w_220_606, w_220_607, w_220_611, w_220_618, w_220_620, w_220_622, w_220_633, w_220_634, w_220_639, w_220_641, w_220_642, w_220_673, w_220_675, w_220_687, w_220_699, w_220_701, w_220_702, w_220_715, w_220_718, w_220_728, w_220_730, w_220_736, w_220_737, w_220_743, w_220_747, w_220_759, w_220_760, w_220_765, w_220_766, w_220_772, w_220_773, w_220_774, w_220_780, w_220_786, w_220_787, w_220_789, w_220_790, w_220_796, w_220_797, w_220_812, w_220_822, w_220_825, w_220_833, w_220_837, w_220_839, w_220_852, w_220_866, w_220_884, w_220_888, w_220_897, w_220_902, w_220_911, w_220_912, w_220_913, w_220_920, w_220_923, w_220_924, w_220_928, w_220_935, w_220_936, w_220_938, w_220_939, w_220_940, w_220_951, w_220_952, w_220_953, w_220_1026, w_220_1050, w_220_1067, w_220_1068, w_220_1078, w_220_1086, w_220_1087, w_220_1089, w_220_1098, w_220_1109, w_220_1124, w_220_1125, w_220_1129, w_220_1132, w_220_1134, w_220_1164, w_220_1174, w_220_1179, w_220_1195, w_220_1208, w_220_1224, w_220_1227, w_220_1232, w_220_1235, w_220_1237, w_220_1246, w_220_1247, w_220_1252, w_220_1255, w_220_1262, w_220_1278, w_220_1280, w_220_1297, w_220_1301, w_220_1314, w_220_1321, w_220_1328, w_220_1333, w_220_1339, w_220_1343, w_220_1348, w_220_1358, w_220_1366, w_220_1375, w_220_1378, w_220_1386, w_220_1400, w_220_1431, w_220_1451, w_220_1456, w_220_1458, w_220_1463, w_220_1468, w_220_1469, w_220_1490, w_220_1499, w_220_1500, w_220_1503, w_220_1504, w_220_1514, w_220_1532, w_220_1547, w_220_1562, w_220_1565, w_220_1579, w_220_1581, w_220_1590, w_220_1604, w_220_1606, w_220_1627, w_220_1630, w_220_1645, w_220_1657, w_220_1673, w_220_1682, w_220_1684, w_220_1687, w_220_1688, w_220_1695, w_220_1704, w_220_1709, w_220_1718, w_220_1727, w_220_1735, w_220_1750, w_220_1784, w_220_1796, w_220_1803, w_220_1804, w_220_1818, w_220_1821, w_220_1828, w_220_1835, w_220_1857, w_220_1860, w_220_1862, w_220_1873, w_220_1886, w_220_1897, w_220_1898, w_220_1909, w_220_1914, w_220_1917, w_220_1926, w_220_1931, w_220_1944, w_220_1946, w_220_1957, w_220_1966, w_220_1993, w_220_2010, w_220_2031, w_220_2035, w_220_2042, w_220_2057, w_220_2062, w_220_2086, w_220_2094, w_220_2095, w_220_2116, w_220_2117, w_220_2128, w_220_2131, w_220_2142, w_220_2143, w_220_2153, w_220_2154, w_220_2156, w_220_2160, w_220_2168, w_220_2170, w_220_2178, w_220_2181, w_220_2189, w_220_2207, w_220_2210, w_220_2212, w_220_2217, w_220_2223, w_220_2228, w_220_2234, w_220_2242, w_220_2248, w_220_2250, w_220_2265, w_220_2301, w_220_2306, w_220_2340, w_220_2351, w_220_2356, w_220_2360, w_220_2362, w_220_2365, w_220_2369, w_220_2370, w_220_2376, w_220_2379, w_220_2389, w_220_2402, w_220_2434, w_220_2441, w_220_2442, w_220_2454, w_220_2456, w_220_2471, w_220_2479, w_220_2489, w_220_2516, w_220_2519, w_220_2529, w_220_2536, w_220_2551, w_220_2560, w_220_2564, w_220_2569, w_220_2572, w_220_2594, w_220_2621, w_220_2634, w_220_2639, w_220_2674, w_220_2680, w_220_2684, w_220_2693, w_220_2698, w_220_2700, w_220_2715, w_220_2721, w_220_2724, w_220_2728, w_220_2738, w_220_2741, w_220_2750, w_220_2761, w_220_2780, w_220_2782, w_220_2792, w_220_2798, w_220_2823, w_220_2835, w_220_2839, w_220_2843, w_220_2844, w_220_2847, w_220_2862, w_220_2864, w_220_2875, w_220_2883, w_220_2890, w_220_2900, w_220_2902, w_220_2908, w_220_2909, w_220_2914, w_220_2939, w_220_2943, w_220_2962, w_220_2965, w_220_2968, w_220_2969, w_220_2979, w_220_2985, w_220_2986, w_220_2989, w_220_2991, w_220_3001, w_220_3021, w_220_3057, w_220_3059, w_220_3066, w_220_3068, w_220_3074, w_220_3076, w_220_3088, w_220_3091, w_220_3102, w_220_3104, w_220_3133, w_220_3143, w_220_3144, w_220_3145, w_220_3148, w_220_3153, w_220_3154, w_220_3159, w_220_3161, w_220_3168, w_220_3171, w_220_3206, w_220_3235, w_220_3248, w_220_3253, w_220_3271, w_220_3276, w_220_3289, w_220_3290, w_220_3302, w_220_3313, w_220_3317, w_220_3321, w_220_3329, w_220_3333, w_220_3340, w_220_3354, w_220_3358, w_220_3372, w_220_3373, w_220_3374, w_220_3388, w_220_3392, w_220_3394, w_220_3398, w_220_3409, w_220_3426, w_220_3444, w_220_3450, w_220_3454, w_220_3470, w_220_3481, w_220_3500, w_220_3509, w_220_3537, w_220_3547, w_220_3578, w_220_3597, w_220_3599, w_220_3601, w_220_3621, w_220_3627, w_220_3628, w_220_3630, w_220_3634, w_220_3636, w_220_3638, w_220_3652, w_220_3653, w_220_3655, w_220_3656, w_220_3676, w_220_3687, w_220_3688, w_220_3690, w_220_3693, w_220_3698, w_220_3713, w_220_3721, w_220_3738, w_220_3740, w_220_3753, w_220_3757, w_220_3769, w_220_3797, w_220_3799, w_220_3804, w_220_3823, w_220_3824, w_220_3828, w_220_3829, w_220_3833, w_220_3850, w_220_3851, w_220_3867, w_220_3877, w_220_3897, w_220_3903, w_220_3906, w_220_3910, w_220_3954, w_220_3957, w_220_3967, w_220_3972, w_220_3983, w_220_3984, w_220_3990, w_220_4014, w_220_4030, w_220_4034, w_220_4035, w_220_4036, w_220_4037, w_220_4038, w_220_4042, w_220_4043, w_220_4044, w_220_4045, w_220_4046, w_220_4047, w_220_4048, w_220_4049, w_220_4050, w_220_4051, w_220_4053;
  wire w_221_000, w_221_024, w_221_025, w_221_027, w_221_028, w_221_033, w_221_048, w_221_052, w_221_053, w_221_054, w_221_057, w_221_058, w_221_059, w_221_061, w_221_069, w_221_072, w_221_076, w_221_089, w_221_091, w_221_097, w_221_101, w_221_105, w_221_110, w_221_116, w_221_118, w_221_121, w_221_124, w_221_138, w_221_142, w_221_148, w_221_149, w_221_161, w_221_175, w_221_178, w_221_186, w_221_187, w_221_188, w_221_190, w_221_191, w_221_200, w_221_207, w_221_209, w_221_213, w_221_214, w_221_217, w_221_220, w_221_221, w_221_223, w_221_229, w_221_241, w_221_249, w_221_259, w_221_261, w_221_267, w_221_273, w_221_284, w_221_285, w_221_289, w_221_290, w_221_296, w_221_301, w_221_314, w_221_323, w_221_343, w_221_347, w_221_348, w_221_349, w_221_350, w_221_355, w_221_360, w_221_362, w_221_364, w_221_369, w_221_370, w_221_372, w_221_374, w_221_375, w_221_380, w_221_382, w_221_385, w_221_389, w_221_391, w_221_394, w_221_395, w_221_398, w_221_401, w_221_414, w_221_418, w_221_423, w_221_425, w_221_434, w_221_444, w_221_448, w_221_454, w_221_456, w_221_459, w_221_462, w_221_465, w_221_472, w_221_484, w_221_485, w_221_492, w_221_495, w_221_503, w_221_504, w_221_507, w_221_509, w_221_514, w_221_524, w_221_534, w_221_546, w_221_551, w_221_554, w_221_559, w_221_560, w_221_561, w_221_565, w_221_568, w_221_585, w_221_592, w_221_599, w_221_600, w_221_601, w_221_602, w_221_603, w_221_604, w_221_608, w_221_621, w_221_627, w_221_631, w_221_640, w_221_643, w_221_646, w_221_651, w_221_666, w_221_675, w_221_678, w_221_687, w_221_695, w_221_717, w_221_718, w_221_722, w_221_726, w_221_730, w_221_735, w_221_739, w_221_740, w_221_743, w_221_750, w_221_754, w_221_761, w_221_771, w_221_772, w_221_783, w_221_788, w_221_791, w_221_792, w_221_794, w_221_795, w_221_796, w_221_805, w_221_807, w_221_810, w_221_814, w_221_816, w_221_819, w_221_821, w_221_822, w_221_826, w_221_829, w_221_830, w_221_835, w_221_836, w_221_841, w_221_845, w_221_849, w_221_855, w_221_864, w_221_868, w_221_871, w_221_873, w_221_874, w_221_877, w_221_879, w_221_882, w_221_886, w_221_896, w_221_909, w_221_910, w_221_914, w_221_916, w_221_918, w_221_922, w_221_924, w_221_929, w_221_941, w_221_942, w_221_952, w_221_954, w_221_955, w_221_962, w_221_970, w_221_977, w_221_995, w_221_1005, w_221_1021, w_221_1026, w_221_1030, w_221_1035, w_221_1038, w_221_1042, w_221_1048, w_221_1054, w_221_1056, w_221_1058, w_221_1059, w_221_1060, w_221_1064, w_221_1067, w_221_1069, w_221_1071, w_221_1075, w_221_1084, w_221_1087, w_221_1089, w_221_1094, w_221_1102, w_221_1110, w_221_1114, w_221_1116, w_221_1117, w_221_1126, w_221_1128, w_221_1130, w_221_1133, w_221_1135, w_221_1136, w_221_1137, w_221_1143, w_221_1150, w_221_1152, w_221_1155, w_221_1156, w_221_1161, w_221_1162, w_221_1169, w_221_1170, w_221_1172, w_221_1178, w_221_1185, w_221_1206, w_221_1210, w_221_1216, w_221_1222, w_221_1228, w_221_1230, w_221_1239, w_221_1250, w_221_1265, w_221_1278, w_221_1281, w_221_1287, w_221_1290, w_221_1291, w_221_1292, w_221_1296, w_221_1301, w_221_1303, w_221_1304, w_221_1307, w_221_1311, w_221_1312, w_221_1318, w_221_1321, w_221_1322, w_221_1330, w_221_1342, w_221_1349, w_221_1357, w_221_1364, w_221_1365, w_221_1366, w_221_1367, w_221_1370, w_221_1376, w_221_1380, w_221_1400, w_221_1406, w_221_1414, w_221_1415, w_221_1426, w_221_1427, w_221_1429, w_221_1432, w_221_1438, w_221_1442, w_221_1444, w_221_1460, w_221_1466, w_221_1469, w_221_1473, w_221_1480, w_221_1483, w_221_1487, w_221_1490, w_221_1497, w_221_1498, w_221_1511, w_221_1514, w_221_1529, w_221_1535, w_221_1544, w_221_1545, w_221_1553, w_221_1575, w_221_1578, w_221_1581, w_221_1583, w_221_1591, w_221_1595, w_221_1605, w_221_1615, w_221_1627, w_221_1642, w_221_1643, w_221_1655, w_221_1658, w_221_1663, w_221_1665, w_221_1669, w_221_1670, w_221_1671, w_221_1681, w_221_1682, w_221_1683, w_221_1691, w_221_1693, w_221_1695, w_221_1702, w_221_1707, w_221_1717, w_221_1718, w_221_1729, w_221_1730, w_221_1734, w_221_1735, w_221_1737, w_221_1761, w_221_1768, w_221_1770, w_221_1779, w_221_1803, w_221_1807, w_221_1813, w_221_1822, w_221_1845, w_221_1851, w_221_1852, w_221_1863, w_221_1864, w_221_1889, w_221_1900, w_221_1914, w_221_1917, w_221_1919, w_221_1922, w_221_1931, w_221_1938, w_221_1945, w_221_1948, w_221_1959, w_221_1975, w_221_1991, w_221_2008, w_221_2009, w_221_2020, w_221_2026, w_221_2031, w_221_2054, w_221_2059, w_221_2075, w_221_2081, w_221_2087, w_221_2089, w_221_2132, w_221_2139, w_221_2144, w_221_2150, w_221_2166, w_221_2174, w_221_2181, w_221_2188, w_221_2202, w_221_2205, w_221_2208, w_221_2212, w_221_2217, w_221_2225, w_221_2232, w_221_2236, w_221_2237, w_221_2242, w_221_2247, w_221_2251, w_221_2254, w_221_2257, w_221_2270, w_221_2311, w_221_2321, w_221_2323, w_221_2328, w_221_2333, w_221_2340, w_221_2359, w_221_2360, w_221_2362, w_221_2364, w_221_2392, w_221_2403, w_221_2405, w_221_2407, w_221_2412, w_221_2423, w_221_2424, w_221_2426, w_221_2431, w_221_2442, w_221_2450, w_221_2465, w_221_2467, w_221_2475, w_221_2485, w_221_2488, w_221_2499, w_221_2502, w_221_2532, w_221_2534, w_221_2537, w_221_2539, w_221_2563, w_221_2579, w_221_2591, w_221_2602, w_221_2610, w_221_2635, w_221_2650, w_221_2655, w_221_2656, w_221_2671, w_221_2683, w_221_2687, w_221_2704, w_221_2711, w_221_2714, w_221_2719, w_221_2726, w_221_2738, w_221_2746, w_221_2783, w_221_2784, w_221_2789, w_221_2796, w_221_2833, w_221_2838, w_221_2845, w_221_2852, w_221_2853, w_221_2855, w_221_2859, w_221_2869, w_221_2875, w_221_2889, w_221_2905, w_221_2916, w_221_2937, w_221_2943, w_221_2961, w_221_2964, w_221_2979, w_221_2983, w_221_2997, w_221_3002, w_221_3007, w_221_3030, w_221_3031, w_221_3039, w_221_3055, w_221_3070, w_221_3110, w_221_3116, w_221_3131, w_221_3155, w_221_3157, w_221_3171, w_221_3173, w_221_3176, w_221_3181, w_221_3190, w_221_3193, w_221_3200, w_221_3205, w_221_3210, w_221_3224, w_221_3228, w_221_3248, w_221_3254, w_221_3255;
  wire w_222_001, w_222_002, w_222_005, w_222_006, w_222_007, w_222_008, w_222_010, w_222_011, w_222_013, w_222_014, w_222_015, w_222_016, w_222_017, w_222_021, w_222_024, w_222_025, w_222_029, w_222_030, w_222_031, w_222_035, w_222_036, w_222_037, w_222_039, w_222_041, w_222_043, w_222_045, w_222_046, w_222_050, w_222_052, w_222_056, w_222_057, w_222_059, w_222_060, w_222_061, w_222_062, w_222_066, w_222_069, w_222_073, w_222_074, w_222_076, w_222_081, w_222_082, w_222_085, w_222_086, w_222_090, w_222_092, w_222_093, w_222_096, w_222_098, w_222_100, w_222_102, w_222_103, w_222_108, w_222_110, w_222_111, w_222_114, w_222_116, w_222_118, w_222_119, w_222_123, w_222_127, w_222_129, w_222_130, w_222_131, w_222_133, w_222_134, w_222_137, w_222_139, w_222_144, w_222_145, w_222_148, w_222_149, w_222_150, w_222_152, w_222_153, w_222_154, w_222_155, w_222_156, w_222_158, w_222_162, w_222_163, w_222_165, w_222_166, w_222_168, w_222_172, w_222_175, w_222_176, w_222_181, w_222_183, w_222_184, w_222_186, w_222_187, w_222_188, w_222_190, w_222_191, w_222_192, w_222_194, w_222_195, w_222_197, w_222_200, w_222_201, w_222_205, w_222_207, w_222_208, w_222_209, w_222_211, w_222_212, w_222_214, w_222_215, w_222_217, w_222_219, w_222_220, w_222_221, w_222_222, w_222_230, w_222_231, w_222_232, w_222_233, w_222_234, w_222_237, w_222_238, w_222_239, w_222_241, w_222_242, w_222_245, w_222_246, w_222_248, w_222_249, w_222_251, w_222_255, w_222_257, w_222_258, w_222_261, w_222_263, w_222_269, w_222_270, w_222_271, w_222_274, w_222_276, w_222_277, w_222_279, w_222_280, w_222_282, w_222_283, w_222_284, w_222_287, w_222_288, w_222_290, w_222_291, w_222_292, w_222_296, w_222_298, w_222_300, w_222_301, w_222_303, w_222_304, w_222_305, w_222_312, w_222_313, w_222_314, w_222_317, w_222_318, w_222_320, w_222_324, w_222_331, w_222_332, w_222_334, w_222_336, w_222_337, w_222_340, w_222_341, w_222_342, w_222_343, w_222_344, w_222_349, w_222_350, w_222_353, w_222_355, w_222_357, w_222_358, w_222_361, w_222_364, w_222_372, w_222_375, w_222_378, w_222_382, w_222_384, w_222_386, w_222_387, w_222_392, w_222_393, w_222_394, w_222_396, w_222_397, w_222_398, w_222_401, w_222_402, w_222_403, w_222_404, w_222_408, w_222_410, w_222_411, w_222_414, w_222_416, w_222_417, w_222_418, w_222_419, w_222_422, w_222_424, w_222_427, w_222_428, w_222_430, w_222_432, w_222_434, w_222_436, w_222_437, w_222_438, w_222_443, w_222_444, w_222_447, w_222_448, w_222_451, w_222_452, w_222_454, w_222_455, w_222_456, w_222_457, w_222_458, w_222_459, w_222_460, w_222_461, w_222_463, w_222_464, w_222_465, w_222_467, w_222_469, w_222_470, w_222_471, w_222_478, w_222_479, w_222_482, w_222_485, w_222_486, w_222_488, w_222_491, w_222_493, w_222_494, w_222_495, w_222_503, w_222_505, w_222_506, w_222_509, w_222_512, w_222_513, w_222_515, w_222_518, w_222_520, w_222_521, w_222_522, w_222_531, w_222_535, w_222_536, w_222_537, w_222_538, w_222_539, w_222_540, w_222_542, w_222_544, w_222_545, w_222_546, w_222_548, w_222_553, w_222_555, w_222_556, w_222_558, w_222_561, w_222_562, w_222_563, w_222_566, w_222_568, w_222_571, w_222_575, w_222_577, w_222_578, w_222_579, w_222_580, w_222_581, w_222_586, w_222_587, w_222_589, w_222_590, w_222_592, w_222_598, w_222_601, w_222_602, w_222_607, w_222_608, w_222_610, w_222_611, w_222_612, w_222_613, w_222_619, w_222_621, w_222_624, w_222_627, w_222_629, w_222_631, w_222_633, w_222_639, w_222_643, w_222_644, w_222_646, w_222_650, w_222_652, w_222_653, w_222_656, w_222_660, w_222_662, w_222_665, w_222_666, w_222_668, w_222_669, w_222_678, w_222_682, w_222_683, w_222_685, w_222_689, w_222_696, w_222_699, w_222_700, w_222_704, w_222_706, w_222_707, w_222_710, w_222_711, w_222_718, w_222_721, w_222_723, w_222_725, w_222_727, w_222_729, w_222_730, w_222_738, w_222_740, w_222_744, w_222_748, w_222_750, w_222_755, w_222_756, w_222_759, w_222_760, w_222_761, w_222_765, w_222_766, w_222_770, w_222_774, w_222_775, w_222_777, w_222_779, w_222_781, w_222_784, w_222_785, w_222_788, w_222_793, w_222_798, w_222_799, w_222_800, w_222_802, w_222_804, w_222_807, w_222_808, w_222_810, w_222_812, w_222_815, w_222_818, w_222_821, w_222_825, w_222_826, w_222_827, w_222_831, w_222_833, w_222_834, w_222_840, w_222_842, w_222_844, w_222_845, w_222_847, w_222_850, w_222_851, w_222_852, w_222_853, w_222_854, w_222_856, w_222_861, w_222_862, w_222_863, w_222_864, w_222_865, w_222_866, w_222_867, w_222_870, w_222_872, w_222_874, w_222_875, w_222_876, w_222_877, w_222_879, w_222_881, w_222_883, w_222_886, w_222_889, w_222_890, w_222_893, w_222_897, w_222_898, w_222_899, w_222_901, w_222_902, w_222_903, w_222_905, w_222_907, w_222_908, w_222_909, w_222_910;
  wire w_223_003, w_223_006, w_223_015, w_223_016, w_223_018, w_223_023, w_223_026, w_223_029, w_223_032, w_223_037, w_223_041, w_223_043, w_223_047, w_223_049, w_223_050, w_223_064, w_223_066, w_223_067, w_223_080, w_223_082, w_223_089, w_223_094, w_223_102, w_223_103, w_223_107, w_223_111, w_223_120, w_223_127, w_223_128, w_223_129, w_223_130, w_223_131, w_223_133, w_223_140, w_223_158, w_223_166, w_223_169, w_223_179, w_223_183, w_223_186, w_223_187, w_223_190, w_223_191, w_223_195, w_223_198, w_223_221, w_223_225, w_223_230, w_223_237, w_223_240, w_223_241, w_223_245, w_223_246, w_223_250, w_223_255, w_223_259, w_223_262, w_223_269, w_223_271, w_223_275, w_223_276, w_223_301, w_223_305, w_223_309, w_223_314, w_223_315, w_223_317, w_223_328, w_223_335, w_223_337, w_223_338, w_223_347, w_223_355, w_223_365, w_223_368, w_223_371, w_223_372, w_223_379, w_223_380, w_223_385, w_223_388, w_223_390, w_223_392, w_223_396, w_223_401, w_223_407, w_223_408, w_223_412, w_223_423, w_223_425, w_223_437, w_223_452, w_223_453, w_223_459, w_223_462, w_223_467, w_223_471, w_223_476, w_223_478, w_223_479, w_223_482, w_223_488, w_223_490, w_223_498, w_223_510, w_223_516, w_223_523, w_223_533, w_223_535, w_223_539, w_223_540, w_223_544, w_223_550, w_223_552, w_223_555, w_223_557, w_223_558, w_223_559, w_223_563, w_223_565, w_223_575, w_223_576, w_223_585, w_223_586, w_223_598, w_223_603, w_223_606, w_223_613, w_223_614, w_223_615, w_223_616, w_223_618, w_223_619, w_223_626, w_223_631, w_223_637, w_223_639, w_223_646, w_223_651, w_223_653, w_223_657, w_223_659, w_223_665, w_223_673, w_223_678, w_223_680, w_223_685, w_223_686, w_223_689, w_223_696, w_223_697, w_223_716, w_223_723, w_223_728, w_223_730, w_223_732, w_223_734, w_223_741, w_223_745, w_223_746, w_223_751, w_223_752, w_223_756, w_223_774, w_223_778, w_223_787, w_223_789, w_223_791, w_223_792, w_223_806, w_223_810, w_223_813, w_223_814, w_223_817, w_223_818, w_223_820, w_223_823, w_223_830, w_223_832, w_223_833, w_223_841, w_223_844, w_223_852, w_223_864, w_223_874, w_223_875, w_223_876, w_223_877, w_223_878, w_223_884, w_223_889, w_223_899, w_223_900, w_223_902, w_223_903, w_223_910, w_223_911, w_223_922, w_223_924, w_223_926, w_223_929, w_223_945, w_223_952, w_223_957, w_223_961, w_223_967, w_223_970, w_223_973, w_223_985, w_223_989, w_223_993, w_223_1009, w_223_1010, w_223_1021, w_223_1023, w_223_1030, w_223_1033, w_223_1036, w_223_1038, w_223_1041, w_223_1060, w_223_1062, w_223_1067, w_223_1073, w_223_1075, w_223_1079, w_223_1089, w_223_1095, w_223_1101, w_223_1114, w_223_1120, w_223_1139, w_223_1148, w_223_1159, w_223_1160, w_223_1164, w_223_1167, w_223_1174, w_223_1180, w_223_1183, w_223_1185, w_223_1190, w_223_1197, w_223_1200, w_223_1205, w_223_1209, w_223_1216, w_223_1217, w_223_1228, w_223_1232, w_223_1237, w_223_1238, w_223_1240, w_223_1245, w_223_1249, w_223_1254, w_223_1256, w_223_1258, w_223_1260, w_223_1264, w_223_1266, w_223_1269, w_223_1274, w_223_1279, w_223_1280, w_223_1281, w_223_1282, w_223_1283, w_223_1287, w_223_1296, w_223_1308, w_223_1310, w_223_1323, w_223_1326, w_223_1330, w_223_1344, w_223_1346, w_223_1347, w_223_1350, w_223_1353, w_223_1355, w_223_1356, w_223_1365, w_223_1367, w_223_1382, w_223_1392, w_223_1401, w_223_1403, w_223_1404, w_223_1410, w_223_1412, w_223_1413, w_223_1415, w_223_1425, w_223_1434, w_223_1438, w_223_1443, w_223_1451, w_223_1452, w_223_1457, w_223_1460, w_223_1461, w_223_1464, w_223_1465, w_223_1472, w_223_1473, w_223_1481, w_223_1485, w_223_1487, w_223_1490, w_223_1491, w_223_1492, w_223_1493, w_223_1494, w_223_1499, w_223_1502, w_223_1504, w_223_1505, w_223_1506, w_223_1507, w_223_1513, w_223_1518, w_223_1523, w_223_1545, w_223_1546, w_223_1549, w_223_1551, w_223_1555, w_223_1557, w_223_1574, w_223_1577, w_223_1579, w_223_1583, w_223_1585, w_223_1589, w_223_1590, w_223_1591, w_223_1592, w_223_1594, w_223_1597, w_223_1598, w_223_1599, w_223_1601, w_223_1603, w_223_1605, w_223_1609, w_223_1613, w_223_1620, w_223_1628, w_223_1638, w_223_1645, w_223_1646, w_223_1651, w_223_1656, w_223_1657, w_223_1664, w_223_1665, w_223_1667, w_223_1673, w_223_1683, w_223_1684, w_223_1691, w_223_1693, w_223_1695, w_223_1699, w_223_1702, w_223_1706, w_223_1709, w_223_1714, w_223_1716, w_223_1721, w_223_1726, w_223_1727, w_223_1730, w_223_1736, w_223_1741, w_223_1743, w_223_1747, w_223_1749, w_223_1750, w_223_1751, w_223_1756, w_223_1759, w_223_1762, w_223_1765, w_223_1772, w_223_1779, w_223_1789, w_223_1798, w_223_1801, w_223_1807, w_223_1808, w_223_1810, w_223_1817, w_223_1824, w_223_1825, w_223_1826, w_223_1827, w_223_1828, w_223_1834, w_223_1836, w_223_1837, w_223_1838, w_223_1840, w_223_1843, w_223_1850, w_223_1851, w_223_1852, w_223_1854, w_223_1856, w_223_1861, w_223_1862, w_223_1866, w_223_1869, w_223_1870, w_223_1872, w_223_1874, w_223_1875, w_223_1885, w_223_1889, w_223_1890, w_223_1891, w_223_1895, w_223_1901, w_223_1902, w_223_1908, w_223_1912, w_223_1919, w_223_1920, w_223_1950, w_223_1952, w_223_1957, w_223_1964, w_223_1972, w_223_1974, w_223_1979, w_223_1985, w_223_1995, w_223_2000, w_223_2008, w_223_2012, w_223_2015, w_223_2016, w_223_2017, w_223_2018, w_223_2021, w_223_2022, w_223_2029, w_223_2030, w_223_2031, w_223_2041, w_223_2050, w_223_2059, w_223_2060, w_223_2077, w_223_2081, w_223_2085, w_223_2086, w_223_2091, w_223_2093, w_223_2095, w_223_2097, w_223_2100, w_223_2107, w_223_2111, w_223_2118, w_223_2124, w_223_2126, w_223_2131, w_223_2142, w_223_2146, w_223_2147, w_223_2148, w_223_2149, w_223_2156, w_223_2158, w_223_2163, w_223_2171, w_223_2172, w_223_2177, w_223_2193, w_223_2197, w_223_2198, w_223_2201, w_223_2207, w_223_2214, w_223_2221, w_223_2244, w_223_2245, w_223_2251, w_223_2252, w_223_2253, w_223_2254, w_223_2261, w_223_2267, w_223_2277, w_223_2278, w_223_2280, w_223_2284, w_223_2285, w_223_2291, w_223_2292, w_223_2295, w_223_2296, w_223_2304, w_223_2313, w_223_2316, w_223_2327, w_223_2331, w_223_2335, w_223_2338, w_223_2339, w_223_2344, w_223_2346, w_223_2353, w_223_2356, w_223_2363, w_223_2364, w_223_2370, w_223_2372, w_223_2376, w_223_2383, w_223_2389, w_223_2392, w_223_2398, w_223_2410, w_223_2422, w_223_2423, w_223_2430, w_223_2433, w_223_2435, w_223_2445, w_223_2452, w_223_2454, w_223_2465, w_223_2476, w_223_2477, w_223_2492, w_223_2495, w_223_2502, w_223_2505, w_223_2507, w_223_2512, w_223_2531, w_223_2535, w_223_2556, w_223_2557, w_223_2576, w_223_2578, w_223_2588, w_223_2589, w_223_2604;
  wire w_224_000, w_224_002, w_224_004, w_224_005, w_224_006, w_224_007, w_224_008, w_224_009, w_224_010, w_224_013, w_224_015, w_224_018, w_224_020, w_224_022, w_224_027, w_224_029, w_224_030, w_224_031, w_224_032, w_224_033, w_224_038, w_224_040, w_224_041, w_224_043, w_224_045, w_224_047, w_224_048, w_224_054, w_224_058, w_224_060, w_224_061, w_224_065, w_224_067, w_224_071, w_224_072, w_224_073, w_224_076, w_224_077, w_224_078, w_224_080, w_224_081, w_224_083, w_224_084, w_224_086, w_224_088, w_224_090, w_224_091, w_224_092, w_224_093, w_224_097, w_224_098, w_224_102, w_224_103, w_224_108, w_224_113, w_224_114, w_224_118, w_224_123, w_224_125, w_224_128, w_224_130, w_224_132, w_224_133, w_224_134, w_224_138, w_224_139, w_224_140, w_224_141, w_224_142, w_224_146, w_224_155, w_224_160, w_224_161, w_224_162, w_224_164, w_224_171, w_224_174, w_224_180, w_224_186, w_224_187, w_224_190, w_224_191, w_224_194, w_224_195, w_224_196, w_224_197, w_224_198, w_224_199, w_224_202, w_224_203, w_224_205, w_224_206, w_224_207, w_224_209, w_224_210, w_224_220, w_224_221, w_224_223, w_224_228, w_224_230, w_224_231, w_224_232, w_224_238, w_224_239, w_224_241, w_224_244, w_224_245, w_224_250, w_224_265, w_224_271, w_224_277, w_224_280, w_224_281, w_224_286, w_224_288, w_224_291, w_224_292, w_224_295, w_224_297, w_224_302, w_224_303, w_224_305, w_224_306, w_224_307, w_224_312, w_224_318, w_224_319, w_224_320, w_224_322, w_224_323, w_224_326, w_224_327, w_224_328, w_224_329, w_224_330, w_224_333, w_224_334, w_224_339, w_224_340, w_224_348, w_224_349, w_224_351, w_224_352, w_224_354, w_224_358, w_224_360, w_224_361, w_224_364, w_224_365, w_224_366, w_224_367, w_224_372, w_224_375, w_224_378, w_224_379, w_224_381, w_224_382, w_224_388, w_224_395, w_224_397, w_224_398, w_224_400, w_224_407, w_224_408, w_224_413, w_224_414, w_224_415, w_224_416, w_224_420, w_224_426, w_224_430, w_224_433, w_224_436, w_224_437, w_224_439, w_224_440, w_224_443, w_224_444, w_224_448, w_224_449, w_224_453, w_224_454, w_224_456, w_224_458, w_224_463, w_224_471, w_224_473, w_224_475, w_224_477, w_224_481, w_224_482, w_224_484, w_224_485, w_224_486, w_224_488, w_224_491, w_224_496, w_224_498, w_224_499, w_224_503, w_224_504, w_224_508, w_224_511, w_224_512, w_224_516, w_224_519, w_224_521, w_224_526, w_224_532, w_224_535, w_224_538, w_224_539, w_224_540, w_224_542, w_224_543, w_224_544, w_224_545, w_224_547, w_224_548, w_224_555, w_224_556, w_224_558, w_224_563, w_224_566, w_224_570, w_224_574, w_224_578, w_224_583, w_224_588, w_224_590, w_224_595, w_224_597, w_224_604, w_224_608, w_224_610, w_224_616, w_224_619, w_224_626, w_224_627, w_224_629, w_224_630, w_224_634, w_224_635, w_224_636, w_224_639, w_224_640, w_224_641, w_224_645, w_224_646, w_224_647, w_224_649, w_224_652, w_224_657, w_224_658, w_224_663, w_224_670, w_224_671, w_224_672, w_224_673, w_224_675, w_224_676, w_224_678, w_224_681, w_224_682, w_224_690, w_224_691, w_224_692, w_224_694, w_224_695, w_224_698, w_224_700, w_224_704, w_224_706, w_224_707, w_224_712, w_224_715, w_224_716, w_224_719, w_224_723, w_224_726, w_224_728, w_224_731, w_224_733, w_224_735, w_224_738, w_224_741, w_224_742, w_224_745, w_224_753, w_224_755, w_224_757, w_224_762, w_224_764, w_224_766, w_224_770, w_224_771, w_224_772, w_224_774, w_224_775, w_224_777, w_224_783, w_224_785, w_224_786, w_224_787, w_224_793, w_224_801, w_224_802, w_224_804, w_224_805, w_224_806, w_224_808, w_224_809, w_224_810, w_224_811, w_224_813, w_224_814, w_224_815, w_224_817, w_224_822, w_224_826, w_224_830, w_224_831, w_224_834, w_224_848, w_224_849, w_224_854, w_224_856, w_224_857, w_224_860, w_224_861, w_224_862, w_224_865, w_224_866, w_224_868, w_224_870, w_224_874, w_224_878, w_224_880, w_224_883, w_224_885, w_224_887, w_224_890, w_224_892, w_224_893, w_224_900, w_224_907, w_224_908, w_224_911, w_224_912, w_224_918, w_224_919, w_224_922, w_224_923, w_224_927, w_224_929, w_224_931, w_224_939, w_224_940, w_224_941, w_224_943, w_224_945, w_224_951, w_224_959, w_224_960, w_224_961, w_224_962, w_224_964, w_224_965, w_224_967, w_224_969, w_224_973, w_224_981, w_224_984, w_224_985, w_224_991, w_224_993, w_224_994, w_224_996, w_224_998, w_224_1001, w_224_1004, w_224_1006, w_224_1007, w_224_1010, w_224_1014, w_224_1018, w_224_1023, w_224_1026, w_224_1027, w_224_1030, w_224_1032, w_224_1037, w_224_1040, w_224_1042, w_224_1045, w_224_1049, w_224_1054, w_224_1056, w_224_1057, w_224_1058, w_224_1059, w_224_1062, w_224_1064, w_224_1065, w_224_1066, w_224_1067, w_224_1072, w_224_1079, w_224_1082, w_224_1084, w_224_1087, w_224_1089, w_224_1091, w_224_1092, w_224_1097, w_224_1100, w_224_1103, w_224_1105, w_224_1106, w_224_1108, w_224_1111, w_224_1112, w_224_1113, w_224_1115, w_224_1117, w_224_1122, w_224_1123, w_224_1130, w_224_1131, w_224_1134, w_224_1139, w_224_1140, w_224_1144, w_224_1145, w_224_1148, w_224_1149, w_224_1151, w_224_1154, w_224_1155, w_224_1158, w_224_1160, w_224_1168, w_224_1176, w_224_1181, w_224_1183, w_224_1189, w_224_1190, w_224_1191, w_224_1193, w_224_1194, w_224_1196, w_224_1197, w_224_1198, w_224_1201, w_224_1202, w_224_1204, w_224_1205, w_224_1206, w_224_1207, w_224_1209, w_224_1210, w_224_1211, w_224_1212, w_224_1214, w_224_1217, w_224_1218, w_224_1219, w_224_1221, w_224_1223, w_224_1224, w_224_1225, w_224_1227;
  wire w_225_000, w_225_002, w_225_005, w_225_006, w_225_008, w_225_009, w_225_010, w_225_011, w_225_012, w_225_018, w_225_019, w_225_021, w_225_023, w_225_025, w_225_027, w_225_029, w_225_030, w_225_031, w_225_038, w_225_039, w_225_040, w_225_041, w_225_042, w_225_043, w_225_044, w_225_046, w_225_048, w_225_050, w_225_051, w_225_054, w_225_058, w_225_059, w_225_060, w_225_061, w_225_063, w_225_065, w_225_067, w_225_068, w_225_071, w_225_073, w_225_077, w_225_079, w_225_081, w_225_082, w_225_083, w_225_085, w_225_091, w_225_093, w_225_096, w_225_098, w_225_099, w_225_101, w_225_102, w_225_103, w_225_104, w_225_105, w_225_108, w_225_110, w_225_112, w_225_113, w_225_114, w_225_115, w_225_116, w_225_117, w_225_120, w_225_121, w_225_122, w_225_123, w_225_124, w_225_125, w_225_127, w_225_130, w_225_132, w_225_134, w_225_136, w_225_140, w_225_141, w_225_146, w_225_147, w_225_151, w_225_152, w_225_153, w_225_154, w_225_157, w_225_158, w_225_160, w_225_167, w_225_168, w_225_169, w_225_171, w_225_172, w_225_179, w_225_182, w_225_184, w_225_185, w_225_186, w_225_188, w_225_198, w_225_200, w_225_201, w_225_205, w_225_208, w_225_209, w_225_210, w_225_212, w_225_215, w_225_216, w_225_219, w_225_220, w_225_226, w_225_230, w_225_231, w_225_232, w_225_233, w_225_237, w_225_241, w_225_248, w_225_249, w_225_250, w_225_252, w_225_253, w_225_254, w_225_256, w_225_260, w_225_261, w_225_262, w_225_263, w_225_265, w_225_267, w_225_268, w_225_269, w_225_272, w_225_276, w_225_277, w_225_278, w_225_280, w_225_281, w_225_282, w_225_284, w_225_286, w_225_287, w_225_289, w_225_290, w_225_293, w_225_295, w_225_298, w_225_299, w_225_300, w_225_301, w_225_302, w_225_307, w_225_309, w_225_310, w_225_315, w_225_316, w_225_317, w_225_318, w_225_320, w_225_321, w_225_325, w_225_327, w_225_329, w_225_330, w_225_331, w_225_334, w_225_335, w_225_340, w_225_341, w_225_342, w_225_343, w_225_345, w_225_346, w_225_348, w_225_350, w_225_351, w_225_353, w_225_354, w_225_361, w_225_362, w_225_363, w_225_365, w_225_367, w_225_370, w_225_371, w_225_372, w_225_374, w_225_375, w_225_376, w_225_377, w_225_379, w_225_380, w_225_381, w_225_382, w_225_383, w_225_386, w_225_387, w_225_388, w_225_389, w_225_390, w_225_391, w_225_392, w_225_394, w_225_395, w_225_397, w_225_398, w_225_400, w_225_404, w_225_405, w_225_408, w_225_411, w_225_412, w_225_417, w_225_422, w_225_428, w_225_429, w_225_430, w_225_432, w_225_433, w_225_435, w_225_436, w_225_437, w_225_442, w_225_443, w_225_444, w_225_446, w_225_448, w_225_449, w_225_450, w_225_452, w_225_453, w_225_454, w_225_455, w_225_456, w_225_457, w_225_458, w_225_459, w_225_461, w_225_463, w_225_464, w_225_465, w_225_466, w_225_469, w_225_470, w_225_471, w_225_472, w_225_473, w_225_474, w_225_476, w_225_477, w_225_480, w_225_482, w_225_489, w_225_494, w_225_495, w_225_497, w_225_498, w_225_499, w_225_500, w_225_504, w_225_508, w_225_510, w_225_513, w_225_514, w_225_515, w_225_516, w_225_518, w_225_519, w_225_520, w_225_522, w_225_524, w_225_525, w_225_526, w_225_527, w_225_529, w_225_532, w_225_535, w_225_537, w_225_541, w_225_542, w_225_544, w_225_545, w_225_548, w_225_549, w_225_550, w_225_551, w_225_555, w_225_557, w_225_563, w_225_564, w_225_566, w_225_567, w_225_569, w_225_570, w_225_574, w_225_575, w_225_576, w_225_579, w_225_580, w_225_581, w_225_582, w_225_584, w_225_587, w_225_593, w_225_596, w_225_598, w_225_599, w_225_600, w_225_603, w_225_608, w_225_611, w_225_612, w_225_613, w_225_614, w_225_617, w_225_618, w_225_619, w_225_622, w_225_628, w_225_630, w_225_636, w_225_637, w_225_640, w_225_643, w_225_646, w_225_648, w_225_649, w_225_652, w_225_657, w_225_661, w_225_662, w_225_663, w_225_664, w_225_665, w_225_667, w_225_668, w_225_671, w_225_672, w_225_673, w_225_678, w_225_681, w_225_682, w_225_684, w_225_686, w_225_689, w_225_691, w_225_692, w_225_694, w_225_700, w_225_701, w_225_702, w_225_703, w_225_704, w_225_706, w_225_709, w_225_710, w_225_716, w_225_717, w_225_718, w_225_720, w_225_721, w_225_724, w_225_726, w_225_728, w_225_729, w_225_730, w_225_733, w_225_736, w_225_739, w_225_740, w_225_742, w_225_743, w_225_747, w_225_752, w_225_753, w_225_755, w_225_758, w_225_764, w_225_766, w_225_767, w_225_768, w_225_769, w_225_774, w_225_776, w_225_777, w_225_778, w_225_781, w_225_782, w_225_786, w_225_787, w_225_790, w_225_791, w_225_796, w_225_801, w_225_802, w_225_803, w_225_805, w_225_808, w_225_810, w_225_811, w_225_813, w_225_815, w_225_817, w_225_818, w_225_820, w_225_821, w_225_824, w_225_828, w_225_829, w_225_830, w_225_831, w_225_834, w_225_835, w_225_838, w_225_840, w_225_841, w_225_842, w_225_843, w_225_845, w_225_847, w_225_848, w_225_851, w_225_852, w_225_855, w_225_857, w_225_859, w_225_861, w_225_862, w_225_864, w_225_867, w_225_868, w_225_870, w_225_873, w_225_877, w_225_879, w_225_881, w_225_894, w_225_895, w_225_900;
  wire w_226_002, w_226_004, w_226_011, w_226_020, w_226_023, w_226_025, w_226_026, w_226_027, w_226_035, w_226_039, w_226_041, w_226_046, w_226_056, w_226_061, w_226_063, w_226_070, w_226_082, w_226_094, w_226_097, w_226_103, w_226_108, w_226_109, w_226_114, w_226_122, w_226_128, w_226_132, w_226_134, w_226_139, w_226_143, w_226_148, w_226_150, w_226_156, w_226_157, w_226_171, w_226_173, w_226_175, w_226_177, w_226_179, w_226_181, w_226_185, w_226_187, w_226_208, w_226_210, w_226_211, w_226_213, w_226_221, w_226_235, w_226_237, w_226_240, w_226_242, w_226_244, w_226_248, w_226_257, w_226_263, w_226_274, w_226_278, w_226_279, w_226_296, w_226_299, w_226_313, w_226_314, w_226_315, w_226_317, w_226_325, w_226_331, w_226_337, w_226_338, w_226_339, w_226_343, w_226_344, w_226_349, w_226_354, w_226_355, w_226_356, w_226_358, w_226_365, w_226_376, w_226_377, w_226_385, w_226_387, w_226_390, w_226_394, w_226_397, w_226_404, w_226_406, w_226_413, w_226_414, w_226_420, w_226_426, w_226_430, w_226_431, w_226_443, w_226_453, w_226_460, w_226_462, w_226_469, w_226_474, w_226_478, w_226_490, w_226_494, w_226_497, w_226_506, w_226_507, w_226_516, w_226_517, w_226_518, w_226_519, w_226_520, w_226_523, w_226_528, w_226_531, w_226_539, w_226_544, w_226_550, w_226_552, w_226_562, w_226_595, w_226_605, w_226_606, w_226_611, w_226_612, w_226_617, w_226_618, w_226_619, w_226_621, w_226_624, w_226_631, w_226_636, w_226_641, w_226_642, w_226_652, w_226_653, w_226_657, w_226_676, w_226_680, w_226_686, w_226_695, w_226_699, w_226_713, w_226_724, w_226_727, w_226_729, w_226_736, w_226_737, w_226_738, w_226_740, w_226_743, w_226_745, w_226_760, w_226_767, w_226_772, w_226_775, w_226_777, w_226_778, w_226_789, w_226_797, w_226_801, w_226_815, w_226_829, w_226_842, w_226_846, w_226_853, w_226_863, w_226_867, w_226_870, w_226_872, w_226_873, w_226_875, w_226_877, w_226_879, w_226_894, w_226_906, w_226_907, w_226_912, w_226_913, w_226_916, w_226_917, w_226_924, w_226_934, w_226_940, w_226_942, w_226_945, w_226_951, w_226_960, w_226_961, w_226_964, w_226_965, w_226_972, w_226_990, w_226_991, w_226_1001, w_226_1003, w_226_1009, w_226_1018, w_226_1027, w_226_1030, w_226_1038, w_226_1040, w_226_1056, w_226_1060, w_226_1068, w_226_1079, w_226_1081, w_226_1082, w_226_1099, w_226_1100, w_226_1105, w_226_1109, w_226_1112, w_226_1133, w_226_1152, w_226_1156, w_226_1158, w_226_1161, w_226_1167, w_226_1169, w_226_1171, w_226_1173, w_226_1180, w_226_1181, w_226_1186, w_226_1187, w_226_1199, w_226_1202, w_226_1206, w_226_1208, w_226_1214, w_226_1216, w_226_1227, w_226_1228, w_226_1232, w_226_1240, w_226_1243, w_226_1245, w_226_1247, w_226_1249, w_226_1253, w_226_1254, w_226_1260, w_226_1267, w_226_1270, w_226_1276, w_226_1290, w_226_1298, w_226_1304, w_226_1310, w_226_1316, w_226_1335, w_226_1340, w_226_1341, w_226_1344, w_226_1348, w_226_1349, w_226_1355, w_226_1361, w_226_1362, w_226_1365, w_226_1367, w_226_1370, w_226_1379, w_226_1381, w_226_1382, w_226_1383, w_226_1387, w_226_1401, w_226_1407, w_226_1408, w_226_1409, w_226_1414, w_226_1415, w_226_1417, w_226_1419, w_226_1421, w_226_1427, w_226_1432, w_226_1444, w_226_1450, w_226_1454, w_226_1467, w_226_1474, w_226_1479, w_226_1500, w_226_1501, w_226_1503, w_226_1511, w_226_1517, w_226_1523, w_226_1528, w_226_1532, w_226_1540, w_226_1547, w_226_1550, w_226_1552, w_226_1574, w_226_1578, w_226_1584, w_226_1585, w_226_1589, w_226_1593, w_226_1597, w_226_1600, w_226_1603, w_226_1611, w_226_1613, w_226_1625, w_226_1628, w_226_1634, w_226_1641, w_226_1647, w_226_1650, w_226_1651, w_226_1653, w_226_1661, w_226_1668, w_226_1669, w_226_1670, w_226_1675, w_226_1681, w_226_1689, w_226_1695, w_226_1702, w_226_1716, w_226_1733, w_226_1754, w_226_1755, w_226_1757, w_226_1763, w_226_1766, w_226_1768, w_226_1776, w_226_1777, w_226_1779, w_226_1780, w_226_1784, w_226_1796, w_226_1806, w_226_1807, w_226_1812, w_226_1816, w_226_1818, w_226_1824, w_226_1828, w_226_1834, w_226_1835, w_226_1836, w_226_1847, w_226_1850, w_226_1867, w_226_1871, w_226_1876, w_226_1882, w_226_1885, w_226_1891, w_226_1892, w_226_1896, w_226_1904, w_226_1907, w_226_1911, w_226_1913, w_226_1916, w_226_1917, w_226_1922, w_226_1925, w_226_1936, w_226_1941, w_226_1952, w_226_1957, w_226_1958, w_226_1970, w_226_1974, w_226_1980, w_226_1988, w_226_1992, w_226_1993, w_226_1998, w_226_2014, w_226_2024, w_226_2031, w_226_2057, w_226_2060, w_226_2073, w_226_2074, w_226_2078, w_226_2082, w_226_2105, w_226_2119, w_226_2121, w_226_2139, w_226_2142, w_226_2153, w_226_2172, w_226_2190, w_226_2196, w_226_2203, w_226_2204, w_226_2216, w_226_2221, w_226_2247, w_226_2250, w_226_2256, w_226_2260, w_226_2271, w_226_2274, w_226_2282, w_226_2284, w_226_2293, w_226_2295, w_226_2300, w_226_2321, w_226_2338, w_226_2349, w_226_2353, w_226_2354, w_226_2356, w_226_2370, w_226_2378, w_226_2381, w_226_2399, w_226_2405, w_226_2422, w_226_2425, w_226_2428, w_226_2461, w_226_2463, w_226_2485, w_226_2488, w_226_2490, w_226_2507, w_226_2514, w_226_2541, w_226_2543, w_226_2552, w_226_2567, w_226_2583, w_226_2590, w_226_2591, w_226_2592, w_226_2596, w_226_2605, w_226_2609, w_226_2611, w_226_2613, w_226_2651, w_226_2665, w_226_2666, w_226_2669, w_226_2671, w_226_2687, w_226_2708, w_226_2726, w_226_2733, w_226_2741, w_226_2744, w_226_2751, w_226_2778, w_226_2784, w_226_2795, w_226_2801, w_226_2807, w_226_2814, w_226_2816, w_226_2827, w_226_2829, w_226_2837, w_226_2841, w_226_2857, w_226_2865, w_226_2866, w_226_2869, w_226_2891, w_226_2903, w_226_2909, w_226_2923, w_226_2944, w_226_2948, w_226_2951, w_226_2957, w_226_2964, w_226_2969, w_226_2975;
  wire w_227_002, w_227_004, w_227_007, w_227_010, w_227_015, w_227_018, w_227_021, w_227_024, w_227_029, w_227_031, w_227_033, w_227_035, w_227_036, w_227_037, w_227_039, w_227_048, w_227_049, w_227_055, w_227_058, w_227_059, w_227_061, w_227_063, w_227_065, w_227_068, w_227_070, w_227_071, w_227_075, w_227_077, w_227_091, w_227_093, w_227_094, w_227_096, w_227_102, w_227_105, w_227_106, w_227_116, w_227_119, w_227_120, w_227_121, w_227_122, w_227_127, w_227_129, w_227_130, w_227_131, w_227_135, w_227_137, w_227_142, w_227_151, w_227_157, w_227_158, w_227_161, w_227_165, w_227_169, w_227_182, w_227_183, w_227_186, w_227_189, w_227_196, w_227_197, w_227_198, w_227_201, w_227_210, w_227_212, w_227_219, w_227_226, w_227_235, w_227_240, w_227_243, w_227_252, w_227_255, w_227_260, w_227_261, w_227_262, w_227_263, w_227_264, w_227_265, w_227_273, w_227_280, w_227_286, w_227_289, w_227_290, w_227_296, w_227_298, w_227_302, w_227_304, w_227_306, w_227_309, w_227_313, w_227_314, w_227_323, w_227_326, w_227_332, w_227_339, w_227_340, w_227_342, w_227_344, w_227_348, w_227_349, w_227_356, w_227_358, w_227_361, w_227_363, w_227_365, w_227_367, w_227_369, w_227_370, w_227_373, w_227_376, w_227_381, w_227_391, w_227_392, w_227_393, w_227_394, w_227_395, w_227_396, w_227_399, w_227_401, w_227_409, w_227_411, w_227_417, w_227_421, w_227_422, w_227_423, w_227_427, w_227_431, w_227_434, w_227_435, w_227_442, w_227_443, w_227_453, w_227_456, w_227_464, w_227_471, w_227_474, w_227_477, w_227_481, w_227_484, w_227_488, w_227_491, w_227_501, w_227_502, w_227_504, w_227_511, w_227_521, w_227_530, w_227_532, w_227_537, w_227_538, w_227_549, w_227_551, w_227_555, w_227_557, w_227_560, w_227_562, w_227_564, w_227_565, w_227_571, w_227_573, w_227_574, w_227_576, w_227_588, w_227_589, w_227_595, w_227_599, w_227_603, w_227_605, w_227_608, w_227_617, w_227_623, w_227_627, w_227_633, w_227_635, w_227_636, w_227_638, w_227_640, w_227_641, w_227_649, w_227_651, w_227_654, w_227_655, w_227_656, w_227_660, w_227_661, w_227_662, w_227_664, w_227_665, w_227_666, w_227_677, w_227_682, w_227_683, w_227_684, w_227_689, w_227_695, w_227_696, w_227_697, w_227_698, w_227_699, w_227_702, w_227_704, w_227_705, w_227_707, w_227_710, w_227_717, w_227_718, w_227_719, w_227_722, w_227_726, w_227_728, w_227_730, w_227_732, w_227_737, w_227_738, w_227_749, w_227_750, w_227_752, w_227_760, w_227_763, w_227_764, w_227_766, w_227_768, w_227_770, w_227_776, w_227_781, w_227_791, w_227_792, w_227_795, w_227_796, w_227_797, w_227_798, w_227_803, w_227_808, w_227_812, w_227_813, w_227_819, w_227_826, w_227_833, w_227_834, w_227_837, w_227_839, w_227_841, w_227_842, w_227_848, w_227_853, w_227_861, w_227_866, w_227_868, w_227_873, w_227_876, w_227_882, w_227_883, w_227_894, w_227_897, w_227_900, w_227_902, w_227_903, w_227_906, w_227_914, w_227_915, w_227_916, w_227_926, w_227_935, w_227_936, w_227_938, w_227_940, w_227_941, w_227_950, w_227_951, w_227_952, w_227_956, w_227_958, w_227_961, w_227_963, w_227_967, w_227_970, w_227_976, w_227_977, w_227_981, w_227_983, w_227_994, w_227_997, w_227_999, w_227_1000, w_227_1005, w_227_1006, w_227_1008, w_227_1010, w_227_1015, w_227_1018, w_227_1019, w_227_1023, w_227_1027, w_227_1035, w_227_1037, w_227_1040, w_227_1041, w_227_1043, w_227_1044, w_227_1046, w_227_1051, w_227_1059, w_227_1061, w_227_1067, w_227_1070, w_227_1071, w_227_1079, w_227_1080, w_227_1081, w_227_1082, w_227_1084, w_227_1087, w_227_1089, w_227_1093, w_227_1094, w_227_1095, w_227_1098, w_227_1113, w_227_1114, w_227_1115, w_227_1116, w_227_1120, w_227_1122, w_227_1123, w_227_1125, w_227_1126, w_227_1134, w_227_1139, w_227_1145, w_227_1150, w_227_1153, w_227_1154, w_227_1155, w_227_1156, w_227_1158, w_227_1160, w_227_1163, w_227_1164, w_227_1165, w_227_1168, w_227_1174, w_227_1177, w_227_1178, w_227_1181, w_227_1187, w_227_1195, w_227_1198, w_227_1200, w_227_1203, w_227_1204, w_227_1208, w_227_1211, w_227_1213, w_227_1215, w_227_1221, w_227_1223, w_227_1232, w_227_1235, w_227_1241, w_227_1261, w_227_1279, w_227_1284, w_227_1289, w_227_1292, w_227_1297, w_227_1299, w_227_1300, w_227_1305, w_227_1306, w_227_1310, w_227_1311, w_227_1313, w_227_1316, w_227_1319, w_227_1337, w_227_1352, w_227_1353, w_227_1362, w_227_1365, w_227_1368, w_227_1383, w_227_1389, w_227_1394, w_227_1395, w_227_1398, w_227_1407, w_227_1410, w_227_1413, w_227_1423, w_227_1426, w_227_1427, w_227_1439, w_227_1447, w_227_1454, w_227_1457, w_227_1467, w_227_1476, w_227_1482, w_227_1484, w_227_1493, w_227_1494, w_227_1501, w_227_1517, w_227_1525, w_227_1526, w_227_1528, w_227_1529, w_227_1531, w_227_1546, w_227_1554, w_227_1556, w_227_1559, w_227_1561, w_227_1574, w_227_1576, w_227_1578, w_227_1584, w_227_1590, w_227_1591, w_227_1599, w_227_1600, w_227_1605, w_227_1608, w_227_1618, w_227_1620, w_227_1623, w_227_1624, w_227_1629, w_227_1630, w_227_1632, w_227_1643, w_227_1647, w_227_1648, w_227_1651, w_227_1656, w_227_1664, w_227_1665, w_227_1674, w_227_1675, w_227_1695, w_227_1698, w_227_1701, w_227_1702, w_227_1708, w_227_1710, w_227_1714, w_227_1718, w_227_1721, w_227_1730, w_227_1731, w_227_1732, w_227_1745, w_227_1749, w_227_1758, w_227_1760, w_227_1770, w_227_1777, w_227_1782, w_227_1784, w_227_1786, w_227_1798, w_227_1802, w_227_1805, w_227_1808, w_227_1810, w_227_1811, w_227_1815, w_227_1824, w_227_1828, w_227_1831, w_227_1843, w_227_1848, w_227_1851, w_227_1857, w_227_1859, w_227_1861, w_227_1862, w_227_1863, w_227_1864;
  wire w_228_001, w_228_003, w_228_005, w_228_007, w_228_008, w_228_010, w_228_013, w_228_015, w_228_018, w_228_019, w_228_021, w_228_023, w_228_031, w_228_034, w_228_040, w_228_042, w_228_044, w_228_047, w_228_049, w_228_051, w_228_057, w_228_058, w_228_060, w_228_063, w_228_065, w_228_067, w_228_068, w_228_074, w_228_080, w_228_081, w_228_084, w_228_086, w_228_088, w_228_090, w_228_091, w_228_092, w_228_093, w_228_094, w_228_095, w_228_098, w_228_107, w_228_108, w_228_109, w_228_111, w_228_112, w_228_113, w_228_114, w_228_116, w_228_117, w_228_120, w_228_122, w_228_124, w_228_131, w_228_133, w_228_134, w_228_135, w_228_136, w_228_137, w_228_140, w_228_142, w_228_146, w_228_147, w_228_148, w_228_149, w_228_151, w_228_153, w_228_154, w_228_157, w_228_159, w_228_160, w_228_161, w_228_163, w_228_169, w_228_171, w_228_175, w_228_177, w_228_178, w_228_180, w_228_181, w_228_182, w_228_184, w_228_185, w_228_189, w_228_190, w_228_195, w_228_197, w_228_198, w_228_199, w_228_200, w_228_202, w_228_203, w_228_205, w_228_206, w_228_209, w_228_210, w_228_211, w_228_213, w_228_214, w_228_215, w_228_216, w_228_217, w_228_225, w_228_228, w_228_231, w_228_232, w_228_235, w_228_238, w_228_240, w_228_243, w_228_244, w_228_246, w_228_250, w_228_253, w_228_254, w_228_255, w_228_256, w_228_257, w_228_259, w_228_263, w_228_264, w_228_265, w_228_266, w_228_269, w_228_273, w_228_275, w_228_276, w_228_281, w_228_283, w_228_284, w_228_286, w_228_288, w_228_289, w_228_290, w_228_291, w_228_293, w_228_302, w_228_305, w_228_308, w_228_309, w_228_311, w_228_316, w_228_317, w_228_324, w_228_329, w_228_330, w_228_338, w_228_339, w_228_340, w_228_341, w_228_346, w_228_349, w_228_350, w_228_351, w_228_352, w_228_353, w_228_355, w_228_357, w_228_358, w_228_359, w_228_364, w_228_365, w_228_370, w_228_382, w_228_386, w_228_387, w_228_388, w_228_391, w_228_395, w_228_396, w_228_397, w_228_398, w_228_400, w_228_401, w_228_402, w_228_403, w_228_405, w_228_416, w_228_419, w_228_420, w_228_423, w_228_426, w_228_435, w_228_436, w_228_439, w_228_440, w_228_442, w_228_443, w_228_445, w_228_446, w_228_448, w_228_450, w_228_452, w_228_455, w_228_457, w_228_458, w_228_460, w_228_461, w_228_463, w_228_468, w_228_471, w_228_472, w_228_475, w_228_476, w_228_480, w_228_481, w_228_484, w_228_487, w_228_494, w_228_498, w_228_501, w_228_507, w_228_508, w_228_511, w_228_513, w_228_515, w_228_521, w_228_526, w_228_529, w_228_533, w_228_540, w_228_543, w_228_544, w_228_545, w_228_546, w_228_552, w_228_553, w_228_555, w_228_559, w_228_561, w_228_563, w_228_568, w_228_569, w_228_574, w_228_577, w_228_578, w_228_579, w_228_584, w_228_588, w_228_590, w_228_591, w_228_592, w_228_593, w_228_594, w_228_595, w_228_598, w_228_606, w_228_610, w_228_616, w_228_624, w_228_626, w_228_628, w_228_631, w_228_637, w_228_638, w_228_640, w_228_642, w_228_644, w_228_647, w_228_648, w_228_653, w_228_654, w_228_655, w_228_657, w_228_658, w_228_659, w_228_660, w_228_661, w_228_665, w_228_668, w_228_669, w_228_670, w_228_672, w_228_677, w_228_680, w_228_685, w_228_686, w_228_690, w_228_695, w_228_698, w_228_699, w_228_701, w_228_703, w_228_705, w_228_710, w_228_711, w_228_712, w_228_713, w_228_715, w_228_717, w_228_718, w_228_723, w_228_727, w_228_729, w_228_735, w_228_739, w_228_746, w_228_748, w_228_749, w_228_752, w_228_754, w_228_760, w_228_765, w_228_772, w_228_776, w_228_777, w_228_779, w_228_780, w_228_781, w_228_782, w_228_786, w_228_797, w_228_798, w_228_800, w_228_805, w_228_806, w_228_810, w_228_811, w_228_816, w_228_818, w_228_822, w_228_823, w_228_830, w_228_832, w_228_841, w_228_842, w_228_845, w_228_846, w_228_849, w_228_850, w_228_851, w_228_855, w_228_856, w_228_865, w_228_869, w_228_870, w_228_873, w_228_875, w_228_876, w_228_877, w_228_878, w_228_880, w_228_882, w_228_888, w_228_892, w_228_896, w_228_897, w_228_899, w_228_901, w_228_904, w_228_905, w_228_913, w_228_916, w_228_917, w_228_918, w_228_919, w_228_923, w_228_929, w_228_930, w_228_934, w_228_939, w_228_948, w_228_950, w_228_952, w_228_953, w_228_956, w_228_957, w_228_959, w_228_960, w_228_963, w_228_964, w_228_971, w_228_976, w_228_981, w_228_986, w_228_987, w_228_992, w_228_993, w_228_994, w_228_995, w_228_997, w_228_998, w_228_1005, w_228_1007, w_228_1010, w_228_1014, w_228_1020, w_228_1022, w_228_1023, w_228_1024, w_228_1033, w_228_1034, w_228_1035, w_228_1036, w_228_1039, w_228_1040, w_228_1041, w_228_1042, w_228_1048, w_228_1052, w_228_1054, w_228_1055, w_228_1056, w_228_1057, w_228_1059, w_228_1060, w_228_1061, w_228_1063, w_228_1066, w_228_1069, w_228_1075, w_228_1076, w_228_1078, w_228_1081, w_228_1084, w_228_1085, w_228_1093, w_228_1096, w_228_1099, w_228_1104, w_228_1107, w_228_1109, w_228_1115, w_228_1118, w_228_1119, w_228_1123, w_228_1127, w_228_1129, w_228_1131, w_228_1137, w_228_1138, w_228_1139;
  wire w_229_010, w_229_017, w_229_026, w_229_042, w_229_052, w_229_061, w_229_062, w_229_065, w_229_067, w_229_069, w_229_079, w_229_082, w_229_101, w_229_106, w_229_109, w_229_112, w_229_116, w_229_120, w_229_123, w_229_126, w_229_131, w_229_137, w_229_138, w_229_140, w_229_143, w_229_150, w_229_153, w_229_167, w_229_180, w_229_183, w_229_188, w_229_191, w_229_200, w_229_204, w_229_205, w_229_207, w_229_218, w_229_233, w_229_237, w_229_241, w_229_243, w_229_253, w_229_255, w_229_260, w_229_263, w_229_268, w_229_276, w_229_278, w_229_280, w_229_288, w_229_291, w_229_294, w_229_297, w_229_298, w_229_306, w_229_308, w_229_309, w_229_312, w_229_313, w_229_314, w_229_317, w_229_323, w_229_324, w_229_330, w_229_333, w_229_339, w_229_340, w_229_348, w_229_351, w_229_352, w_229_368, w_229_370, w_229_373, w_229_376, w_229_379, w_229_384, w_229_391, w_229_394, w_229_401, w_229_405, w_229_414, w_229_424, w_229_433, w_229_437, w_229_441, w_229_442, w_229_446, w_229_448, w_229_449, w_229_453, w_229_456, w_229_458, w_229_462, w_229_465, w_229_482, w_229_500, w_229_501, w_229_502, w_229_508, w_229_510, w_229_513, w_229_516, w_229_528, w_229_551, w_229_552, w_229_553, w_229_556, w_229_562, w_229_569, w_229_572, w_229_573, w_229_578, w_229_585, w_229_594, w_229_597, w_229_598, w_229_599, w_229_603, w_229_609, w_229_611, w_229_612, w_229_618, w_229_621, w_229_625, w_229_630, w_229_633, w_229_639, w_229_643, w_229_647, w_229_648, w_229_649, w_229_655, w_229_656, w_229_669, w_229_670, w_229_671, w_229_672, w_229_675, w_229_686, w_229_689, w_229_695, w_229_699, w_229_700, w_229_702, w_229_708, w_229_714, w_229_717, w_229_731, w_229_736, w_229_738, w_229_740, w_229_743, w_229_744, w_229_750, w_229_753, w_229_756, w_229_757, w_229_761, w_229_765, w_229_783, w_229_787, w_229_796, w_229_798, w_229_800, w_229_808, w_229_809, w_229_810, w_229_831, w_229_832, w_229_834, w_229_840, w_229_841, w_229_842, w_229_848, w_229_853, w_229_857, w_229_860, w_229_871, w_229_872, w_229_874, w_229_879, w_229_881, w_229_882, w_229_883, w_229_885, w_229_900, w_229_903, w_229_905, w_229_915, w_229_926, w_229_927, w_229_933, w_229_942, w_229_948, w_229_956, w_229_970, w_229_973, w_229_979, w_229_981, w_229_992, w_229_998, w_229_1001, w_229_1010, w_229_1015, w_229_1024, w_229_1026, w_229_1030, w_229_1037, w_229_1051, w_229_1059, w_229_1063, w_229_1073, w_229_1075, w_229_1082, w_229_1086, w_229_1096, w_229_1098, w_229_1102, w_229_1108, w_229_1112, w_229_1113, w_229_1120, w_229_1123, w_229_1128, w_229_1141, w_229_1158, w_229_1162, w_229_1164, w_229_1165, w_229_1170, w_229_1194, w_229_1195, w_229_1208, w_229_1213, w_229_1214, w_229_1215, w_229_1216, w_229_1219, w_229_1222, w_229_1228, w_229_1230, w_229_1238, w_229_1249, w_229_1252, w_229_1253, w_229_1256, w_229_1257, w_229_1285, w_229_1306, w_229_1308, w_229_1316, w_229_1347, w_229_1373, w_229_1379, w_229_1380, w_229_1381, w_229_1383, w_229_1391, w_229_1406, w_229_1412, w_229_1422, w_229_1426, w_229_1437, w_229_1438, w_229_1463, w_229_1481, w_229_1483, w_229_1492, w_229_1501, w_229_1504, w_229_1508, w_229_1509, w_229_1524, w_229_1525, w_229_1527, w_229_1530, w_229_1531, w_229_1561, w_229_1578, w_229_1586, w_229_1591, w_229_1602, w_229_1603, w_229_1607, w_229_1611, w_229_1620, w_229_1628, w_229_1641, w_229_1646, w_229_1658, w_229_1690, w_229_1702, w_229_1720, w_229_1727, w_229_1730, w_229_1735, w_229_1736, w_229_1741, w_229_1753, w_229_1756, w_229_1770, w_229_1791, w_229_1798, w_229_1803, w_229_1827, w_229_1828, w_229_1860, w_229_1862, w_229_1869, w_229_1875, w_229_1884, w_229_1887, w_229_1892, w_229_1898, w_229_1917, w_229_1928, w_229_1932, w_229_1935, w_229_1958, w_229_1959, w_229_1963, w_229_1976, w_229_1980, w_229_1986, w_229_2004, w_229_2014, w_229_2033, w_229_2049, w_229_2089, w_229_2093, w_229_2099, w_229_2107, w_229_2116, w_229_2117, w_229_2126, w_229_2147, w_229_2156, w_229_2183, w_229_2200, w_229_2223, w_229_2278, w_229_2283, w_229_2285, w_229_2286, w_229_2288, w_229_2290, w_229_2295, w_229_2315, w_229_2316, w_229_2330, w_229_2333, w_229_2343, w_229_2350, w_229_2365, w_229_2366, w_229_2373, w_229_2385, w_229_2387, w_229_2390, w_229_2396, w_229_2398, w_229_2420, w_229_2431, w_229_2479, w_229_2483, w_229_2508, w_229_2530, w_229_2548, w_229_2550, w_229_2558, w_229_2563, w_229_2573, w_229_2575, w_229_2583, w_229_2584, w_229_2586, w_229_2598, w_229_2651, w_229_2652, w_229_2653, w_229_2664, w_229_2678, w_229_2683, w_229_2704, w_229_2722, w_229_2723, w_229_2741, w_229_2763, w_229_2766, w_229_2783, w_229_2793, w_229_2795, w_229_2799, w_229_2804, w_229_2820, w_229_2825, w_229_2833, w_229_2834, w_229_2838, w_229_2840, w_229_2848, w_229_2862, w_229_2863, w_229_2877, w_229_2890, w_229_2904, w_229_2917, w_229_2924, w_229_2942, w_229_2949, w_229_2953, w_229_2954, w_229_2967, w_229_2969, w_229_2977, w_229_2983, w_229_2987, w_229_3000, w_229_3032, w_229_3037, w_229_3050, w_229_3051, w_229_3054, w_229_3058, w_229_3063, w_229_3083, w_229_3086, w_229_3090, w_229_3104, w_229_3113, w_229_3114, w_229_3132, w_229_3137, w_229_3144, w_229_3159, w_229_3166, w_229_3178, w_229_3196, w_229_3198, w_229_3212, w_229_3217, w_229_3220, w_229_3230, w_229_3239, w_229_3242, w_229_3253, w_229_3255, w_229_3264, w_229_3265, w_229_3269, w_229_3276, w_229_3293, w_229_3302, w_229_3312, w_229_3316, w_229_3349, w_229_3350, w_229_3353, w_229_3354, w_229_3370, w_229_3373, w_229_3376, w_229_3380, w_229_3381, w_229_3419, w_229_3421, w_229_3425, w_229_3435, w_229_3441, w_229_3454, w_229_3459, w_229_3460, w_229_3462, w_229_3492, w_229_3496, w_229_3498, w_229_3500, w_229_3505, w_229_3513, w_229_3523, w_229_3527, w_229_3531, w_229_3536, w_229_3563, w_229_3571, w_229_3573, w_229_3593, w_229_3599, w_229_3600, w_229_3606, w_229_3609, w_229_3613, w_229_3620, w_229_3636, w_229_3649, w_229_3659, w_229_3696, w_229_3698, w_229_3725, w_229_3730, w_229_3736, w_229_3813, w_229_3818, w_229_3827, w_229_3830, w_229_3847, w_229_3851, w_229_3855, w_229_3858, w_229_3860, w_229_3861;
  wire w_230_013, w_230_015, w_230_016, w_230_022, w_230_028, w_230_031, w_230_036, w_230_043, w_230_050, w_230_051, w_230_054, w_230_058, w_230_059, w_230_060, w_230_064, w_230_065, w_230_068, w_230_070, w_230_072, w_230_098, w_230_103, w_230_105, w_230_107, w_230_111, w_230_113, w_230_116, w_230_124, w_230_128, w_230_134, w_230_138, w_230_139, w_230_144, w_230_145, w_230_146, w_230_147, w_230_148, w_230_158, w_230_160, w_230_161, w_230_162, w_230_178, w_230_195, w_230_196, w_230_197, w_230_199, w_230_207, w_230_208, w_230_210, w_230_220, w_230_224, w_230_228, w_230_230, w_230_233, w_230_244, w_230_252, w_230_255, w_230_258, w_230_260, w_230_263, w_230_266, w_230_267, w_230_272, w_230_276, w_230_277, w_230_279, w_230_280, w_230_291, w_230_294, w_230_295, w_230_296, w_230_302, w_230_304, w_230_312, w_230_317, w_230_319, w_230_321, w_230_327, w_230_332, w_230_338, w_230_345, w_230_346, w_230_352, w_230_357, w_230_360, w_230_362, w_230_372, w_230_379, w_230_381, w_230_385, w_230_388, w_230_392, w_230_396, w_230_400, w_230_403, w_230_414, w_230_424, w_230_427, w_230_430, w_230_433, w_230_436, w_230_439, w_230_446, w_230_455, w_230_463, w_230_466, w_230_467, w_230_475, w_230_488, w_230_496, w_230_504, w_230_505, w_230_510, w_230_512, w_230_519, w_230_524, w_230_535, w_230_558, w_230_571, w_230_576, w_230_581, w_230_584, w_230_587, w_230_594, w_230_597, w_230_605, w_230_609, w_230_613, w_230_624, w_230_627, w_230_633, w_230_634, w_230_635, w_230_638, w_230_639, w_230_646, w_230_647, w_230_648, w_230_650, w_230_653, w_230_660, w_230_672, w_230_675, w_230_678, w_230_680, w_230_682, w_230_703, w_230_704, w_230_705, w_230_706, w_230_715, w_230_721, w_230_722, w_230_727, w_230_743, w_230_749, w_230_760, w_230_768, w_230_778, w_230_780, w_230_785, w_230_795, w_230_827, w_230_844, w_230_845, w_230_853, w_230_857, w_230_862, w_230_875, w_230_884, w_230_893, w_230_905, w_230_919, w_230_920, w_230_931, w_230_939, w_230_943, w_230_950, w_230_957, w_230_962, w_230_976, w_230_995, w_230_1011, w_230_1022, w_230_1026, w_230_1032, w_230_1039, w_230_1049, w_230_1055, w_230_1058, w_230_1070, w_230_1071, w_230_1094, w_230_1100, w_230_1119, w_230_1134, w_230_1136, w_230_1140, w_230_1141, w_230_1147, w_230_1152, w_230_1166, w_230_1173, w_230_1180, w_230_1191, w_230_1203, w_230_1204, w_230_1205, w_230_1214, w_230_1215, w_230_1219, w_230_1232, w_230_1234, w_230_1255, w_230_1283, w_230_1295, w_230_1302, w_230_1310, w_230_1327, w_230_1329, w_230_1351, w_230_1356, w_230_1364, w_230_1367, w_230_1379, w_230_1385, w_230_1389, w_230_1407, w_230_1416, w_230_1431, w_230_1438, w_230_1442, w_230_1446, w_230_1460, w_230_1465, w_230_1470, w_230_1483, w_230_1485, w_230_1492, w_230_1494, w_230_1497, w_230_1499, w_230_1520, w_230_1530, w_230_1532, w_230_1543, w_230_1552, w_230_1571, w_230_1574, w_230_1580, w_230_1594, w_230_1597, w_230_1623, w_230_1648, w_230_1653, w_230_1658, w_230_1661, w_230_1663, w_230_1681, w_230_1683, w_230_1691, w_230_1701, w_230_1704, w_230_1705, w_230_1708, w_230_1728, w_230_1735, w_230_1741, w_230_1750, w_230_1757, w_230_1759, w_230_1760, w_230_1763, w_230_1765, w_230_1767, w_230_1776, w_230_1778, w_230_1789, w_230_1819, w_230_1835, w_230_1847, w_230_1849, w_230_1854, w_230_1856, w_230_1876, w_230_1877, w_230_1884, w_230_1889, w_230_1898, w_230_1910, w_230_1948, w_230_1966, w_230_1976, w_230_1989, w_230_2015, w_230_2020, w_230_2038, w_230_2070, w_230_2071, w_230_2074, w_230_2091, w_230_2092, w_230_2099, w_230_2102, w_230_2109, w_230_2122, w_230_2182, w_230_2184, w_230_2191, w_230_2193, w_230_2198, w_230_2199, w_230_2202, w_230_2211, w_230_2240, w_230_2253, w_230_2266, w_230_2290, w_230_2301, w_230_2316, w_230_2321, w_230_2327, w_230_2336, w_230_2337, w_230_2367, w_230_2368, w_230_2385, w_230_2389, w_230_2399, w_230_2406, w_230_2407, w_230_2408, w_230_2411, w_230_2413, w_230_2438, w_230_2458, w_230_2479, w_230_2500, w_230_2513, w_230_2514, w_230_2550, w_230_2553, w_230_2564, w_230_2565, w_230_2568, w_230_2572, w_230_2576, w_230_2586, w_230_2597, w_230_2605, w_230_2608, w_230_2610, w_230_2611, w_230_2619, w_230_2623, w_230_2631, w_230_2638, w_230_2644, w_230_2653, w_230_2673, w_230_2684, w_230_2692, w_230_2699, w_230_2707, w_230_2710, w_230_2714, w_230_2727, w_230_2728, w_230_2740, w_230_2742, w_230_2746, w_230_2773, w_230_2778, w_230_2786, w_230_2799, w_230_2808, w_230_2816, w_230_2817, w_230_2824, w_230_2829, w_230_2838, w_230_2848, w_230_2877, w_230_2878, w_230_2885, w_230_2897, w_230_2902, w_230_2903, w_230_2904, w_230_2907, w_230_2922, w_230_2933, w_230_2946, w_230_2949, w_230_2956, w_230_2957, w_230_2961, w_230_2968, w_230_2971, w_230_3000, w_230_3009, w_230_3020, w_230_3026, w_230_3028, w_230_3034, w_230_3036, w_230_3040, w_230_3041, w_230_3056, w_230_3061, w_230_3074, w_230_3078, w_230_3080, w_230_3100, w_230_3116, w_230_3121, w_230_3126, w_230_3133, w_230_3167, w_230_3169, w_230_3186, w_230_3206, w_230_3210, w_230_3214, w_230_3217, w_230_3218, w_230_3224, w_230_3232, w_230_3239, w_230_3248, w_230_3251, w_230_3254, w_230_3265, w_230_3268, w_230_3271, w_230_3276, w_230_3281, w_230_3298, w_230_3307, w_230_3309, w_230_3316, w_230_3346, w_230_3352, w_230_3354, w_230_3360, w_230_3368, w_230_3372, w_230_3379, w_230_3393, w_230_3412, w_230_3438, w_230_3447, w_230_3452, w_230_3459, w_230_3461, w_230_3462, w_230_3469, w_230_3485, w_230_3489, w_230_3490, w_230_3496, w_230_3497, w_230_3500, w_230_3503, w_230_3528, w_230_3533, w_230_3542, w_230_3544, w_230_3545, w_230_3572, w_230_3592, w_230_3594, w_230_3613, w_230_3615, w_230_3620, w_230_3651, w_230_3663, w_230_3665, w_230_3674, w_230_3693, w_230_3698, w_230_3701, w_230_3718, w_230_3720, w_230_3730, w_230_3737, w_230_3756, w_230_3770, w_230_3784, w_230_3785, w_230_3793, w_230_3811, w_230_3832, w_230_3858, w_230_3862, w_230_3867, w_230_3909, w_230_3914, w_230_3916, w_230_3937, w_230_3946, w_230_3947, w_230_3949, w_230_3951, w_230_3954, w_230_3956, w_230_3960, w_230_3963, w_230_3968, w_230_3969, w_230_3976, w_230_3988, w_230_4011, w_230_4012, w_230_4023, w_230_4029, w_230_4037, w_230_4049, w_230_4052, w_230_4058, w_230_4060, w_230_4067, w_230_4070, w_230_4075, w_230_4085, w_230_4087, w_230_4093, w_230_4103, w_230_4118, w_230_4130, w_230_4160, w_230_4176, w_230_4177, w_230_4188, w_230_4194, w_230_4216, w_230_4223, w_230_4228, w_230_4239, w_230_4243, w_230_4252, w_230_4261, w_230_4271, w_230_4272, w_230_4273, w_230_4274, w_230_4275, w_230_4277, w_230_4279, w_230_4280, w_230_4281, w_230_4282, w_230_4283, w_230_4284, w_230_4285, w_230_4286, w_230_4288, w_230_4290, w_230_4291, w_230_4292, w_230_4293, w_230_4295, w_230_4297, w_230_4298, w_230_4299, w_230_4300, w_230_4301, w_230_4302, w_230_4303, w_230_4304, w_230_4306;
  wire w_231_009, w_231_010, w_231_022, w_231_024, w_231_029, w_231_034, w_231_035, w_231_036, w_231_040, w_231_044, w_231_045, w_231_050, w_231_052, w_231_055, w_231_056, w_231_063, w_231_065, w_231_070, w_231_073, w_231_077, w_231_078, w_231_081, w_231_083, w_231_088, w_231_090, w_231_091, w_231_095, w_231_098, w_231_110, w_231_113, w_231_114, w_231_124, w_231_127, w_231_130, w_231_133, w_231_140, w_231_141, w_231_143, w_231_154, w_231_156, w_231_160, w_231_162, w_231_165, w_231_177, w_231_188, w_231_189, w_231_190, w_231_197, w_231_198, w_231_199, w_231_211, w_231_217, w_231_221, w_231_224, w_231_227, w_231_239, w_231_242, w_231_244, w_231_245, w_231_248, w_231_249, w_231_253, w_231_254, w_231_261, w_231_262, w_231_268, w_231_272, w_231_278, w_231_294, w_231_299, w_231_300, w_231_309, w_231_310, w_231_313, w_231_320, w_231_321, w_231_322, w_231_323, w_231_330, w_231_332, w_231_338, w_231_342, w_231_346, w_231_350, w_231_352, w_231_353, w_231_354, w_231_355, w_231_356, w_231_358, w_231_360, w_231_373, w_231_383, w_231_384, w_231_391, w_231_397, w_231_400, w_231_405, w_231_414, w_231_416, w_231_420, w_231_422, w_231_424, w_231_425, w_231_432, w_231_433, w_231_435, w_231_437, w_231_449, w_231_466, w_231_467, w_231_483, w_231_486, w_231_487, w_231_489, w_231_492, w_231_508, w_231_511, w_231_512, w_231_516, w_231_525, w_231_530, w_231_533, w_231_536, w_231_539, w_231_542, w_231_563, w_231_574, w_231_576, w_231_583, w_231_584, w_231_585, w_231_586, w_231_591, w_231_592, w_231_605, w_231_606, w_231_609, w_231_628, w_231_632, w_231_635, w_231_643, w_231_646, w_231_650, w_231_651, w_231_657, w_231_664, w_231_665, w_231_669, w_231_675, w_231_676, w_231_677, w_231_682, w_231_688, w_231_689, w_231_690, w_231_691, w_231_697, w_231_698, w_231_702, w_231_705, w_231_718, w_231_720, w_231_730, w_231_741, w_231_747, w_231_752, w_231_755, w_231_762, w_231_765, w_231_766, w_231_780, w_231_788, w_231_792, w_231_793, w_231_794, w_231_797, w_231_801, w_231_806, w_231_821, w_231_825, w_231_826, w_231_830, w_231_836, w_231_840, w_231_841, w_231_848, w_231_857, w_231_858, w_231_862, w_231_865, w_231_868, w_231_870, w_231_871, w_231_875, w_231_883, w_231_887, w_231_891, w_231_895, w_231_899, w_231_903, w_231_910, w_231_929, w_231_932, w_231_933, w_231_950, w_231_953, w_231_954, w_231_956, w_231_967, w_231_972, w_231_974, w_231_975, w_231_976, w_231_979, w_231_986, w_231_987, w_231_999, w_231_1000, w_231_1013, w_231_1021, w_231_1023, w_231_1025, w_231_1026, w_231_1027, w_231_1030, w_231_1040, w_231_1042, w_231_1045, w_231_1046, w_231_1064, w_231_1072, w_231_1086, w_231_1090, w_231_1093, w_231_1097, w_231_1101, w_231_1104, w_231_1107, w_231_1108, w_231_1117, w_231_1125, w_231_1131, w_231_1139, w_231_1142, w_231_1157, w_231_1159, w_231_1163, w_231_1167, w_231_1176, w_231_1181, w_231_1188, w_231_1195, w_231_1200, w_231_1208, w_231_1212, w_231_1219, w_231_1223, w_231_1224, w_231_1234, w_231_1238, w_231_1241, w_231_1243, w_231_1244, w_231_1251, w_231_1258, w_231_1263, w_231_1275, w_231_1286, w_231_1288, w_231_1291, w_231_1295, w_231_1298, w_231_1307, w_231_1312, w_231_1319, w_231_1320, w_231_1326, w_231_1331, w_231_1332, w_231_1334, w_231_1338, w_231_1346, w_231_1347, w_231_1348, w_231_1354, w_231_1357, w_231_1358, w_231_1361, w_231_1370, w_231_1371, w_231_1373, w_231_1376, w_231_1377, w_231_1392, w_231_1395, w_231_1397, w_231_1403, w_231_1405, w_231_1406, w_231_1409, w_231_1414, w_231_1421, w_231_1422, w_231_1423, w_231_1428, w_231_1432, w_231_1436, w_231_1442, w_231_1446, w_231_1451, w_231_1459, w_231_1460, w_231_1464, w_231_1470, w_231_1472, w_231_1473, w_231_1475, w_231_1478, w_231_1482, w_231_1484, w_231_1486, w_231_1487, w_231_1489, w_231_1492, w_231_1497, w_231_1500, w_231_1504, w_231_1516, w_231_1532, w_231_1537, w_231_1544, w_231_1546, w_231_1554, w_231_1558, w_231_1561, w_231_1573, w_231_1580, w_231_1588, w_231_1590, w_231_1591, w_231_1603, w_231_1615, w_231_1616, w_231_1618, w_231_1622, w_231_1626, w_231_1633, w_231_1639, w_231_1640, w_231_1645, w_231_1647, w_231_1662, w_231_1671, w_231_1675, w_231_1682, w_231_1690, w_231_1701, w_231_1708, w_231_1712, w_231_1714, w_231_1719, w_231_1726, w_231_1732, w_231_1740, w_231_1757, w_231_1758, w_231_1764, w_231_1766, w_231_1767, w_231_1778, w_231_1779, w_231_1789, w_231_1790, w_231_1794, w_231_1798, w_231_1800, w_231_1803, w_231_1806, w_231_1809, w_231_1811, w_231_1826, w_231_1828, w_231_1833, w_231_1834, w_231_1839, w_231_1841, w_231_1844, w_231_1849, w_231_1852, w_231_1853, w_231_1860, w_231_1864, w_231_1866, w_231_1873, w_231_1877, w_231_1900, w_231_1917, w_231_1919, w_231_1920, w_231_1922, w_231_1924, w_231_1931, w_231_1933, w_231_1938, w_231_1941, w_231_1949, w_231_1952, w_231_1954, w_231_1955, w_231_1957, w_231_1959, w_231_1960, w_231_1972, w_231_1973, w_231_1975, w_231_1980, w_231_1986, w_231_1995, w_231_1998, w_231_1999, w_231_2000, w_231_2006, w_231_2019, w_231_2024, w_231_2044, w_231_2051, w_231_2056, w_231_2058, w_231_2062, w_231_2064, w_231_2065, w_231_2068, w_231_2072, w_231_2074, w_231_2075, w_231_2081, w_231_2092, w_231_2093, w_231_2106, w_231_2109, w_231_2110, w_231_2112, w_231_2132, w_231_2135, w_231_2138, w_231_2140, w_231_2141, w_231_2152, w_231_2159, w_231_2175, w_231_2177, w_231_2178, w_231_2199, w_231_2201, w_231_2203, w_231_2206, w_231_2207, w_231_2212, w_231_2218, w_231_2223, w_231_2230, w_231_2231, w_231_2233, w_231_2239, w_231_2246, w_231_2253, w_231_2257, w_231_2268, w_231_2273, w_231_2274, w_231_2276, w_231_2283, w_231_2284, w_231_2287, w_231_2298, w_231_2299, w_231_2300, w_231_2304, w_231_2305, w_231_2313, w_231_2317, w_231_2321, w_231_2323, w_231_2328, w_231_2333, w_231_2348, w_231_2349, w_231_2362, w_231_2373, w_231_2376, w_231_2381, w_231_2382, w_231_2386, w_231_2393, w_231_2438, w_231_2461, w_231_2471, w_231_2474, w_231_2481, w_231_2486, w_231_2497, w_231_2502, w_231_2504, w_231_2505, w_231_2518, w_231_2536, w_231_2540, w_231_2556, w_231_2565, w_231_2601, w_231_2610, w_231_2613, w_231_2629, w_231_2640, w_231_2641, w_231_2642, w_231_2658;
  wire w_232_002, w_232_004, w_232_010, w_232_011, w_232_013, w_232_023, w_232_026, w_232_032, w_232_039, w_232_042, w_232_050, w_232_052, w_232_054, w_232_057, w_232_067, w_232_072, w_232_082, w_232_094, w_232_095, w_232_100, w_232_109, w_232_117, w_232_124, w_232_125, w_232_127, w_232_130, w_232_133, w_232_134, w_232_135, w_232_138, w_232_143, w_232_147, w_232_149, w_232_151, w_232_153, w_232_154, w_232_157, w_232_158, w_232_159, w_232_161, w_232_167, w_232_178, w_232_179, w_232_181, w_232_188, w_232_197, w_232_201, w_232_202, w_232_205, w_232_208, w_232_211, w_232_214, w_232_215, w_232_216, w_232_219, w_232_225, w_232_229, w_232_231, w_232_236, w_232_238, w_232_240, w_232_249, w_232_254, w_232_262, w_232_265, w_232_273, w_232_282, w_232_283, w_232_284, w_232_285, w_232_291, w_232_292, w_232_296, w_232_303, w_232_310, w_232_311, w_232_315, w_232_320, w_232_322, w_232_326, w_232_328, w_232_330, w_232_331, w_232_335, w_232_336, w_232_339, w_232_340, w_232_341, w_232_343, w_232_344, w_232_346, w_232_349, w_232_354, w_232_355, w_232_361, w_232_362, w_232_366, w_232_370, w_232_371, w_232_379, w_232_386, w_232_390, w_232_391, w_232_392, w_232_395, w_232_399, w_232_402, w_232_403, w_232_405, w_232_409, w_232_417, w_232_419, w_232_420, w_232_427, w_232_429, w_232_431, w_232_433, w_232_434, w_232_436, w_232_438, w_232_439, w_232_440, w_232_442, w_232_443, w_232_444, w_232_447, w_232_449, w_232_455, w_232_460, w_232_461, w_232_463, w_232_465, w_232_468, w_232_472, w_232_480, w_232_482, w_232_483, w_232_484, w_232_486, w_232_487, w_232_488, w_232_489, w_232_490, w_232_491, w_232_494, w_232_497, w_232_502, w_232_504, w_232_508, w_232_510, w_232_516, w_232_518, w_232_525, w_232_529, w_232_531, w_232_532, w_232_534, w_232_535, w_232_542, w_232_544, w_232_550, w_232_552, w_232_556, w_232_557, w_232_560, w_232_562, w_232_563, w_232_564, w_232_565, w_232_566, w_232_567, w_232_569, w_232_570, w_232_573, w_232_576, w_232_577, w_232_579, w_232_580, w_232_582, w_232_584, w_232_590, w_232_592, w_232_595, w_232_603, w_232_604, w_232_610, w_232_616, w_232_620, w_232_621, w_232_627, w_232_632, w_232_641, w_232_642, w_232_651, w_232_655, w_232_658, w_232_664, w_232_668, w_232_670, w_232_671, w_232_673, w_232_674, w_232_676, w_232_684, w_232_688, w_232_690, w_232_700, w_232_701, w_232_712, w_232_713, w_232_714, w_232_716, w_232_724, w_232_730, w_232_738, w_232_739, w_232_741, w_232_744, w_232_746, w_232_747, w_232_750, w_232_751, w_232_754, w_232_756, w_232_757, w_232_761, w_232_767, w_232_769, w_232_770, w_232_771, w_232_772, w_232_773, w_232_774, w_232_775, w_232_789, w_232_792, w_232_793, w_232_802, w_232_807, w_232_808, w_232_809, w_232_812, w_232_820, w_232_821, w_232_822, w_232_832, w_232_833, w_232_834, w_232_846, w_232_850, w_232_852, w_232_853, w_232_857, w_232_859, w_232_860, w_232_877, w_232_891, w_232_898, w_232_901, w_232_903, w_232_917, w_232_920, w_232_924, w_232_925, w_232_926, w_232_932, w_232_934, w_232_937, w_232_939, w_232_955, w_232_957, w_232_958, w_232_959, w_232_966, w_232_972, w_232_973, w_232_983, w_232_990, w_232_994, w_232_997, w_232_998, w_232_1002, w_232_1003, w_232_1004, w_232_1006, w_232_1020, w_232_1022, w_232_1029, w_232_1032, w_232_1038, w_232_1043, w_232_1046, w_232_1054, w_232_1058, w_232_1059, w_232_1060, w_232_1063, w_232_1074, w_232_1077, w_232_1078, w_232_1088, w_232_1092, w_232_1094, w_232_1103, w_232_1106, w_232_1114, w_232_1116, w_232_1119, w_232_1125, w_232_1131, w_232_1135, w_232_1136, w_232_1139, w_232_1140, w_232_1144, w_232_1145, w_232_1146, w_232_1161, w_232_1165, w_232_1178, w_232_1180, w_232_1188, w_232_1189, w_232_1192, w_232_1194, w_232_1195, w_232_1197, w_232_1201, w_232_1203, w_232_1210, w_232_1225, w_232_1233, w_232_1238, w_232_1244, w_232_1250, w_232_1256, w_232_1257, w_232_1259, w_232_1261, w_232_1262, w_232_1263, w_232_1266, w_232_1267, w_232_1275, w_232_1282, w_232_1292, w_232_1296, w_232_1299, w_232_1303, w_232_1304, w_232_1314, w_232_1315, w_232_1325, w_232_1332, w_232_1334, w_232_1346, w_232_1353, w_232_1354, w_232_1360, w_232_1361, w_232_1373, w_232_1374, w_232_1391, w_232_1406, w_232_1411, w_232_1412, w_232_1423, w_232_1429, w_232_1433, w_232_1437, w_232_1442, w_232_1450, w_232_1454, w_232_1460, w_232_1462, w_232_1463, w_232_1468, w_232_1475, w_232_1483, w_232_1484, w_232_1490, w_232_1497, w_232_1503, w_232_1515, w_232_1521, w_232_1525, w_232_1526, w_232_1527, w_232_1528, w_232_1530, w_232_1544, w_232_1550, w_232_1565, w_232_1569, w_232_1570, w_232_1573, w_232_1577, w_232_1582, w_232_1594, w_232_1600, w_232_1602, w_232_1603, w_232_1605, w_232_1606, w_232_1607, w_232_1625, w_232_1631, w_232_1635, w_232_1637, w_232_1639, w_232_1644, w_232_1645, w_232_1653, w_232_1654, w_232_1668, w_232_1689, w_232_1691, w_232_1692, w_232_1718, w_232_1719, w_232_1723, w_232_1739, w_232_1741, w_232_1746, w_232_1748, w_232_1749, w_232_1759, w_232_1762, w_232_1764, w_232_1767, w_232_1769, w_232_1782, w_232_1790, w_232_1798, w_232_1800, w_232_1802, w_232_1803, w_232_1806, w_232_1809, w_232_1811, w_232_1827, w_232_1832, w_232_1835, w_232_1854, w_232_1859, w_232_1861, w_232_1862, w_232_1868, w_232_1869, w_232_1876, w_232_1879, w_232_1882, w_232_1883, w_232_1885, w_232_1897, w_232_1899, w_232_1900, w_232_1903, w_232_1905, w_232_1914, w_232_1924, w_232_1928, w_232_1930, w_232_1931, w_232_1934, w_232_1939, w_232_1943, w_232_1950, w_232_1963, w_232_1964, w_232_1965, w_232_1966, w_232_1967, w_232_1968, w_232_1969, w_232_1970, w_232_1974, w_232_1975, w_232_1976, w_232_1978;
  wire w_233_008, w_233_011, w_233_013, w_233_018, w_233_019, w_233_021, w_233_023, w_233_027, w_233_028, w_233_029, w_233_036, w_233_040, w_233_041, w_233_049, w_233_053, w_233_066, w_233_070, w_233_072, w_233_076, w_233_080, w_233_081, w_233_084, w_233_089, w_233_090, w_233_093, w_233_098, w_233_099, w_233_105, w_233_108, w_233_114, w_233_122, w_233_124, w_233_129, w_233_131, w_233_132, w_233_135, w_233_138, w_233_145, w_233_146, w_233_147, w_233_148, w_233_155, w_233_165, w_233_171, w_233_173, w_233_174, w_233_176, w_233_177, w_233_179, w_233_181, w_233_184, w_233_185, w_233_187, w_233_191, w_233_194, w_233_197, w_233_198, w_233_199, w_233_207, w_233_208, w_233_211, w_233_214, w_233_219, w_233_221, w_233_223, w_233_225, w_233_227, w_233_230, w_233_232, w_233_237, w_233_239, w_233_242, w_233_243, w_233_252, w_233_254, w_233_260, w_233_262, w_233_267, w_233_269, w_233_278, w_233_281, w_233_285, w_233_288, w_233_290, w_233_291, w_233_295, w_233_307, w_233_312, w_233_314, w_233_319, w_233_320, w_233_321, w_233_322, w_233_323, w_233_327, w_233_328, w_233_329, w_233_330, w_233_333, w_233_338, w_233_339, w_233_340, w_233_348, w_233_360, w_233_364, w_233_365, w_233_374, w_233_375, w_233_380, w_233_382, w_233_389, w_233_398, w_233_401, w_233_402, w_233_405, w_233_417, w_233_418, w_233_419, w_233_420, w_233_423, w_233_427, w_233_432, w_233_433, w_233_434, w_233_437, w_233_441, w_233_445, w_233_446, w_233_447, w_233_455, w_233_459, w_233_462, w_233_463, w_233_467, w_233_471, w_233_473, w_233_478, w_233_481, w_233_491, w_233_506, w_233_508, w_233_509, w_233_520, w_233_522, w_233_524, w_233_526, w_233_528, w_233_532, w_233_535, w_233_536, w_233_543, w_233_544, w_233_548, w_233_549, w_233_550, w_233_557, w_233_565, w_233_566, w_233_573, w_233_581, w_233_592, w_233_593, w_233_606, w_233_611, w_233_617, w_233_618, w_233_622, w_233_625, w_233_627, w_233_628, w_233_630, w_233_633, w_233_636, w_233_645, w_233_648, w_233_651, w_233_652, w_233_653, w_233_654, w_233_660, w_233_676, w_233_681, w_233_682, w_233_686, w_233_688, w_233_691, w_233_695, w_233_696, w_233_698, w_233_707, w_233_711, w_233_716, w_233_723, w_233_726, w_233_730, w_233_733, w_233_735, w_233_740, w_233_745, w_233_751, w_233_767, w_233_768, w_233_773, w_233_775, w_233_780, w_233_795, w_233_799, w_233_804, w_233_806, w_233_808, w_233_809, w_233_813, w_233_816, w_233_817, w_233_821, w_233_822, w_233_841, w_233_843, w_233_844, w_233_852, w_233_858, w_233_860, w_233_868, w_233_873, w_233_884, w_233_885, w_233_890, w_233_894, w_233_898, w_233_906, w_233_918, w_233_940, w_233_945, w_233_960, w_233_962, w_233_967, w_233_970, w_233_972, w_233_976, w_233_979, w_233_980, w_233_983, w_233_986, w_233_992, w_233_995, w_233_996, w_233_1006, w_233_1008, w_233_1011, w_233_1014, w_233_1016, w_233_1024, w_233_1026, w_233_1029, w_233_1045, w_233_1064, w_233_1065, w_233_1070, w_233_1073, w_233_1078, w_233_1079, w_233_1088, w_233_1091, w_233_1092, w_233_1094, w_233_1102, w_233_1103, w_233_1106, w_233_1111, w_233_1114, w_233_1119, w_233_1129, w_233_1137, w_233_1138, w_233_1139, w_233_1142, w_233_1144, w_233_1151, w_233_1155, w_233_1156, w_233_1157, w_233_1164, w_233_1172, w_233_1173, w_233_1174, w_233_1178, w_233_1186, w_233_1195, w_233_1201, w_233_1202, w_233_1203, w_233_1213, w_233_1216, w_233_1217, w_233_1221, w_233_1228, w_233_1231, w_233_1243, w_233_1256, w_233_1262, w_233_1267, w_233_1270, w_233_1273, w_233_1284, w_233_1287, w_233_1288, w_233_1289, w_233_1300, w_233_1304, w_233_1311, w_233_1316, w_233_1325, w_233_1326, w_233_1328, w_233_1330, w_233_1331, w_233_1341, w_233_1348, w_233_1351, w_233_1353, w_233_1375, w_233_1376, w_233_1377, w_233_1378, w_233_1392, w_233_1393, w_233_1395, w_233_1400, w_233_1402, w_233_1406, w_233_1407, w_233_1410, w_233_1412, w_233_1415, w_233_1427, w_233_1433, w_233_1434, w_233_1448, w_233_1460, w_233_1464, w_233_1475, w_233_1485, w_233_1495, w_233_1515, w_233_1517, w_233_1522, w_233_1524, w_233_1534, w_233_1535, w_233_1537, w_233_1550, w_233_1553, w_233_1554, w_233_1558, w_233_1570, w_233_1576, w_233_1584, w_233_1589, w_233_1593, w_233_1597, w_233_1599, w_233_1601, w_233_1604, w_233_1615, w_233_1619, w_233_1627, w_233_1629, w_233_1639, w_233_1641, w_233_1645, w_233_1649, w_233_1650, w_233_1653, w_233_1658, w_233_1666, w_233_1674, w_233_1676, w_233_1681, w_233_1682, w_233_1692, w_233_1697, w_233_1699, w_233_1700, w_233_1704, w_233_1705, w_233_1709, w_233_1714, w_233_1725, w_233_1734, w_233_1736, w_233_1748, w_233_1753, w_233_1759, w_233_1763, w_233_1771, w_233_1787, w_233_1788, w_233_1806, w_233_1808, w_233_1810, w_233_1817, w_233_1819, w_233_1824, w_233_1831, w_233_1834, w_233_1835, w_233_1842, w_233_1843, w_233_1847, w_233_1851, w_233_1858, w_233_1866, w_233_1868, w_233_1871, w_233_1873, w_233_1875, w_233_1878, w_233_1882, w_233_1888, w_233_1894, w_233_1901, w_233_1906, w_233_1912, w_233_1914, w_233_1924, w_233_1931, w_233_1935, w_233_1945, w_233_1954, w_233_1960, w_233_1963, w_233_1969, w_233_1971, w_233_1981, w_233_1984, w_233_1993, w_233_2001, w_233_2002, w_233_2004, w_233_2007, w_233_2009, w_233_2010, w_233_2011, w_233_2018, w_233_2030, w_233_2034, w_233_2035, w_233_2038, w_233_2047, w_233_2049, w_233_2050, w_233_2053, w_233_2054, w_233_2063, w_233_2064, w_233_2070, w_233_2071, w_233_2076, w_233_2078, w_233_2080, w_233_2084, w_233_2110, w_233_2114, w_233_2115, w_233_2127, w_233_2129, w_233_2140, w_233_2144, w_233_2152, w_233_2157, w_233_2158, w_233_2162, w_233_2167, w_233_2169, w_233_2172, w_233_2176, w_233_2183, w_233_2196, w_233_2197, w_233_2202, w_233_2204, w_233_2215, w_233_2217, w_233_2237, w_233_2239, w_233_2240, w_233_2242, w_233_2244, w_233_2246, w_233_2250, w_233_2259, w_233_2260, w_233_2261, w_233_2262, w_233_2263, w_233_2264, w_233_2265, w_233_2266, w_233_2267, w_233_2268, w_233_2272, w_233_2273, w_233_2274, w_233_2275, w_233_2276, w_233_2277, w_233_2278, w_233_2279, w_233_2280, w_233_2281, w_233_2282, w_233_2283, w_233_2285;
  wire w_234_006, w_234_007, w_234_012, w_234_013, w_234_019, w_234_020, w_234_022, w_234_025, w_234_027, w_234_030, w_234_031, w_234_032, w_234_044, w_234_045, w_234_050, w_234_055, w_234_056, w_234_063, w_234_065, w_234_069, w_234_072, w_234_079, w_234_081, w_234_088, w_234_095, w_234_108, w_234_123, w_234_124, w_234_137, w_234_139, w_234_140, w_234_142, w_234_148, w_234_152, w_234_164, w_234_165, w_234_166, w_234_173, w_234_175, w_234_189, w_234_193, w_234_194, w_234_208, w_234_213, w_234_223, w_234_224, w_234_226, w_234_229, w_234_236, w_234_238, w_234_249, w_234_250, w_234_252, w_234_256, w_234_264, w_234_265, w_234_268, w_234_269, w_234_294, w_234_295, w_234_297, w_234_301, w_234_303, w_234_311, w_234_314, w_234_325, w_234_327, w_234_337, w_234_342, w_234_343, w_234_347, w_234_358, w_234_377, w_234_383, w_234_389, w_234_390, w_234_391, w_234_392, w_234_394, w_234_397, w_234_399, w_234_404, w_234_405, w_234_408, w_234_410, w_234_411, w_234_414, w_234_415, w_234_417, w_234_433, w_234_440, w_234_441, w_234_447, w_234_455, w_234_460, w_234_465, w_234_467, w_234_476, w_234_485, w_234_486, w_234_489, w_234_490, w_234_491, w_234_497, w_234_503, w_234_504, w_234_506, w_234_513, w_234_518, w_234_519, w_234_524, w_234_532, w_234_533, w_234_540, w_234_543, w_234_546, w_234_554, w_234_559, w_234_561, w_234_572, w_234_575, w_234_577, w_234_589, w_234_592, w_234_598, w_234_600, w_234_601, w_234_607, w_234_608, w_234_609, w_234_618, w_234_620, w_234_622, w_234_627, w_234_631, w_234_634, w_234_635, w_234_637, w_234_638, w_234_639, w_234_642, w_234_644, w_234_646, w_234_651, w_234_656, w_234_663, w_234_673, w_234_679, w_234_684, w_234_686, w_234_695, w_234_698, w_234_699, w_234_700, w_234_704, w_234_707, w_234_709, w_234_710, w_234_718, w_234_723, w_234_733, w_234_737, w_234_742, w_234_743, w_234_745, w_234_749, w_234_750, w_234_760, w_234_764, w_234_767, w_234_772, w_234_776, w_234_779, w_234_788, w_234_806, w_234_813, w_234_814, w_234_815, w_234_820, w_234_827, w_234_833, w_234_854, w_234_855, w_234_864, w_234_870, w_234_876, w_234_878, w_234_884, w_234_885, w_234_890, w_234_907, w_234_913, w_234_920, w_234_944, w_234_945, w_234_953, w_234_957, w_234_968, w_234_970, w_234_971, w_234_976, w_234_985, w_234_990, w_234_991, w_234_992, w_234_993, w_234_1008, w_234_1031, w_234_1032, w_234_1034, w_234_1041, w_234_1043, w_234_1044, w_234_1048, w_234_1061, w_234_1065, w_234_1073, w_234_1080, w_234_1096, w_234_1098, w_234_1103, w_234_1106, w_234_1114, w_234_1116, w_234_1122, w_234_1123, w_234_1134, w_234_1159, w_234_1162, w_234_1166, w_234_1170, w_234_1174, w_234_1182, w_234_1188, w_234_1189, w_234_1201, w_234_1220, w_234_1231, w_234_1235, w_234_1237, w_234_1254, w_234_1257, w_234_1259, w_234_1262, w_234_1265, w_234_1266, w_234_1267, w_234_1278, w_234_1289, w_234_1293, w_234_1298, w_234_1303, w_234_1304, w_234_1305, w_234_1309, w_234_1314, w_234_1329, w_234_1333, w_234_1336, w_234_1340, w_234_1349, w_234_1367, w_234_1368, w_234_1369, w_234_1372, w_234_1379, w_234_1383, w_234_1386, w_234_1387, w_234_1389, w_234_1395, w_234_1418, w_234_1419, w_234_1426, w_234_1436, w_234_1454, w_234_1487, w_234_1505, w_234_1506, w_234_1509, w_234_1518, w_234_1530, w_234_1539, w_234_1540, w_234_1561, w_234_1590, w_234_1591, w_234_1596, w_234_1619, w_234_1634, w_234_1645, w_234_1666, w_234_1710, w_234_1715, w_234_1726, w_234_1730, w_234_1734, w_234_1749, w_234_1750, w_234_1763, w_234_1768, w_234_1773, w_234_1776, w_234_1802, w_234_1813, w_234_1827, w_234_1837, w_234_1838, w_234_1842, w_234_1844, w_234_1853, w_234_1866, w_234_1869, w_234_1878, w_234_1885, w_234_1900, w_234_1901, w_234_1903, w_234_1920, w_234_1928, w_234_1951, w_234_1952, w_234_1965, w_234_1970, w_234_1980, w_234_1987, w_234_1997, w_234_2002, w_234_2004, w_234_2017, w_234_2019, w_234_2023, w_234_2029, w_234_2030, w_234_2054, w_234_2059, w_234_2064, w_234_2079, w_234_2086, w_234_2099, w_234_2101, w_234_2104, w_234_2133, w_234_2174, w_234_2177, w_234_2183, w_234_2187, w_234_2188, w_234_2191, w_234_2217, w_234_2222, w_234_2223, w_234_2247, w_234_2254, w_234_2258, w_234_2261, w_234_2265, w_234_2269, w_234_2274, w_234_2300, w_234_2305, w_234_2311, w_234_2329, w_234_2330, w_234_2332, w_234_2363, w_234_2368, w_234_2378, w_234_2381, w_234_2392, w_234_2397, w_234_2410, w_234_2412, w_234_2414, w_234_2422, w_234_2429, w_234_2444, w_234_2457, w_234_2466, w_234_2504, w_234_2506, w_234_2552, w_234_2567, w_234_2585, w_234_2586, w_234_2588, w_234_2598, w_234_2610, w_234_2645, w_234_2651, w_234_2690, w_234_2702, w_234_2705, w_234_2757, w_234_2770, w_234_2783, w_234_2789, w_234_2799, w_234_2802, w_234_2828, w_234_2833, w_234_2836, w_234_2839, w_234_2862, w_234_2876, w_234_2877, w_234_2880, w_234_2893, w_234_2908, w_234_2932, w_234_2955, w_234_2963, w_234_2965, w_234_2973, w_234_2974, w_234_2985, w_234_2986, w_234_2988, w_234_2994, w_234_3003, w_234_3020, w_234_3030, w_234_3035, w_234_3045, w_234_3059, w_234_3060, w_234_3072, w_234_3089, w_234_3091, w_234_3094, w_234_3121, w_234_3127, w_234_3131, w_234_3139, w_234_3167, w_234_3168, w_234_3176, w_234_3180, w_234_3198, w_234_3202, w_234_3204, w_234_3214, w_234_3217, w_234_3218, w_234_3243, w_234_3245, w_234_3252, w_234_3257, w_234_3258, w_234_3262, w_234_3269, w_234_3275, w_234_3278, w_234_3279, w_234_3285, w_234_3287, w_234_3292, w_234_3296, w_234_3306, w_234_3319, w_234_3321, w_234_3326, w_234_3330, w_234_3338, w_234_3348, w_234_3367, w_234_3373, w_234_3387, w_234_3399, w_234_3409, w_234_3426, w_234_3427, w_234_3429, w_234_3442, w_234_3452, w_234_3453, w_234_3472, w_234_3476, w_234_3502, w_234_3508, w_234_3511, w_234_3514, w_234_3524, w_234_3536, w_234_3545, w_234_3571, w_234_3575, w_234_3579, w_234_3588, w_234_3592, w_234_3604, w_234_3605, w_234_3606, w_234_3608, w_234_3610, w_234_3611, w_234_3612, w_234_3613, w_234_3614, w_234_3615, w_234_3616, w_234_3617, w_234_3618, w_234_3619, w_234_3620, w_234_3621, w_234_3623;
  wire w_235_001, w_235_002, w_235_006, w_235_007, w_235_008, w_235_009, w_235_011, w_235_012, w_235_013, w_235_014, w_235_015, w_235_016, w_235_017, w_235_018, w_235_019, w_235_020, w_235_021, w_235_022, w_235_023, w_235_024, w_235_026, w_235_027, w_235_028, w_235_029, w_235_030, w_235_031, w_235_032, w_235_033, w_235_034, w_235_035, w_235_037, w_235_038, w_235_040, w_235_041, w_235_042, w_235_044, w_235_045, w_235_046, w_235_047, w_235_048, w_235_050, w_235_053, w_235_054, w_235_056, w_235_057, w_235_059, w_235_060, w_235_061, w_235_062, w_235_063, w_235_064, w_235_066, w_235_070, w_235_071, w_235_072, w_235_073, w_235_074, w_235_075, w_235_076, w_235_077, w_235_079, w_235_080, w_235_083, w_235_084, w_235_085, w_235_086, w_235_088, w_235_089, w_235_090, w_235_091, w_235_092, w_235_093, w_235_094, w_235_095, w_235_096, w_235_097, w_235_099, w_235_100, w_235_101, w_235_103, w_235_104, w_235_105, w_235_107, w_235_108, w_235_109, w_235_111, w_235_112, w_235_114, w_235_115, w_235_116, w_235_118, w_235_119, w_235_120, w_235_121, w_235_122, w_235_123, w_235_125, w_235_126, w_235_127, w_235_128, w_235_129, w_235_131, w_235_132, w_235_133, w_235_134, w_235_136, w_235_137, w_235_138, w_235_139, w_235_140, w_235_141, w_235_142, w_235_143, w_235_144, w_235_145, w_235_146, w_235_147, w_235_148, w_235_149, w_235_150, w_235_151, w_235_152, w_235_153, w_235_155, w_235_156, w_235_157, w_235_158, w_235_159, w_235_160, w_235_161, w_235_162, w_235_163, w_235_164, w_235_165, w_235_166, w_235_168, w_235_169, w_235_170, w_235_171, w_235_172, w_235_174, w_235_175, w_235_176, w_235_178, w_235_179, w_235_182, w_235_183, w_235_187, w_235_188, w_235_189, w_235_191, w_235_192, w_235_193, w_235_194, w_235_196, w_235_197, w_235_198, w_235_200, w_235_201, w_235_202, w_235_203, w_235_204, w_235_206, w_235_207, w_235_210, w_235_211, w_235_213, w_235_214, w_235_217, w_235_218, w_235_219, w_235_221, w_235_222, w_235_223, w_235_224, w_235_225, w_235_227, w_235_229, w_235_230, w_235_231, w_235_232, w_235_233, w_235_235, w_235_237, w_235_238, w_235_239, w_235_240, w_235_241, w_235_242, w_235_243, w_235_244, w_235_245, w_235_246, w_235_247, w_235_248, w_235_250, w_235_251, w_235_252, w_235_253, w_235_254, w_235_255, w_235_256, w_235_257, w_235_259, w_235_260, w_235_261, w_235_262, w_235_263, w_235_264, w_235_267, w_235_268, w_235_269, w_235_270, w_235_271, w_235_272, w_235_273, w_235_274, w_235_275, w_235_276, w_235_277, w_235_278, w_235_282, w_235_284, w_235_286, w_235_287, w_235_288, w_235_289, w_235_291, w_235_292, w_235_293, w_235_295, w_235_296, w_235_297, w_235_299, w_235_302, w_235_303, w_235_305, w_235_306, w_235_307, w_235_308, w_235_309, w_235_310, w_235_311, w_235_312, w_235_314, w_235_315, w_235_316, w_235_317, w_235_318, w_235_320, w_235_321, w_235_322, w_235_323, w_235_324, w_235_326, w_235_327, w_235_328, w_235_329, w_235_330, w_235_335, w_235_336, w_235_338, w_235_339, w_235_341, w_235_343, w_235_344, w_235_345, w_235_346, w_235_347, w_235_349, w_235_350, w_235_351, w_235_353, w_235_354, w_235_355, w_235_356, w_235_358, w_235_359, w_235_360, w_235_363, w_235_365;
  wire w_236_004, w_236_005, w_236_010, w_236_014, w_236_017, w_236_018, w_236_029, w_236_030, w_236_031, w_236_032, w_236_036, w_236_038, w_236_040, w_236_046, w_236_048, w_236_049, w_236_051, w_236_053, w_236_054, w_236_055, w_236_057, w_236_059, w_236_061, w_236_062, w_236_064, w_236_068, w_236_070, w_236_071, w_236_074, w_236_075, w_236_080, w_236_083, w_236_084, w_236_087, w_236_090, w_236_091, w_236_093, w_236_094, w_236_100, w_236_107, w_236_113, w_236_115, w_236_117, w_236_118, w_236_120, w_236_121, w_236_132, w_236_135, w_236_136, w_236_137, w_236_141, w_236_143, w_236_146, w_236_156, w_236_158, w_236_164, w_236_177, w_236_180, w_236_181, w_236_184, w_236_188, w_236_194, w_236_203, w_236_207, w_236_209, w_236_213, w_236_215, w_236_218, w_236_219, w_236_220, w_236_221, w_236_229, w_236_232, w_236_233, w_236_234, w_236_237, w_236_239, w_236_242, w_236_246, w_236_259, w_236_260, w_236_262, w_236_266, w_236_268, w_236_269, w_236_272, w_236_273, w_236_278, w_236_291, w_236_297, w_236_301, w_236_303, w_236_306, w_236_308, w_236_315, w_236_316, w_236_318, w_236_319, w_236_320, w_236_322, w_236_331, w_236_333, w_236_338, w_236_343, w_236_354, w_236_356, w_236_362, w_236_363, w_236_364, w_236_368, w_236_370, w_236_371, w_236_374, w_236_379, w_236_386, w_236_390, w_236_396, w_236_401, w_236_404, w_236_405, w_236_412, w_236_413, w_236_414, w_236_417, w_236_418, w_236_427, w_236_428, w_236_429, w_236_432, w_236_433, w_236_440, w_236_441, w_236_442, w_236_449, w_236_450, w_236_451, w_236_454, w_236_462, w_236_465, w_236_466, w_236_470, w_236_489, w_236_491, w_236_494, w_236_495, w_236_502, w_236_506, w_236_508, w_236_514, w_236_515, w_236_516, w_236_518, w_236_520, w_236_524, w_236_525, w_236_529, w_236_531, w_236_534, w_236_535, w_236_536, w_236_544, w_236_545, w_236_546, w_236_558, w_236_565, w_236_568, w_236_569, w_236_573, w_236_578, w_236_579, w_236_581, w_236_584, w_236_585, w_236_587, w_236_597, w_236_598, w_236_602, w_236_603, w_236_604, w_236_610, w_236_611, w_236_613, w_236_619, w_236_622, w_236_623, w_236_624, w_236_625, w_236_628, w_236_631, w_236_632, w_236_634, w_236_635, w_236_636, w_236_638, w_236_639, w_236_641, w_236_645, w_236_646, w_236_649, w_236_651, w_236_653, w_236_655, w_236_660, w_236_665, w_236_671, w_236_673, w_236_675, w_236_676, w_236_677, w_236_686, w_236_687, w_236_693, w_236_694, w_236_695, w_236_699, w_236_711, w_236_712, w_236_716, w_236_718, w_236_719, w_236_720, w_236_721, w_236_727, w_236_728, w_236_729, w_236_730, w_236_732, w_236_742, w_236_744, w_236_750, w_236_752, w_236_753, w_236_762, w_236_763, w_236_770, w_236_779, w_236_781, w_236_788, w_236_790, w_236_793, w_236_798, w_236_807, w_236_811, w_236_812, w_236_818, w_236_822, w_236_823, w_236_827, w_236_828, w_236_830, w_236_832, w_236_838, w_236_840, w_236_848, w_236_855, w_236_856, w_236_859, w_236_861, w_236_863, w_236_868, w_236_874, w_236_875, w_236_879, w_236_889, w_236_892, w_236_894, w_236_895, w_236_896, w_236_898, w_236_899, w_236_901, w_236_904, w_236_905, w_236_913, w_236_915, w_236_919, w_236_922, w_236_929, w_236_936, w_236_945, w_236_948, w_236_952, w_236_953, w_236_963, w_236_968, w_236_969, w_236_970, w_236_972, w_236_974, w_236_983, w_236_988, w_236_995, w_236_997, w_236_1000, w_236_1001, w_236_1004, w_236_1012, w_236_1015, w_236_1016, w_236_1018, w_236_1025, w_236_1028, w_236_1030, w_236_1031, w_236_1036, w_236_1043, w_236_1047, w_236_1049, w_236_1053, w_236_1054, w_236_1055, w_236_1060, w_236_1061, w_236_1063, w_236_1068, w_236_1069, w_236_1074, w_236_1083, w_236_1089, w_236_1090, w_236_1097, w_236_1103, w_236_1104, w_236_1105, w_236_1109, w_236_1117, w_236_1122, w_236_1123, w_236_1125, w_236_1130, w_236_1132, w_236_1133, w_236_1135, w_236_1137, w_236_1145, w_236_1151, w_236_1159, w_236_1160, w_236_1161, w_236_1163, w_236_1164, w_236_1170, w_236_1173, w_236_1174, w_236_1175, w_236_1189, w_236_1191, w_236_1192, w_236_1193, w_236_1195, w_236_1198, w_236_1203, w_236_1207, w_236_1209, w_236_1212, w_236_1227, w_236_1228, w_236_1229, w_236_1233, w_236_1240, w_236_1243, w_236_1251, w_236_1260, w_236_1262, w_236_1269, w_236_1270, w_236_1276, w_236_1284, w_236_1286, w_236_1289, w_236_1292, w_236_1294, w_236_1296, w_236_1300, w_236_1308, w_236_1310, w_236_1311, w_236_1318, w_236_1319, w_236_1322, w_236_1327, w_236_1342, w_236_1350, w_236_1354, w_236_1358, w_236_1359, w_236_1360, w_236_1363, w_236_1367, w_236_1369, w_236_1372, w_236_1373, w_236_1376, w_236_1377, w_236_1378, w_236_1381, w_236_1384, w_236_1387, w_236_1388, w_236_1391, w_236_1392, w_236_1396, w_236_1398, w_236_1407, w_236_1408, w_236_1409, w_236_1412, w_236_1417, w_236_1421, w_236_1423, w_236_1426, w_236_1433, w_236_1434, w_236_1441, w_236_1443, w_236_1444, w_236_1447, w_236_1448, w_236_1451, w_236_1456, w_236_1457, w_236_1462, w_236_1463, w_236_1467, w_236_1474, w_236_1477, w_236_1480, w_236_1481, w_236_1484, w_236_1488, w_236_1489, w_236_1490, w_236_1491, w_236_1496, w_236_1503, w_236_1505, w_236_1506, w_236_1507, w_236_1509, w_236_1514, w_236_1517, w_236_1523, w_236_1526, w_236_1529, w_236_1530, w_236_1531, w_236_1532, w_236_1534, w_236_1535, w_236_1547, w_236_1548, w_236_1549, w_236_1550, w_236_1554, w_236_1555, w_236_1556, w_236_1565, w_236_1567, w_236_1574, w_236_1575, w_236_1577, w_236_1578, w_236_1579, w_236_1582, w_236_1583, w_236_1586, w_236_1591, w_236_1594, w_236_1597, w_236_1598, w_236_1603, w_236_1605, w_236_1612, w_236_1621, w_236_1624, w_236_1626, w_236_1630, w_236_1632, w_236_1634;
  wire w_237_006, w_237_015, w_237_017, w_237_028, w_237_030, w_237_037, w_237_043, w_237_044, w_237_045, w_237_052, w_237_053, w_237_069, w_237_071, w_237_072, w_237_074, w_237_078, w_237_081, w_237_086, w_237_092, w_237_094, w_237_095, w_237_098, w_237_100, w_237_108, w_237_111, w_237_113, w_237_114, w_237_116, w_237_118, w_237_126, w_237_131, w_237_146, w_237_147, w_237_176, w_237_183, w_237_185, w_237_188, w_237_191, w_237_205, w_237_208, w_237_221, w_237_228, w_237_230, w_237_235, w_237_239, w_237_246, w_237_257, w_237_274, w_237_283, w_237_288, w_237_292, w_237_330, w_237_332, w_237_334, w_237_346, w_237_354, w_237_358, w_237_370, w_237_378, w_237_403, w_237_404, w_237_410, w_237_413, w_237_414, w_237_421, w_237_464, w_237_475, w_237_482, w_237_502, w_237_506, w_237_513, w_237_526, w_237_558, w_237_574, w_237_580, w_237_582, w_237_588, w_237_589, w_237_603, w_237_647, w_237_653, w_237_662, w_237_666, w_237_668, w_237_674, w_237_692, w_237_696, w_237_712, w_237_720, w_237_731, w_237_742, w_237_744, w_237_746, w_237_751, w_237_757, w_237_766, w_237_770, w_237_783, w_237_786, w_237_795, w_237_798, w_237_806, w_237_808, w_237_818, w_237_822, w_237_844, w_237_850, w_237_890, w_237_895, w_237_904, w_237_913, w_237_916, w_237_917, w_237_934, w_237_935, w_237_936, w_237_938, w_237_950, w_237_955, w_237_981, w_237_994, w_237_1010, w_237_1012, w_237_1018, w_237_1019, w_237_1028, w_237_1043, w_237_1044, w_237_1058, w_237_1084, w_237_1090, w_237_1096, w_237_1098, w_237_1104, w_237_1108, w_237_1118, w_237_1127, w_237_1134, w_237_1135, w_237_1148, w_237_1154, w_237_1162, w_237_1188, w_237_1192, w_237_1213, w_237_1215, w_237_1219, w_237_1220, w_237_1250, w_237_1254, w_237_1258, w_237_1287, w_237_1311, w_237_1318, w_237_1326, w_237_1330, w_237_1337, w_237_1338, w_237_1371, w_237_1387, w_237_1399, w_237_1416, w_237_1442, w_237_1446, w_237_1462, w_237_1466, w_237_1481, w_237_1490, w_237_1491, w_237_1495, w_237_1501, w_237_1505, w_237_1515, w_237_1516, w_237_1517, w_237_1518, w_237_1521, w_237_1549, w_237_1552, w_237_1555, w_237_1563, w_237_1564, w_237_1566, w_237_1575, w_237_1580, w_237_1596, w_237_1603, w_237_1605, w_237_1627, w_237_1636, w_237_1641, w_237_1664, w_237_1669, w_237_1693, w_237_1699, w_237_1716, w_237_1718, w_237_1723, w_237_1727, w_237_1729, w_237_1733, w_237_1759, w_237_1763, w_237_1783, w_237_1784, w_237_1803, w_237_1822, w_237_1839, w_237_1856, w_237_1861, w_237_1867, w_237_1868, w_237_1882, w_237_1886, w_237_1889, w_237_1899, w_237_1916, w_237_1928, w_237_1942, w_237_1943, w_237_1946, w_237_1953, w_237_1958, w_237_1960, w_237_1971, w_237_2017, w_237_2031, w_237_2045, w_237_2053, w_237_2064, w_237_2073, w_237_2080, w_237_2082, w_237_2087, w_237_2091, w_237_2109, w_237_2122, w_237_2129, w_237_2143, w_237_2210, w_237_2213, w_237_2222, w_237_2224, w_237_2239, w_237_2248, w_237_2249, w_237_2255, w_237_2257, w_237_2262, w_237_2292, w_237_2309, w_237_2311, w_237_2312, w_237_2314, w_237_2357, w_237_2363, w_237_2369, w_237_2386, w_237_2399, w_237_2404, w_237_2405, w_237_2412, w_237_2414, w_237_2426, w_237_2427, w_237_2431, w_237_2444, w_237_2453, w_237_2465, w_237_2482, w_237_2484, w_237_2491, w_237_2531, w_237_2544, w_237_2552, w_237_2576, w_237_2592, w_237_2601, w_237_2609, w_237_2610, w_237_2611, w_237_2627, w_237_2633, w_237_2651, w_237_2663, w_237_2673, w_237_2678, w_237_2688, w_237_2706, w_237_2718, w_237_2723, w_237_2725, w_237_2728, w_237_2729, w_237_2733, w_237_2741, w_237_2743, w_237_2766, w_237_2775, w_237_2779, w_237_2781, w_237_2790, w_237_2800, w_237_2812, w_237_2818, w_237_2825, w_237_2840, w_237_2845, w_237_2847, w_237_2851, w_237_2852, w_237_2861, w_237_2866, w_237_2870, w_237_2879, w_237_2880, w_237_2883, w_237_2907, w_237_2911, w_237_2914, w_237_2924, w_237_2929, w_237_2940, w_237_2946, w_237_2948, w_237_2968, w_237_2971, w_237_2986, w_237_2989, w_237_2999, w_237_3015, w_237_3025, w_237_3033, w_237_3043, w_237_3046, w_237_3066, w_237_3069, w_237_3074, w_237_3084, w_237_3097, w_237_3098, w_237_3101, w_237_3107, w_237_3108, w_237_3136, w_237_3147, w_237_3149, w_237_3152, w_237_3155, w_237_3171, w_237_3176, w_237_3182, w_237_3192, w_237_3195, w_237_3228, w_237_3232, w_237_3249, w_237_3263, w_237_3266, w_237_3267, w_237_3273, w_237_3281, w_237_3285, w_237_3286, w_237_3289, w_237_3316, w_237_3325, w_237_3337, w_237_3342, w_237_3349, w_237_3351, w_237_3360, w_237_3373, w_237_3399, w_237_3404, w_237_3421, w_237_3429, w_237_3434, w_237_3442, w_237_3469, w_237_3472, w_237_3491, w_237_3492, w_237_3494, w_237_3496, w_237_3505, w_237_3510, w_237_3512, w_237_3516, w_237_3524, w_237_3556, w_237_3560, w_237_3563, w_237_3583, w_237_3584, w_237_3592, w_237_3597, w_237_3599, w_237_3610, w_237_3615, w_237_3619, w_237_3625, w_237_3635, w_237_3648, w_237_3671, w_237_3675, w_237_3678, w_237_3687, w_237_3688, w_237_3693, w_237_3703, w_237_3712, w_237_3740, w_237_3747, w_237_3766, w_237_3794, w_237_3801, w_237_3819, w_237_3821, w_237_3831, w_237_3833, w_237_3839, w_237_3843, w_237_3861, w_237_3865, w_237_3879, w_237_3890, w_237_3895, w_237_3912, w_237_3924, w_237_3953, w_237_3960, w_237_3965, w_237_3968, w_237_3980, w_237_3986, w_237_3997, w_237_4010, w_237_4023, w_237_4033, w_237_4034, w_237_4036, w_237_4038, w_237_4052, w_237_4054, w_237_4058, w_237_4062, w_237_4075, w_237_4078, w_237_4100, w_237_4103, w_237_4110, w_237_4118, w_237_4122, w_237_4127, w_237_4136, w_237_4183, w_237_4192, w_237_4202, w_237_4211, w_237_4215, w_237_4224, w_237_4239, w_237_4257, w_237_4265, w_237_4268, w_237_4284, w_237_4286, w_237_4292, w_237_4294, w_237_4303, w_237_4313, w_237_4321, w_237_4328, w_237_4329, w_237_4335, w_237_4345, w_237_4347, w_237_4354, w_237_4369, w_237_4375, w_237_4408, w_237_4414, w_237_4415, w_237_4425, w_237_4428, w_237_4452, w_237_4455, w_237_4461, w_237_4485, w_237_4493, w_237_4510, w_237_4528, w_237_4531, w_237_4537, w_237_4542, w_237_4547, w_237_4550, w_237_4594, w_237_4599, w_237_4620, w_237_4625, w_237_4640, w_237_4661, w_237_4667, w_237_4669, w_237_4670, w_237_4671, w_237_4681, w_237_4689, w_237_4694, w_237_4698, w_237_4721, w_237_4728, w_237_4729, w_237_4732, w_237_4737, w_237_4744, w_237_4747, w_237_4767, w_237_4787, w_237_4791, w_237_4796, w_237_4801, w_237_4812, w_237_4836, w_237_4839, w_237_4847, w_237_4854, w_237_4855, w_237_4868, w_237_4882, w_237_4883, w_237_4884, w_237_4885;
  wire w_238_000, w_238_001, w_238_002, w_238_003, w_238_004, w_238_005, w_238_007, w_238_008, w_238_009, w_238_010, w_238_011, w_238_012, w_238_013, w_238_015, w_238_016, w_238_017, w_238_019, w_238_020, w_238_021, w_238_023, w_238_024, w_238_025, w_238_027, w_238_028, w_238_029, w_238_030, w_238_031, w_238_032, w_238_033, w_238_034, w_238_035, w_238_036, w_238_037, w_238_038, w_238_039, w_238_040, w_238_041, w_238_042, w_238_043, w_238_044, w_238_045, w_238_046, w_238_047, w_238_048, w_238_049, w_238_050, w_238_051, w_238_052, w_238_053, w_238_054, w_238_055, w_238_056, w_238_057, w_238_058, w_238_059, w_238_060, w_238_061, w_238_062, w_238_064, w_238_065, w_238_067, w_238_068, w_238_070, w_238_071, w_238_072, w_238_073, w_238_074, w_238_075, w_238_076, w_238_077, w_238_078, w_238_079, w_238_080, w_238_081, w_238_082, w_238_083, w_238_084, w_238_085, w_238_086, w_238_087, w_238_088, w_238_089, w_238_090, w_238_091, w_238_092, w_238_093, w_238_094, w_238_095, w_238_096, w_238_097, w_238_099, w_238_101, w_238_102, w_238_103, w_238_104, w_238_105, w_238_106, w_238_107, w_238_108, w_238_109, w_238_110, w_238_111, w_238_112, w_238_113, w_238_114, w_238_115, w_238_116, w_238_117, w_238_120, w_238_121, w_238_122, w_238_123, w_238_124, w_238_125, w_238_126, w_238_127, w_238_128, w_238_130, w_238_131, w_238_132, w_238_133, w_238_134, w_238_135, w_238_137, w_238_139, w_238_140, w_238_141, w_238_142, w_238_143, w_238_144, w_238_145, w_238_146, w_238_147, w_238_149, w_238_150, w_238_151, w_238_153, w_238_154, w_238_155, w_238_156, w_238_157, w_238_158, w_238_159, w_238_160, w_238_161, w_238_162, w_238_163, w_238_164, w_238_165, w_238_166, w_238_167, w_238_168, w_238_169, w_238_170, w_238_171, w_238_172, w_238_173, w_238_174, w_238_175, w_238_176, w_238_177, w_238_178, w_238_179, w_238_180, w_238_181, w_238_183, w_238_184, w_238_185, w_238_186, w_238_187, w_238_189, w_238_190, w_238_191, w_238_192, w_238_194, w_238_195, w_238_196, w_238_197, w_238_198, w_238_199, w_238_200, w_238_201, w_238_202, w_238_204, w_238_205, w_238_206, w_238_207, w_238_208, w_238_209, w_238_210, w_238_211, w_238_212, w_238_213, w_238_215, w_238_216, w_238_219, w_238_220, w_238_221, w_238_222, w_238_224, w_238_225, w_238_226, w_238_227, w_238_228, w_238_229, w_238_230, w_238_234, w_238_235, w_238_236, w_238_237, w_238_238, w_238_239, w_238_240, w_238_241, w_238_243;
  wire w_239_001, w_239_005, w_239_019, w_239_027, w_239_055, w_239_056, w_239_061, w_239_067, w_239_070, w_239_080, w_239_081, w_239_085, w_239_091, w_239_105, w_239_108, w_239_110, w_239_117, w_239_119, w_239_121, w_239_122, w_239_127, w_239_133, w_239_141, w_239_145, w_239_148, w_239_149, w_239_153, w_239_154, w_239_155, w_239_159, w_239_160, w_239_161, w_239_168, w_239_169, w_239_175, w_239_178, w_239_185, w_239_186, w_239_187, w_239_188, w_239_195, w_239_205, w_239_206, w_239_212, w_239_220, w_239_221, w_239_248, w_239_252, w_239_254, w_239_264, w_239_270, w_239_274, w_239_278, w_239_285, w_239_291, w_239_294, w_239_305, w_239_314, w_239_320, w_239_324, w_239_326, w_239_334, w_239_336, w_239_346, w_239_351, w_239_353, w_239_367, w_239_371, w_239_376, w_239_389, w_239_391, w_239_396, w_239_403, w_239_409, w_239_410, w_239_416, w_239_417, w_239_424, w_239_426, w_239_438, w_239_449, w_239_458, w_239_462, w_239_463, w_239_471, w_239_475, w_239_478, w_239_480, w_239_484, w_239_496, w_239_502, w_239_504, w_239_509, w_239_521, w_239_532, w_239_545, w_239_549, w_239_550, w_239_551, w_239_569, w_239_576, w_239_583, w_239_589, w_239_595, w_239_597, w_239_602, w_239_607, w_239_612, w_239_620, w_239_622, w_239_624, w_239_629, w_239_635, w_239_640, w_239_647, w_239_650, w_239_656, w_239_657, w_239_661, w_239_664, w_239_666, w_239_668, w_239_672, w_239_673, w_239_674, w_239_685, w_239_686, w_239_704, w_239_712, w_239_719, w_239_720, w_239_725, w_239_728, w_239_729, w_239_731, w_239_738, w_239_743, w_239_749, w_239_754, w_239_768, w_239_777, w_239_779, w_239_785, w_239_790, w_239_792, w_239_794, w_239_796, w_239_799, w_239_808, w_239_818, w_239_819, w_239_828, w_239_832, w_239_837, w_239_839, w_239_843, w_239_847, w_239_850, w_239_851, w_239_853, w_239_862, w_239_870, w_239_876, w_239_884, w_239_889, w_239_898, w_239_900, w_239_904, w_239_909, w_239_910, w_239_922, w_239_923, w_239_927, w_239_931, w_239_934, w_239_948, w_239_951, w_239_957, w_239_958, w_239_962, w_239_964, w_239_970, w_239_977, w_239_978, w_239_980, w_239_989, w_239_996, w_239_998, w_239_999, w_239_1009, w_239_1016, w_239_1028, w_239_1034, w_239_1035, w_239_1036, w_239_1037, w_239_1044, w_239_1054, w_239_1065, w_239_1079, w_239_1084, w_239_1089, w_239_1091, w_239_1094, w_239_1096, w_239_1098, w_239_1100, w_239_1105, w_239_1115, w_239_1119, w_239_1121, w_239_1133, w_239_1136, w_239_1138, w_239_1142, w_239_1143, w_239_1148, w_239_1150, w_239_1162, w_239_1163, w_239_1167, w_239_1170, w_239_1176, w_239_1178, w_239_1181, w_239_1199, w_239_1202, w_239_1204, w_239_1205, w_239_1209, w_239_1216, w_239_1225, w_239_1241, w_239_1261, w_239_1275, w_239_1278, w_239_1294, w_239_1296, w_239_1302, w_239_1305, w_239_1310, w_239_1315, w_239_1316, w_239_1336, w_239_1340, w_239_1366, w_239_1377, w_239_1381, w_239_1383, w_239_1398, w_239_1402, w_239_1425, w_239_1429, w_239_1436, w_239_1448, w_239_1457, w_239_1463, w_239_1469, w_239_1476, w_239_1483, w_239_1492, w_239_1505, w_239_1518, w_239_1519, w_239_1526, w_239_1538, w_239_1547, w_239_1548, w_239_1552, w_239_1559, w_239_1564, w_239_1565, w_239_1575, w_239_1576, w_239_1599, w_239_1624, w_239_1625, w_239_1632, w_239_1634, w_239_1638, w_239_1670, w_239_1685, w_239_1693, w_239_1699, w_239_1707, w_239_1715, w_239_1717, w_239_1726, w_239_1732, w_239_1737, w_239_1739, w_239_1769, w_239_1774, w_239_1776, w_239_1787, w_239_1791, w_239_1802, w_239_1803, w_239_1805, w_239_1820, w_239_1822, w_239_1834, w_239_1855, w_239_1856, w_239_1858, w_239_1870, w_239_1885, w_239_1905, w_239_1929, w_239_1931, w_239_1939, w_239_1944, w_239_1950, w_239_1962, w_239_1973, w_239_1988, w_239_2002, w_239_2011, w_239_2075, w_239_2087, w_239_2105, w_239_2116, w_239_2122, w_239_2127, w_239_2132, w_239_2140, w_239_2147, w_239_2153, w_239_2173, w_239_2176, w_239_2182, w_239_2192, w_239_2202, w_239_2208, w_239_2219, w_239_2223, w_239_2232, w_239_2238, w_239_2249, w_239_2263, w_239_2266, w_239_2268, w_239_2276, w_239_2281, w_239_2310, w_239_2311, w_239_2336, w_239_2371, w_239_2382, w_239_2384, w_239_2387, w_239_2388, w_239_2390, w_239_2406, w_239_2407, w_239_2410, w_239_2416, w_239_2418, w_239_2422, w_239_2424, w_239_2427, w_239_2429, w_239_2435, w_239_2440, w_239_2451, w_239_2471, w_239_2476, w_239_2478, w_239_2493, w_239_2529, w_239_2534, w_239_2544, w_239_2545, w_239_2549, w_239_2554, w_239_2632, w_239_2638, w_239_2657, w_239_2659, w_239_2679, w_239_2688, w_239_2691, w_239_2708, w_239_2712, w_239_2716, w_239_2717, w_239_2733, w_239_2735, w_239_2746, w_239_2764, w_239_2769, w_239_2777, w_239_2779, w_239_2812, w_239_2821, w_239_2830, w_239_2833, w_239_2844, w_239_2856, w_239_2871, w_239_2886, w_239_2903, w_239_2905, w_239_2913, w_239_2954, w_239_2956, w_239_2978, w_239_3011, w_239_3015, w_239_3052, w_239_3056, w_239_3067, w_239_3068, w_239_3094, w_239_3098, w_239_3102, w_239_3131, w_239_3132, w_239_3134, w_239_3168, w_239_3169, w_239_3175, w_239_3188, w_239_3191, w_239_3200, w_239_3210, w_239_3213, w_239_3241, w_239_3247, w_239_3257, w_239_3272, w_239_3280, w_239_3286, w_239_3299, w_239_3309, w_239_3317, w_239_3318, w_239_3322, w_239_3328, w_239_3332, w_239_3360, w_239_3361, w_239_3377, w_239_3378, w_239_3397, w_239_3407, w_239_3409, w_239_3414, w_239_3424, w_239_3426, w_239_3427, w_239_3429, w_239_3434, w_239_3444, w_239_3445, w_239_3450, w_239_3455, w_239_3456, w_239_3463, w_239_3470, w_239_3473, w_239_3478, w_239_3483, w_239_3487, w_239_3492, w_239_3506, w_239_3514, w_239_3521, w_239_3535, w_239_3547, w_239_3549, w_239_3552, w_239_3559, w_239_3563, w_239_3568, w_239_3569, w_239_3575, w_239_3576, w_239_3578, w_239_3595, w_239_3598, w_239_3603, w_239_3611, w_239_3620, w_239_3630, w_239_3649, w_239_3654, w_239_3670, w_239_3671;
  wire w_240_003, w_240_014, w_240_017, w_240_018, w_240_025, w_240_026, w_240_027, w_240_029, w_240_051, w_240_053, w_240_054, w_240_077, w_240_080, w_240_083, w_240_086, w_240_091, w_240_094, w_240_112, w_240_128, w_240_131, w_240_136, w_240_139, w_240_145, w_240_152, w_240_161, w_240_162, w_240_165, w_240_166, w_240_169, w_240_170, w_240_173, w_240_174, w_240_176, w_240_178, w_240_181, w_240_187, w_240_191, w_240_198, w_240_199, w_240_203, w_240_209, w_240_218, w_240_219, w_240_231, w_240_232, w_240_233, w_240_236, w_240_257, w_240_258, w_240_268, w_240_269, w_240_289, w_240_292, w_240_293, w_240_295, w_240_297, w_240_304, w_240_317, w_240_323, w_240_328, w_240_332, w_240_358, w_240_365, w_240_367, w_240_368, w_240_376, w_240_381, w_240_386, w_240_396, w_240_398, w_240_400, w_240_406, w_240_410, w_240_428, w_240_438, w_240_449, w_240_459, w_240_461, w_240_464, w_240_473, w_240_488, w_240_491, w_240_500, w_240_501, w_240_502, w_240_505, w_240_508, w_240_515, w_240_526, w_240_532, w_240_534, w_240_536, w_240_537, w_240_543, w_240_564, w_240_569, w_240_571, w_240_575, w_240_583, w_240_591, w_240_593, w_240_596, w_240_601, w_240_613, w_240_614, w_240_616, w_240_621, w_240_622, w_240_625, w_240_629, w_240_631, w_240_636, w_240_652, w_240_656, w_240_658, w_240_659, w_240_676, w_240_689, w_240_696, w_240_698, w_240_726, w_240_738, w_240_749, w_240_776, w_240_777, w_240_780, w_240_795, w_240_814, w_240_853, w_240_856, w_240_862, w_240_883, w_240_896, w_240_897, w_240_900, w_240_924, w_240_940, w_240_946, w_240_947, w_240_967, w_240_972, w_240_981, w_240_989, w_240_1003, w_240_1008, w_240_1011, w_240_1034, w_240_1035, w_240_1038, w_240_1043, w_240_1049, w_240_1057, w_240_1075, w_240_1085, w_240_1086, w_240_1114, w_240_1120, w_240_1127, w_240_1143, w_240_1148, w_240_1150, w_240_1162, w_240_1189, w_240_1201, w_240_1202, w_240_1221, w_240_1224, w_240_1250, w_240_1264, w_240_1269, w_240_1272, w_240_1290, w_240_1291, w_240_1293, w_240_1313, w_240_1314, w_240_1349, w_240_1375, w_240_1388, w_240_1400, w_240_1410, w_240_1448, w_240_1451, w_240_1490, w_240_1507, w_240_1510, w_240_1512, w_240_1514, w_240_1515, w_240_1517, w_240_1524, w_240_1529, w_240_1530, w_240_1542, w_240_1552, w_240_1589, w_240_1606, w_240_1626, w_240_1631, w_240_1647, w_240_1661, w_240_1681, w_240_1688, w_240_1693, w_240_1708, w_240_1730, w_240_1735, w_240_1754, w_240_1757, w_240_1760, w_240_1762, w_240_1771, w_240_1773, w_240_1775, w_240_1799, w_240_1800, w_240_1835, w_240_1860, w_240_1873, w_240_1877, w_240_1897, w_240_1904, w_240_1914, w_240_1933, w_240_1935, w_240_1943, w_240_1957, w_240_1970, w_240_1971, w_240_1990, w_240_1993, w_240_2002, w_240_2004, w_240_2006, w_240_2026, w_240_2028, w_240_2039, w_240_2046, w_240_2047, w_240_2059, w_240_2082, w_240_2089, w_240_2093, w_240_2097, w_240_2105, w_240_2116, w_240_2143, w_240_2157, w_240_2161, w_240_2165, w_240_2189, w_240_2200, w_240_2235, w_240_2251, w_240_2257, w_240_2262, w_240_2275, w_240_2285, w_240_2286, w_240_2293, w_240_2303, w_240_2338, w_240_2341, w_240_2349, w_240_2354, w_240_2357, w_240_2358, w_240_2362, w_240_2390, w_240_2401, w_240_2426, w_240_2427, w_240_2442, w_240_2447, w_240_2463, w_240_2472, w_240_2485, w_240_2495, w_240_2504, w_240_2505, w_240_2516, w_240_2523, w_240_2527, w_240_2538, w_240_2544, w_240_2548, w_240_2553, w_240_2575, w_240_2586, w_240_2630, w_240_2649, w_240_2665, w_240_2677, w_240_2682, w_240_2683, w_240_2694, w_240_2697, w_240_2700, w_240_2705, w_240_2706, w_240_2729, w_240_2740, w_240_2743, w_240_2746, w_240_2758, w_240_2786, w_240_2795, w_240_2796, w_240_2811, w_240_2826, w_240_2839, w_240_2846, w_240_2848, w_240_2849, w_240_2850, w_240_2858, w_240_2864, w_240_2865, w_240_2877, w_240_2905, w_240_2908, w_240_2926, w_240_2946, w_240_2951, w_240_2956, w_240_2962, w_240_2974, w_240_2978, w_240_2982, w_240_2985, w_240_2986, w_240_3000, w_240_3016, w_240_3028, w_240_3035, w_240_3038, w_240_3045, w_240_3048, w_240_3050, w_240_3052, w_240_3056, w_240_3061, w_240_3068, w_240_3071, w_240_3073, w_240_3077, w_240_3090, w_240_3093, w_240_3098, w_240_3116, w_240_3121, w_240_3122, w_240_3125, w_240_3126, w_240_3131, w_240_3137, w_240_3139, w_240_3140, w_240_3165, w_240_3183, w_240_3189, w_240_3193, w_240_3208, w_240_3210, w_240_3230, w_240_3256, w_240_3283, w_240_3295, w_240_3299, w_240_3300, w_240_3304, w_240_3314, w_240_3322, w_240_3376, w_240_3384, w_240_3387, w_240_3396, w_240_3404, w_240_3431, w_240_3439, w_240_3446, w_240_3468, w_240_3471, w_240_3473, w_240_3487, w_240_3507, w_240_3511, w_240_3516, w_240_3518, w_240_3529, w_240_3536, w_240_3562, w_240_3563, w_240_3573, w_240_3600, w_240_3613, w_240_3618, w_240_3625, w_240_3633, w_240_3635, w_240_3674, w_240_3684, w_240_3688, w_240_3696, w_240_3704, w_240_3712, w_240_3734, w_240_3735, w_240_3738, w_240_3773, w_240_3786, w_240_3787, w_240_3813, w_240_3820, w_240_3831, w_240_3836, w_240_3875, w_240_3883, w_240_3905, w_240_3911, w_240_3916, w_240_3917, w_240_3918, w_240_3920, w_240_3950, w_240_3966, w_240_3974, w_240_3981, w_240_4021, w_240_4037, w_240_4058, w_240_4084, w_240_4085, w_240_4087, w_240_4088, w_240_4103, w_240_4112, w_240_4125, w_240_4127, w_240_4129, w_240_4147, w_240_4151, w_240_4161, w_240_4167, w_240_4170, w_240_4184, w_240_4195, w_240_4206, w_240_4208, w_240_4209, w_240_4213, w_240_4221, w_240_4224, w_240_4247, w_240_4266, w_240_4272, w_240_4275, w_240_4293, w_240_4294, w_240_4295, w_240_4296, w_240_4297, w_240_4298, w_240_4299, w_240_4300, w_240_4301, w_240_4302, w_240_4306, w_240_4307, w_240_4308, w_240_4309, w_240_4310, w_240_4311, w_240_4312, w_240_4313, w_240_4314, w_240_4315, w_240_4316, w_240_4317, w_240_4319;
  wire w_241_006, w_241_011, w_241_033, w_241_035, w_241_038, w_241_041, w_241_054, w_241_055, w_241_061, w_241_069, w_241_071, w_241_073, w_241_077, w_241_078, w_241_082, w_241_087, w_241_091, w_241_107, w_241_111, w_241_119, w_241_120, w_241_123, w_241_127, w_241_137, w_241_143, w_241_145, w_241_146, w_241_153, w_241_154, w_241_164, w_241_167, w_241_172, w_241_176, w_241_182, w_241_187, w_241_197, w_241_198, w_241_200, w_241_208, w_241_213, w_241_229, w_241_242, w_241_245, w_241_250, w_241_252, w_241_258, w_241_260, w_241_261, w_241_262, w_241_277, w_241_278, w_241_279, w_241_283, w_241_297, w_241_301, w_241_302, w_241_303, w_241_306, w_241_308, w_241_311, w_241_318, w_241_320, w_241_325, w_241_327, w_241_335, w_241_336, w_241_339, w_241_347, w_241_352, w_241_359, w_241_369, w_241_381, w_241_395, w_241_400, w_241_401, w_241_403, w_241_426, w_241_428, w_241_431, w_241_434, w_241_438, w_241_442, w_241_444, w_241_450, w_241_451, w_241_456, w_241_458, w_241_461, w_241_464, w_241_469, w_241_478, w_241_489, w_241_496, w_241_497, w_241_498, w_241_503, w_241_509, w_241_511, w_241_521, w_241_528, w_241_545, w_241_546, w_241_553, w_241_555, w_241_558, w_241_560, w_241_569, w_241_577, w_241_581, w_241_587, w_241_596, w_241_610, w_241_621, w_241_635, w_241_653, w_241_657, w_241_660, w_241_663, w_241_665, w_241_666, w_241_667, w_241_671, w_241_679, w_241_682, w_241_683, w_241_685, w_241_688, w_241_697, w_241_702, w_241_704, w_241_709, w_241_721, w_241_722, w_241_728, w_241_730, w_241_744, w_241_747, w_241_753, w_241_754, w_241_756, w_241_762, w_241_773, w_241_776, w_241_777, w_241_781, w_241_786, w_241_789, w_241_790, w_241_800, w_241_805, w_241_808, w_241_815, w_241_820, w_241_835, w_241_837, w_241_839, w_241_843, w_241_849, w_241_851, w_241_852, w_241_855, w_241_861, w_241_869, w_241_875, w_241_880, w_241_895, w_241_896, w_241_901, w_241_908, w_241_909, w_241_914, w_241_915, w_241_926, w_241_939, w_241_943, w_241_947, w_241_951, w_241_955, w_241_971, w_241_976, w_241_977, w_241_981, w_241_989, w_241_994, w_241_996, w_241_999, w_241_1002, w_241_1006, w_241_1007, w_241_1008, w_241_1009, w_241_1010, w_241_1016, w_241_1017, w_241_1024, w_241_1034, w_241_1035, w_241_1040, w_241_1044, w_241_1051, w_241_1055, w_241_1056, w_241_1061, w_241_1062, w_241_1064, w_241_1067, w_241_1071, w_241_1079, w_241_1081, w_241_1106, w_241_1107, w_241_1109, w_241_1110, w_241_1111, w_241_1119, w_241_1126, w_241_1130, w_241_1131, w_241_1135, w_241_1136, w_241_1138, w_241_1143, w_241_1145, w_241_1147, w_241_1155, w_241_1165, w_241_1170, w_241_1174, w_241_1177, w_241_1184, w_241_1186, w_241_1187, w_241_1189, w_241_1195, w_241_1199, w_241_1204, w_241_1213, w_241_1215, w_241_1222, w_241_1229, w_241_1230, w_241_1231, w_241_1234, w_241_1242, w_241_1244, w_241_1252, w_241_1258, w_241_1266, w_241_1268, w_241_1271, w_241_1277, w_241_1279, w_241_1282, w_241_1284, w_241_1289, w_241_1290, w_241_1291, w_241_1298, w_241_1299, w_241_1315, w_241_1319, w_241_1320, w_241_1326, w_241_1336, w_241_1338, w_241_1339, w_241_1346, w_241_1351, w_241_1354, w_241_1361, w_241_1366, w_241_1368, w_241_1373, w_241_1379, w_241_1387, w_241_1400, w_241_1418, w_241_1429, w_241_1431, w_241_1433, w_241_1435, w_241_1439, w_241_1451, w_241_1465, w_241_1469, w_241_1479, w_241_1482, w_241_1485, w_241_1486, w_241_1499, w_241_1501, w_241_1507, w_241_1508, w_241_1518, w_241_1521, w_241_1524, w_241_1532, w_241_1533, w_241_1538, w_241_1543, w_241_1548, w_241_1556, w_241_1557, w_241_1558, w_241_1575, w_241_1581, w_241_1586, w_241_1601, w_241_1602, w_241_1604, w_241_1607, w_241_1608, w_241_1628, w_241_1629, w_241_1648, w_241_1651, w_241_1655, w_241_1665, w_241_1678, w_241_1679, w_241_1680, w_241_1681, w_241_1684, w_241_1695, w_241_1706, w_241_1707, w_241_1709, w_241_1728, w_241_1742, w_241_1745, w_241_1754, w_241_1759, w_241_1760, w_241_1763, w_241_1772, w_241_1779, w_241_1782, w_241_1788, w_241_1795, w_241_1798, w_241_1800, w_241_1801, w_241_1812, w_241_1823, w_241_1824, w_241_1828, w_241_1830, w_241_1831, w_241_1846, w_241_1855, w_241_1862, w_241_1863, w_241_1872, w_241_1888, w_241_1899, w_241_1906, w_241_1925, w_241_1933, w_241_1935, w_241_1941, w_241_1946, w_241_1948, w_241_1953, w_241_1963, w_241_1967, w_241_1968, w_241_1974, w_241_1975, w_241_1987, w_241_2007, w_241_2012, w_241_2017, w_241_2021, w_241_2025, w_241_2034, w_241_2037, w_241_2050, w_241_2066, w_241_2079, w_241_2092, w_241_2093, w_241_2114, w_241_2115, w_241_2116, w_241_2120, w_241_2130, w_241_2138, w_241_2142, w_241_2152, w_241_2155, w_241_2170, w_241_2174, w_241_2182, w_241_2190, w_241_2194, w_241_2203, w_241_2225, w_241_2230, w_241_2235, w_241_2246, w_241_2255, w_241_2268, w_241_2271, w_241_2273, w_241_2275, w_241_2289, w_241_2292, w_241_2298, w_241_2327, w_241_2337, w_241_2376, w_241_2383, w_241_2387, w_241_2400, w_241_2431, w_241_2432, w_241_2434, w_241_2448, w_241_2449, w_241_2466, w_241_2467, w_241_2474, w_241_2480, w_241_2483, w_241_2487, w_241_2489, w_241_2490, w_241_2492, w_241_2496, w_241_2529, w_241_2542, w_241_2554, w_241_2597, w_241_2599, w_241_2610, w_241_2613, w_241_2625, w_241_2629, w_241_2641, w_241_2645, w_241_2695, w_241_2701, w_241_2709, w_241_2716, w_241_2732, w_241_2749, w_241_2761, w_241_2765, w_241_2769, w_241_2778, w_241_2782, w_241_2796, w_241_2801, w_241_2803, w_241_2812, w_241_2817, w_241_2820, w_241_2825, w_241_2833, w_241_2841, w_241_2853, w_241_2858, w_241_2870, w_241_2874, w_241_2883, w_241_2892, w_241_2915, w_241_2963, w_241_2967, w_241_2970, w_241_2975, w_241_2989, w_241_2997, w_241_2999, w_241_3014, w_241_3015, w_241_3023, w_241_3033, w_241_3050, w_241_3066, w_241_3067, w_241_3070, w_241_3071, w_241_3102, w_241_3121, w_241_3126, w_241_3130, w_241_3131, w_241_3132, w_241_3133, w_241_3134, w_241_3135, w_241_3136, w_241_3137, w_241_3141, w_241_3142, w_241_3143, w_241_3144, w_241_3145, w_241_3146, w_241_3147, w_241_3148, w_241_3149, w_241_3150, w_241_3151, w_241_3152, w_241_3154;
  wire w_242_005, w_242_016, w_242_024, w_242_036, w_242_042, w_242_043, w_242_044, w_242_049, w_242_050, w_242_054, w_242_058, w_242_069, w_242_073, w_242_074, w_242_076, w_242_089, w_242_090, w_242_091, w_242_094, w_242_099, w_242_103, w_242_119, w_242_122, w_242_124, w_242_126, w_242_129, w_242_132, w_242_134, w_242_135, w_242_142, w_242_145, w_242_151, w_242_155, w_242_159, w_242_161, w_242_165, w_242_172, w_242_176, w_242_183, w_242_188, w_242_189, w_242_192, w_242_194, w_242_198, w_242_201, w_242_208, w_242_210, w_242_211, w_242_212, w_242_226, w_242_227, w_242_236, w_242_253, w_242_254, w_242_255, w_242_258, w_242_260, w_242_262, w_242_267, w_242_275, w_242_278, w_242_284, w_242_286, w_242_303, w_242_308, w_242_312, w_242_313, w_242_315, w_242_323, w_242_330, w_242_334, w_242_338, w_242_351, w_242_364, w_242_365, w_242_369, w_242_377, w_242_378, w_242_379, w_242_382, w_242_387, w_242_397, w_242_404, w_242_406, w_242_416, w_242_418, w_242_423, w_242_428, w_242_429, w_242_432, w_242_454, w_242_456, w_242_462, w_242_470, w_242_471, w_242_472, w_242_485, w_242_489, w_242_491, w_242_499, w_242_502, w_242_505, w_242_509, w_242_510, w_242_512, w_242_519, w_242_524, w_242_545, w_242_550, w_242_552, w_242_555, w_242_559, w_242_560, w_242_566, w_242_586, w_242_592, w_242_595, w_242_607, w_242_619, w_242_621, w_242_623, w_242_632, w_242_633, w_242_636, w_242_647, w_242_648, w_242_652, w_242_658, w_242_667, w_242_669, w_242_673, w_242_681, w_242_686, w_242_688, w_242_698, w_242_699, w_242_700, w_242_720, w_242_724, w_242_740, w_242_743, w_242_746, w_242_747, w_242_749, w_242_754, w_242_761, w_242_770, w_242_775, w_242_778, w_242_786, w_242_813, w_242_819, w_242_825, w_242_832, w_242_833, w_242_837, w_242_838, w_242_850, w_242_854, w_242_866, w_242_874, w_242_876, w_242_880, w_242_895, w_242_898, w_242_904, w_242_908, w_242_911, w_242_912, w_242_915, w_242_917, w_242_918, w_242_920, w_242_925, w_242_932, w_242_941, w_242_942, w_242_944, w_242_959, w_242_968, w_242_977, w_242_979, w_242_982, w_242_984, w_242_985, w_242_992, w_242_996, w_242_1001, w_242_1009, w_242_1010, w_242_1039, w_242_1043, w_242_1045, w_242_1053, w_242_1058, w_242_1063, w_242_1067, w_242_1068, w_242_1072, w_242_1074, w_242_1094, w_242_1095, w_242_1096, w_242_1106, w_242_1109, w_242_1111, w_242_1117, w_242_1119, w_242_1121, w_242_1122, w_242_1123, w_242_1133, w_242_1135, w_242_1136, w_242_1141, w_242_1146, w_242_1147, w_242_1148, w_242_1149, w_242_1152, w_242_1160, w_242_1165, w_242_1171, w_242_1180, w_242_1182, w_242_1185, w_242_1187, w_242_1188, w_242_1194, w_242_1196, w_242_1197, w_242_1212, w_242_1214, w_242_1218, w_242_1224, w_242_1225, w_242_1226, w_242_1228, w_242_1230, w_242_1232, w_242_1234, w_242_1235, w_242_1252, w_242_1267, w_242_1268, w_242_1270, w_242_1272, w_242_1282, w_242_1290, w_242_1323, w_242_1352, w_242_1353, w_242_1365, w_242_1366, w_242_1394, w_242_1398, w_242_1409, w_242_1463, w_242_1468, w_242_1477, w_242_1482, w_242_1483, w_242_1484, w_242_1495, w_242_1498, w_242_1506, w_242_1516, w_242_1519, w_242_1528, w_242_1565, w_242_1578, w_242_1586, w_242_1589, w_242_1595, w_242_1610, w_242_1621, w_242_1630, w_242_1633, w_242_1640, w_242_1655, w_242_1662, w_242_1671, w_242_1672, w_242_1687, w_242_1698, w_242_1702, w_242_1711, w_242_1731, w_242_1737, w_242_1741, w_242_1751, w_242_1768, w_242_1784, w_242_1796, w_242_1821, w_242_1822, w_242_1823, w_242_1849, w_242_1850, w_242_1862, w_242_1863, w_242_1881, w_242_1888, w_242_1894, w_242_1896, w_242_1907, w_242_1944, w_242_1956, w_242_1965, w_242_1968, w_242_1970, w_242_1975, w_242_1977, w_242_1997, w_242_2008, w_242_2027, w_242_2038, w_242_2057, w_242_2065, w_242_2081, w_242_2092, w_242_2098, w_242_2100, w_242_2101, w_242_2105, w_242_2106, w_242_2108, w_242_2118, w_242_2151, w_242_2157, w_242_2162, w_242_2167, w_242_2170, w_242_2171, w_242_2177, w_242_2193, w_242_2219, w_242_2230, w_242_2247, w_242_2248, w_242_2274, w_242_2276, w_242_2280, w_242_2287, w_242_2288, w_242_2292, w_242_2298, w_242_2317, w_242_2318, w_242_2337, w_242_2346, w_242_2358, w_242_2363, w_242_2366, w_242_2367, w_242_2374, w_242_2375, w_242_2378, w_242_2390, w_242_2440, w_242_2453, w_242_2456, w_242_2458, w_242_2468, w_242_2474, w_242_2494, w_242_2512, w_242_2514, w_242_2517, w_242_2528, w_242_2534, w_242_2535, w_242_2562, w_242_2574, w_242_2590, w_242_2595, w_242_2598, w_242_2600, w_242_2612, w_242_2615, w_242_2621, w_242_2629, w_242_2632, w_242_2646, w_242_2674, w_242_2699, w_242_2703, w_242_2704, w_242_2711, w_242_2718, w_242_2723, w_242_2731, w_242_2733, w_242_2753, w_242_2756, w_242_2774, w_242_2786, w_242_2804, w_242_2819, w_242_2828, w_242_2830, w_242_2836, w_242_2843, w_242_2855, w_242_2859, w_242_2862, w_242_2863, w_242_2872, w_242_2874, w_242_2876, w_242_2877, w_242_2878, w_242_2879, w_242_2894, w_242_2936, w_242_2937, w_242_2943, w_242_2945, w_242_2958, w_242_2960, w_242_2967, w_242_2974, w_242_2984, w_242_2992, w_242_2995, w_242_2997, w_242_3002, w_242_3004, w_242_3011, w_242_3017, w_242_3019, w_242_3040, w_242_3055, w_242_3081, w_242_3089, w_242_3105, w_242_3106, w_242_3117, w_242_3150, w_242_3165, w_242_3182, w_242_3195, w_242_3220, w_242_3223, w_242_3226, w_242_3228, w_242_3230, w_242_3236, w_242_3248, w_242_3253, w_242_3258, w_242_3270, w_242_3281, w_242_3296, w_242_3300, w_242_3323, w_242_3329, w_242_3339, w_242_3349, w_242_3373, w_242_3379, w_242_3394, w_242_3403, w_242_3436, w_242_3441, w_242_3451, w_242_3454, w_242_3475, w_242_3482, w_242_3493, w_242_3496, w_242_3504, w_242_3513, w_242_3524, w_242_3537, w_242_3549, w_242_3550, w_242_3561, w_242_3564, w_242_3570, w_242_3587, w_242_3614, w_242_3618, w_242_3631, w_242_3632, w_242_3636, w_242_3644, w_242_3649, w_242_3663, w_242_3668, w_242_3674, w_242_3675, w_242_3681, w_242_3683, w_242_3686, w_242_3691, w_242_3707, w_242_3713, w_242_3714, w_242_3717, w_242_3727, w_242_3729, w_242_3736, w_242_3740, w_242_3742;
  wire w_243_003, w_243_004, w_243_005, w_243_008, w_243_013, w_243_015, w_243_022, w_243_028, w_243_052, w_243_054, w_243_055, w_243_057, w_243_059, w_243_063, w_243_065, w_243_067, w_243_092, w_243_094, w_243_096, w_243_098, w_243_101, w_243_104, w_243_108, w_243_110, w_243_114, w_243_115, w_243_124, w_243_136, w_243_140, w_243_143, w_243_144, w_243_145, w_243_149, w_243_161, w_243_167, w_243_169, w_243_184, w_243_192, w_243_194, w_243_195, w_243_213, w_243_214, w_243_223, w_243_224, w_243_227, w_243_228, w_243_233, w_243_236, w_243_242, w_243_250, w_243_257, w_243_265, w_243_270, w_243_274, w_243_277, w_243_283, w_243_284, w_243_295, w_243_296, w_243_300, w_243_305, w_243_307, w_243_308, w_243_311, w_243_315, w_243_317, w_243_325, w_243_327, w_243_332, w_243_342, w_243_346, w_243_347, w_243_349, w_243_352, w_243_357, w_243_359, w_243_374, w_243_376, w_243_377, w_243_381, w_243_382, w_243_387, w_243_388, w_243_400, w_243_413, w_243_417, w_243_418, w_243_422, w_243_429, w_243_434, w_243_440, w_243_447, w_243_449, w_243_456, w_243_458, w_243_463, w_243_464, w_243_477, w_243_487, w_243_490, w_243_497, w_243_505, w_243_510, w_243_534, w_243_537, w_243_546, w_243_553, w_243_561, w_243_566, w_243_567, w_243_570, w_243_577, w_243_584, w_243_593, w_243_594, w_243_602, w_243_603, w_243_604, w_243_609, w_243_610, w_243_612, w_243_616, w_243_620, w_243_622, w_243_623, w_243_626, w_243_643, w_243_645, w_243_650, w_243_655, w_243_656, w_243_660, w_243_665, w_243_667, w_243_668, w_243_673, w_243_684, w_243_687, w_243_702, w_243_706, w_243_714, w_243_715, w_243_722, w_243_731, w_243_733, w_243_745, w_243_751, w_243_766, w_243_767, w_243_768, w_243_777, w_243_784, w_243_785, w_243_788, w_243_789, w_243_791, w_243_792, w_243_793, w_243_798, w_243_803, w_243_821, w_243_826, w_243_830, w_243_838, w_243_842, w_243_843, w_243_845, w_243_847, w_243_851, w_243_852, w_243_858, w_243_859, w_243_863, w_243_865, w_243_878, w_243_887, w_243_892, w_243_898, w_243_904, w_243_908, w_243_917, w_243_940, w_243_942, w_243_943, w_243_955, w_243_959, w_243_960, w_243_967, w_243_982, w_243_989, w_243_999, w_243_1015, w_243_1017, w_243_1019, w_243_1028, w_243_1029, w_243_1030, w_243_1033, w_243_1036, w_243_1043, w_243_1044, w_243_1053, w_243_1060, w_243_1085, w_243_1086, w_243_1091, w_243_1092, w_243_1100, w_243_1101, w_243_1114, w_243_1128, w_243_1142, w_243_1161, w_243_1165, w_243_1177, w_243_1178, w_243_1184, w_243_1193, w_243_1211, w_243_1226, w_243_1227, w_243_1234, w_243_1235, w_243_1240, w_243_1241, w_243_1245, w_243_1251, w_243_1257, w_243_1258, w_243_1270, w_243_1284, w_243_1285, w_243_1286, w_243_1289, w_243_1292, w_243_1294, w_243_1295, w_243_1297, w_243_1301, w_243_1303, w_243_1305, w_243_1321, w_243_1326, w_243_1330, w_243_1332, w_243_1333, w_243_1340, w_243_1344, w_243_1354, w_243_1356, w_243_1358, w_243_1366, w_243_1369, w_243_1376, w_243_1381, w_243_1382, w_243_1394, w_243_1396, w_243_1405, w_243_1413, w_243_1416, w_243_1418, w_243_1421, w_243_1423, w_243_1424, w_243_1427, w_243_1429, w_243_1432, w_243_1434, w_243_1443, w_243_1457, w_243_1460, w_243_1477, w_243_1479, w_243_1489, w_243_1495, w_243_1498, w_243_1502, w_243_1504, w_243_1515, w_243_1521, w_243_1524, w_243_1528, w_243_1531, w_243_1535, w_243_1551, w_243_1557, w_243_1563, w_243_1566, w_243_1567, w_243_1569, w_243_1574, w_243_1579, w_243_1584, w_243_1588, w_243_1591, w_243_1594, w_243_1606, w_243_1609, w_243_1611, w_243_1637, w_243_1641, w_243_1650, w_243_1659, w_243_1665, w_243_1670, w_243_1678, w_243_1696, w_243_1711, w_243_1725, w_243_1728, w_243_1732, w_243_1736, w_243_1770, w_243_1783, w_243_1787, w_243_1796, w_243_1801, w_243_1820, w_243_1823, w_243_1830, w_243_1835, w_243_1842, w_243_1892, w_243_1894, w_243_1898, w_243_1904, w_243_1907, w_243_1918, w_243_1922, w_243_1940, w_243_1975, w_243_1987, w_243_1990, w_243_2001, w_243_2010, w_243_2011, w_243_2034, w_243_2045, w_243_2046, w_243_2058, w_243_2066, w_243_2135, w_243_2137, w_243_2168, w_243_2183, w_243_2195, w_243_2205, w_243_2218, w_243_2220, w_243_2226, w_243_2235, w_243_2236, w_243_2239, w_243_2257, w_243_2260, w_243_2270, w_243_2320, w_243_2325, w_243_2330, w_243_2341, w_243_2345, w_243_2356, w_243_2369, w_243_2405, w_243_2408, w_243_2420, w_243_2429, w_243_2432, w_243_2447, w_243_2449, w_243_2473, w_243_2499, w_243_2518, w_243_2527, w_243_2532, w_243_2538, w_243_2556, w_243_2560, w_243_2561, w_243_2583, w_243_2589, w_243_2590, w_243_2611, w_243_2625, w_243_2626, w_243_2657, w_243_2660, w_243_2669, w_243_2680, w_243_2694, w_243_2724, w_243_2736, w_243_2739, w_243_2751, w_243_2791, w_243_2811, w_243_2815, w_243_2818, w_243_2819, w_243_2822, w_243_2826, w_243_2846, w_243_2865, w_243_2876, w_243_2891, w_243_2900, w_243_2903, w_243_2945, w_243_2947, w_243_2968, w_243_2974, w_243_2985, w_243_2995, w_243_3000, w_243_3007, w_243_3011, w_243_3012, w_243_3016, w_243_3018, w_243_3019, w_243_3024, w_243_3027, w_243_3037, w_243_3042, w_243_3048, w_243_3049, w_243_3066, w_243_3068, w_243_3073, w_243_3075, w_243_3086, w_243_3100, w_243_3108, w_243_3114, w_243_3134, w_243_3149, w_243_3166, w_243_3188, w_243_3194, w_243_3210, w_243_3218, w_243_3220, w_243_3221, w_243_3233, w_243_3252, w_243_3257, w_243_3264, w_243_3268, w_243_3280, w_243_3306, w_243_3315, w_243_3323, w_243_3328, w_243_3350;
  wire w_244_000, w_244_002, w_244_006, w_244_017, w_244_037, w_244_038, w_244_039, w_244_047, w_244_049, w_244_050, w_244_052, w_244_054, w_244_060, w_244_065, w_244_067, w_244_069, w_244_073, w_244_076, w_244_085, w_244_088, w_244_098, w_244_100, w_244_101, w_244_104, w_244_110, w_244_125, w_244_135, w_244_145, w_244_147, w_244_150, w_244_157, w_244_159, w_244_165, w_244_166, w_244_171, w_244_174, w_244_189, w_244_196, w_244_199, w_244_201, w_244_206, w_244_211, w_244_214, w_244_219, w_244_226, w_244_229, w_244_236, w_244_247, w_244_250, w_244_251, w_244_252, w_244_256, w_244_261, w_244_262, w_244_267, w_244_274, w_244_276, w_244_281, w_244_282, w_244_283, w_244_300, w_244_311, w_244_313, w_244_321, w_244_323, w_244_327, w_244_331, w_244_338, w_244_340, w_244_348, w_244_349, w_244_351, w_244_354, w_244_355, w_244_359, w_244_361, w_244_363, w_244_371, w_244_379, w_244_385, w_244_390, w_244_391, w_244_392, w_244_393, w_244_403, w_244_409, w_244_419, w_244_420, w_244_425, w_244_435, w_244_436, w_244_439, w_244_440, w_244_448, w_244_459, w_244_460, w_244_482, w_244_486, w_244_508, w_244_510, w_244_511, w_244_513, w_244_519, w_244_551, w_244_555, w_244_556, w_244_563, w_244_564, w_244_567, w_244_568, w_244_576, w_244_586, w_244_592, w_244_611, w_244_625, w_244_630, w_244_633, w_244_636, w_244_637, w_244_648, w_244_654, w_244_671, w_244_673, w_244_678, w_244_680, w_244_688, w_244_698, w_244_703, w_244_723, w_244_734, w_244_736, w_244_743, w_244_750, w_244_752, w_244_760, w_244_762, w_244_772, w_244_793, w_244_795, w_244_802, w_244_810, w_244_830, w_244_833, w_244_840, w_244_845, w_244_848, w_244_850, w_244_861, w_244_872, w_244_875, w_244_877, w_244_881, w_244_882, w_244_886, w_244_887, w_244_890, w_244_902, w_244_903, w_244_905, w_244_907, w_244_912, w_244_923, w_244_924, w_244_941, w_244_957, w_244_962, w_244_970, w_244_971, w_244_973, w_244_976, w_244_978, w_244_982, w_244_985, w_244_994, w_244_996, w_244_1001, w_244_1007, w_244_1010, w_244_1018, w_244_1023, w_244_1026, w_244_1027, w_244_1028, w_244_1036, w_244_1037, w_244_1044, w_244_1055, w_244_1056, w_244_1058, w_244_1063, w_244_1069, w_244_1070, w_244_1071, w_244_1081, w_244_1087, w_244_1089, w_244_1090, w_244_1094, w_244_1107, w_244_1111, w_244_1112, w_244_1113, w_244_1114, w_244_1119, w_244_1129, w_244_1131, w_244_1133, w_244_1160, w_244_1166, w_244_1167, w_244_1169, w_244_1174, w_244_1178, w_244_1195, w_244_1205, w_244_1215, w_244_1232, w_244_1233, w_244_1240, w_244_1242, w_244_1243, w_244_1244, w_244_1256, w_244_1260, w_244_1265, w_244_1271, w_244_1280, w_244_1292, w_244_1295, w_244_1297, w_244_1310, w_244_1313, w_244_1316, w_244_1323, w_244_1334, w_244_1335, w_244_1336, w_244_1338, w_244_1349, w_244_1362, w_244_1366, w_244_1370, w_244_1374, w_244_1375, w_244_1389, w_244_1403, w_244_1405, w_244_1417, w_244_1418, w_244_1435, w_244_1441, w_244_1442, w_244_1457, w_244_1458, w_244_1459, w_244_1460, w_244_1463, w_244_1482, w_244_1485, w_244_1493, w_244_1496, w_244_1498, w_244_1512, w_244_1521, w_244_1525, w_244_1541, w_244_1544, w_244_1549, w_244_1552, w_244_1561, w_244_1592, w_244_1593, w_244_1601, w_244_1602, w_244_1610, w_244_1616, w_244_1621, w_244_1628, w_244_1629, w_244_1640, w_244_1653, w_244_1662, w_244_1665, w_244_1670, w_244_1673, w_244_1680, w_244_1690, w_244_1695, w_244_1700, w_244_1705, w_244_1711, w_244_1722, w_244_1727, w_244_1730, w_244_1732, w_244_1735, w_244_1740, w_244_1744, w_244_1746, w_244_1765, w_244_1777, w_244_1783, w_244_1786, w_244_1789, w_244_1799, w_244_1803, w_244_1817, w_244_1821, w_244_1823, w_244_1825, w_244_1837, w_244_1840, w_244_1845, w_244_1848, w_244_1863, w_244_1864, w_244_1867, w_244_1872, w_244_1873, w_244_1889, w_244_1890, w_244_1894, w_244_1895, w_244_1899, w_244_1900, w_244_1909, w_244_1913, w_244_1914, w_244_1915, w_244_1921, w_244_1923, w_244_1935, w_244_1940, w_244_1951, w_244_1952, w_244_1953, w_244_1960, w_244_1965, w_244_1966, w_244_1969, w_244_1975, w_244_1977, w_244_1981, w_244_1987, w_244_1993, w_244_2009, w_244_2010, w_244_2018, w_244_2020, w_244_2023, w_244_2024, w_244_2026, w_244_2028, w_244_2033, w_244_2041, w_244_2059, w_244_2063, w_244_2066, w_244_2079, w_244_2085, w_244_2094, w_244_2095, w_244_2112, w_244_2114, w_244_2126, w_244_2127, w_244_2135, w_244_2137, w_244_2150, w_244_2159, w_244_2167, w_244_2185, w_244_2192, w_244_2209, w_244_2210, w_244_2215, w_244_2217, w_244_2231, w_244_2252, w_244_2264, w_244_2265, w_244_2266, w_244_2270, w_244_2271, w_244_2277, w_244_2278, w_244_2283, w_244_2287, w_244_2289, w_244_2293, w_244_2297, w_244_2298, w_244_2301, w_244_2304, w_244_2314, w_244_2320, w_244_2323, w_244_2327, w_244_2339, w_244_2340, w_244_2346, w_244_2351, w_244_2355, w_244_2357, w_244_2361, w_244_2362, w_244_2369, w_244_2371, w_244_2384, w_244_2398, w_244_2402, w_244_2408, w_244_2409, w_244_2413, w_244_2419, w_244_2420, w_244_2423, w_244_2428, w_244_2429, w_244_2430, w_244_2442, w_244_2443, w_244_2450, w_244_2455, w_244_2485, w_244_2492, w_244_2499, w_244_2504;
  wire w_245_002, w_245_007, w_245_008, w_245_009, w_245_011, w_245_013, w_245_015, w_245_016, w_245_017, w_245_018, w_245_019, w_245_020, w_245_022, w_245_023, w_245_025, w_245_028, w_245_029, w_245_030, w_245_031, w_245_038, w_245_041, w_245_044, w_245_046, w_245_048, w_245_049, w_245_050, w_245_051, w_245_054, w_245_055, w_245_060, w_245_062, w_245_065, w_245_066, w_245_067, w_245_068, w_245_069, w_245_074, w_245_076, w_245_077, w_245_078, w_245_080, w_245_081, w_245_082, w_245_085, w_245_087, w_245_088, w_245_094, w_245_099, w_245_101, w_245_103, w_245_106, w_245_107, w_245_108, w_245_109, w_245_112, w_245_113, w_245_114, w_245_116, w_245_117, w_245_119, w_245_120, w_245_121, w_245_122, w_245_125, w_245_126, w_245_127, w_245_128, w_245_132, w_245_133, w_245_136, w_245_139, w_245_141, w_245_144, w_245_145, w_245_146, w_245_148, w_245_154, w_245_157, w_245_158, w_245_160, w_245_161, w_245_163, w_245_164, w_245_165, w_245_166, w_245_168, w_245_169, w_245_170, w_245_172, w_245_176, w_245_177, w_245_180, w_245_181, w_245_185, w_245_186, w_245_192, w_245_193, w_245_196, w_245_198, w_245_199, w_245_200, w_245_201, w_245_202, w_245_203, w_245_204, w_245_207, w_245_208, w_245_209, w_245_210, w_245_211, w_245_213, w_245_214, w_245_216, w_245_222, w_245_224, w_245_228, w_245_229, w_245_233, w_245_234, w_245_235, w_245_237, w_245_241, w_245_243, w_245_244, w_245_245, w_245_248, w_245_249, w_245_250, w_245_252, w_245_254, w_245_257, w_245_260, w_245_262, w_245_263, w_245_264, w_245_266, w_245_267, w_245_270, w_245_271, w_245_274, w_245_277, w_245_280, w_245_281, w_245_282, w_245_286, w_245_287, w_245_289, w_245_290, w_245_291, w_245_293, w_245_296, w_245_297, w_245_298, w_245_299, w_245_301, w_245_303, w_245_305, w_245_307, w_245_308, w_245_310, w_245_311, w_245_315, w_245_316, w_245_317, w_245_319, w_245_321, w_245_322, w_245_323, w_245_325, w_245_326, w_245_327, w_245_330, w_245_333, w_245_334, w_245_337, w_245_338, w_245_339, w_245_340, w_245_344, w_245_347, w_245_350, w_245_354, w_245_355, w_245_356, w_245_357, w_245_359, w_245_361, w_245_362, w_245_363, w_245_364, w_245_367, w_245_368, w_245_369, w_245_370, w_245_371, w_245_374, w_245_376, w_245_378, w_245_380, w_245_381, w_245_382, w_245_383, w_245_384, w_245_385, w_245_387, w_245_388, w_245_391, w_245_392, w_245_393, w_245_398, w_245_399, w_245_405, w_245_406, w_245_407, w_245_408, w_245_410, w_245_411, w_245_412, w_245_413, w_245_416, w_245_417, w_245_418, w_245_422, w_245_423, w_245_424, w_245_426, w_245_427, w_245_428, w_245_432, w_245_433, w_245_434, w_245_436, w_245_437, w_245_438, w_245_440, w_245_443, w_245_444, w_245_448, w_245_449, w_245_453, w_245_454, w_245_455, w_245_457, w_245_459, w_245_460, w_245_461, w_245_462, w_245_465, w_245_466, w_245_467, w_245_469, w_245_473, w_245_475, w_245_477, w_245_480, w_245_481, w_245_483, w_245_485, w_245_486, w_245_487, w_245_488, w_245_490, w_245_491, w_245_492, w_245_493, w_245_494, w_245_497, w_245_499, w_245_500, w_245_502, w_245_503, w_245_504, w_245_505, w_245_507, w_245_508, w_245_509, w_245_513, w_245_516, w_245_517, w_245_518, w_245_519, w_245_520, w_245_521, w_245_522, w_245_523, w_245_525, w_245_527, w_245_528, w_245_529, w_245_530, w_245_531, w_245_532, w_245_535, w_245_538, w_245_542, w_245_544, w_245_545, w_245_549, w_245_554, w_245_556, w_245_557, w_245_560, w_245_561, w_245_562, w_245_564, w_245_565, w_245_566, w_245_570, w_245_572, w_245_573, w_245_574, w_245_575, w_245_576, w_245_579, w_245_581, w_245_582, w_245_584, w_245_585, w_245_590, w_245_592, w_245_593, w_245_595, w_245_596, w_245_597, w_245_600, w_245_601, w_245_603, w_245_605, w_245_606, w_245_607, w_245_610, w_245_612, w_245_614, w_245_615, w_245_618, w_245_619, w_245_620, w_245_621, w_245_622, w_245_623;
  wire w_246_000, w_246_001, w_246_004, w_246_005, w_246_006, w_246_008, w_246_010, w_246_011, w_246_012, w_246_015, w_246_016, w_246_018, w_246_022, w_246_026, w_246_027, w_246_028, w_246_030, w_246_032, w_246_033, w_246_034, w_246_036, w_246_040, w_246_043, w_246_048, w_246_050, w_246_051, w_246_054, w_246_055, w_246_056, w_246_058, w_246_060, w_246_061, w_246_062, w_246_063, w_246_064, w_246_067, w_246_068, w_246_071, w_246_073, w_246_075, w_246_076, w_246_077, w_246_078, w_246_082, w_246_083, w_246_086, w_246_087, w_246_088, w_246_089, w_246_091, w_246_092, w_246_094, w_246_095, w_246_099, w_246_100, w_246_101, w_246_102, w_246_103, w_246_104, w_246_107, w_246_108, w_246_110, w_246_113, w_246_116, w_246_118, w_246_119, w_246_120, w_246_122, w_246_125, w_246_127, w_246_128, w_246_130, w_246_135, w_246_138, w_246_141, w_246_142, w_246_143, w_246_144, w_246_147, w_246_149, w_246_150, w_246_153, w_246_155, w_246_156, w_246_158, w_246_161, w_246_162, w_246_163, w_246_164, w_246_166, w_246_167, w_246_168, w_246_171, w_246_175, w_246_178, w_246_180, w_246_184, w_246_188, w_246_192, w_246_195, w_246_197, w_246_198, w_246_204, w_246_208, w_246_213, w_246_216, w_246_217, w_246_219, w_246_220, w_246_221, w_246_224, w_246_225, w_246_226, w_246_227, w_246_228, w_246_234, w_246_236, w_246_237, w_246_238, w_246_239, w_246_241, w_246_242, w_246_243, w_246_244, w_246_246, w_246_248, w_246_250, w_246_251, w_246_252, w_246_253, w_246_255, w_246_256, w_246_257, w_246_258, w_246_262, w_246_263, w_246_264, w_246_265, w_246_266, w_246_267, w_246_271, w_246_277, w_246_278, w_246_280, w_246_281, w_246_287, w_246_288, w_246_292, w_246_293, w_246_296, w_246_298, w_246_300, w_246_302, w_246_304, w_246_305, w_246_307, w_246_309, w_246_311, w_246_312, w_246_313, w_246_316, w_246_319, w_246_325, w_246_326, w_246_329, w_246_330, w_246_331, w_246_334, w_246_336, w_246_337, w_246_339, w_246_341, w_246_342, w_246_344, w_246_345, w_246_346, w_246_349, w_246_351, w_246_353, w_246_355, w_246_356, w_246_358, w_246_359, w_246_360, w_246_366, w_246_367, w_246_368, w_246_370, w_246_371, w_246_373, w_246_375, w_246_376, w_246_378, w_246_380, w_246_383, w_246_384, w_246_386, w_246_388, w_246_389, w_246_391, w_246_392, w_246_394, w_246_397, w_246_398, w_246_401, w_246_402, w_246_404, w_246_406, w_246_409, w_246_410, w_246_411, w_246_414, w_246_416, w_246_419, w_246_420, w_246_421, w_246_423, w_246_425, w_246_427, w_246_428, w_246_432, w_246_435, w_246_436, w_246_437, w_246_438, w_246_440, w_246_441, w_246_442, w_246_443, w_246_444, w_246_446, w_246_448, w_246_449, w_246_452, w_246_455, w_246_456, w_246_459, w_246_462, w_246_463, w_246_464, w_246_465, w_246_468, w_246_470, w_246_471, w_246_473, w_246_474, w_246_475, w_246_477, w_246_481, w_246_484, w_246_485, w_246_486, w_246_490, w_246_492, w_246_493, w_246_494, w_246_495, w_246_498, w_246_499, w_246_504, w_246_507, w_246_512, w_246_515, w_246_516, w_246_518, w_246_519, w_246_520, w_246_522, w_246_525, w_246_526, w_246_531, w_246_532, w_246_534, w_246_535, w_246_536, w_246_538, w_246_539, w_246_541, w_246_542, w_246_544, w_246_545, w_246_547, w_246_548, w_246_549, w_246_551, w_246_552, w_246_553, w_246_554, w_246_555, w_246_556, w_246_557, w_246_558, w_246_559, w_246_561, w_246_563, w_246_565, w_246_566, w_246_568, w_246_571, w_246_575, w_246_576, w_246_577, w_246_580, w_246_581, w_246_582, w_246_583, w_246_586, w_246_588, w_246_593, w_246_595, w_246_598, w_246_599, w_246_600, w_246_602, w_246_603, w_246_604, w_246_606, w_246_607, w_246_608, w_246_611, w_246_612, w_246_614, w_246_616, w_246_617, w_246_618, w_246_619, w_246_620, w_246_623, w_246_624, w_246_627, w_246_628, w_246_631, w_246_633, w_246_636, w_246_638, w_246_641, w_246_642, w_246_644, w_246_645, w_246_646, w_246_647, w_246_648, w_246_650, w_246_652, w_246_658, w_246_660, w_246_661, w_246_662, w_246_664, w_246_665, w_246_666, w_246_670, w_246_672, w_246_673, w_246_674, w_246_676;
  wire w_247_005, w_247_008, w_247_011, w_247_015, w_247_031, w_247_036, w_247_043, w_247_054, w_247_059, w_247_063, w_247_069, w_247_075, w_247_081, w_247_097, w_247_098, w_247_105, w_247_106, w_247_107, w_247_110, w_247_112, w_247_116, w_247_134, w_247_146, w_247_149, w_247_150, w_247_155, w_247_158, w_247_162, w_247_163, w_247_165, w_247_169, w_247_177, w_247_181, w_247_183, w_247_186, w_247_194, w_247_199, w_247_212, w_247_216, w_247_217, w_247_239, w_247_240, w_247_242, w_247_248, w_247_250, w_247_252, w_247_254, w_247_261, w_247_264, w_247_265, w_247_273, w_247_278, w_247_287, w_247_289, w_247_292, w_247_295, w_247_301, w_247_322, w_247_331, w_247_337, w_247_343, w_247_349, w_247_358, w_247_362, w_247_371, w_247_374, w_247_378, w_247_389, w_247_395, w_247_397, w_247_402, w_247_404, w_247_410, w_247_412, w_247_417, w_247_420, w_247_421, w_247_431, w_247_433, w_247_450, w_247_458, w_247_461, w_247_462, w_247_471, w_247_476, w_247_481, w_247_492, w_247_494, w_247_495, w_247_498, w_247_500, w_247_501, w_247_507, w_247_510, w_247_513, w_247_516, w_247_521, w_247_528, w_247_538, w_247_548, w_247_554, w_247_560, w_247_569, w_247_570, w_247_574, w_247_578, w_247_580, w_247_582, w_247_584, w_247_586, w_247_595, w_247_600, w_247_604, w_247_608, w_247_624, w_247_635, w_247_642, w_247_644, w_247_648, w_247_649, w_247_666, w_247_671, w_247_673, w_247_677, w_247_689, w_247_707, w_247_732, w_247_741, w_247_745, w_247_748, w_247_751, w_247_761, w_247_773, w_247_774, w_247_776, w_247_782, w_247_815, w_247_821, w_247_846, w_247_851, w_247_854, w_247_857, w_247_868, w_247_884, w_247_894, w_247_896, w_247_950, w_247_972, w_247_997, w_247_1007, w_247_1009, w_247_1052, w_247_1089, w_247_1094, w_247_1095, w_247_1107, w_247_1108, w_247_1121, w_247_1125, w_247_1133, w_247_1155, w_247_1174, w_247_1187, w_247_1194, w_247_1201, w_247_1209, w_247_1216, w_247_1231, w_247_1238, w_247_1241, w_247_1245, w_247_1268, w_247_1269, w_247_1291, w_247_1292, w_247_1297, w_247_1313, w_247_1315, w_247_1339, w_247_1343, w_247_1371, w_247_1373, w_247_1381, w_247_1393, w_247_1397, w_247_1429, w_247_1433, w_247_1434, w_247_1449, w_247_1452, w_247_1469, w_247_1486, w_247_1490, w_247_1498, w_247_1504, w_247_1509, w_247_1517, w_247_1556, w_247_1560, w_247_1596, w_247_1597, w_247_1614, w_247_1618, w_247_1620, w_247_1627, w_247_1629, w_247_1645, w_247_1653, w_247_1664, w_247_1672, w_247_1673, w_247_1689, w_247_1700, w_247_1709, w_247_1711, w_247_1736, w_247_1740, w_247_1758, w_247_1761, w_247_1767, w_247_1770, w_247_1782, w_247_1788, w_247_1800, w_247_1802, w_247_1824, w_247_1827, w_247_1835, w_247_1836, w_247_1854, w_247_1868, w_247_1892, w_247_1894, w_247_1898, w_247_1905, w_247_1925, w_247_1928, w_247_1929, w_247_1960, w_247_1967, w_247_1969, w_247_1976, w_247_1980, w_247_1986, w_247_1990, w_247_1997, w_247_2006, w_247_2013, w_247_2029, w_247_2030, w_247_2040, w_247_2042, w_247_2047, w_247_2058, w_247_2079, w_247_2081, w_247_2087, w_247_2099, w_247_2104, w_247_2110, w_247_2111, w_247_2113, w_247_2124, w_247_2142, w_247_2146, w_247_2153, w_247_2189, w_247_2216, w_247_2222, w_247_2229, w_247_2235, w_247_2242, w_247_2266, w_247_2272, w_247_2289, w_247_2297, w_247_2301, w_247_2303, w_247_2306, w_247_2310, w_247_2320, w_247_2342, w_247_2361, w_247_2364, w_247_2371, w_247_2379, w_247_2418, w_247_2441, w_247_2456, w_247_2478, w_247_2496, w_247_2500, w_247_2513, w_247_2531, w_247_2576, w_247_2603, w_247_2605, w_247_2608, w_247_2609, w_247_2635, w_247_2643, w_247_2654, w_247_2668, w_247_2677, w_247_2722, w_247_2755, w_247_2783, w_247_2799, w_247_2801, w_247_2811, w_247_2813, w_247_2819, w_247_2831, w_247_2832, w_247_2835, w_247_2840, w_247_2843, w_247_2880, w_247_2900, w_247_2925, w_247_2926, w_247_2934, w_247_2949, w_247_2952, w_247_2961, w_247_2963, w_247_2964, w_247_2971, w_247_2981, w_247_2985, w_247_2987, w_247_2990, w_247_2991, w_247_2993, w_247_2999, w_247_3016, w_247_3024, w_247_3028, w_247_3031, w_247_3045, w_247_3049, w_247_3054, w_247_3070, w_247_3075, w_247_3077, w_247_3078, w_247_3097, w_247_3101, w_247_3131, w_247_3166, w_247_3169, w_247_3190, w_247_3192, w_247_3199, w_247_3220, w_247_3224, w_247_3227, w_247_3240, w_247_3241, w_247_3254, w_247_3264, w_247_3266, w_247_3274, w_247_3279, w_247_3302, w_247_3318, w_247_3325, w_247_3331, w_247_3341, w_247_3343, w_247_3347, w_247_3364, w_247_3371, w_247_3375, w_247_3378, w_247_3388, w_247_3389, w_247_3393, w_247_3396, w_247_3402, w_247_3426, w_247_3428, w_247_3482, w_247_3490, w_247_3496, w_247_3519, w_247_3525, w_247_3565, w_247_3574, w_247_3585, w_247_3587, w_247_3588, w_247_3598, w_247_3600, w_247_3601, w_247_3630, w_247_3637, w_247_3665, w_247_3681, w_247_3685, w_247_3689, w_247_3691, w_247_3708, w_247_3722, w_247_3747, w_247_3755, w_247_3756, w_247_3766, w_247_3771, w_247_3775, w_247_3782, w_247_3789, w_247_3814, w_247_3816, w_247_3821, w_247_3823, w_247_3840, w_247_3841, w_247_3845, w_247_3850, w_247_3852, w_247_3869, w_247_3871, w_247_3884, w_247_3885, w_247_3892, w_247_3893, w_247_3894, w_247_3927, w_247_3933, w_247_3955, w_247_3957, w_247_3958, w_247_3961, w_247_3987, w_247_4004, w_247_4008, w_247_4012, w_247_4016, w_247_4019, w_247_4022, w_247_4034, w_247_4057, w_247_4061, w_247_4069, w_247_4075, w_247_4078, w_247_4083, w_247_4095, w_247_4117, w_247_4122, w_247_4126, w_247_4135, w_247_4136, w_247_4144, w_247_4156, w_247_4158, w_247_4163, w_247_4184, w_247_4187, w_247_4190, w_247_4225, w_247_4272, w_247_4273, w_247_4288;
  wire w_248_005, w_248_006, w_248_012, w_248_020, w_248_021, w_248_031, w_248_041, w_248_051, w_248_054, w_248_060, w_248_067, w_248_068, w_248_074, w_248_099, w_248_105, w_248_115, w_248_121, w_248_131, w_248_136, w_248_144, w_248_145, w_248_154, w_248_171, w_248_172, w_248_173, w_248_176, w_248_177, w_248_180, w_248_185, w_248_193, w_248_196, w_248_205, w_248_217, w_248_218, w_248_221, w_248_230, w_248_237, w_248_239, w_248_240, w_248_242, w_248_251, w_248_252, w_248_253, w_248_259, w_248_282, w_248_303, w_248_304, w_248_316, w_248_318, w_248_341, w_248_343, w_248_344, w_248_348, w_248_349, w_248_374, w_248_375, w_248_377, w_248_393, w_248_400, w_248_402, w_248_403, w_248_404, w_248_415, w_248_419, w_248_421, w_248_422, w_248_430, w_248_435, w_248_438, w_248_450, w_248_452, w_248_457, w_248_472, w_248_482, w_248_493, w_248_497, w_248_503, w_248_505, w_248_506, w_248_515, w_248_530, w_248_532, w_248_533, w_248_535, w_248_537, w_248_538, w_248_553, w_248_557, w_248_563, w_248_570, w_248_578, w_248_580, w_248_582, w_248_584, w_248_597, w_248_606, w_248_607, w_248_609, w_248_610, w_248_614, w_248_616, w_248_619, w_248_623, w_248_625, w_248_634, w_248_638, w_248_639, w_248_641, w_248_642, w_248_643, w_248_644, w_248_645, w_248_647, w_248_650, w_248_668, w_248_670, w_248_674, w_248_678, w_248_683, w_248_691, w_248_693, w_248_707, w_248_717, w_248_718, w_248_722, w_248_725, w_248_749, w_248_751, w_248_760, w_248_766, w_248_769, w_248_774, w_248_782, w_248_786, w_248_788, w_248_795, w_248_796, w_248_798, w_248_799, w_248_805, w_248_808, w_248_810, w_248_818, w_248_827, w_248_832, w_248_835, w_248_852, w_248_859, w_248_866, w_248_867, w_248_877, w_248_885, w_248_887, w_248_888, w_248_890, w_248_900, w_248_909, w_248_912, w_248_915, w_248_919, w_248_929, w_248_954, w_248_956, w_248_963, w_248_968, w_248_980, w_248_986, w_248_990, w_248_995, w_248_997, w_248_1002, w_248_1003, w_248_1011, w_248_1013, w_248_1021, w_248_1025, w_248_1029, w_248_1032, w_248_1044, w_248_1050, w_248_1053, w_248_1055, w_248_1056, w_248_1085, w_248_1087, w_248_1101, w_248_1103, w_248_1109, w_248_1113, w_248_1114, w_248_1119, w_248_1120, w_248_1129, w_248_1141, w_248_1142, w_248_1143, w_248_1150, w_248_1161, w_248_1162, w_248_1163, w_248_1165, w_248_1167, w_248_1168, w_248_1171, w_248_1180, w_248_1182, w_248_1184, w_248_1185, w_248_1187, w_248_1193, w_248_1195, w_248_1199, w_248_1206, w_248_1207, w_248_1215, w_248_1217, w_248_1226, w_248_1227, w_248_1229, w_248_1230, w_248_1232, w_248_1245, w_248_1246, w_248_1250, w_248_1251, w_248_1254, w_248_1257, w_248_1272, w_248_1275, w_248_1276, w_248_1282, w_248_1294, w_248_1296, w_248_1301, w_248_1307, w_248_1314, w_248_1315, w_248_1318, w_248_1320, w_248_1329, w_248_1330, w_248_1331, w_248_1333, w_248_1340, w_248_1345, w_248_1346, w_248_1352, w_248_1354, w_248_1356, w_248_1357, w_248_1359, w_248_1361, w_248_1362, w_248_1364, w_248_1366, w_248_1380, w_248_1385, w_248_1395, w_248_1400, w_248_1411, w_248_1426, w_248_1429, w_248_1430, w_248_1436, w_248_1441, w_248_1453, w_248_1456, w_248_1457, w_248_1464, w_248_1465, w_248_1471, w_248_1474, w_248_1479, w_248_1490, w_248_1492, w_248_1497, w_248_1499, w_248_1511, w_248_1512, w_248_1515, w_248_1523, w_248_1525, w_248_1527, w_248_1533, w_248_1538, w_248_1540, w_248_1542, w_248_1543, w_248_1546, w_248_1556, w_248_1557, w_248_1562, w_248_1563, w_248_1571, w_248_1574, w_248_1582, w_248_1593, w_248_1596, w_248_1598, w_248_1601, w_248_1627, w_248_1641, w_248_1650, w_248_1664, w_248_1665, w_248_1667, w_248_1671, w_248_1677, w_248_1695, w_248_1698, w_248_1714, w_248_1718, w_248_1719, w_248_1722, w_248_1725, w_248_1729, w_248_1736, w_248_1740, w_248_1743, w_248_1744, w_248_1757, w_248_1772, w_248_1773, w_248_1780, w_248_1782, w_248_1783, w_248_1791, w_248_1799, w_248_1816, w_248_1829, w_248_1835, w_248_1848, w_248_1852, w_248_1861, w_248_1862, w_248_1867, w_248_1885, w_248_1906, w_248_1915, w_248_1934, w_248_1935, w_248_1941, w_248_1956, w_248_1966, w_248_1969, w_248_1971, w_248_1976, w_248_1998, w_248_2035, w_248_2037, w_248_2045, w_248_2047, w_248_2049, w_248_2051, w_248_2069, w_248_2072, w_248_2079, w_248_2104, w_248_2112, w_248_2125, w_248_2137, w_248_2152, w_248_2171, w_248_2189, w_248_2220, w_248_2229, w_248_2247, w_248_2263, w_248_2273, w_248_2299, w_248_2308, w_248_2318, w_248_2324, w_248_2332, w_248_2359, w_248_2364, w_248_2375, w_248_2377, w_248_2395, w_248_2401, w_248_2409, w_248_2421, w_248_2422, w_248_2423, w_248_2430, w_248_2450, w_248_2461, w_248_2474, w_248_2478, w_248_2481, w_248_2488, w_248_2493, w_248_2496, w_248_2526, w_248_2551, w_248_2565, w_248_2566, w_248_2567, w_248_2582, w_248_2590, w_248_2602, w_248_2615, w_248_2619, w_248_2622, w_248_2628, w_248_2641, w_248_2645, w_248_2649, w_248_2657, w_248_2672, w_248_2677, w_248_2697, w_248_2698, w_248_2721, w_248_2760, w_248_2765, w_248_2774, w_248_2784, w_248_2791, w_248_2809, w_248_2824, w_248_2854, w_248_2882, w_248_2888, w_248_2903, w_248_2919, w_248_2929, w_248_2937, w_248_2948, w_248_2965, w_248_2973, w_248_2974, w_248_3023, w_248_3051, w_248_3055, w_248_3070, w_248_3081, w_248_3083, w_248_3094, w_248_3095, w_248_3111, w_248_3113, w_248_3128, w_248_3132, w_248_3141, w_248_3146, w_248_3164, w_248_3171, w_248_3174, w_248_3179, w_248_3190, w_248_3192, w_248_3198;
  wire w_249_001, w_249_007, w_249_009, w_249_011, w_249_013, w_249_018, w_249_021, w_249_023, w_249_024, w_249_025, w_249_033, w_249_035, w_249_047, w_249_048, w_249_050, w_249_051, w_249_060, w_249_063, w_249_071, w_249_076, w_249_079, w_249_087, w_249_095, w_249_106, w_249_109, w_249_111, w_249_123, w_249_126, w_249_128, w_249_131, w_249_137, w_249_140, w_249_144, w_249_149, w_249_153, w_249_160, w_249_174, w_249_179, w_249_187, w_249_188, w_249_189, w_249_202, w_249_205, w_249_216, w_249_219, w_249_222, w_249_223, w_249_228, w_249_229, w_249_234, w_249_235, w_249_245, w_249_255, w_249_256, w_249_263, w_249_264, w_249_273, w_249_274, w_249_277, w_249_280, w_249_281, w_249_282, w_249_295, w_249_304, w_249_306, w_249_313, w_249_322, w_249_326, w_249_333, w_249_334, w_249_352, w_249_355, w_249_356, w_249_360, w_249_376, w_249_381, w_249_384, w_249_389, w_249_396, w_249_407, w_249_416, w_249_423, w_249_424, w_249_439, w_249_441, w_249_443, w_249_446, w_249_452, w_249_456, w_249_458, w_249_460, w_249_461, w_249_481, w_249_483, w_249_491, w_249_496, w_249_499, w_249_502, w_249_518, w_249_522, w_249_526, w_249_539, w_249_543, w_249_553, w_249_555, w_249_565, w_249_568, w_249_580, w_249_586, w_249_588, w_249_589, w_249_590, w_249_592, w_249_601, w_249_613, w_249_614, w_249_622, w_249_623, w_249_624, w_249_628, w_249_634, w_249_635, w_249_645, w_249_646, w_249_656, w_249_659, w_249_663, w_249_667, w_249_669, w_249_683, w_249_685, w_249_702, w_249_714, w_249_717, w_249_719, w_249_724, w_249_731, w_249_737, w_249_747, w_249_761, w_249_763, w_249_765, w_249_772, w_249_779, w_249_793, w_249_801, w_249_803, w_249_805, w_249_813, w_249_814, w_249_824, w_249_827, w_249_838, w_249_846, w_249_849, w_249_856, w_249_864, w_249_865, w_249_868, w_249_871, w_249_872, w_249_885, w_249_888, w_249_899, w_249_904, w_249_905, w_249_908, w_249_922, w_249_927, w_249_932, w_249_934, w_249_937, w_249_940, w_249_941, w_249_948, w_249_953, w_249_954, w_249_962, w_249_966, w_249_969, w_249_970, w_249_973, w_249_974, w_249_986, w_249_990, w_249_991, w_249_992, w_249_993, w_249_998, w_249_1003, w_249_1011, w_249_1015, w_249_1018, w_249_1022, w_249_1027, w_249_1030, w_249_1034, w_249_1036, w_249_1039, w_249_1042, w_249_1044, w_249_1050, w_249_1051, w_249_1060, w_249_1061, w_249_1064, w_249_1068, w_249_1072, w_249_1095, w_249_1112, w_249_1125, w_249_1132, w_249_1134, w_249_1150, w_249_1155, w_249_1158, w_249_1159, w_249_1161, w_249_1167, w_249_1192, w_249_1193, w_249_1194, w_249_1195, w_249_1196, w_249_1199, w_249_1202, w_249_1206, w_249_1208, w_249_1210, w_249_1213, w_249_1218, w_249_1219, w_249_1222, w_249_1234, w_249_1250, w_249_1259, w_249_1262, w_249_1266, w_249_1267, w_249_1275, w_249_1285, w_249_1286, w_249_1288, w_249_1291, w_249_1293, w_249_1298, w_249_1302, w_249_1315, w_249_1316, w_249_1317, w_249_1322, w_249_1324, w_249_1343, w_249_1345, w_249_1349, w_249_1353, w_249_1355, w_249_1357, w_249_1362, w_249_1371, w_249_1383, w_249_1384, w_249_1385, w_249_1394, w_249_1416, w_249_1421, w_249_1428, w_249_1429, w_249_1431, w_249_1433, w_249_1434, w_249_1438, w_249_1449, w_249_1452, w_249_1469, w_249_1478, w_249_1484, w_249_1497, w_249_1504, w_249_1505, w_249_1513, w_249_1518, w_249_1520, w_249_1538, w_249_1551, w_249_1556, w_249_1564, w_249_1565, w_249_1567, w_249_1572, w_249_1574, w_249_1575, w_249_1581, w_249_1584, w_249_1586, w_249_1596, w_249_1600, w_249_1604, w_249_1608, w_249_1614, w_249_1618, w_249_1620, w_249_1628, w_249_1634, w_249_1642, w_249_1645, w_249_1646, w_249_1662, w_249_1666, w_249_1668, w_249_1673, w_249_1674, w_249_1686, w_249_1689, w_249_1691, w_249_1700, w_249_1705, w_249_1706, w_249_1711, w_249_1712, w_249_1713, w_249_1716, w_249_1726, w_249_1738, w_249_1745, w_249_1748, w_249_1751, w_249_1783, w_249_1787, w_249_1790, w_249_1798, w_249_1799, w_249_1800, w_249_1803, w_249_1813, w_249_1819, w_249_1823, w_249_1828, w_249_1845, w_249_1846, w_249_1850, w_249_1851, w_249_1852, w_249_1871, w_249_1882, w_249_1886, w_249_1891, w_249_1910, w_249_1913, w_249_1920, w_249_1934, w_249_1952, w_249_1970, w_249_1972, w_249_1975, w_249_1991, w_249_1994, w_249_2009, w_249_2014, w_249_2016, w_249_2030, w_249_2033, w_249_2042, w_249_2051, w_249_2054, w_249_2060, w_249_2072, w_249_2076, w_249_2084, w_249_2091, w_249_2093, w_249_2109, w_249_2115, w_249_2180, w_249_2183, w_249_2190, w_249_2205, w_249_2209, w_249_2218, w_249_2219, w_249_2225, w_249_2229, w_249_2237, w_249_2245, w_249_2256, w_249_2257, w_249_2265, w_249_2271, w_249_2289, w_249_2294, w_249_2296, w_249_2308, w_249_2314, w_249_2316, w_249_2347, w_249_2366, w_249_2384, w_249_2389, w_249_2398, w_249_2402, w_249_2407, w_249_2414, w_249_2422, w_249_2437, w_249_2443, w_249_2449, w_249_2458, w_249_2469, w_249_2478, w_249_2493, w_249_2497, w_249_2501, w_249_2504, w_249_2528, w_249_2540, w_249_2571, w_249_2572, w_249_2573, w_249_2575, w_249_2600, w_249_2616, w_249_2624, w_249_2627, w_249_2636, w_249_2644, w_249_2651, w_249_2656, w_249_2661, w_249_2686, w_249_2695, w_249_2716, w_249_2720, w_249_2729, w_249_2737, w_249_2740, w_249_2745, w_249_2762, w_249_2778, w_249_2780, w_249_2788, w_249_2803, w_249_2804, w_249_2829, w_249_2830, w_249_2836, w_249_2857, w_249_2859, w_249_2890, w_249_2907, w_249_2910, w_249_2928, w_249_2929, w_249_2948, w_249_2966, w_249_2967, w_249_2973, w_249_2978, w_249_3032, w_249_3037, w_249_3065, w_249_3071, w_249_3081, w_249_3093, w_249_3112, w_249_3122, w_249_3124, w_249_3130, w_249_3133, w_249_3149, w_249_3151, w_249_3156, w_249_3166, w_249_3177, w_249_3178, w_249_3179, w_249_3180, w_249_3181, w_249_3182, w_249_3183, w_249_3184, w_249_3188, w_249_3189, w_249_3190, w_249_3192;
  wire w_250_001, w_250_003, w_250_004, w_250_006, w_250_007, w_250_009, w_250_010, w_250_011, w_250_012, w_250_013, w_250_014, w_250_015, w_250_016, w_250_018, w_250_019, w_250_020, w_250_021, w_250_022, w_250_023, w_250_024, w_250_025, w_250_026, w_250_027, w_250_028, w_250_029, w_250_030, w_250_031, w_250_032, w_250_033, w_250_034, w_250_035, w_250_037, w_250_039, w_250_040, w_250_043, w_250_044, w_250_045, w_250_046, w_250_048, w_250_049, w_250_051, w_250_052, w_250_054, w_250_055, w_250_056, w_250_058, w_250_060, w_250_065, w_250_066, w_250_067, w_250_068, w_250_069, w_250_070, w_250_072, w_250_074, w_250_075, w_250_076, w_250_077, w_250_078, w_250_079, w_250_080, w_250_081, w_250_082, w_250_083, w_250_084, w_250_085, w_250_087, w_250_088, w_250_089, w_250_090, w_250_093, w_250_094, w_250_096, w_250_100, w_250_101, w_250_105, w_250_106, w_250_107, w_250_108, w_250_110, w_250_111, w_250_112, w_250_113, w_250_115, w_250_116, w_250_117, w_250_119, w_250_120, w_250_121, w_250_123, w_250_127, w_250_128, w_250_130, w_250_132, w_250_133, w_250_134, w_250_135, w_250_136, w_250_139, w_250_141, w_250_142, w_250_144, w_250_145, w_250_146, w_250_148, w_250_149, w_250_150, w_250_151, w_250_152, w_250_154, w_250_155, w_250_156, w_250_157, w_250_158, w_250_159, w_250_160, w_250_161, w_250_163, w_250_166, w_250_168, w_250_169, w_250_170, w_250_171, w_250_172, w_250_173, w_250_174, w_250_175, w_250_176, w_250_177, w_250_178, w_250_180, w_250_181, w_250_182, w_250_183, w_250_184, w_250_185, w_250_186, w_250_187, w_250_188, w_250_189, w_250_191, w_250_193, w_250_196, w_250_198, w_250_199, w_250_200, w_250_202, w_250_203, w_250_204, w_250_205, w_250_206, w_250_207, w_250_208, w_250_209, w_250_210, w_250_212, w_250_213, w_250_214, w_250_215, w_250_216, w_250_217, w_250_218, w_250_219, w_250_220, w_250_222, w_250_223, w_250_224, w_250_227, w_250_228, w_250_229, w_250_230, w_250_231, w_250_232, w_250_234, w_250_236, w_250_238, w_250_239, w_250_241, w_250_244, w_250_245, w_250_247, w_250_248, w_250_249, w_250_251, w_250_252, w_250_253, w_250_256, w_250_257, w_250_258, w_250_259, w_250_260, w_250_261, w_250_262, w_250_263, w_250_264, w_250_265, w_250_266, w_250_267, w_250_269, w_250_271, w_250_272, w_250_273, w_250_274, w_250_275, w_250_276, w_250_278, w_250_279, w_250_281, w_250_282, w_250_283, w_250_284, w_250_285, w_250_286, w_250_287, w_250_289, w_250_291, w_250_294, w_250_295, w_250_296, w_250_298, w_250_299, w_250_300, w_250_301, w_250_302, w_250_303, w_250_304, w_250_306, w_250_307, w_250_308, w_250_310, w_250_311, w_250_312, w_250_314, w_250_315, w_250_319, w_250_320, w_250_323, w_250_324, w_250_326, w_250_329, w_250_330, w_250_332, w_250_333, w_250_334, w_250_335, w_250_336, w_250_337, w_250_338, w_250_339, w_250_341, w_250_342, w_250_343, w_250_344, w_250_345, w_250_349, w_250_350, w_250_351, w_250_352, w_250_354, w_250_356, w_250_357, w_250_359, w_250_361, w_250_362, w_250_363, w_250_364, w_250_365, w_250_366, w_250_367, w_250_369, w_250_370, w_250_371, w_250_374, w_250_375, w_250_376, w_250_377, w_250_378, w_250_379, w_250_380;
  wire w_251_001, w_251_007, w_251_008, w_251_012, w_251_013, w_251_019, w_251_023, w_251_027, w_251_032, w_251_034, w_251_036, w_251_037, w_251_043, w_251_044, w_251_045, w_251_046, w_251_047, w_251_048, w_251_052, w_251_054, w_251_055, w_251_056, w_251_058, w_251_062, w_251_063, w_251_065, w_251_074, w_251_084, w_251_096, w_251_099, w_251_100, w_251_102, w_251_109, w_251_112, w_251_114, w_251_116, w_251_118, w_251_119, w_251_121, w_251_123, w_251_135, w_251_137, w_251_138, w_251_146, w_251_150, w_251_152, w_251_155, w_251_157, w_251_161, w_251_163, w_251_167, w_251_173, w_251_176, w_251_180, w_251_181, w_251_184, w_251_185, w_251_192, w_251_199, w_251_203, w_251_208, w_251_213, w_251_218, w_251_227, w_251_229, w_251_232, w_251_237, w_251_244, w_251_249, w_251_253, w_251_258, w_251_263, w_251_265, w_251_270, w_251_273, w_251_274, w_251_286, w_251_287, w_251_289, w_251_299, w_251_303, w_251_310, w_251_318, w_251_322, w_251_324, w_251_332, w_251_333, w_251_338, w_251_341, w_251_346, w_251_351, w_251_359, w_251_374, w_251_378, w_251_385, w_251_388, w_251_390, w_251_394, w_251_397, w_251_400, w_251_407, w_251_418, w_251_420, w_251_422, w_251_423, w_251_426, w_251_428, w_251_434, w_251_440, w_251_447, w_251_449, w_251_458, w_251_465, w_251_469, w_251_472, w_251_473, w_251_482, w_251_490, w_251_492, w_251_497, w_251_501, w_251_511, w_251_521, w_251_537, w_251_551, w_251_552, w_251_563, w_251_566, w_251_583, w_251_584, w_251_613, w_251_650, w_251_653, w_251_667, w_251_682, w_251_684, w_251_685, w_251_687, w_251_696, w_251_703, w_251_704, w_251_706, w_251_709, w_251_713, w_251_722, w_251_724, w_251_725, w_251_726, w_251_751, w_251_753, w_251_755, w_251_762, w_251_781, w_251_782, w_251_785, w_251_789, w_251_793, w_251_800, w_251_801, w_251_823, w_251_825, w_251_830, w_251_840, w_251_843, w_251_846, w_251_853, w_251_856, w_251_862, w_251_865, w_251_872, w_251_875, w_251_878, w_251_879, w_251_880, w_251_881, w_251_882, w_251_884, w_251_887, w_251_888, w_251_893, w_251_915, w_251_926, w_251_930, w_251_932, w_251_935, w_251_942, w_251_944, w_251_954, w_251_959, w_251_962, w_251_968, w_251_984, w_251_992, w_251_994, w_251_998, w_251_1001, w_251_1006, w_251_1030, w_251_1035, w_251_1041, w_251_1047, w_251_1051, w_251_1054, w_251_1063, w_251_1075, w_251_1079, w_251_1080, w_251_1093, w_251_1099, w_251_1102, w_251_1110, w_251_1111, w_251_1125, w_251_1136, w_251_1144, w_251_1146, w_251_1154, w_251_1173, w_251_1177, w_251_1178, w_251_1185, w_251_1187, w_251_1190, w_251_1191, w_251_1194, w_251_1199, w_251_1202, w_251_1219, w_251_1228, w_251_1233, w_251_1248, w_251_1271, w_251_1272, w_251_1273, w_251_1289, w_251_1291, w_251_1298, w_251_1301, w_251_1302, w_251_1305, w_251_1306, w_251_1308, w_251_1311, w_251_1314, w_251_1316, w_251_1319, w_251_1324, w_251_1325, w_251_1332, w_251_1346, w_251_1353, w_251_1367, w_251_1376, w_251_1378, w_251_1383, w_251_1394, w_251_1398, w_251_1406, w_251_1423, w_251_1424, w_251_1426, w_251_1437, w_251_1438, w_251_1440, w_251_1444, w_251_1452, w_251_1454, w_251_1455, w_251_1456, w_251_1461, w_251_1476, w_251_1479, w_251_1480, w_251_1490, w_251_1505, w_251_1511, w_251_1512, w_251_1522, w_251_1532, w_251_1541, w_251_1542, w_251_1543, w_251_1544, w_251_1552, w_251_1560, w_251_1570, w_251_1573, w_251_1574, w_251_1577, w_251_1590, w_251_1601, w_251_1602, w_251_1605, w_251_1608, w_251_1625, w_251_1631, w_251_1634, w_251_1638, w_251_1641, w_251_1648, w_251_1651, w_251_1657, w_251_1665, w_251_1674, w_251_1684, w_251_1706, w_251_1711, w_251_1716, w_251_1724, w_251_1731, w_251_1736, w_251_1747, w_251_1753, w_251_1755, w_251_1768, w_251_1774, w_251_1778, w_251_1794, w_251_1797, w_251_1798, w_251_1807, w_251_1813, w_251_1817, w_251_1822, w_251_1826, w_251_1827, w_251_1849, w_251_1853, w_251_1861, w_251_1867, w_251_1877, w_251_1882, w_251_1889, w_251_1895, w_251_1899, w_251_1903, w_251_1905, w_251_1911, w_251_1916, w_251_1918, w_251_1937, w_251_1944, w_251_1963, w_251_1976, w_251_1997, w_251_2003, w_251_2009, w_251_2010, w_251_2013, w_251_2015, w_251_2016, w_251_2024, w_251_2026, w_251_2028, w_251_2030, w_251_2037, w_251_2041, w_251_2044, w_251_2046, w_251_2049, w_251_2053, w_251_2058, w_251_2072, w_251_2074, w_251_2076, w_251_2083, w_251_2084, w_251_2086, w_251_2104, w_251_2114, w_251_2115, w_251_2129, w_251_2133, w_251_2136, w_251_2140, w_251_2141, w_251_2146, w_251_2147, w_251_2154, w_251_2157, w_251_2161, w_251_2162, w_251_2163, w_251_2164, w_251_2172, w_251_2176, w_251_2177, w_251_2179, w_251_2182, w_251_2186, w_251_2188, w_251_2207, w_251_2210, w_251_2231, w_251_2232, w_251_2242, w_251_2244, w_251_2245, w_251_2246, w_251_2248, w_251_2250, w_251_2262, w_251_2264, w_251_2266, w_251_2277, w_251_2280, w_251_2284, w_251_2285, w_251_2288, w_251_2290, w_251_2291, w_251_2295, w_251_2301, w_251_2306, w_251_2318, w_251_2322, w_251_2324, w_251_2328, w_251_2351, w_251_2358, w_251_2369, w_251_2373, w_251_2375, w_251_2398, w_251_2404, w_251_2407, w_251_2416, w_251_2417, w_251_2425, w_251_2428, w_251_2431, w_251_2432, w_251_2433, w_251_2434, w_251_2435, w_251_2436;
  wire w_252_005, w_252_006, w_252_009, w_252_010, w_252_012, w_252_023, w_252_033, w_252_056, w_252_057, w_252_058, w_252_060, w_252_062, w_252_067, w_252_070, w_252_074, w_252_078, w_252_081, w_252_082, w_252_102, w_252_109, w_252_111, w_252_112, w_252_124, w_252_141, w_252_145, w_252_154, w_252_155, w_252_165, w_252_169, w_252_174, w_252_180, w_252_182, w_252_191, w_252_193, w_252_195, w_252_211, w_252_213, w_252_214, w_252_216, w_252_226, w_252_233, w_252_234, w_252_237, w_252_239, w_252_256, w_252_275, w_252_282, w_252_296, w_252_298, w_252_312, w_252_313, w_252_319, w_252_326, w_252_327, w_252_336, w_252_346, w_252_351, w_252_359, w_252_363, w_252_366, w_252_386, w_252_390, w_252_397, w_252_401, w_252_409, w_252_411, w_252_413, w_252_415, w_252_423, w_252_426, w_252_431, w_252_432, w_252_435, w_252_443, w_252_452, w_252_454, w_252_459, w_252_464, w_252_470, w_252_473, w_252_477, w_252_480, w_252_483, w_252_492, w_252_495, w_252_496, w_252_512, w_252_515, w_252_520, w_252_536, w_252_541, w_252_544, w_252_559, w_252_567, w_252_574, w_252_577, w_252_583, w_252_586, w_252_593, w_252_596, w_252_600, w_252_603, w_252_604, w_252_606, w_252_609, w_252_615, w_252_616, w_252_617, w_252_618, w_252_622, w_252_623, w_252_624, w_252_650, w_252_659, w_252_668, w_252_674, w_252_676, w_252_681, w_252_682, w_252_686, w_252_689, w_252_696, w_252_702, w_252_706, w_252_707, w_252_712, w_252_715, w_252_717, w_252_721, w_252_724, w_252_727, w_252_736, w_252_739, w_252_745, w_252_749, w_252_760, w_252_764, w_252_766, w_252_767, w_252_773, w_252_775, w_252_778, w_252_779, w_252_780, w_252_785, w_252_790, w_252_792, w_252_795, w_252_797, w_252_806, w_252_819, w_252_824, w_252_825, w_252_855, w_252_860, w_252_865, w_252_872, w_252_876, w_252_883, w_252_884, w_252_885, w_252_902, w_252_904, w_252_906, w_252_910, w_252_919, w_252_926, w_252_929, w_252_937, w_252_957, w_252_968, w_252_976, w_252_978, w_252_985, w_252_991, w_252_993, w_252_994, w_252_998, w_252_1006, w_252_1009, w_252_1025, w_252_1029, w_252_1031, w_252_1040, w_252_1051, w_252_1052, w_252_1053, w_252_1054, w_252_1056, w_252_1057, w_252_1065, w_252_1074, w_252_1075, w_252_1081, w_252_1084, w_252_1089, w_252_1097, w_252_1105, w_252_1107, w_252_1115, w_252_1119, w_252_1121, w_252_1124, w_252_1135, w_252_1138, w_252_1142, w_252_1143, w_252_1144, w_252_1147, w_252_1149, w_252_1157, w_252_1160, w_252_1164, w_252_1166, w_252_1174, w_252_1175, w_252_1179, w_252_1186, w_252_1191, w_252_1195, w_252_1196, w_252_1199, w_252_1200, w_252_1204, w_252_1205, w_252_1222, w_252_1224, w_252_1226, w_252_1239, w_252_1240, w_252_1250, w_252_1270, w_252_1273, w_252_1274, w_252_1277, w_252_1280, w_252_1286, w_252_1301, w_252_1304, w_252_1319, w_252_1329, w_252_1331, w_252_1334, w_252_1340, w_252_1352, w_252_1356, w_252_1367, w_252_1368, w_252_1370, w_252_1387, w_252_1389, w_252_1390, w_252_1391, w_252_1392, w_252_1395, w_252_1396, w_252_1400, w_252_1402, w_252_1405, w_252_1413, w_252_1421, w_252_1432, w_252_1433, w_252_1438, w_252_1449, w_252_1450, w_252_1466, w_252_1470, w_252_1472, w_252_1475, w_252_1476, w_252_1481, w_252_1483, w_252_1506, w_252_1523, w_252_1525, w_252_1530, w_252_1539, w_252_1552, w_252_1553, w_252_1554, w_252_1555, w_252_1558, w_252_1586, w_252_1594, w_252_1597, w_252_1606, w_252_1614, w_252_1621, w_252_1630, w_252_1632, w_252_1633, w_252_1634, w_252_1637, w_252_1642, w_252_1651, w_252_1661, w_252_1665, w_252_1669, w_252_1681, w_252_1686, w_252_1689, w_252_1696, w_252_1703, w_252_1704, w_252_1706, w_252_1720, w_252_1722, w_252_1723, w_252_1725, w_252_1733, w_252_1735, w_252_1770, w_252_1774, w_252_1785, w_252_1804, w_252_1805, w_252_1807, w_252_1813, w_252_1815, w_252_1823, w_252_1830, w_252_1834, w_252_1835, w_252_1838, w_252_1850, w_252_1853, w_252_1890, w_252_1892, w_252_1896, w_252_1897, w_252_1898, w_252_1901, w_252_1905, w_252_1911, w_252_1912, w_252_1913, w_252_1915, w_252_1919, w_252_1928, w_252_1929, w_252_1942, w_252_1945, w_252_1947, w_252_1955, w_252_1969, w_252_1974, w_252_1994, w_252_1995, w_252_2000, w_252_2008, w_252_2019, w_252_2025, w_252_2030, w_252_2035, w_252_2048, w_252_2049, w_252_2061, w_252_2066, w_252_2071, w_252_2072, w_252_2074, w_252_2075, w_252_2081, w_252_2084, w_252_2086, w_252_2092, w_252_2094, w_252_2095, w_252_2098, w_252_2103, w_252_2105, w_252_2108, w_252_2113, w_252_2115, w_252_2118, w_252_2121, w_252_2124, w_252_2126, w_252_2127, w_252_2129, w_252_2131, w_252_2137, w_252_2138, w_252_2144, w_252_2148, w_252_2160, w_252_2161, w_252_2165, w_252_2166, w_252_2170, w_252_2178, w_252_2179, w_252_2182, w_252_2187, w_252_2197, w_252_2202, w_252_2203, w_252_2205, w_252_2207, w_252_2209, w_252_2211, w_252_2216, w_252_2222, w_252_2224, w_252_2226, w_252_2228, w_252_2235, w_252_2237, w_252_2238, w_252_2243, w_252_2245, w_252_2247, w_252_2276, w_252_2277, w_252_2279, w_252_2282, w_252_2287, w_252_2291, w_252_2299, w_252_2300, w_252_2307, w_252_2313, w_252_2314, w_252_2321, w_252_2329, w_252_2334, w_252_2339, w_252_2340, w_252_2355, w_252_2360, w_252_2362, w_252_2365, w_252_2385, w_252_2388, w_252_2391, w_252_2394, w_252_2397, w_252_2408, w_252_2413, w_252_2414, w_252_2417, w_252_2419, w_252_2423, w_252_2430, w_252_2432, w_252_2450, w_252_2456, w_252_2460, w_252_2462, w_252_2480, w_252_2493, w_252_2501, w_252_2502, w_252_2519, w_252_2523, w_252_2532, w_252_2537, w_252_2552, w_252_2555, w_252_2564, w_252_2565, w_252_2569;
  wire w_253_003, w_253_007, w_253_022, w_253_023, w_253_043, w_253_045, w_253_048, w_253_051, w_253_059, w_253_062, w_253_074, w_253_084, w_253_087, w_253_090, w_253_095, w_253_100, w_253_105, w_253_122, w_253_134, w_253_142, w_253_149, w_253_162, w_253_166, w_253_171, w_253_183, w_253_196, w_253_210, w_253_215, w_253_216, w_253_220, w_253_226, w_253_227, w_253_232, w_253_252, w_253_253, w_253_265, w_253_267, w_253_269, w_253_272, w_253_279, w_253_287, w_253_313, w_253_314, w_253_316, w_253_327, w_253_332, w_253_334, w_253_342, w_253_344, w_253_351, w_253_352, w_253_353, w_253_355, w_253_363, w_253_366, w_253_368, w_253_369, w_253_372, w_253_379, w_253_381, w_253_382, w_253_383, w_253_390, w_253_395, w_253_399, w_253_400, w_253_405, w_253_411, w_253_419, w_253_424, w_253_427, w_253_428, w_253_429, w_253_431, w_253_442, w_253_443, w_253_445, w_253_449, w_253_472, w_253_477, w_253_479, w_253_482, w_253_484, w_253_495, w_253_501, w_253_502, w_253_506, w_253_519, w_253_524, w_253_525, w_253_536, w_253_537, w_253_539, w_253_549, w_253_562, w_253_567, w_253_568, w_253_573, w_253_574, w_253_586, w_253_598, w_253_607, w_253_610, w_253_615, w_253_617, w_253_628, w_253_636, w_253_639, w_253_642, w_253_644, w_253_649, w_253_651, w_253_669, w_253_672, w_253_682, w_253_689, w_253_690, w_253_692, w_253_697, w_253_700, w_253_704, w_253_706, w_253_710, w_253_722, w_253_725, w_253_731, w_253_733, w_253_735, w_253_736, w_253_740, w_253_756, w_253_761, w_253_771, w_253_775, w_253_776, w_253_797, w_253_798, w_253_803, w_253_815, w_253_816, w_253_843, w_253_846, w_253_851, w_253_856, w_253_858, w_253_861, w_253_883, w_253_886, w_253_902, w_253_909, w_253_925, w_253_926, w_253_934, w_253_943, w_253_944, w_253_946, w_253_956, w_253_971, w_253_974, w_253_981, w_253_989, w_253_994, w_253_1002, w_253_1011, w_253_1012, w_253_1014, w_253_1016, w_253_1017, w_253_1018, w_253_1021, w_253_1029, w_253_1035, w_253_1036, w_253_1042, w_253_1046, w_253_1048, w_253_1052, w_253_1053, w_253_1056, w_253_1066, w_253_1068, w_253_1076, w_253_1087, w_253_1100, w_253_1103, w_253_1105, w_253_1107, w_253_1111, w_253_1122, w_253_1125, w_253_1134, w_253_1139, w_253_1143, w_253_1149, w_253_1151, w_253_1155, w_253_1157, w_253_1158, w_253_1165, w_253_1181, w_253_1182, w_253_1185, w_253_1200, w_253_1202, w_253_1232, w_253_1256, w_253_1259, w_253_1276, w_253_1282, w_253_1287, w_253_1310, w_253_1315, w_253_1319, w_253_1326, w_253_1333, w_253_1340, w_253_1343, w_253_1346, w_253_1352, w_253_1354, w_253_1360, w_253_1373, w_253_1375, w_253_1377, w_253_1382, w_253_1396, w_253_1400, w_253_1406, w_253_1413, w_253_1427, w_253_1429, w_253_1434, w_253_1438, w_253_1439, w_253_1440, w_253_1449, w_253_1454, w_253_1464, w_253_1468, w_253_1482, w_253_1484, w_253_1506, w_253_1518, w_253_1521, w_253_1544, w_253_1547, w_253_1548, w_253_1560, w_253_1576, w_253_1578, w_253_1589, w_253_1591, w_253_1597, w_253_1600, w_253_1603, w_253_1604, w_253_1615, w_253_1647, w_253_1660, w_253_1681, w_253_1683, w_253_1689, w_253_1690, w_253_1705, w_253_1729, w_253_1733, w_253_1737, w_253_1739, w_253_1744, w_253_1752, w_253_1756, w_253_1759, w_253_1769, w_253_1770, w_253_1774, w_253_1779, w_253_1782, w_253_1794, w_253_1832, w_253_1845, w_253_1854, w_253_1858, w_253_1879, w_253_1897, w_253_1911, w_253_1915, w_253_1917, w_253_1921, w_253_1925, w_253_1956, w_253_1991, w_253_1996, w_253_1999, w_253_2015, w_253_2030, w_253_2047, w_253_2048, w_253_2057, w_253_2058, w_253_2065, w_253_2074, w_253_2088, w_253_2092, w_253_2101, w_253_2135, w_253_2140, w_253_2142, w_253_2162, w_253_2176, w_253_2181, w_253_2191, w_253_2194, w_253_2210, w_253_2213, w_253_2227, w_253_2243, w_253_2253, w_253_2258, w_253_2265, w_253_2305, w_253_2310, w_253_2334, w_253_2344, w_253_2360, w_253_2368, w_253_2369, w_253_2387, w_253_2397, w_253_2407, w_253_2409, w_253_2410, w_253_2413, w_253_2417, w_253_2428, w_253_2430, w_253_2434, w_253_2446, w_253_2456, w_253_2458, w_253_2462, w_253_2476, w_253_2477, w_253_2483, w_253_2498, w_253_2499, w_253_2503, w_253_2505, w_253_2506, w_253_2511, w_253_2530, w_253_2533, w_253_2537, w_253_2540, w_253_2548, w_253_2575, w_253_2581, w_253_2599, w_253_2601, w_253_2602, w_253_2624, w_253_2631, w_253_2652, w_253_2653, w_253_2654, w_253_2666, w_253_2673, w_253_2676, w_253_2687, w_253_2725, w_253_2741, w_253_2752, w_253_2756, w_253_2758, w_253_2760, w_253_2772, w_253_2787, w_253_2789, w_253_2792, w_253_2797, w_253_2800, w_253_2808, w_253_2816, w_253_2831, w_253_2861, w_253_2872, w_253_2877, w_253_2885, w_253_2889, w_253_2892, w_253_2895, w_253_2897, w_253_2910, w_253_2914, w_253_2933, w_253_2939, w_253_2961, w_253_2966, w_253_2976, w_253_2978, w_253_2982, w_253_2994, w_253_3005, w_253_3023, w_253_3028, w_253_3072, w_253_3084, w_253_3090, w_253_3092, w_253_3098, w_253_3105, w_253_3107, w_253_3110, w_253_3117, w_253_3118, w_253_3128, w_253_3154, w_253_3167, w_253_3177, w_253_3179, w_253_3188, w_253_3189, w_253_3192, w_253_3195, w_253_3196, w_253_3202, w_253_3205, w_253_3220, w_253_3228, w_253_3229, w_253_3242, w_253_3248, w_253_3255, w_253_3257, w_253_3271, w_253_3284, w_253_3302, w_253_3311, w_253_3313, w_253_3323, w_253_3335, w_253_3336, w_253_3358, w_253_3380, w_253_3390, w_253_3404, w_253_3412, w_253_3427, w_253_3431, w_253_3445, w_253_3449, w_253_3467, w_253_3473, w_253_3483, w_253_3484, w_253_3498, w_253_3512, w_253_3532, w_253_3536, w_253_3540, w_253_3548, w_253_3554, w_253_3555, w_253_3567, w_253_3581, w_253_3583, w_253_3587, w_253_3592, w_253_3594, w_253_3608, w_253_3610, w_253_3617, w_253_3637, w_253_3644, w_253_3665, w_253_3669, w_253_3685, w_253_3686, w_253_3690, w_253_3722, w_253_3723, w_253_3750, w_253_3762, w_253_3766, w_253_3786, w_253_3801, w_253_3810, w_253_3811, w_253_3832, w_253_3833, w_253_3834, w_253_3836;
  wire w_254_012, w_254_018, w_254_021, w_254_032, w_254_034, w_254_036, w_254_045, w_254_051, w_254_052, w_254_054, w_254_056, w_254_066, w_254_070, w_254_077, w_254_078, w_254_080, w_254_095, w_254_097, w_254_116, w_254_119, w_254_134, w_254_137, w_254_142, w_254_147, w_254_148, w_254_149, w_254_155, w_254_164, w_254_171, w_254_173, w_254_194, w_254_198, w_254_208, w_254_210, w_254_216, w_254_217, w_254_220, w_254_233, w_254_239, w_254_245, w_254_247, w_254_249, w_254_252, w_254_260, w_254_261, w_254_267, w_254_275, w_254_278, w_254_283, w_254_293, w_254_294, w_254_297, w_254_306, w_254_309, w_254_315, w_254_320, w_254_324, w_254_329, w_254_334, w_254_343, w_254_351, w_254_352, w_254_360, w_254_367, w_254_374, w_254_378, w_254_383, w_254_385, w_254_387, w_254_390, w_254_392, w_254_401, w_254_402, w_254_409, w_254_426, w_254_431, w_254_436, w_254_446, w_254_452, w_254_459, w_254_461, w_254_474, w_254_476, w_254_478, w_254_482, w_254_483, w_254_503, w_254_508, w_254_509, w_254_514, w_254_523, w_254_527, w_254_529, w_254_541, w_254_554, w_254_556, w_254_557, w_254_560, w_254_561, w_254_562, w_254_567, w_254_571, w_254_573, w_254_579, w_254_586, w_254_587, w_254_590, w_254_594, w_254_616, w_254_618, w_254_640, w_254_641, w_254_643, w_254_646, w_254_647, w_254_658, w_254_660, w_254_670, w_254_686, w_254_690, w_254_692, w_254_693, w_254_709, w_254_715, w_254_718, w_254_719, w_254_723, w_254_726, w_254_744, w_254_745, w_254_750, w_254_753, w_254_755, w_254_756, w_254_765, w_254_770, w_254_777, w_254_788, w_254_789, w_254_790, w_254_793, w_254_794, w_254_817, w_254_821, w_254_823, w_254_833, w_254_837, w_254_851, w_254_854, w_254_856, w_254_860, w_254_863, w_254_870, w_254_873, w_254_882, w_254_896, w_254_898, w_254_905, w_254_910, w_254_926, w_254_931, w_254_951, w_254_964, w_254_969, w_254_972, w_254_974, w_254_983, w_254_988, w_254_992, w_254_993, w_254_995, w_254_996, w_254_1023, w_254_1025, w_254_1033, w_254_1034, w_254_1036, w_254_1037, w_254_1052, w_254_1062, w_254_1087, w_254_1089, w_254_1110, w_254_1112, w_254_1114, w_254_1122, w_254_1124, w_254_1125, w_254_1137, w_254_1147, w_254_1154, w_254_1155, w_254_1177, w_254_1188, w_254_1193, w_254_1194, w_254_1200, w_254_1202, w_254_1205, w_254_1210, w_254_1230, w_254_1240, w_254_1243, w_254_1251, w_254_1252, w_254_1272, w_254_1275, w_254_1278, w_254_1287, w_254_1304, w_254_1312, w_254_1316, w_254_1318, w_254_1323, w_254_1329, w_254_1331, w_254_1339, w_254_1344, w_254_1350, w_254_1351, w_254_1354, w_254_1362, w_254_1378, w_254_1395, w_254_1396, w_254_1398, w_254_1428, w_254_1429, w_254_1447, w_254_1451, w_254_1460, w_254_1467, w_254_1479, w_254_1510, w_254_1513, w_254_1520, w_254_1529, w_254_1535, w_254_1551, w_254_1567, w_254_1570, w_254_1576, w_254_1593, w_254_1631, w_254_1635, w_254_1649, w_254_1661, w_254_1685, w_254_1698, w_254_1700, w_254_1701, w_254_1705, w_254_1711, w_254_1734, w_254_1743, w_254_1749, w_254_1773, w_254_1775, w_254_1781, w_254_1786, w_254_1789, w_254_1800, w_254_1812, w_254_1822, w_254_1835, w_254_1843, w_254_1847, w_254_1854, w_254_1865, w_254_1875, w_254_1882, w_254_1884, w_254_1897, w_254_1916, w_254_1920, w_254_1958, w_254_1959, w_254_1982, w_254_1992, w_254_1993, w_254_1994, w_254_2006, w_254_2018, w_254_2024, w_254_2031, w_254_2032, w_254_2033, w_254_2047, w_254_2062, w_254_2066, w_254_2083, w_254_2087, w_254_2095, w_254_2100, w_254_2114, w_254_2140, w_254_2154, w_254_2171, w_254_2196, w_254_2201, w_254_2220, w_254_2226, w_254_2228, w_254_2229, w_254_2239, w_254_2240, w_254_2254, w_254_2263, w_254_2271, w_254_2285, w_254_2288, w_254_2293, w_254_2304, w_254_2307, w_254_2310, w_254_2321, w_254_2323, w_254_2328, w_254_2330, w_254_2339, w_254_2351, w_254_2363, w_254_2402, w_254_2406, w_254_2413, w_254_2416, w_254_2422, w_254_2426, w_254_2432, w_254_2437, w_254_2446, w_254_2471, w_254_2485, w_254_2488, w_254_2520, w_254_2524, w_254_2534, w_254_2539, w_254_2547, w_254_2548, w_254_2554, w_254_2562, w_254_2567, w_254_2569, w_254_2573, w_254_2588, w_254_2589, w_254_2592, w_254_2600, w_254_2616, w_254_2633, w_254_2670, w_254_2674, w_254_2677, w_254_2679, w_254_2686, w_254_2687, w_254_2700, w_254_2741, w_254_2747, w_254_2748, w_254_2759, w_254_2764, w_254_2768, w_254_2790, w_254_2818, w_254_2830, w_254_2832, w_254_2847, w_254_2849, w_254_2851, w_254_2852, w_254_2865, w_254_2867, w_254_2874, w_254_2880, w_254_2891, w_254_2894, w_254_2909, w_254_2916, w_254_2923, w_254_2929, w_254_2934, w_254_2957, w_254_2962, w_254_2974, w_254_2987, w_254_2990, w_254_3006, w_254_3021, w_254_3024, w_254_3028, w_254_3035, w_254_3037, w_254_3097, w_254_3108, w_254_3115, w_254_3125, w_254_3133, w_254_3140, w_254_3149, w_254_3186, w_254_3187, w_254_3215, w_254_3227, w_254_3228, w_254_3230, w_254_3233, w_254_3247, w_254_3249, w_254_3280, w_254_3290, w_254_3300, w_254_3351, w_254_3356, w_254_3358, w_254_3362, w_254_3364, w_254_3393, w_254_3409, w_254_3430, w_254_3431, w_254_3460, w_254_3465, w_254_3481, w_254_3486, w_254_3495, w_254_3519, w_254_3526, w_254_3539, w_254_3546, w_254_3549, w_254_3565, w_254_3567, w_254_3581, w_254_3582, w_254_3589, w_254_3596, w_254_3598, w_254_3599, w_254_3600, w_254_3601, w_254_3602, w_254_3603, w_254_3604, w_254_3605, w_254_3606, w_254_3607, w_254_3611, w_254_3612, w_254_3613, w_254_3614, w_254_3615, w_254_3616, w_254_3617, w_254_3618, w_254_3619, w_254_3620, w_254_3622;
  wire w_255_002, w_255_010, w_255_021, w_255_023, w_255_024, w_255_034, w_255_036, w_255_040, w_255_041, w_255_046, w_255_047, w_255_050, w_255_051, w_255_052, w_255_054, w_255_057, w_255_061, w_255_064, w_255_065, w_255_066, w_255_067, w_255_070, w_255_071, w_255_072, w_255_073, w_255_077, w_255_085, w_255_090, w_255_091, w_255_096, w_255_098, w_255_100, w_255_106, w_255_110, w_255_111, w_255_115, w_255_117, w_255_118, w_255_123, w_255_126, w_255_127, w_255_130, w_255_131, w_255_133, w_255_136, w_255_153, w_255_161, w_255_162, w_255_166, w_255_167, w_255_169, w_255_171, w_255_172, w_255_179, w_255_180, w_255_181, w_255_194, w_255_198, w_255_200, w_255_201, w_255_206, w_255_218, w_255_220, w_255_226, w_255_227, w_255_228, w_255_231, w_255_232, w_255_238, w_255_244, w_255_248, w_255_249, w_255_251, w_255_252, w_255_253, w_255_259, w_255_266, w_255_268, w_255_274, w_255_275, w_255_278, w_255_281, w_255_283, w_255_284, w_255_291, w_255_294, w_255_296, w_255_305, w_255_312, w_255_313, w_255_317, w_255_324, w_255_325, w_255_326, w_255_331, w_255_337, w_255_339, w_255_340, w_255_342, w_255_346, w_255_350, w_255_352, w_255_357, w_255_358, w_255_359, w_255_360, w_255_362, w_255_365, w_255_368, w_255_369, w_255_373, w_255_382, w_255_383, w_255_387, w_255_389, w_255_391, w_255_394, w_255_396, w_255_397, w_255_402, w_255_403, w_255_406, w_255_414, w_255_416, w_255_418, w_255_424, w_255_427, w_255_428, w_255_429, w_255_430, w_255_431, w_255_437, w_255_438, w_255_443, w_255_445, w_255_448, w_255_452, w_255_453, w_255_455, w_255_456, w_255_457, w_255_458, w_255_459, w_255_461, w_255_464, w_255_472, w_255_478, w_255_486, w_255_489, w_255_496, w_255_501, w_255_504, w_255_505, w_255_508, w_255_514, w_255_515, w_255_519, w_255_521, w_255_523, w_255_525, w_255_526, w_255_529, w_255_535, w_255_540, w_255_543, w_255_545, w_255_562, w_255_565, w_255_569, w_255_574, w_255_575, w_255_576, w_255_578, w_255_581, w_255_582, w_255_586, w_255_588, w_255_591, w_255_593, w_255_599, w_255_604, w_255_605, w_255_608, w_255_609, w_255_610, w_255_615, w_255_619, w_255_620, w_255_624, w_255_626, w_255_629, w_255_630, w_255_632, w_255_633, w_255_637, w_255_641, w_255_643, w_255_644, w_255_650, w_255_654, w_255_656, w_255_663, w_255_665, w_255_677, w_255_678, w_255_679, w_255_701, w_255_714, w_255_717, w_255_719, w_255_726, w_255_729, w_255_736, w_255_739, w_255_741, w_255_742, w_255_743, w_255_745, w_255_746, w_255_751, w_255_752, w_255_754, w_255_757, w_255_759, w_255_760, w_255_765, w_255_768, w_255_769, w_255_771, w_255_775, w_255_779, w_255_781, w_255_785, w_255_788, w_255_791, w_255_792, w_255_796, w_255_797, w_255_798, w_255_799, w_255_800, w_255_802, w_255_804, w_255_807, w_255_808, w_255_810, w_255_814, w_255_819, w_255_823, w_255_825, w_255_829, w_255_837, w_255_840, w_255_841, w_255_842, w_255_843, w_255_845, w_255_850, w_255_853, w_255_862, w_255_863, w_255_864, w_255_866, w_255_867, w_255_869, w_255_876, w_255_877, w_255_879, w_255_896, w_255_897, w_255_898, w_255_905, w_255_910, w_255_912, w_255_914, w_255_921, w_255_923, w_255_926, w_255_928, w_255_929, w_255_931, w_255_934, w_255_936, w_255_937, w_255_944, w_255_946, w_255_947, w_255_956, w_255_965, w_255_976, w_255_987, w_255_994, w_255_1006, w_255_1018, w_255_1021, w_255_1023, w_255_1028, w_255_1029, w_255_1032, w_255_1033, w_255_1039, w_255_1043, w_255_1054, w_255_1055, w_255_1058, w_255_1063, w_255_1067, w_255_1078, w_255_1084, w_255_1092, w_255_1093, w_255_1094, w_255_1101, w_255_1103, w_255_1105, w_255_1106, w_255_1107, w_255_1108, w_255_1112, w_255_1117, w_255_1121, w_255_1122, w_255_1123, w_255_1124, w_255_1131, w_255_1136, w_255_1138, w_255_1146, w_255_1151, w_255_1152, w_255_1154, w_255_1157, w_255_1160, w_255_1162, w_255_1163, w_255_1168, w_255_1171, w_255_1173, w_255_1175, w_255_1178, w_255_1187, w_255_1189, w_255_1190, w_255_1194, w_255_1197, w_255_1200, w_255_1201, w_255_1202, w_255_1209, w_255_1210, w_255_1211, w_255_1218, w_255_1220, w_255_1221, w_255_1226, w_255_1227, w_255_1235, w_255_1241, w_255_1242, w_255_1245, w_255_1248, w_255_1252, w_255_1253, w_255_1257, w_255_1260, w_255_1263, w_255_1271, w_255_1272, w_255_1274, w_255_1278, w_255_1280, w_255_1281, w_255_1282, w_255_1283, w_255_1286, w_255_1292, w_255_1302, w_255_1306, w_255_1310, w_255_1317, w_255_1321, w_255_1325, w_255_1328, w_255_1329, w_255_1331, w_255_1332, w_255_1339, w_255_1340, w_255_1344, w_255_1345, w_255_1346, w_255_1350, w_255_1352, w_255_1353, w_255_1359, w_255_1363, w_255_1370, w_255_1372, w_255_1373, w_255_1374, w_255_1375, w_255_1378, w_255_1386, w_255_1387, w_255_1388, w_255_1389, w_255_1390, w_255_1391, w_255_1392, w_255_1393, w_255_1394, w_255_1398, w_255_1399, w_255_1400, w_255_1401, w_255_1402, w_255_1403, w_255_1404, w_255_1405, w_255_1406, w_255_1408;
  wire w_256_015, w_256_021, w_256_031, w_256_039, w_256_043, w_256_044, w_256_050, w_256_053, w_256_058, w_256_062, w_256_068, w_256_076, w_256_078, w_256_085, w_256_093, w_256_097, w_256_098, w_256_104, w_256_106, w_256_112, w_256_113, w_256_114, w_256_115, w_256_123, w_256_125, w_256_126, w_256_135, w_256_140, w_256_146, w_256_147, w_256_150, w_256_151, w_256_153, w_256_161, w_256_164, w_256_167, w_256_168, w_256_174, w_256_178, w_256_179, w_256_180, w_256_184, w_256_187, w_256_192, w_256_195, w_256_197, w_256_201, w_256_205, w_256_212, w_256_218, w_256_219, w_256_220, w_256_221, w_256_226, w_256_228, w_256_230, w_256_237, w_256_241, w_256_243, w_256_249, w_256_255, w_256_261, w_256_262, w_256_274, w_256_278, w_256_280, w_256_285, w_256_286, w_256_287, w_256_292, w_256_302, w_256_303, w_256_309, w_256_312, w_256_314, w_256_316, w_256_320, w_256_331, w_256_341, w_256_357, w_256_368, w_256_373, w_256_374, w_256_382, w_256_383, w_256_387, w_256_388, w_256_389, w_256_393, w_256_394, w_256_396, w_256_407, w_256_416, w_256_417, w_256_418, w_256_432, w_256_435, w_256_443, w_256_446, w_256_450, w_256_451, w_256_468, w_256_473, w_256_486, w_256_487, w_256_492, w_256_493, w_256_497, w_256_501, w_256_502, w_256_503, w_256_508, w_256_511, w_256_525, w_256_527, w_256_530, w_256_534, w_256_544, w_256_549, w_256_551, w_256_554, w_256_562, w_256_568, w_256_569, w_256_571, w_256_573, w_256_574, w_256_575, w_256_576, w_256_581, w_256_590, w_256_601, w_256_602, w_256_608, w_256_611, w_256_622, w_256_625, w_256_626, w_256_635, w_256_644, w_256_647, w_256_650, w_256_651, w_256_652, w_256_658, w_256_660, w_256_668, w_256_674, w_256_682, w_256_683, w_256_691, w_256_693, w_256_694, w_256_696, w_256_704, w_256_705, w_256_706, w_256_715, w_256_717, w_256_719, w_256_722, w_256_734, w_256_740, w_256_741, w_256_752, w_256_755, w_256_763, w_256_780, w_256_785, w_256_798, w_256_805, w_256_809, w_256_814, w_256_817, w_256_825, w_256_828, w_256_832, w_256_842, w_256_864, w_256_866, w_256_868, w_256_883, w_256_894, w_256_902, w_256_903, w_256_925, w_256_927, w_256_929, w_256_955, w_256_959, w_256_962, w_256_971, w_256_980, w_256_990, w_256_992, w_256_1000, w_256_1002, w_256_1005, w_256_1008, w_256_1035, w_256_1043, w_256_1045, w_256_1047, w_256_1054, w_256_1058, w_256_1065, w_256_1068, w_256_1071, w_256_1073, w_256_1074, w_256_1075, w_256_1076, w_256_1092, w_256_1099, w_256_1109, w_256_1113, w_256_1120, w_256_1131, w_256_1138, w_256_1147, w_256_1150, w_256_1158, w_256_1168, w_256_1169, w_256_1176, w_256_1193, w_256_1198, w_256_1206, w_256_1244, w_256_1252, w_256_1258, w_256_1260, w_256_1264, w_256_1269, w_256_1271, w_256_1275, w_256_1277, w_256_1279, w_256_1288, w_256_1296, w_256_1303, w_256_1309, w_256_1319, w_256_1328, w_256_1330, w_256_1332, w_256_1333, w_256_1334, w_256_1336, w_256_1358, w_256_1361, w_256_1374, w_256_1387, w_256_1388, w_256_1397, w_256_1406, w_256_1407, w_256_1411, w_256_1414, w_256_1421, w_256_1423, w_256_1426, w_256_1427, w_256_1432, w_256_1433, w_256_1439, w_256_1442, w_256_1446, w_256_1455, w_256_1461, w_256_1463, w_256_1466, w_256_1467, w_256_1472, w_256_1484, w_256_1488, w_256_1489, w_256_1492, w_256_1496, w_256_1499, w_256_1510, w_256_1518, w_256_1520, w_256_1525, w_256_1528, w_256_1529, w_256_1552, w_256_1561, w_256_1562, w_256_1568, w_256_1570, w_256_1573, w_256_1575, w_256_1599, w_256_1601, w_256_1605, w_256_1606, w_256_1607, w_256_1612, w_256_1625, w_256_1639, w_256_1646, w_256_1647, w_256_1649, w_256_1663, w_256_1664, w_256_1673, w_256_1681, w_256_1682, w_256_1683, w_256_1703, w_256_1705, w_256_1707, w_256_1711, w_256_1712, w_256_1720, w_256_1725, w_256_1726, w_256_1731, w_256_1735, w_256_1736, w_256_1748, w_256_1753, w_256_1756, w_256_1758, w_256_1761, w_256_1773, w_256_1775, w_256_1782, w_256_1795, w_256_1798, w_256_1800, w_256_1805, w_256_1809, w_256_1824, w_256_1825, w_256_1830, w_256_1831, w_256_1836, w_256_1844, w_256_1846, w_256_1847, w_256_1853, w_256_1864, w_256_1877, w_256_1878, w_256_1911, w_256_1913, w_256_1914, w_256_1917, w_256_1927, w_256_1936, w_256_1937, w_256_1947, w_256_1949, w_256_1950, w_256_1959, w_256_1986, w_256_1995, w_256_2004, w_256_2007, w_256_2020, w_256_2023, w_256_2028, w_256_2031, w_256_2038, w_256_2042, w_256_2044, w_256_2059, w_256_2060, w_256_2072, w_256_2073, w_256_2081, w_256_2083, w_256_2088, w_256_2101;
  wire w_257_000, w_257_001, w_257_002, w_257_003, w_257_004, w_257_005, w_257_006, w_257_007, w_257_008, w_257_009, w_257_010, w_257_011, w_257_012, w_257_013, w_257_014, w_257_015, w_257_016, w_257_017, w_257_019, w_257_021, w_257_023, w_257_024, w_257_025, w_257_026, w_257_027, w_257_028, w_257_029, w_257_030, w_257_031, w_257_032, w_257_033, w_257_034, w_257_035, w_257_036, w_257_037, w_257_038, w_257_039, w_257_040, w_257_041, w_257_042, w_257_043, w_257_044, w_257_045, w_257_046, w_257_047, w_257_048, w_257_049, w_257_050, w_257_051, w_257_052, w_257_053, w_257_054, w_257_055, w_257_056, w_257_057, w_257_058, w_257_059, w_257_060, w_257_061, w_257_062, w_257_063, w_257_064, w_257_065, w_257_067, w_257_068, w_257_069, w_257_070, w_257_071, w_257_072, w_257_073, w_257_074, w_257_075, w_257_076, w_257_077, w_257_078, w_257_079, w_257_080, w_257_081, w_257_082, w_257_083, w_257_084, w_257_085, w_257_086, w_257_087, w_257_088, w_257_089, w_257_090, w_257_091, w_257_092, w_257_093, w_257_094, w_257_095, w_257_096, w_257_097, w_257_098, w_257_099, w_257_100, w_257_101, w_257_102, w_257_103, w_257_104, w_257_105, w_257_106, w_257_107, w_257_108, w_257_109, w_257_110, w_257_111, w_257_112, w_257_113, w_257_114, w_257_115, w_257_116, w_257_117, w_257_119, w_257_120, w_257_121, w_257_122, w_257_123, w_257_124, w_257_125, w_257_127, w_257_129, w_257_131, w_257_132, w_257_133, w_257_135, w_257_136, w_257_137, w_257_138, w_257_139, w_257_140, w_257_141, w_257_142, w_257_143, w_257_144, w_257_145, w_257_147, w_257_148, w_257_149, w_257_151, w_257_152, w_257_153, w_257_154, w_257_156, w_257_157, w_257_158, w_257_159, w_257_160, w_257_161, w_257_163, w_257_165, w_257_167, w_257_168, w_257_169, w_257_170, w_257_171, w_257_172, w_257_173, w_257_174, w_257_175, w_257_176, w_257_178, w_257_179, w_257_180, w_257_181, w_257_182, w_257_183, w_257_184, w_257_185, w_257_186, w_257_188, w_257_189;
  wire w_258_006, w_258_009, w_258_015, w_258_044, w_258_046, w_258_047, w_258_054, w_258_059, w_258_060, w_258_064, w_258_071, w_258_092, w_258_094, w_258_101, w_258_109, w_258_111, w_258_115, w_258_119, w_258_122, w_258_123, w_258_125, w_258_131, w_258_134, w_258_136, w_258_151, w_258_152, w_258_158, w_258_159, w_258_167, w_258_170, w_258_177, w_258_179, w_258_197, w_258_203, w_258_207, w_258_215, w_258_221, w_258_231, w_258_247, w_258_262, w_258_263, w_258_265, w_258_266, w_258_273, w_258_274, w_258_285, w_258_288, w_258_293, w_258_298, w_258_302, w_258_318, w_258_321, w_258_330, w_258_333, w_258_335, w_258_343, w_258_345, w_258_362, w_258_371, w_258_384, w_258_385, w_258_386, w_258_394, w_258_401, w_258_404, w_258_424, w_258_427, w_258_428, w_258_429, w_258_443, w_258_449, w_258_452, w_258_456, w_258_470, w_258_482, w_258_483, w_258_516, w_258_518, w_258_519, w_258_520, w_258_528, w_258_529, w_258_531, w_258_532, w_258_536, w_258_541, w_258_543, w_258_545, w_258_553, w_258_554, w_258_561, w_258_562, w_258_563, w_258_571, w_258_603, w_258_606, w_258_608, w_258_615, w_258_618, w_258_623, w_258_625, w_258_627, w_258_628, w_258_635, w_258_638, w_258_642, w_258_645, w_258_653, w_258_663, w_258_685, w_258_687, w_258_692, w_258_707, w_258_708, w_258_709, w_258_712, w_258_716, w_258_732, w_258_740, w_258_742, w_258_743, w_258_746, w_258_748, w_258_750, w_258_773, w_258_774, w_258_775, w_258_786, w_258_799, w_258_803, w_258_807, w_258_809, w_258_811, w_258_813, w_258_815, w_258_825, w_258_835, w_258_839, w_258_841, w_258_847, w_258_848, w_258_854, w_258_856, w_258_857, w_258_861, w_258_863, w_258_867, w_258_873, w_258_880, w_258_898, w_258_900, w_258_902, w_258_908, w_258_912, w_258_932, w_258_938, w_258_943, w_258_945, w_258_956, w_258_959, w_258_965, w_258_969, w_258_975, w_258_976, w_258_977, w_258_996, w_258_1000, w_258_1005, w_258_1007, w_258_1009, w_258_1014, w_258_1017, w_258_1018, w_258_1028, w_258_1049, w_258_1056, w_258_1063, w_258_1075, w_258_1082, w_258_1087, w_258_1092, w_258_1094, w_258_1111, w_258_1130, w_258_1138, w_258_1142, w_258_1152, w_258_1157, w_258_1158, w_258_1160, w_258_1165, w_258_1170, w_258_1175, w_258_1178, w_258_1186, w_258_1195, w_258_1205, w_258_1207, w_258_1208, w_258_1213, w_258_1217, w_258_1227, w_258_1231, w_258_1234, w_258_1238, w_258_1253, w_258_1254, w_258_1265, w_258_1274, w_258_1283, w_258_1284, w_258_1289, w_258_1290, w_258_1300, w_258_1304, w_258_1305, w_258_1309, w_258_1320, w_258_1325, w_258_1333, w_258_1346, w_258_1349, w_258_1350, w_258_1361, w_258_1364, w_258_1379, w_258_1384, w_258_1385, w_258_1408, w_258_1409, w_258_1421, w_258_1428, w_258_1431, w_258_1442, w_258_1449, w_258_1473, w_258_1481, w_258_1485, w_258_1486, w_258_1487, w_258_1492, w_258_1495, w_258_1496, w_258_1502, w_258_1505, w_258_1507, w_258_1511, w_258_1515, w_258_1518, w_258_1527, w_258_1534, w_258_1549, w_258_1550, w_258_1562, w_258_1564, w_258_1566, w_258_1573, w_258_1576, w_258_1577, w_258_1581, w_258_1586, w_258_1589, w_258_1591, w_258_1595, w_258_1601, w_258_1619, w_258_1627, w_258_1635, w_258_1642, w_258_1644, w_258_1645, w_258_1650, w_258_1659, w_258_1660, w_258_1673, w_258_1675, w_258_1677, w_258_1678, w_258_1680, w_258_1689, w_258_1699, w_258_1703, w_258_1705, w_258_1715, w_258_1725, w_258_1736, w_258_1739, w_258_1742, w_258_1743, w_258_1744, w_258_1752, w_258_1757, w_258_1761, w_258_1774, w_258_1777, w_258_1783, w_258_1784, w_258_1799, w_258_1800, w_258_1802, w_258_1812, w_258_1814, w_258_1819, w_258_1827, w_258_1829, w_258_1841, w_258_1844, w_258_1847, w_258_1849, w_258_1856, w_258_1859, w_258_1865, w_258_1870, w_258_1874, w_258_1877, w_258_1878, w_258_1880, w_258_1884, w_258_1894, w_258_1896, w_258_1906, w_258_1909, w_258_1914, w_258_1917, w_258_1920, w_258_1921, w_258_1926, w_258_1930, w_258_1936, w_258_1946, w_258_1950, w_258_1958, w_258_1959, w_258_1969, w_258_1971, w_258_1972, w_258_1987, w_258_1988, w_258_1990, w_258_1998, w_258_2004, w_258_2005, w_258_2008, w_258_2009, w_258_2010, w_258_2014, w_258_2017, w_258_2034, w_258_2048, w_258_2049, w_258_2051, w_258_2058, w_258_2060, w_258_2063, w_258_2089, w_258_2093, w_258_2097, w_258_2105, w_258_2114, w_258_2116, w_258_2119, w_258_2122, w_258_2128, w_258_2135, w_258_2136, w_258_2144, w_258_2146, w_258_2149, w_258_2151, w_258_2155, w_258_2172, w_258_2176, w_258_2178, w_258_2184, w_258_2187, w_258_2188, w_258_2191, w_258_2192, w_258_2204, w_258_2207, w_258_2218, w_258_2220, w_258_2221, w_258_2224, w_258_2231, w_258_2237, w_258_2241, w_258_2246, w_258_2252, w_258_2257, w_258_2272, w_258_2275, w_258_2279, w_258_2285, w_258_2287, w_258_2302, w_258_2306, w_258_2309, w_258_2318, w_258_2323, w_258_2343, w_258_2349, w_258_2354, w_258_2361, w_258_2362, w_258_2363, w_258_2368, w_258_2382, w_258_2384, w_258_2399, w_258_2402, w_258_2410, w_258_2424, w_258_2427, w_258_2442, w_258_2463, w_258_2482, w_258_2489, w_258_2491, w_258_2516, w_258_2528, w_258_2598, w_258_2603, w_258_2605, w_258_2620;
  wire w_259_004, w_259_008, w_259_009, w_259_011, w_259_016, w_259_018, w_259_023, w_259_024, w_259_025, w_259_029, w_259_030, w_259_035, w_259_037, w_259_040, w_259_045, w_259_046, w_259_057, w_259_062, w_259_063, w_259_066, w_259_067, w_259_072, w_259_079, w_259_081, w_259_082, w_259_085, w_259_089, w_259_092, w_259_094, w_259_095, w_259_099, w_259_101, w_259_104, w_259_106, w_259_107, w_259_108, w_259_110, w_259_113, w_259_114, w_259_117, w_259_123, w_259_124, w_259_127, w_259_129, w_259_130, w_259_134, w_259_136, w_259_140, w_259_142, w_259_144, w_259_148, w_259_149, w_259_153, w_259_156, w_259_157, w_259_158, w_259_161, w_259_163, w_259_164, w_259_165, w_259_169, w_259_174, w_259_178, w_259_180, w_259_181, w_259_184, w_259_185, w_259_187, w_259_188, w_259_189, w_259_190, w_259_192, w_259_194, w_259_195, w_259_197, w_259_198, w_259_202, w_259_204, w_259_206, w_259_208, w_259_210, w_259_214, w_259_215, w_259_219, w_259_220, w_259_225, w_259_227, w_259_232, w_259_236, w_259_238, w_259_239, w_259_241, w_259_242, w_259_243, w_259_244, w_259_248, w_259_250, w_259_251, w_259_252, w_259_255, w_259_259, w_259_260, w_259_263, w_259_264, w_259_269, w_259_270, w_259_271, w_259_272, w_259_275, w_259_278, w_259_281, w_259_282, w_259_284, w_259_289, w_259_291, w_259_292, w_259_293, w_259_300, w_259_303, w_259_304, w_259_310, w_259_313, w_259_316, w_259_319, w_259_320, w_259_322, w_259_326, w_259_328, w_259_329, w_259_336, w_259_337, w_259_339, w_259_340, w_259_342, w_259_346, w_259_349, w_259_353, w_259_354, w_259_355, w_259_357, w_259_360, w_259_366, w_259_367, w_259_370, w_259_374, w_259_375, w_259_376, w_259_378, w_259_379, w_259_387, w_259_390, w_259_392, w_259_393, w_259_397, w_259_399, w_259_400, w_259_401, w_259_402, w_259_403, w_259_405, w_259_411, w_259_412, w_259_413, w_259_415, w_259_418, w_259_429, w_259_433, w_259_435, w_259_438, w_259_440, w_259_441, w_259_442, w_259_443, w_259_445, w_259_446, w_259_447, w_259_449, w_259_450, w_259_451, w_259_459, w_259_460, w_259_463, w_259_465, w_259_466, w_259_472, w_259_474, w_259_475, w_259_476, w_259_478, w_259_480, w_259_481, w_259_482, w_259_483, w_259_496, w_259_497, w_259_500, w_259_502, w_259_506, w_259_515, w_259_516, w_259_519, w_259_522, w_259_524, w_259_529, w_259_530, w_259_534, w_259_536, w_259_538, w_259_539, w_259_541, w_259_544, w_259_546, w_259_547, w_259_551, w_259_553, w_259_555, w_259_557, w_259_563, w_259_565, w_259_566, w_259_569, w_259_570, w_259_571, w_259_573, w_259_574, w_259_575, w_259_578, w_259_591, w_259_597, w_259_600, w_259_602, w_259_603, w_259_604, w_259_607, w_259_608, w_259_610, w_259_612, w_259_614, w_259_617, w_259_619, w_259_620, w_259_621, w_259_622, w_259_626, w_259_634, w_259_639, w_259_641, w_259_642, w_259_643, w_259_644, w_259_645, w_259_647, w_259_653, w_259_654, w_259_656, w_259_668, w_259_675, w_259_677, w_259_680, w_259_682, w_259_683, w_259_685, w_259_688, w_259_693, w_259_697, w_259_698, w_259_703, w_259_705, w_259_706, w_259_709, w_259_717, w_259_718, w_259_723, w_259_724, w_259_725, w_259_730, w_259_732, w_259_738, w_259_740, w_259_742, w_259_747, w_259_749, w_259_754, w_259_758, w_259_762, w_259_764, w_259_770, w_259_773, w_259_776, w_259_777, w_259_778, w_259_779, w_259_782, w_259_785, w_259_788, w_259_789, w_259_791, w_259_796, w_259_797, w_259_800, w_259_808, w_259_811, w_259_812, w_259_815, w_259_816, w_259_824, w_259_825, w_259_826, w_259_827, w_259_828, w_259_829, w_259_834, w_259_836, w_259_838, w_259_848, w_259_850, w_259_854, w_259_857, w_259_861, w_259_863, w_259_868, w_259_870, w_259_876, w_259_881, w_259_882, w_259_886, w_259_888, w_259_889, w_259_891, w_259_893, w_259_894, w_259_895, w_259_897, w_259_898, w_259_901, w_259_904, w_259_906, w_259_907, w_259_908, w_259_910, w_259_914, w_259_917, w_259_918, w_259_921, w_259_925, w_259_927, w_259_929, w_259_933, w_259_941, w_259_943, w_259_945, w_259_946, w_259_949, w_259_951, w_259_954, w_259_955, w_259_957, w_259_959, w_259_961, w_259_962, w_259_963, w_259_965, w_259_966, w_259_969, w_259_971, w_259_974, w_259_979, w_259_983, w_259_988, w_259_989, w_259_991, w_259_992, w_259_995, w_259_996;
  wire w_260_000, w_260_001, w_260_002, w_260_006, w_260_012, w_260_020, w_260_026, w_260_027, w_260_028, w_260_029, w_260_030, w_260_034, w_260_035, w_260_040, w_260_045, w_260_058, w_260_059, w_260_061, w_260_065, w_260_066, w_260_072, w_260_074, w_260_080, w_260_087, w_260_088, w_260_096, w_260_097, w_260_106, w_260_112, w_260_124, w_260_126, w_260_127, w_260_130, w_260_132, w_260_136, w_260_137, w_260_146, w_260_148, w_260_151, w_260_158, w_260_161, w_260_164, w_260_167, w_260_168, w_260_175, w_260_178, w_260_183, w_260_184, w_260_185, w_260_191, w_260_193, w_260_194, w_260_199, w_260_202, w_260_205, w_260_217, w_260_220, w_260_227, w_260_231, w_260_236, w_260_241, w_260_246, w_260_249, w_260_254, w_260_261, w_260_282, w_260_288, w_260_292, w_260_300, w_260_303, w_260_306, w_260_311, w_260_319, w_260_322, w_260_326, w_260_329, w_260_340, w_260_341, w_260_342, w_260_351, w_260_353, w_260_354, w_260_357, w_260_362, w_260_367, w_260_370, w_260_381, w_260_382, w_260_385, w_260_388, w_260_391, w_260_409, w_260_410, w_260_414, w_260_422, w_260_425, w_260_426, w_260_433, w_260_435, w_260_440, w_260_443, w_260_445, w_260_446, w_260_450, w_260_455, w_260_463, w_260_464, w_260_468, w_260_469, w_260_472, w_260_475, w_260_482, w_260_484, w_260_488, w_260_495, w_260_499, w_260_522, w_260_529, w_260_534, w_260_535, w_260_536, w_260_537, w_260_544, w_260_545, w_260_550, w_260_553, w_260_554, w_260_556, w_260_559, w_260_560, w_260_564, w_260_567, w_260_568, w_260_569, w_260_571, w_260_575, w_260_580, w_260_582, w_260_588, w_260_592, w_260_602, w_260_609, w_260_620, w_260_623, w_260_624, w_260_632, w_260_635, w_260_637, w_260_645, w_260_648, w_260_660, w_260_666, w_260_668, w_260_672, w_260_674, w_260_675, w_260_676, w_260_678, w_260_691, w_260_694, w_260_695, w_260_704, w_260_707, w_260_715, w_260_717, w_260_718, w_260_724, w_260_733, w_260_751, w_260_765, w_260_769, w_260_771, w_260_778, w_260_783, w_260_785, w_260_796, w_260_797, w_260_801, w_260_802, w_260_804, w_260_805, w_260_815, w_260_818, w_260_828, w_260_829, w_260_830, w_260_835, w_260_872, w_260_873, w_260_877, w_260_884, w_260_896, w_260_909, w_260_920, w_260_925, w_260_935, w_260_937, w_260_942, w_260_943, w_260_947, w_260_951, w_260_955, w_260_968, w_260_977, w_260_982, w_260_984, w_260_991, w_260_993, w_260_995, w_260_1017, w_260_1020, w_260_1030, w_260_1032, w_260_1035, w_260_1040, w_260_1043, w_260_1044, w_260_1051, w_260_1053, w_260_1056, w_260_1068, w_260_1072, w_260_1073, w_260_1079, w_260_1083, w_260_1095, w_260_1107, w_260_1109, w_260_1116, w_260_1122, w_260_1124, w_260_1125, w_260_1129, w_260_1137, w_260_1139, w_260_1149, w_260_1156, w_260_1163, w_260_1164, w_260_1176, w_260_1188, w_260_1193, w_260_1205, w_260_1206, w_260_1208, w_260_1212, w_260_1213, w_260_1218, w_260_1221, w_260_1229, w_260_1231, w_260_1233, w_260_1241, w_260_1242, w_260_1247, w_260_1258, w_260_1259, w_260_1262, w_260_1265, w_260_1272, w_260_1277, w_260_1280, w_260_1281, w_260_1285, w_260_1286, w_260_1293, w_260_1306, w_260_1316, w_260_1318, w_260_1327, w_260_1332, w_260_1335, w_260_1343, w_260_1344, w_260_1351, w_260_1368, w_260_1369, w_260_1375, w_260_1376, w_260_1379, w_260_1381, w_260_1386, w_260_1405, w_260_1408, w_260_1414, w_260_1416, w_260_1429, w_260_1434, w_260_1437, w_260_1438, w_260_1440, w_260_1443, w_260_1461, w_260_1465, w_260_1466, w_260_1467, w_260_1471, w_260_1482, w_260_1484, w_260_1493, w_260_1494, w_260_1497, w_260_1517, w_260_1526, w_260_1537, w_260_1544, w_260_1548, w_260_1556, w_260_1563, w_260_1566, w_260_1567, w_260_1569, w_260_1581, w_260_1587, w_260_1595, w_260_1597, w_260_1598, w_260_1599, w_260_1609, w_260_1611, w_260_1616, w_260_1622, w_260_1626, w_260_1628, w_260_1638, w_260_1662, w_260_1667, w_260_1675, w_260_1681, w_260_1686, w_260_1691, w_260_1694, w_260_1710, w_260_1717, w_260_1721, w_260_1736, w_260_1737, w_260_1753, w_260_1755, w_260_1768, w_260_1773, w_260_1775, w_260_1777, w_260_1779, w_260_1782, w_260_1789, w_260_1793, w_260_1797, w_260_1802, w_260_1808, w_260_1810, w_260_1829, w_260_1847, w_260_1852, w_260_1858, w_260_1870, w_260_1873, w_260_1874, w_260_1883, w_260_1886, w_260_1896, w_260_1902, w_260_1905, w_260_1906, w_260_1914, w_260_1917, w_260_1922, w_260_1925, w_260_1926, w_260_1928, w_260_1933, w_260_1936, w_260_1958, w_260_1969, w_260_1977, w_260_1986, w_260_1988, w_260_1994, w_260_1995, w_260_1996, w_260_2016, w_260_2019, w_260_2027, w_260_2030, w_260_2035, w_260_2039, w_260_2042, w_260_2054, w_260_2060, w_260_2065, w_260_2067, w_260_2077, w_260_2078, w_260_2085, w_260_2093, w_260_2099, w_260_2101, w_260_2107, w_260_2108;
  wire w_261_001, w_261_006, w_261_010, w_261_011, w_261_012, w_261_013, w_261_014, w_261_016, w_261_018, w_261_020, w_261_022, w_261_023, w_261_025, w_261_027, w_261_028, w_261_029, w_261_030, w_261_031, w_261_033, w_261_034, w_261_037, w_261_041, w_261_048, w_261_050, w_261_055, w_261_056, w_261_057, w_261_061, w_261_062, w_261_068, w_261_069, w_261_070, w_261_071, w_261_072, w_261_073, w_261_074, w_261_075, w_261_077, w_261_078, w_261_081, w_261_082, w_261_088, w_261_095, w_261_098, w_261_100, w_261_101, w_261_103, w_261_107, w_261_108, w_261_110, w_261_112, w_261_113, w_261_114, w_261_115, w_261_120, w_261_125, w_261_132, w_261_133, w_261_136, w_261_145, w_261_146, w_261_148, w_261_153, w_261_154, w_261_155, w_261_156, w_261_157, w_261_166, w_261_167, w_261_168, w_261_169, w_261_170, w_261_171, w_261_172, w_261_174, w_261_177, w_261_178, w_261_179, w_261_180, w_261_185, w_261_187, w_261_190, w_261_192, w_261_193, w_261_195, w_261_198, w_261_199, w_261_201, w_261_202, w_261_203, w_261_205, w_261_206, w_261_207, w_261_208, w_261_209, w_261_210, w_261_211, w_261_213, w_261_215, w_261_217, w_261_220, w_261_221, w_261_226, w_261_229, w_261_231, w_261_232, w_261_234, w_261_242, w_261_250, w_261_251, w_261_252, w_261_260, w_261_262, w_261_263, w_261_267, w_261_270, w_261_272, w_261_274, w_261_275, w_261_276, w_261_278, w_261_282, w_261_284, w_261_289, w_261_291, w_261_292, w_261_295, w_261_298, w_261_304, w_261_306, w_261_307, w_261_308, w_261_311, w_261_315, w_261_316, w_261_317, w_261_325, w_261_329, w_261_334, w_261_338, w_261_340, w_261_343, w_261_345, w_261_351, w_261_354, w_261_355, w_261_357, w_261_361, w_261_365, w_261_366, w_261_374, w_261_376, w_261_379, w_261_380, w_261_381, w_261_382, w_261_384, w_261_388, w_261_400, w_261_407, w_261_409, w_261_411, w_261_413, w_261_415, w_261_418, w_261_419, w_261_420, w_261_421, w_261_423, w_261_428, w_261_430, w_261_432, w_261_434, w_261_435, w_261_436, w_261_437, w_261_438, w_261_440, w_261_442, w_261_448, w_261_451, w_261_455, w_261_458, w_261_460, w_261_461, w_261_462, w_261_463, w_261_464, w_261_466, w_261_468, w_261_469, w_261_476, w_261_478, w_261_480, w_261_481, w_261_483, w_261_487, w_261_490, w_261_494, w_261_495, w_261_496, w_261_497, w_261_498, w_261_499, w_261_500, w_261_501, w_261_504, w_261_505, w_261_506, w_261_508, w_261_511, w_261_514, w_261_515, w_261_518, w_261_519, w_261_520, w_261_522, w_261_529, w_261_538, w_261_544, w_261_545, w_261_548, w_261_550, w_261_551, w_261_553, w_261_556, w_261_560, w_261_562, w_261_564, w_261_565, w_261_566, w_261_569, w_261_574, w_261_576, w_261_584, w_261_587, w_261_591, w_261_592, w_261_595, w_261_600, w_261_603, w_261_604, w_261_608, w_261_612, w_261_613, w_261_614, w_261_617, w_261_618, w_261_619, w_261_620, w_261_623, w_261_624, w_261_626, w_261_631, w_261_643, w_261_644, w_261_647, w_261_650, w_261_653, w_261_654, w_261_655, w_261_656, w_261_657, w_261_659, w_261_662, w_261_664, w_261_666, w_261_667, w_261_677, w_261_679, w_261_683, w_261_684, w_261_685, w_261_689, w_261_700, w_261_701, w_261_705, w_261_708, w_261_712, w_261_713, w_261_714, w_261_715, w_261_718, w_261_719, w_261_723, w_261_724, w_261_731, w_261_734, w_261_738, w_261_743, w_261_745, w_261_746, w_261_750, w_261_752, w_261_755, w_261_757, w_261_759, w_261_760, w_261_761, w_261_763, w_261_775, w_261_776, w_261_778, w_261_780, w_261_783, w_261_785, w_261_793, w_261_794, w_261_797, w_261_800, w_261_808, w_261_812, w_261_816, w_261_826, w_261_828, w_261_830, w_261_832, w_261_833, w_261_836, w_261_839, w_261_840, w_261_842, w_261_844, w_261_845, w_261_849, w_261_851, w_261_852, w_261_856, w_261_862, w_261_864, w_261_867, w_261_869, w_261_870, w_261_871, w_261_881, w_261_882, w_261_884, w_261_888, w_261_889, w_261_891, w_261_894, w_261_896, w_261_899, w_261_903, w_261_904, w_261_909, w_261_911, w_261_914, w_261_923, w_261_925, w_261_936, w_261_940, w_261_942;
  wire w_262_000, w_262_002, w_262_003, w_262_004, w_262_015, w_262_020, w_262_022, w_262_051, w_262_062, w_262_077, w_262_080, w_262_087, w_262_111, w_262_113, w_262_116, w_262_124, w_262_125, w_262_129, w_262_130, w_262_135, w_262_138, w_262_146, w_262_147, w_262_149, w_262_169, w_262_172, w_262_176, w_262_179, w_262_182, w_262_190, w_262_192, w_262_197, w_262_199, w_262_200, w_262_210, w_262_214, w_262_215, w_262_220, w_262_228, w_262_240, w_262_242, w_262_243, w_262_246, w_262_249, w_262_253, w_262_259, w_262_260, w_262_264, w_262_265, w_262_268, w_262_273, w_262_276, w_262_282, w_262_288, w_262_289, w_262_291, w_262_316, w_262_319, w_262_320, w_262_321, w_262_324, w_262_328, w_262_332, w_262_334, w_262_348, w_262_355, w_262_364, w_262_375, w_262_389, w_262_397, w_262_407, w_262_412, w_262_416, w_262_418, w_262_421, w_262_422, w_262_423, w_262_428, w_262_437, w_262_442, w_262_445, w_262_455, w_262_483, w_262_494, w_262_495, w_262_500, w_262_501, w_262_517, w_262_518, w_262_519, w_262_531, w_262_536, w_262_538, w_262_543, w_262_544, w_262_550, w_262_562, w_262_564, w_262_569, w_262_578, w_262_579, w_262_586, w_262_588, w_262_591, w_262_595, w_262_601, w_262_627, w_262_636, w_262_643, w_262_644, w_262_645, w_262_649, w_262_653, w_262_656, w_262_664, w_262_665, w_262_673, w_262_677, w_262_680, w_262_687, w_262_688, w_262_696, w_262_700, w_262_704, w_262_712, w_262_723, w_262_736, w_262_746, w_262_751, w_262_756, w_262_758, w_262_760, w_262_771, w_262_787, w_262_789, w_262_791, w_262_800, w_262_801, w_262_808, w_262_811, w_262_815, w_262_816, w_262_830, w_262_841, w_262_846, w_262_867, w_262_874, w_262_883, w_262_884, w_262_896, w_262_901, w_262_902, w_262_909, w_262_912, w_262_914, w_262_924, w_262_937, w_262_941, w_262_945, w_262_953, w_262_963, w_262_969, w_262_979, w_262_1001, w_262_1010, w_262_1028, w_262_1035, w_262_1057, w_262_1063, w_262_1119, w_262_1126, w_262_1130, w_262_1139, w_262_1145, w_262_1151, w_262_1153, w_262_1166, w_262_1171, w_262_1207, w_262_1233, w_262_1247, w_262_1249, w_262_1251, w_262_1263, w_262_1269, w_262_1279, w_262_1285, w_262_1288, w_262_1291, w_262_1319, w_262_1333, w_262_1356, w_262_1371, w_262_1400, w_262_1401, w_262_1430, w_262_1433, w_262_1447, w_262_1452, w_262_1469, w_262_1473, w_262_1503, w_262_1548, w_262_1568, w_262_1571, w_262_1591, w_262_1592, w_262_1596, w_262_1604, w_262_1609, w_262_1611, w_262_1619, w_262_1651, w_262_1661, w_262_1669, w_262_1676, w_262_1686, w_262_1692, w_262_1710, w_262_1724, w_262_1730, w_262_1745, w_262_1769, w_262_1780, w_262_1781, w_262_1785, w_262_1792, w_262_1794, w_262_1805, w_262_1806, w_262_1808, w_262_1852, w_262_1855, w_262_1859, w_262_1861, w_262_1876, w_262_1885, w_262_1899, w_262_1900, w_262_1903, w_262_1926, w_262_1947, w_262_1960, w_262_1982, w_262_1983, w_262_1993, w_262_1999, w_262_2004, w_262_2015, w_262_2021, w_262_2039, w_262_2042, w_262_2043, w_262_2045, w_262_2058, w_262_2061, w_262_2066, w_262_2075, w_262_2080, w_262_2096, w_262_2104, w_262_2117, w_262_2141, w_262_2144, w_262_2148, w_262_2154, w_262_2185, w_262_2191, w_262_2215, w_262_2218, w_262_2222, w_262_2226, w_262_2238, w_262_2253, w_262_2258, w_262_2261, w_262_2266, w_262_2281, w_262_2296, w_262_2299, w_262_2302, w_262_2308, w_262_2319, w_262_2322, w_262_2340, w_262_2342, w_262_2373, w_262_2378, w_262_2381, w_262_2388, w_262_2407, w_262_2440, w_262_2442, w_262_2449, w_262_2460, w_262_2461, w_262_2468, w_262_2472, w_262_2479, w_262_2491, w_262_2504, w_262_2512, w_262_2518, w_262_2519, w_262_2526, w_262_2551, w_262_2553, w_262_2569, w_262_2572, w_262_2578, w_262_2581, w_262_2588, w_262_2615, w_262_2628, w_262_2638, w_262_2639, w_262_2646, w_262_2675, w_262_2679, w_262_2683, w_262_2688, w_262_2689, w_262_2721, w_262_2724, w_262_2730, w_262_2738, w_262_2743, w_262_2757, w_262_2759, w_262_2772, w_262_2774, w_262_2778, w_262_2793, w_262_2798, w_262_2817, w_262_2822, w_262_2823, w_262_2836, w_262_2840, w_262_2857, w_262_2885, w_262_2891, w_262_2899, w_262_2919, w_262_2931, w_262_2951, w_262_2959, w_262_2976, w_262_2980, w_262_2981, w_262_2998, w_262_3008, w_262_3042, w_262_3054, w_262_3072, w_262_3090, w_262_3095, w_262_3111, w_262_3129, w_262_3132, w_262_3135, w_262_3170, w_262_3182, w_262_3189, w_262_3272, w_262_3284, w_262_3296, w_262_3303, w_262_3337, w_262_3357, w_262_3387, w_262_3396, w_262_3400, w_262_3401, w_262_3403, w_262_3405, w_262_3418, w_262_3421, w_262_3430, w_262_3444, w_262_3445, w_262_3449, w_262_3450, w_262_3465, w_262_3483, w_262_3487, w_262_3496, w_262_3535, w_262_3537, w_262_3562, w_262_3592, w_262_3599, w_262_3607, w_262_3634, w_262_3641, w_262_3659, w_262_3660, w_262_3680, w_262_3683, w_262_3684, w_262_3701, w_262_3705, w_262_3730, w_262_3740, w_262_3745, w_262_3746, w_262_3755, w_262_3756, w_262_3766, w_262_3792, w_262_3793, w_262_3796, w_262_3802, w_262_3804, w_262_3823, w_262_3829, w_262_3831, w_262_3840, w_262_3845, w_262_3848, w_262_3861, w_262_3884, w_262_3898, w_262_3924, w_262_3936, w_262_3949, w_262_3955, w_262_3989, w_262_3992, w_262_4018, w_262_4020, w_262_4024, w_262_4026;
  wire w_263_000, w_263_002, w_263_003, w_263_007, w_263_008, w_263_011, w_263_014, w_263_015, w_263_016, w_263_018, w_263_019, w_263_020, w_263_021, w_263_023, w_263_024, w_263_025, w_263_027, w_263_028, w_263_029, w_263_034, w_263_035, w_263_037, w_263_038, w_263_040, w_263_041, w_263_042, w_263_043, w_263_044, w_263_046, w_263_048, w_263_053, w_263_055, w_263_059, w_263_060, w_263_063, w_263_066, w_263_069, w_263_070, w_263_073, w_263_074, w_263_075, w_263_076, w_263_077, w_263_078, w_263_080, w_263_082, w_263_083, w_263_084, w_263_085, w_263_087, w_263_089, w_263_090, w_263_091, w_263_094, w_263_096, w_263_100, w_263_103, w_263_104, w_263_106, w_263_108, w_263_110, w_263_111, w_263_112, w_263_113, w_263_115, w_263_116, w_263_117, w_263_118, w_263_119, w_263_121, w_263_125, w_263_126, w_263_130, w_263_133, w_263_135, w_263_136, w_263_138, w_263_139, w_263_142, w_263_144, w_263_146, w_263_147, w_263_148, w_263_150, w_263_152, w_263_153, w_263_154, w_263_158, w_263_159, w_263_161, w_263_162, w_263_165, w_263_166, w_263_168, w_263_171, w_263_174, w_263_175, w_263_176, w_263_178, w_263_179, w_263_180, w_263_182, w_263_184, w_263_186, w_263_187, w_263_191, w_263_192, w_263_193, w_263_194, w_263_195, w_263_196, w_263_200, w_263_201, w_263_203, w_263_204, w_263_205, w_263_206, w_263_207, w_263_208, w_263_209, w_263_210, w_263_213, w_263_215, w_263_216, w_263_217, w_263_218, w_263_219, w_263_220, w_263_222, w_263_223, w_263_224, w_263_227, w_263_228, w_263_229, w_263_232, w_263_233, w_263_236, w_263_237, w_263_240, w_263_242, w_263_243, w_263_244, w_263_245, w_263_246, w_263_247, w_263_250, w_263_251, w_263_252, w_263_255, w_263_258, w_263_260, w_263_262, w_263_263, w_263_265, w_263_267, w_263_268, w_263_269, w_263_271, w_263_273, w_263_275, w_263_277, w_263_280, w_263_282, w_263_283, w_263_287, w_263_290, w_263_291, w_263_293, w_263_294, w_263_295, w_263_296, w_263_297, w_263_303, w_263_304, w_263_307, w_263_308, w_263_310, w_263_311, w_263_312, w_263_313, w_263_314, w_263_315, w_263_316, w_263_319, w_263_321, w_263_323, w_263_327, w_263_328, w_263_330, w_263_332, w_263_334, w_263_335, w_263_336, w_263_338, w_263_340, w_263_343, w_263_345, w_263_346, w_263_347, w_263_348, w_263_349, w_263_350, w_263_353, w_263_354, w_263_356, w_263_357, w_263_359, w_263_360, w_263_361, w_263_362, w_263_363, w_263_367, w_263_368, w_263_370, w_263_371, w_263_372, w_263_373, w_263_374, w_263_375, w_263_376, w_263_377, w_263_378, w_263_379, w_263_380, w_263_382, w_263_383, w_263_384, w_263_386, w_263_387, w_263_388, w_263_389, w_263_390, w_263_392, w_263_393, w_263_394, w_263_396, w_263_397, w_263_399, w_263_401, w_263_402, w_263_406, w_263_408, w_263_410, w_263_411, w_263_412, w_263_413, w_263_417, w_263_419, w_263_420, w_263_424, w_263_430, w_263_433, w_263_434, w_263_435, w_263_436, w_263_437, w_263_442, w_263_444, w_263_447, w_263_448, w_263_449, w_263_451, w_263_454, w_263_455, w_263_457, w_263_459, w_263_460, w_263_461, w_263_463, w_263_464, w_263_466, w_263_469, w_263_470, w_263_472, w_263_478, w_263_479, w_263_480, w_263_485, w_263_486, w_263_488, w_263_490, w_263_491, w_263_492, w_263_493, w_263_494, w_263_495, w_263_498, w_263_499, w_263_500, w_263_501, w_263_503, w_263_504, w_263_507, w_263_508, w_263_510, w_263_513, w_263_514, w_263_515, w_263_516, w_263_518, w_263_523, w_263_524, w_263_525, w_263_526, w_263_527, w_263_529, w_263_533, w_263_535, w_263_536, w_263_537, w_263_539, w_263_540, w_263_542, w_263_546, w_263_547, w_263_548, w_263_551, w_263_552, w_263_554, w_263_556, w_263_557, w_263_561, w_263_562, w_263_563, w_263_566, w_263_567, w_263_570, w_263_571, w_263_572, w_263_574, w_263_576, w_263_577, w_263_579, w_263_580, w_263_581, w_263_582, w_263_583, w_263_584, w_263_585, w_263_586, w_263_587, w_263_588, w_263_589;
  wire w_264_000, w_264_002, w_264_005, w_264_006, w_264_007, w_264_010, w_264_013, w_264_014, w_264_018, w_264_019, w_264_020, w_264_025, w_264_026, w_264_027, w_264_031, w_264_032, w_264_039, w_264_043, w_264_045, w_264_048, w_264_049, w_264_051, w_264_067, w_264_075, w_264_079, w_264_085, w_264_091, w_264_094, w_264_096, w_264_099, w_264_102, w_264_103, w_264_104, w_264_108, w_264_116, w_264_121, w_264_130, w_264_131, w_264_132, w_264_135, w_264_139, w_264_143, w_264_163, w_264_166, w_264_168, w_264_177, w_264_182, w_264_190, w_264_193, w_264_196, w_264_199, w_264_207, w_264_211, w_264_213, w_264_216, w_264_218, w_264_226, w_264_231, w_264_240, w_264_243, w_264_247, w_264_254, w_264_257, w_264_260, w_264_267, w_264_272, w_264_273, w_264_279, w_264_283, w_264_290, w_264_293, w_264_297, w_264_299, w_264_301, w_264_307, w_264_310, w_264_314, w_264_320, w_264_321, w_264_323, w_264_325, w_264_333, w_264_344, w_264_345, w_264_348, w_264_359, w_264_365, w_264_370, w_264_371, w_264_374, w_264_377, w_264_395, w_264_400, w_264_408, w_264_410, w_264_414, w_264_416, w_264_417, w_264_419, w_264_427, w_264_428, w_264_432, w_264_444, w_264_446, w_264_447, w_264_448, w_264_465, w_264_467, w_264_468, w_264_470, w_264_471, w_264_476, w_264_478, w_264_482, w_264_483, w_264_486, w_264_495, w_264_496, w_264_497, w_264_501, w_264_503, w_264_504, w_264_505, w_264_508, w_264_515, w_264_519, w_264_521, w_264_527, w_264_534, w_264_536, w_264_537, w_264_540, w_264_545, w_264_555, w_264_559, w_264_560, w_264_569, w_264_573, w_264_575, w_264_578, w_264_581, w_264_585, w_264_586, w_264_602, w_264_611, w_264_614, w_264_622, w_264_625, w_264_632, w_264_634, w_264_637, w_264_643, w_264_649, w_264_657, w_264_663, w_264_669, w_264_678, w_264_679, w_264_680, w_264_681, w_264_688, w_264_691, w_264_692, w_264_699, w_264_700, w_264_706, w_264_717, w_264_721, w_264_725, w_264_726, w_264_730, w_264_735, w_264_747, w_264_748, w_264_752, w_264_753, w_264_754, w_264_755, w_264_757, w_264_760, w_264_763, w_264_768, w_264_772, w_264_778, w_264_781, w_264_787, w_264_788, w_264_793, w_264_797, w_264_802, w_264_812, w_264_813, w_264_815, w_264_817, w_264_818, w_264_819, w_264_820, w_264_825, w_264_826, w_264_831, w_264_834, w_264_836, w_264_837, w_264_840, w_264_843, w_264_849, w_264_859, w_264_865, w_264_867, w_264_868, w_264_869, w_264_872, w_264_880, w_264_883, w_264_884, w_264_895, w_264_896, w_264_904, w_264_907, w_264_909, w_264_910, w_264_915, w_264_922, w_264_925, w_264_926, w_264_927, w_264_938, w_264_946, w_264_951, w_264_955, w_264_957, w_264_959, w_264_966, w_264_970, w_264_973, w_264_974, w_264_977, w_264_978, w_264_984, w_264_985, w_264_991, w_264_1002, w_264_1004, w_264_1008, w_264_1010, w_264_1014, w_264_1016, w_264_1020, w_264_1022, w_264_1031, w_264_1038, w_264_1045, w_264_1047, w_264_1062, w_264_1067, w_264_1068, w_264_1070, w_264_1079, w_264_1080, w_264_1083, w_264_1086, w_264_1088, w_264_1090, w_264_1092, w_264_1095, w_264_1109, w_264_1113, w_264_1122, w_264_1130, w_264_1136, w_264_1144, w_264_1147, w_264_1150, w_264_1153, w_264_1156, w_264_1160, w_264_1161, w_264_1162, w_264_1164, w_264_1167, w_264_1168, w_264_1170, w_264_1171, w_264_1188, w_264_1196, w_264_1206, w_264_1212, w_264_1214, w_264_1219, w_264_1222, w_264_1223, w_264_1227, w_264_1228, w_264_1242, w_264_1246, w_264_1249, w_264_1258, w_264_1264, w_264_1265, w_264_1266, w_264_1267, w_264_1280, w_264_1283, w_264_1284, w_264_1292, w_264_1300, w_264_1302, w_264_1315, w_264_1319, w_264_1327, w_264_1332, w_264_1342, w_264_1344, w_264_1347, w_264_1356, w_264_1362, w_264_1364, w_264_1365, w_264_1371, w_264_1372, w_264_1373, w_264_1375, w_264_1376, w_264_1378, w_264_1380, w_264_1382, w_264_1387, w_264_1390, w_264_1394, w_264_1401, w_264_1406, w_264_1413, w_264_1415, w_264_1417, w_264_1418, w_264_1420, w_264_1423, w_264_1434, w_264_1435, w_264_1436, w_264_1437, w_264_1444, w_264_1446, w_264_1449, w_264_1454, w_264_1455, w_264_1460, w_264_1466, w_264_1472, w_264_1478, w_264_1486, w_264_1493, w_264_1497, w_264_1500, w_264_1503, w_264_1506, w_264_1511, w_264_1516, w_264_1518, w_264_1519, w_264_1520, w_264_1526, w_264_1539, w_264_1548, w_264_1555, w_264_1556, w_264_1568, w_264_1569, w_264_1578, w_264_1580, w_264_1581, w_264_1588, w_264_1593, w_264_1595, w_264_1604, w_264_1606, w_264_1617, w_264_1624, w_264_1631, w_264_1634, w_264_1637, w_264_1647, w_264_1649, w_264_1654, w_264_1661, w_264_1676, w_264_1683, w_264_1685, w_264_1687, w_264_1688, w_264_1692, w_264_1696, w_264_1704, w_264_1706, w_264_1715, w_264_1717, w_264_1723, w_264_1725, w_264_1735, w_264_1738, w_264_1746, w_264_1753, w_264_1755, w_264_1764, w_264_1765, w_264_1770, w_264_1771, w_264_1772, w_264_1773, w_264_1774, w_264_1775, w_264_1779, w_264_1780, w_264_1781, w_264_1782, w_264_1783, w_264_1784, w_264_1785, w_264_1786, w_264_1787, w_264_1788, w_264_1790;
  wire w_265_000, w_265_002, w_265_005, w_265_006, w_265_007, w_265_010, w_265_011, w_265_016, w_265_018, w_265_020, w_265_021, w_265_024, w_265_026, w_265_027, w_265_029, w_265_033, w_265_034, w_265_036, w_265_037, w_265_038, w_265_039, w_265_041, w_265_042, w_265_043, w_265_045, w_265_046, w_265_047, w_265_048, w_265_051, w_265_052, w_265_055, w_265_056, w_265_060, w_265_063, w_265_066, w_265_067, w_265_071, w_265_072, w_265_073, w_265_074, w_265_075, w_265_077, w_265_080, w_265_082, w_265_086, w_265_087, w_265_089, w_265_090, w_265_091, w_265_093, w_265_095, w_265_101, w_265_104, w_265_107, w_265_108, w_265_109, w_265_110, w_265_113, w_265_118, w_265_121, w_265_123, w_265_124, w_265_126, w_265_131, w_265_132, w_265_133, w_265_134, w_265_137, w_265_141, w_265_142, w_265_144, w_265_148, w_265_149, w_265_150, w_265_152, w_265_153, w_265_154, w_265_155, w_265_157, w_265_158, w_265_159, w_265_162, w_265_163, w_265_165, w_265_167, w_265_178, w_265_179, w_265_182, w_265_183, w_265_186, w_265_188, w_265_195, w_265_196, w_265_201, w_265_202, w_265_203, w_265_211, w_265_215, w_265_216, w_265_217, w_265_221, w_265_222, w_265_225, w_265_227, w_265_228, w_265_230, w_265_231, w_265_233, w_265_234, w_265_235, w_265_237, w_265_242, w_265_243, w_265_251, w_265_252, w_265_255, w_265_257, w_265_258, w_265_260, w_265_261, w_265_262, w_265_266, w_265_267, w_265_269, w_265_272, w_265_275, w_265_277, w_265_279, w_265_283, w_265_287, w_265_289, w_265_290, w_265_292, w_265_293, w_265_300, w_265_301, w_265_303, w_265_306, w_265_309, w_265_313, w_265_314, w_265_318, w_265_321, w_265_323, w_265_327, w_265_330, w_265_331, w_265_335, w_265_342, w_265_344, w_265_345, w_265_350, w_265_354, w_265_355, w_265_356, w_265_357, w_265_358, w_265_361, w_265_362, w_265_363, w_265_366, w_265_367, w_265_369, w_265_370, w_265_375, w_265_380, w_265_383, w_265_388, w_265_392, w_265_393, w_265_394, w_265_399, w_265_400, w_265_401, w_265_403, w_265_405, w_265_407, w_265_409, w_265_410, w_265_411, w_265_412, w_265_413, w_265_414, w_265_416, w_265_417, w_265_418, w_265_419, w_265_420, w_265_421, w_265_423, w_265_428, w_265_431, w_265_432, w_265_433, w_265_438, w_265_440, w_265_442, w_265_443, w_265_449, w_265_451, w_265_452, w_265_453, w_265_455, w_265_460, w_265_463, w_265_468, w_265_469, w_265_471, w_265_473, w_265_474, w_265_475, w_265_477, w_265_481, w_265_484, w_265_485, w_265_486, w_265_487, w_265_488, w_265_493, w_265_495, w_265_496, w_265_497, w_265_499, w_265_500, w_265_503, w_265_504, w_265_505, w_265_507, w_265_513, w_265_516, w_265_525, w_265_526, w_265_527, w_265_536, w_265_537, w_265_538, w_265_540, w_265_545, w_265_547, w_265_548, w_265_550, w_265_551, w_265_553, w_265_555, w_265_556, w_265_560, w_265_561, w_265_564, w_265_566, w_265_568, w_265_570, w_265_577, w_265_578, w_265_579, w_265_580, w_265_583, w_265_584, w_265_585, w_265_586, w_265_588, w_265_593, w_265_597, w_265_598, w_265_600, w_265_603, w_265_604, w_265_609, w_265_610, w_265_613, w_265_615, w_265_616, w_265_618, w_265_619, w_265_630, w_265_631, w_265_632, w_265_635, w_265_637, w_265_643, w_265_645, w_265_654, w_265_659, w_265_660, w_265_663, w_265_664, w_265_667, w_265_668, w_265_669, w_265_674, w_265_679, w_265_680, w_265_681, w_265_682, w_265_685, w_265_686, w_265_691, w_265_692, w_265_693, w_265_697, w_265_700, w_265_708, w_265_709, w_265_710, w_265_711, w_265_714, w_265_716, w_265_719, w_265_724, w_265_726, w_265_727, w_265_728, w_265_731, w_265_732, w_265_735, w_265_736, w_265_737, w_265_739, w_265_746, w_265_747, w_265_748, w_265_752, w_265_756, w_265_757, w_265_760, w_265_761, w_265_768, w_265_770, w_265_771, w_265_773, w_265_775, w_265_776, w_265_777, w_265_778, w_265_779, w_265_780, w_265_781, w_265_782, w_265_783, w_265_784, w_265_786, w_265_787, w_265_790, w_265_791, w_265_792, w_265_794, w_265_796, w_265_801, w_265_803, w_265_806, w_265_812, w_265_814, w_265_816, w_265_817, w_265_818, w_265_819, w_265_820, w_265_821, w_265_822, w_265_823, w_265_824, w_265_825, w_265_829, w_265_830, w_265_831, w_265_832, w_265_833, w_265_834, w_265_835, w_265_837;
  wire w_266_001, w_266_007, w_266_009, w_266_038, w_266_040, w_266_041, w_266_047, w_266_074, w_266_079, w_266_086, w_266_090, w_266_095, w_266_105, w_266_153, w_266_158, w_266_188, w_266_194, w_266_196, w_266_208, w_266_214, w_266_227, w_266_239, w_266_277, w_266_281, w_266_291, w_266_305, w_266_317, w_266_327, w_266_340, w_266_346, w_266_381, w_266_407, w_266_411, w_266_414, w_266_465, w_266_468, w_266_487, w_266_508, w_266_512, w_266_536, w_266_544, w_266_554, w_266_562, w_266_565, w_266_571, w_266_581, w_266_597, w_266_599, w_266_603, w_266_616, w_266_618, w_266_628, w_266_664, w_266_668, w_266_686, w_266_719, w_266_724, w_266_742, w_266_745, w_266_750, w_266_753, w_266_763, w_266_788, w_266_791, w_266_814, w_266_818, w_266_821, w_266_825, w_266_846, w_266_858, w_266_862, w_266_901, w_266_906, w_266_933, w_266_938, w_266_955, w_266_959, w_266_965, w_266_966, w_266_975, w_266_979, w_266_980, w_266_983, w_266_998, w_266_1007, w_266_1049, w_266_1053, w_266_1055, w_266_1079, w_266_1097, w_266_1120, w_266_1149, w_266_1151, w_266_1169, w_266_1172, w_266_1184, w_266_1192, w_266_1196, w_266_1198, w_266_1220, w_266_1228, w_266_1239, w_266_1247, w_266_1281, w_266_1295, w_266_1304, w_266_1326, w_266_1337, w_266_1356, w_266_1377, w_266_1378, w_266_1389, w_266_1414, w_266_1423, w_266_1430, w_266_1453, w_266_1465, w_266_1489, w_266_1492, w_266_1503, w_266_1514, w_266_1519, w_266_1520, w_266_1521, w_266_1526, w_266_1529, w_266_1535, w_266_1536, w_266_1549, w_266_1562, w_266_1581, w_266_1593, w_266_1599, w_266_1605, w_266_1637, w_266_1653, w_266_1667, w_266_1670, w_266_1700, w_266_1709, w_266_1715, w_266_1721, w_266_1741, w_266_1751, w_266_1752, w_266_1770, w_266_1777, w_266_1784, w_266_1808, w_266_1824, w_266_1837, w_266_1840, w_266_1848, w_266_1851, w_266_1902, w_266_1913, w_266_1924, w_266_1942, w_266_1945, w_266_1947, w_266_1950, w_266_1991, w_266_1996, w_266_1997, w_266_2000, w_266_2002, w_266_2012, w_266_2029, w_266_2047, w_266_2052, w_266_2060, w_266_2066, w_266_2091, w_266_2097, w_266_2099, w_266_2101, w_266_2104, w_266_2119, w_266_2134, w_266_2141, w_266_2146, w_266_2157, w_266_2189, w_266_2255, w_266_2267, w_266_2281, w_266_2286, w_266_2314, w_266_2332, w_266_2333, w_266_2346, w_266_2357, w_266_2360, w_266_2361, w_266_2373, w_266_2392, w_266_2398, w_266_2411, w_266_2431, w_266_2451, w_266_2475, w_266_2478, w_266_2497, w_266_2498, w_266_2499, w_266_2508, w_266_2517, w_266_2526, w_266_2529, w_266_2537, w_266_2588, w_266_2590, w_266_2598, w_266_2600, w_266_2609, w_266_2617, w_266_2631, w_266_2632, w_266_2655, w_266_2670, w_266_2671, w_266_2672, w_266_2681, w_266_2699, w_266_2708, w_266_2742, w_266_2750, w_266_2760, w_266_2763, w_266_2768, w_266_2780, w_266_2781, w_266_2797, w_266_2804, w_266_2832, w_266_2843, w_266_2851, w_266_2864, w_266_2878, w_266_2889, w_266_2897, w_266_2898, w_266_2914, w_266_2929, w_266_2933, w_266_2942, w_266_2971, w_266_2975, w_266_2998, w_266_3000, w_266_3003, w_266_3006, w_266_3012, w_266_3016, w_266_3028, w_266_3047, w_266_3050, w_266_3053, w_266_3058, w_266_3084, w_266_3088, w_266_3089, w_266_3102, w_266_3132, w_266_3136, w_266_3141, w_266_3156, w_266_3159, w_266_3160, w_266_3168, w_266_3170, w_266_3176, w_266_3186, w_266_3199, w_266_3242, w_266_3250, w_266_3253, w_266_3272, w_266_3281, w_266_3284, w_266_3286, w_266_3299, w_266_3305, w_266_3324, w_266_3328, w_266_3343, w_266_3347, w_266_3348, w_266_3351, w_266_3357, w_266_3364, w_266_3417, w_266_3427, w_266_3437, w_266_3439, w_266_3441, w_266_3450, w_266_3471, w_266_3474, w_266_3477, w_266_3479, w_266_3480, w_266_3490, w_266_3493, w_266_3505, w_266_3507, w_266_3512, w_266_3516, w_266_3519, w_266_3529, w_266_3533, w_266_3562, w_266_3589, w_266_3609, w_266_3613, w_266_3626, w_266_3628, w_266_3642, w_266_3650, w_266_3665, w_266_3669, w_266_3676, w_266_3696, w_266_3706, w_266_3710, w_266_3742, w_266_3743, w_266_3760, w_266_3773, w_266_3805, w_266_3815, w_266_3818, w_266_3837, w_266_3860, w_266_3861, w_266_3881, w_266_3882, w_266_3903, w_266_3909, w_266_3916, w_266_3929, w_266_3951, w_266_3959, w_266_3990, w_266_4003, w_266_4015, w_266_4019, w_266_4024, w_266_4035, w_266_4051, w_266_4053, w_266_4056, w_266_4062, w_266_4063, w_266_4069, w_266_4081, w_266_4090, w_266_4100, w_266_4104, w_266_4108, w_266_4113, w_266_4127, w_266_4146, w_266_4162, w_266_4175, w_266_4176, w_266_4214, w_266_4230, w_266_4244, w_266_4282, w_266_4286, w_266_4293, w_266_4303, w_266_4307, w_266_4339, w_266_4343, w_266_4348, w_266_4379, w_266_4394, w_266_4408, w_266_4423, w_266_4449, w_266_4469, w_266_4484, w_266_4507, w_266_4512, w_266_4515, w_266_4530, w_266_4532, w_266_4537, w_266_4539, w_266_4546, w_266_4549, w_266_4567, w_266_4570, w_266_4593, w_266_4596, w_266_4607, w_266_4631, w_266_4643, w_266_4647, w_266_4656, w_266_4663, w_266_4678, w_266_4685, w_266_4686, w_266_4699, w_266_4720, w_266_4730, w_266_4751, w_266_4756, w_266_4764, w_266_4773, w_266_4781, w_266_4789, w_266_4808, w_266_4817, w_266_4826, w_266_4829, w_266_4839, w_266_4862, w_266_4879, w_266_4881, w_266_4890, w_266_4891, w_266_4932, w_266_4933, w_266_4936, w_266_4947, w_266_4970, w_266_4979;
  wire w_267_010, w_267_012, w_267_013, w_267_026, w_267_036, w_267_043, w_267_050, w_267_060, w_267_067, w_267_071, w_267_079, w_267_080, w_267_081, w_267_083, w_267_088, w_267_107, w_267_115, w_267_119, w_267_124, w_267_126, w_267_135, w_267_149, w_267_158, w_267_167, w_267_169, w_267_194, w_267_199, w_267_211, w_267_214, w_267_221, w_267_225, w_267_228, w_267_242, w_267_248, w_267_249, w_267_254, w_267_255, w_267_265, w_267_267, w_267_278, w_267_283, w_267_291, w_267_294, w_267_305, w_267_308, w_267_315, w_267_321, w_267_338, w_267_349, w_267_351, w_267_358, w_267_375, w_267_380, w_267_410, w_267_423, w_267_440, w_267_441, w_267_446, w_267_461, w_267_466, w_267_491, w_267_496, w_267_498, w_267_499, w_267_520, w_267_524, w_267_528, w_267_531, w_267_532, w_267_535, w_267_575, w_267_591, w_267_636, w_267_639, w_267_646, w_267_665, w_267_667, w_267_668, w_267_690, w_267_696, w_267_711, w_267_733, w_267_747, w_267_758, w_267_780, w_267_799, w_267_800, w_267_824, w_267_840, w_267_858, w_267_892, w_267_899, w_267_907, w_267_911, w_267_912, w_267_923, w_267_959, w_267_977, w_267_1009, w_267_1066, w_267_1074, w_267_1083, w_267_1092, w_267_1094, w_267_1101, w_267_1102, w_267_1103, w_267_1115, w_267_1125, w_267_1131, w_267_1142, w_267_1150, w_267_1170, w_267_1177, w_267_1186, w_267_1188, w_267_1213, w_267_1217, w_267_1236, w_267_1263, w_267_1285, w_267_1343, w_267_1357, w_267_1376, w_267_1380, w_267_1399, w_267_1416, w_267_1423, w_267_1438, w_267_1440, w_267_1475, w_267_1476, w_267_1497, w_267_1513, w_267_1524, w_267_1540, w_267_1547, w_267_1558, w_267_1567, w_267_1573, w_267_1608, w_267_1626, w_267_1631, w_267_1665, w_267_1667, w_267_1676, w_267_1696, w_267_1702, w_267_1703, w_267_1704, w_267_1722, w_267_1758, w_267_1762, w_267_1769, w_267_1783, w_267_1819, w_267_1838, w_267_1850, w_267_1858, w_267_1865, w_267_1870, w_267_1871, w_267_1881, w_267_1892, w_267_1898, w_267_1913, w_267_1940, w_267_1943, w_267_1962, w_267_1964, w_267_1975, w_267_2000, w_267_2003, w_267_2016, w_267_2020, w_267_2021, w_267_2039, w_267_2043, w_267_2064, w_267_2069, w_267_2085, w_267_2086, w_267_2092, w_267_2117, w_267_2123, w_267_2125, w_267_2137, w_267_2156, w_267_2173, w_267_2178, w_267_2185, w_267_2189, w_267_2219, w_267_2227, w_267_2234, w_267_2238, w_267_2254, w_267_2267, w_267_2280, w_267_2282, w_267_2292, w_267_2299, w_267_2309, w_267_2319, w_267_2324, w_267_2330, w_267_2348, w_267_2358, w_267_2361, w_267_2366, w_267_2386, w_267_2397, w_267_2405, w_267_2409, w_267_2419, w_267_2424, w_267_2437, w_267_2442, w_267_2460, w_267_2463, w_267_2464, w_267_2467, w_267_2474, w_267_2481, w_267_2492, w_267_2494, w_267_2502, w_267_2509, w_267_2521, w_267_2528, w_267_2544, w_267_2562, w_267_2569, w_267_2570, w_267_2572, w_267_2601, w_267_2630, w_267_2651, w_267_2658, w_267_2664, w_267_2684, w_267_2688, w_267_2696, w_267_2701, w_267_2708, w_267_2711, w_267_2712, w_267_2721, w_267_2724, w_267_2729, w_267_2748, w_267_2752, w_267_2754, w_267_2756, w_267_2782, w_267_2806, w_267_2807, w_267_2808, w_267_2810, w_267_2823, w_267_2846, w_267_2857, w_267_2860, w_267_2868, w_267_2883, w_267_2896, w_267_2898, w_267_2912, w_267_2914, w_267_2917, w_267_2920, w_267_2944, w_267_2946, w_267_2963, w_267_2968, w_267_2988, w_267_3035, w_267_3038, w_267_3063, w_267_3066, w_267_3091, w_267_3101, w_267_3113, w_267_3116, w_267_3205, w_267_3206, w_267_3221, w_267_3249, w_267_3252, w_267_3290, w_267_3295, w_267_3297, w_267_3303, w_267_3312, w_267_3364, w_267_3386, w_267_3387, w_267_3398, w_267_3406, w_267_3408, w_267_3439, w_267_3445, w_267_3471, w_267_3473, w_267_3476, w_267_3489, w_267_3494, w_267_3507, w_267_3519, w_267_3520, w_267_3548, w_267_3558, w_267_3562, w_267_3564, w_267_3568, w_267_3572, w_267_3577, w_267_3592, w_267_3600, w_267_3654, w_267_3663, w_267_3666, w_267_3673, w_267_3674, w_267_3675, w_267_3697, w_267_3703, w_267_3707, w_267_3728, w_267_3746, w_267_3756, w_267_3759, w_267_3769, w_267_3778, w_267_3785, w_267_3794, w_267_3800, w_267_3807, w_267_3836, w_267_3849, w_267_3852, w_267_3865, w_267_3869, w_267_3873, w_267_3877, w_267_3887, w_267_3927, w_267_3928, w_267_3937, w_267_3938, w_267_3946, w_267_3950, w_267_3961, w_267_3967, w_267_3969, w_267_3980, w_267_4013, w_267_4022, w_267_4045, w_267_4055, w_267_4067, w_267_4073, w_267_4081, w_267_4084, w_267_4097, w_267_4098, w_267_4110, w_267_4119, w_267_4146, w_267_4153, w_267_4154, w_267_4215, w_267_4253, w_267_4256, w_267_4283, w_267_4288, w_267_4309, w_267_4331, w_267_4335, w_267_4340, w_267_4355, w_267_4356, w_267_4357, w_267_4368, w_267_4369, w_267_4375, w_267_4381, w_267_4390, w_267_4404, w_267_4419, w_267_4435, w_267_4441, w_267_4479, w_267_4488, w_267_4493, w_267_4497, w_267_4504, w_267_4510, w_267_4513, w_267_4516, w_267_4519, w_267_4524, w_267_4544, w_267_4545, w_267_4631, w_267_4641, w_267_4647, w_267_4668, w_267_4670, w_267_4676, w_267_4681, w_267_4686, w_267_4692;
  wire w_268_002, w_268_003, w_268_005, w_268_006, w_268_008, w_268_017, w_268_020, w_268_021, w_268_023, w_268_024, w_268_025, w_268_028, w_268_029, w_268_032, w_268_036, w_268_037, w_268_040, w_268_042, w_268_046, w_268_051, w_268_054, w_268_055, w_268_059, w_268_064, w_268_068, w_268_071, w_268_072, w_268_073, w_268_074, w_268_076, w_268_077, w_268_078, w_268_082, w_268_083, w_268_091, w_268_092, w_268_103, w_268_104, w_268_106, w_268_111, w_268_112, w_268_119, w_268_121, w_268_125, w_268_128, w_268_132, w_268_136, w_268_137, w_268_140, w_268_142, w_268_146, w_268_148, w_268_154, w_268_155, w_268_157, w_268_158, w_268_164, w_268_168, w_268_170, w_268_172, w_268_179, w_268_182, w_268_183, w_268_185, w_268_191, w_268_194, w_268_197, w_268_199, w_268_207, w_268_210, w_268_211, w_268_213, w_268_214, w_268_218, w_268_219, w_268_226, w_268_227, w_268_232, w_268_244, w_268_246, w_268_249, w_268_255, w_268_259, w_268_261, w_268_268, w_268_272, w_268_278, w_268_279, w_268_282, w_268_285, w_268_297, w_268_300, w_268_301, w_268_302, w_268_306, w_268_311, w_268_317, w_268_318, w_268_323, w_268_327, w_268_328, w_268_329, w_268_333, w_268_335, w_268_338, w_268_342, w_268_348, w_268_350, w_268_351, w_268_356, w_268_358, w_268_359, w_268_375, w_268_379, w_268_381, w_268_383, w_268_385, w_268_404, w_268_409, w_268_412, w_268_422, w_268_424, w_268_429, w_268_432, w_268_434, w_268_435, w_268_439, w_268_444, w_268_447, w_268_449, w_268_452, w_268_456, w_268_467, w_268_472, w_268_473, w_268_477, w_268_478, w_268_479, w_268_483, w_268_486, w_268_488, w_268_492, w_268_507, w_268_510, w_268_516, w_268_521, w_268_525, w_268_531, w_268_534, w_268_537, w_268_546, w_268_547, w_268_551, w_268_555, w_268_557, w_268_566, w_268_569, w_268_571, w_268_575, w_268_576, w_268_587, w_268_589, w_268_594, w_268_617, w_268_622, w_268_636, w_268_638, w_268_640, w_268_644, w_268_651, w_268_656, w_268_658, w_268_659, w_268_660, w_268_665, w_268_671, w_268_672, w_268_679, w_268_685, w_268_689, w_268_693, w_268_696, w_268_699, w_268_700, w_268_705, w_268_706, w_268_715, w_268_722, w_268_725, w_268_739, w_268_740, w_268_742, w_268_744, w_268_748, w_268_753, w_268_756, w_268_760, w_268_767, w_268_768, w_268_770, w_268_775, w_268_776, w_268_783, w_268_792, w_268_793, w_268_795, w_268_802, w_268_805, w_268_807, w_268_811, w_268_815, w_268_816, w_268_818, w_268_820, w_268_823, w_268_834, w_268_842, w_268_843, w_268_845, w_268_852, w_268_857, w_268_861, w_268_865, w_268_875, w_268_878, w_268_879, w_268_880, w_268_882, w_268_888, w_268_889, w_268_891, w_268_893, w_268_897, w_268_899, w_268_902, w_268_903, w_268_909, w_268_910, w_268_918, w_268_919, w_268_926, w_268_928, w_268_929, w_268_931, w_268_932, w_268_937, w_268_938, w_268_942, w_268_947, w_268_949, w_268_951, w_268_952, w_268_955, w_268_958, w_268_964, w_268_965, w_268_973, w_268_976, w_268_977, w_268_979, w_268_982, w_268_986, w_268_997, w_268_999, w_268_1020, w_268_1028, w_268_1030, w_268_1031, w_268_1041, w_268_1051, w_268_1053, w_268_1055, w_268_1057, w_268_1058, w_268_1060, w_268_1062, w_268_1063, w_268_1066, w_268_1077, w_268_1078, w_268_1081, w_268_1083, w_268_1090, w_268_1096, w_268_1107, w_268_1109, w_268_1111, w_268_1119, w_268_1121, w_268_1128, w_268_1129, w_268_1131, w_268_1133, w_268_1136, w_268_1139, w_268_1140, w_268_1141, w_268_1142, w_268_1147, w_268_1153, w_268_1156, w_268_1159, w_268_1165, w_268_1166, w_268_1167, w_268_1168, w_268_1172, w_268_1173, w_268_1184, w_268_1193, w_268_1217, w_268_1224, w_268_1228, w_268_1231, w_268_1235, w_268_1236, w_268_1237, w_268_1249, w_268_1262, w_268_1266, w_268_1270, w_268_1283, w_268_1292, w_268_1294, w_268_1299, w_268_1302, w_268_1304, w_268_1305, w_268_1317, w_268_1327, w_268_1329, w_268_1331, w_268_1332, w_268_1333, w_268_1334, w_268_1337, w_268_1341, w_268_1347, w_268_1350, w_268_1351, w_268_1352, w_268_1368, w_268_1369, w_268_1373, w_268_1378, w_268_1388, w_268_1395, w_268_1404, w_268_1408, w_268_1409, w_268_1411, w_268_1412, w_268_1414, w_268_1415, w_268_1416, w_268_1419, w_268_1425, w_268_1431, w_268_1432, w_268_1436, w_268_1449, w_268_1450, w_268_1458, w_268_1462, w_268_1464, w_268_1467, w_268_1468, w_268_1476, w_268_1479, w_268_1482, w_268_1491, w_268_1494, w_268_1501, w_268_1503, w_268_1504, w_268_1506, w_268_1507, w_268_1508, w_268_1517;
  wire w_269_000, w_269_005, w_269_014, w_269_015, w_269_022, w_269_029, w_269_033, w_269_034, w_269_035, w_269_041, w_269_062, w_269_065, w_269_066, w_269_073, w_269_088, w_269_090, w_269_095, w_269_099, w_269_103, w_269_106, w_269_124, w_269_125, w_269_133, w_269_138, w_269_147, w_269_161, w_269_162, w_269_163, w_269_166, w_269_170, w_269_194, w_269_203, w_269_221, w_269_228, w_269_234, w_269_245, w_269_246, w_269_268, w_269_269, w_269_272, w_269_304, w_269_308, w_269_311, w_269_312, w_269_321, w_269_323, w_269_330, w_269_331, w_269_334, w_269_336, w_269_337, w_269_343, w_269_347, w_269_351, w_269_356, w_269_366, w_269_369, w_269_372, w_269_391, w_269_396, w_269_397, w_269_406, w_269_417, w_269_420, w_269_429, w_269_431, w_269_436, w_269_441, w_269_461, w_269_485, w_269_491, w_269_497, w_269_499, w_269_501, w_269_508, w_269_535, w_269_540, w_269_547, w_269_553, w_269_555, w_269_558, w_269_563, w_269_566, w_269_569, w_269_576, w_269_592, w_269_603, w_269_605, w_269_640, w_269_645, w_269_646, w_269_662, w_269_666, w_269_667, w_269_675, w_269_686, w_269_690, w_269_691, w_269_694, w_269_697, w_269_759, w_269_767, w_269_771, w_269_773, w_269_776, w_269_790, w_269_800, w_269_807, w_269_809, w_269_812, w_269_820, w_269_826, w_269_827, w_269_835, w_269_838, w_269_845, w_269_846, w_269_851, w_269_870, w_269_879, w_269_883, w_269_893, w_269_895, w_269_923, w_269_934, w_269_936, w_269_939, w_269_947, w_269_950, w_269_951, w_269_965, w_269_966, w_269_968, w_269_969, w_269_976, w_269_980, w_269_984, w_269_993, w_269_1014, w_269_1017, w_269_1021, w_269_1024, w_269_1031, w_269_1038, w_269_1040, w_269_1051, w_269_1053, w_269_1054, w_269_1067, w_269_1081, w_269_1082, w_269_1100, w_269_1103, w_269_1113, w_269_1118, w_269_1122, w_269_1123, w_269_1143, w_269_1150, w_269_1151, w_269_1174, w_269_1181, w_269_1197, w_269_1200, w_269_1204, w_269_1205, w_269_1221, w_269_1223, w_269_1229, w_269_1232, w_269_1239, w_269_1248, w_269_1256, w_269_1268, w_269_1269, w_269_1275, w_269_1279, w_269_1301, w_269_1304, w_269_1305, w_269_1308, w_269_1319, w_269_1320, w_269_1329, w_269_1334, w_269_1348, w_269_1350, w_269_1351, w_269_1353, w_269_1357, w_269_1372, w_269_1380, w_269_1398, w_269_1404, w_269_1410, w_269_1432, w_269_1458, w_269_1467, w_269_1469, w_269_1477, w_269_1486, w_269_1489, w_269_1510, w_269_1513, w_269_1518, w_269_1525, w_269_1527, w_269_1531, w_269_1544, w_269_1550, w_269_1566, w_269_1568, w_269_1572, w_269_1579, w_269_1591, w_269_1593, w_269_1625, w_269_1630, w_269_1632, w_269_1633, w_269_1636, w_269_1643, w_269_1656, w_269_1660, w_269_1664, w_269_1676, w_269_1710, w_269_1711, w_269_1712, w_269_1715, w_269_1722, w_269_1733, w_269_1739, w_269_1741, w_269_1744, w_269_1747, w_269_1761, w_269_1769, w_269_1770, w_269_1793, w_269_1806, w_269_1808, w_269_1817, w_269_1818, w_269_1821, w_269_1823, w_269_1824, w_269_1832, w_269_1833, w_269_1836, w_269_1844, w_269_1852, w_269_1862, w_269_1865, w_269_1867, w_269_1872, w_269_1881, w_269_1895, w_269_1909, w_269_1917, w_269_1921, w_269_1922, w_269_1925, w_269_1927, w_269_1928, w_269_1933, w_269_1944, w_269_1949, w_269_1950, w_269_1958, w_269_1959, w_269_1965, w_269_1969, w_269_1975, w_269_1989, w_269_1993, w_269_2004, w_269_2007, w_269_2045, w_269_2056, w_269_2062, w_269_2076, w_269_2094, w_269_2110, w_269_2117, w_269_2124, w_269_2132, w_269_2137, w_269_2143, w_269_2149, w_269_2162, w_269_2191, w_269_2210, w_269_2215, w_269_2217, w_269_2238, w_269_2250, w_269_2260, w_269_2263, w_269_2286, w_269_2291, w_269_2305, w_269_2308, w_269_2314, w_269_2316, w_269_2337, w_269_2339, w_269_2363, w_269_2367, w_269_2373, w_269_2392, w_269_2397, w_269_2400, w_269_2425, w_269_2429, w_269_2454, w_269_2482, w_269_2497, w_269_2521, w_269_2540, w_269_2542, w_269_2575, w_269_2620, w_269_2653, w_269_2654, w_269_2667, w_269_2690, w_269_2695, w_269_2708, w_269_2710, w_269_2732, w_269_2746, w_269_2759, w_269_2762, w_269_2769, w_269_2798, w_269_2814, w_269_2819, w_269_2839, w_269_2850, w_269_2854, w_269_2855, w_269_2866, w_269_2873, w_269_2881, w_269_2890, w_269_2894, w_269_2903, w_269_2910, w_269_2912, w_269_2922, w_269_2952, w_269_2958, w_269_2959, w_269_2960, w_269_2961, w_269_2962, w_269_2964;
  wire w_270_012, w_270_016, w_270_025, w_270_027, w_270_038, w_270_059, w_270_066, w_270_069, w_270_072, w_270_077, w_270_092, w_270_114, w_270_116, w_270_130, w_270_132, w_270_136, w_270_157, w_270_163, w_270_164, w_270_180, w_270_197, w_270_200, w_270_206, w_270_210, w_270_212, w_270_223, w_270_226, w_270_236, w_270_240, w_270_243, w_270_254, w_270_256, w_270_258, w_270_261, w_270_263, w_270_266, w_270_278, w_270_279, w_270_282, w_270_283, w_270_288, w_270_292, w_270_306, w_270_308, w_270_313, w_270_314, w_270_318, w_270_320, w_270_322, w_270_323, w_270_336, w_270_339, w_270_341, w_270_358, w_270_362, w_270_366, w_270_368, w_270_373, w_270_376, w_270_380, w_270_383, w_270_389, w_270_397, w_270_401, w_270_405, w_270_422, w_270_424, w_270_433, w_270_439, w_270_442, w_270_455, w_270_457, w_270_461, w_270_464, w_270_467, w_270_468, w_270_473, w_270_481, w_270_486, w_270_493, w_270_494, w_270_516, w_270_518, w_270_519, w_270_523, w_270_524, w_270_539, w_270_541, w_270_553, w_270_555, w_270_567, w_270_569, w_270_572, w_270_576, w_270_577, w_270_581, w_270_590, w_270_591, w_270_592, w_270_596, w_270_609, w_270_620, w_270_622, w_270_629, w_270_634, w_270_649, w_270_652, w_270_661, w_270_670, w_270_674, w_270_678, w_270_683, w_270_691, w_270_692, w_270_700, w_270_701, w_270_707, w_270_710, w_270_714, w_270_741, w_270_743, w_270_746, w_270_747, w_270_756, w_270_759, w_270_766, w_270_774, w_270_776, w_270_777, w_270_778, w_270_785, w_270_789, w_270_790, w_270_792, w_270_794, w_270_800, w_270_802, w_270_804, w_270_806, w_270_816, w_270_830, w_270_834, w_270_836, w_270_837, w_270_838, w_270_844, w_270_845, w_270_848, w_270_860, w_270_861, w_270_871, w_270_878, w_270_902, w_270_907, w_270_912, w_270_917, w_270_923, w_270_928, w_270_929, w_270_930, w_270_941, w_270_942, w_270_944, w_270_946, w_270_958, w_270_959, w_270_986, w_270_1012, w_270_1017, w_270_1025, w_270_1032, w_270_1043, w_270_1047, w_270_1056, w_270_1061, w_270_1062, w_270_1067, w_270_1077, w_270_1081, w_270_1083, w_270_1088, w_270_1090, w_270_1091, w_270_1095, w_270_1104, w_270_1106, w_270_1107, w_270_1108, w_270_1117, w_270_1125, w_270_1132, w_270_1142, w_270_1173, w_270_1174, w_270_1185, w_270_1188, w_270_1190, w_270_1191, w_270_1192, w_270_1197, w_270_1214, w_270_1216, w_270_1217, w_270_1223, w_270_1225, w_270_1231, w_270_1234, w_270_1240, w_270_1252, w_270_1255, w_270_1256, w_270_1263, w_270_1271, w_270_1274, w_270_1286, w_270_1290, w_270_1294, w_270_1298, w_270_1305, w_270_1309, w_270_1312, w_270_1313, w_270_1317, w_270_1324, w_270_1325, w_270_1330, w_270_1331, w_270_1333, w_270_1337, w_270_1339, w_270_1343, w_270_1344, w_270_1346, w_270_1352, w_270_1353, w_270_1362, w_270_1366, w_270_1367, w_270_1369, w_270_1371, w_270_1388, w_270_1397, w_270_1401, w_270_1406, w_270_1420, w_270_1422, w_270_1423, w_270_1432, w_270_1433, w_270_1435, w_270_1438, w_270_1439, w_270_1441, w_270_1457, w_270_1471, w_270_1472, w_270_1473, w_270_1474, w_270_1489, w_270_1493, w_270_1509, w_270_1510, w_270_1524, w_270_1530, w_270_1538, w_270_1539, w_270_1542, w_270_1550, w_270_1556, w_270_1561, w_270_1562, w_270_1569, w_270_1584, w_270_1591, w_270_1592, w_270_1599, w_270_1607, w_270_1613, w_270_1615, w_270_1622, w_270_1623, w_270_1633, w_270_1645, w_270_1647, w_270_1657, w_270_1659, w_270_1660, w_270_1661, w_270_1665, w_270_1666, w_270_1684, w_270_1687, w_270_1701, w_270_1707, w_270_1718, w_270_1721, w_270_1725, w_270_1727, w_270_1735, w_270_1739, w_270_1754, w_270_1757, w_270_1761, w_270_1762, w_270_1768, w_270_1769, w_270_1774, w_270_1775, w_270_1782, w_270_1784, w_270_1789, w_270_1796, w_270_1801, w_270_1803, w_270_1814, w_270_1819, w_270_1822, w_270_1826, w_270_1828, w_270_1831, w_270_1843, w_270_1849, w_270_1851, w_270_1861, w_270_1875, w_270_1877, w_270_1887, w_270_1889, w_270_1901, w_270_1915, w_270_1918, w_270_1947, w_270_1952, w_270_1954, w_270_1955, w_270_1965, w_270_1975, w_270_1979, w_270_1981, w_270_1982, w_270_1991, w_270_2000, w_270_2001, w_270_2003, w_270_2022, w_270_2030, w_270_2044, w_270_2051, w_270_2065, w_270_2076, w_270_2090, w_270_2094, w_270_2098, w_270_2119, w_270_2125, w_270_2136, w_270_2144, w_270_2146, w_270_2148, w_270_2166, w_270_2175, w_270_2177, w_270_2178, w_270_2179, w_270_2180, w_270_2187, w_270_2195, w_270_2197, w_270_2198, w_270_2200, w_270_2205, w_270_2208, w_270_2210, w_270_2212, w_270_2227, w_270_2238, w_270_2250, w_270_2255, w_270_2258, w_270_2269, w_270_2271, w_270_2277, w_270_2284, w_270_2287, w_270_2288, w_270_2301, w_270_2302, w_270_2309, w_270_2315, w_270_2367, w_270_2404, w_270_2405, w_270_2406, w_270_2414, w_270_2426, w_270_2468, w_270_2474, w_270_2478, w_270_2483, w_270_2495, w_270_2518, w_270_2521, w_270_2532, w_270_2533, w_270_2534, w_270_2568, w_270_2573, w_270_2594, w_270_2597, w_270_2611, w_270_2612, w_270_2633, w_270_2647, w_270_2649, w_270_2653, w_270_2662, w_270_2663, w_270_2664, w_270_2665, w_270_2666, w_270_2667, w_270_2668, w_270_2669, w_270_2670, w_270_2671, w_270_2672, w_270_2674, w_270_2676, w_270_2677, w_270_2678, w_270_2679, w_270_2680, w_270_2681, w_270_2682, w_270_2683, w_270_2685;
  wire w_271_006, w_271_008, w_271_022, w_271_024, w_271_027, w_271_031, w_271_037, w_271_038, w_271_045, w_271_046, w_271_053, w_271_058, w_271_059, w_271_064, w_271_072, w_271_073, w_271_081, w_271_092, w_271_093, w_271_097, w_271_107, w_271_111, w_271_112, w_271_123, w_271_129, w_271_134, w_271_147, w_271_150, w_271_151, w_271_155, w_271_166, w_271_171, w_271_175, w_271_176, w_271_180, w_271_184, w_271_194, w_271_204, w_271_206, w_271_208, w_271_221, w_271_222, w_271_228, w_271_237, w_271_238, w_271_239, w_271_263, w_271_264, w_271_266, w_271_267, w_271_271, w_271_272, w_271_276, w_271_280, w_271_284, w_271_286, w_271_291, w_271_293, w_271_294, w_271_301, w_271_307, w_271_309, w_271_310, w_271_313, w_271_340, w_271_345, w_271_356, w_271_363, w_271_364, w_271_373, w_271_375, w_271_376, w_271_389, w_271_391, w_271_396, w_271_403, w_271_410, w_271_421, w_271_434, w_271_437, w_271_441, w_271_446, w_271_453, w_271_456, w_271_457, w_271_462, w_271_472, w_271_474, w_271_477, w_271_486, w_271_519, w_271_545, w_271_547, w_271_550, w_271_565, w_271_574, w_271_575, w_271_578, w_271_581, w_271_582, w_271_589, w_271_597, w_271_609, w_271_617, w_271_618, w_271_623, w_271_628, w_271_633, w_271_635, w_271_638, w_271_640, w_271_643, w_271_648, w_271_660, w_271_661, w_271_663, w_271_671, w_271_673, w_271_685, w_271_687, w_271_693, w_271_703, w_271_712, w_271_716, w_271_729, w_271_731, w_271_740, w_271_742, w_271_749, w_271_753, w_271_763, w_271_765, w_271_776, w_271_783, w_271_786, w_271_798, w_271_811, w_271_813, w_271_818, w_271_834, w_271_836, w_271_839, w_271_841, w_271_847, w_271_852, w_271_860, w_271_867, w_271_868, w_271_876, w_271_880, w_271_883, w_271_893, w_271_901, w_271_917, w_271_929, w_271_934, w_271_948, w_271_970, w_271_986, w_271_990, w_271_1036, w_271_1049, w_271_1058, w_271_1060, w_271_1075, w_271_1087, w_271_1092, w_271_1095, w_271_1110, w_271_1115, w_271_1133, w_271_1153, w_271_1156, w_271_1160, w_271_1176, w_271_1187, w_271_1199, w_271_1225, w_271_1257, w_271_1262, w_271_1294, w_271_1298, w_271_1314, w_271_1316, w_271_1326, w_271_1356, w_271_1360, w_271_1367, w_271_1371, w_271_1382, w_271_1392, w_271_1425, w_271_1472, w_271_1475, w_271_1482, w_271_1530, w_271_1541, w_271_1558, w_271_1559, w_271_1563, w_271_1570, w_271_1609, w_271_1617, w_271_1624, w_271_1673, w_271_1685, w_271_1686, w_271_1689, w_271_1697, w_271_1710, w_271_1715, w_271_1717, w_271_1718, w_271_1724, w_271_1754, w_271_1793, w_271_1803, w_271_1836, w_271_1837, w_271_1848, w_271_1851, w_271_1873, w_271_1881, w_271_1910, w_271_1915, w_271_1919, w_271_1937, w_271_1941, w_271_1961, w_271_1966, w_271_1988, w_271_1997, w_271_2004, w_271_2010, w_271_2026, w_271_2028, w_271_2030, w_271_2047, w_271_2061, w_271_2063, w_271_2081, w_271_2095, w_271_2099, w_271_2116, w_271_2126, w_271_2137, w_271_2141, w_271_2161, w_271_2168, w_271_2169, w_271_2177, w_271_2184, w_271_2193, w_271_2209, w_271_2224, w_271_2247, w_271_2250, w_271_2256, w_271_2257, w_271_2263, w_271_2273, w_271_2285, w_271_2294, w_271_2303, w_271_2322, w_271_2372, w_271_2374, w_271_2395, w_271_2399, w_271_2400, w_271_2417, w_271_2448, w_271_2462, w_271_2492, w_271_2497, w_271_2504, w_271_2507, w_271_2527, w_271_2529, w_271_2532, w_271_2551, w_271_2574, w_271_2615, w_271_2628, w_271_2650, w_271_2654, w_271_2658, w_271_2659, w_271_2662, w_271_2684, w_271_2690, w_271_2729, w_271_2735, w_271_2738, w_271_2742, w_271_2748, w_271_2771, w_271_2778, w_271_2782, w_271_2783, w_271_2788, w_271_2790, w_271_2794, w_271_2798, w_271_2802, w_271_2804, w_271_2806, w_271_2832, w_271_2836, w_271_2861, w_271_2866, w_271_2872, w_271_2885, w_271_2887, w_271_2895, w_271_2899, w_271_2919, w_271_2955, w_271_2978, w_271_2979, w_271_2986, w_271_2987, w_271_3021, w_271_3030, w_271_3036, w_271_3058, w_271_3071, w_271_3089, w_271_3096, w_271_3132, w_271_3136, w_271_3145, w_271_3161, w_271_3162, w_271_3190, w_271_3207, w_271_3208, w_271_3212, w_271_3223, w_271_3242, w_271_3271, w_271_3278, w_271_3283, w_271_3285, w_271_3299, w_271_3303, w_271_3315, w_271_3317, w_271_3320, w_271_3337, w_271_3343, w_271_3344, w_271_3385, w_271_3387, w_271_3393, w_271_3407, w_271_3417, w_271_3421, w_271_3437, w_271_3444, w_271_3450, w_271_3462, w_271_3463, w_271_3469, w_271_3474, w_271_3486, w_271_3489, w_271_3498, w_271_3499, w_271_3509, w_271_3517, w_271_3531, w_271_3550, w_271_3570, w_271_3584, w_271_3592, w_271_3594, w_271_3603, w_271_3636, w_271_3652, w_271_3660, w_271_3664, w_271_3672, w_271_3696, w_271_3698, w_271_3717, w_271_3724, w_271_3744, w_271_3750, w_271_3756, w_271_3767, w_271_3779, w_271_3781, w_271_3799, w_271_3807, w_271_3808, w_271_3822, w_271_3833, w_271_3844, w_271_3852, w_271_3860, w_271_3869, w_271_3892, w_271_3894, w_271_3896, w_271_3897, w_271_3903, w_271_3911, w_271_3925, w_271_3928, w_271_3931, w_271_3942, w_271_3956, w_271_3958, w_271_3986, w_271_3990, w_271_3991, w_271_3999, w_271_4081;
  wire w_272_000, w_272_001, w_272_002, w_272_003, w_272_004, w_272_005, w_272_006, w_272_007, w_272_008, w_272_009, w_272_010, w_272_011, w_272_012, w_272_013, w_272_014, w_272_015, w_272_016, w_272_017, w_272_018, w_272_019, w_272_020, w_272_021, w_272_022, w_272_023, w_272_024, w_272_025, w_272_026, w_272_027, w_272_028, w_272_029, w_272_030, w_272_031, w_272_032, w_272_033, w_272_034, w_272_035, w_272_036, w_272_037, w_272_038, w_272_039, w_272_041, w_272_042, w_272_043, w_272_044, w_272_045, w_272_046, w_272_047, w_272_048, w_272_049, w_272_050, w_272_051, w_272_052, w_272_053, w_272_054, w_272_055, w_272_056, w_272_057, w_272_058, w_272_059, w_272_061, w_272_062, w_272_063, w_272_064, w_272_065, w_272_066, w_272_067, w_272_068, w_272_069, w_272_070, w_272_071, w_272_072, w_272_073, w_272_074, w_272_075, w_272_076, w_272_077, w_272_078, w_272_079, w_272_080, w_272_082, w_272_083, w_272_084, w_272_086, w_272_087, w_272_088, w_272_089, w_272_090, w_272_091, w_272_092, w_272_093, w_272_094, w_272_095, w_272_096, w_272_097, w_272_098, w_272_099, w_272_100, w_272_101, w_272_102, w_272_103, w_272_104, w_272_105, w_272_106, w_272_107, w_272_108, w_272_109, w_272_110, w_272_111, w_272_112, w_272_113, w_272_114, w_272_115, w_272_116, w_272_117, w_272_118, w_272_119, w_272_120, w_272_121, w_272_122, w_272_123, w_272_125, w_272_126, w_272_127, w_272_128, w_272_129, w_272_130, w_272_131, w_272_132, w_272_133, w_272_134, w_272_136, w_272_137, w_272_138, w_272_139, w_272_140, w_272_141, w_272_142, w_272_143, w_272_144, w_272_145, w_272_146;
  wire w_273_000, w_273_005, w_273_006, w_273_007, w_273_009, w_273_012, w_273_015, w_273_018, w_273_019, w_273_020, w_273_023, w_273_024, w_273_025, w_273_028, w_273_030, w_273_033, w_273_039, w_273_040, w_273_042, w_273_044, w_273_045, w_273_047, w_273_048, w_273_049, w_273_050, w_273_053, w_273_054, w_273_056, w_273_062, w_273_064, w_273_065, w_273_066, w_273_067, w_273_068, w_273_069, w_273_070, w_273_071, w_273_076, w_273_079, w_273_085, w_273_091, w_273_096, w_273_099, w_273_101, w_273_103, w_273_104, w_273_105, w_273_107, w_273_109, w_273_111, w_273_114, w_273_116, w_273_121, w_273_124, w_273_125, w_273_127, w_273_128, w_273_135, w_273_138, w_273_139, w_273_147, w_273_149, w_273_151, w_273_160, w_273_162, w_273_163, w_273_167, w_273_168, w_273_170, w_273_174, w_273_175, w_273_178, w_273_180, w_273_181, w_273_184, w_273_185, w_273_187, w_273_188, w_273_191, w_273_192, w_273_195, w_273_196, w_273_197, w_273_201, w_273_202, w_273_206, w_273_209, w_273_211, w_273_212, w_273_213, w_273_214, w_273_217, w_273_219, w_273_220, w_273_222, w_273_224, w_273_225, w_273_227, w_273_229, w_273_230, w_273_231, w_273_237, w_273_239, w_273_240, w_273_241, w_273_242, w_273_243, w_273_246, w_273_250, w_273_252, w_273_255, w_273_257, w_273_258, w_273_259, w_273_260, w_273_261, w_273_262, w_273_266, w_273_267, w_273_269, w_273_270, w_273_271, w_273_272, w_273_273, w_273_276, w_273_278, w_273_279, w_273_283, w_273_284, w_273_287, w_273_290, w_273_291, w_273_292, w_273_294, w_273_295, w_273_297, w_273_301, w_273_304, w_273_305, w_273_309, w_273_310, w_273_314, w_273_315, w_273_317, w_273_318, w_273_319, w_273_321, w_273_323, w_273_327, w_273_331, w_273_332, w_273_340, w_273_341, w_273_342, w_273_346, w_273_347, w_273_349, w_273_354, w_273_360, w_273_361, w_273_365, w_273_368, w_273_369, w_273_371, w_273_372, w_273_379, w_273_380, w_273_381, w_273_382, w_273_385, w_273_386, w_273_387, w_273_388, w_273_391, w_273_398, w_273_401, w_273_402, w_273_405, w_273_406, w_273_409, w_273_410, w_273_416, w_273_418, w_273_419, w_273_420, w_273_421, w_273_422, w_273_426, w_273_428, w_273_439, w_273_440, w_273_441, w_273_442, w_273_443, w_273_444, w_273_452, w_273_454, w_273_455, w_273_465, w_273_466, w_273_468, w_273_471, w_273_472, w_273_474, w_273_475, w_273_476, w_273_478, w_273_484, w_273_486, w_273_487, w_273_488, w_273_489, w_273_490, w_273_491, w_273_492, w_273_495, w_273_499, w_273_501, w_273_502, w_273_503, w_273_506, w_273_507, w_273_510, w_273_514, w_273_521, w_273_523, w_273_527, w_273_529, w_273_530, w_273_533, w_273_535, w_273_537, w_273_539, w_273_540, w_273_541, w_273_543, w_273_549, w_273_551, w_273_552, w_273_556, w_273_557, w_273_560, w_273_561, w_273_563, w_273_565, w_273_567, w_273_573, w_273_574, w_273_578, w_273_579, w_273_581, w_273_583, w_273_585, w_273_589, w_273_590, w_273_591, w_273_594, w_273_601, w_273_603, w_273_604, w_273_607, w_273_610, w_273_619, w_273_621, w_273_623, w_273_626, w_273_627, w_273_628, w_273_632, w_273_635, w_273_636, w_273_639, w_273_640, w_273_645, w_273_646, w_273_651, w_273_652, w_273_656, w_273_657, w_273_658, w_273_659, w_273_662, w_273_666, w_273_668, w_273_671, w_273_673, w_273_676, w_273_677, w_273_681, w_273_684, w_273_685, w_273_689, w_273_690, w_273_693, w_273_699, w_273_700, w_273_701, w_273_702, w_273_704, w_273_705, w_273_707, w_273_708, w_273_710, w_273_711, w_273_712, w_273_713, w_273_715, w_273_718, w_273_719, w_273_721, w_273_726, w_273_727, w_273_733, w_273_734, w_273_736, w_273_738, w_273_739, w_273_740, w_273_741;
  wire w_274_009, w_274_014, w_274_024, w_274_033, w_274_043, w_274_044, w_274_071, w_274_088, w_274_092, w_274_093, w_274_097, w_274_101, w_274_104, w_274_105, w_274_108, w_274_114, w_274_119, w_274_131, w_274_132, w_274_134, w_274_136, w_274_145, w_274_150, w_274_161, w_274_166, w_274_168, w_274_171, w_274_196, w_274_201, w_274_203, w_274_204, w_274_207, w_274_220, w_274_234, w_274_236, w_274_247, w_274_253, w_274_255, w_274_270, w_274_276, w_274_308, w_274_320, w_274_327, w_274_329, w_274_330, w_274_334, w_274_346, w_274_353, w_274_359, w_274_360, w_274_369, w_274_371, w_274_380, w_274_393, w_274_394, w_274_395, w_274_396, w_274_398, w_274_401, w_274_405, w_274_406, w_274_408, w_274_416, w_274_428, w_274_434, w_274_438, w_274_444, w_274_446, w_274_458, w_274_464, w_274_477, w_274_484, w_274_488, w_274_492, w_274_501, w_274_506, w_274_507, w_274_510, w_274_524, w_274_525, w_274_529, w_274_535, w_274_536, w_274_548, w_274_573, w_274_588, w_274_607, w_274_609, w_274_615, w_274_617, w_274_626, w_274_632, w_274_633, w_274_634, w_274_638, w_274_644, w_274_646, w_274_661, w_274_666, w_274_667, w_274_679, w_274_685, w_274_693, w_274_711, w_274_717, w_274_721, w_274_726, w_274_737, w_274_750, w_274_754, w_274_760, w_274_764, w_274_774, w_274_784, w_274_789, w_274_815, w_274_816, w_274_818, w_274_831, w_274_834, w_274_837, w_274_844, w_274_858, w_274_859, w_274_871, w_274_875, w_274_879, w_274_889, w_274_893, w_274_913, w_274_914, w_274_919, w_274_929, w_274_937, w_274_948, w_274_951, w_274_952, w_274_960, w_274_969, w_274_986, w_274_989, w_274_994, w_274_1004, w_274_1007, w_274_1034, w_274_1040, w_274_1044, w_274_1051, w_274_1055, w_274_1058, w_274_1062, w_274_1068, w_274_1073, w_274_1097, w_274_1103, w_274_1107, w_274_1112, w_274_1113, w_274_1119, w_274_1122, w_274_1132, w_274_1140, w_274_1142, w_274_1153, w_274_1158, w_274_1159, w_274_1160, w_274_1162, w_274_1172, w_274_1174, w_274_1177, w_274_1187, w_274_1191, w_274_1199, w_274_1202, w_274_1233, w_274_1240, w_274_1241, w_274_1257, w_274_1263, w_274_1267, w_274_1275, w_274_1282, w_274_1283, w_274_1286, w_274_1289, w_274_1290, w_274_1293, w_274_1295, w_274_1299, w_274_1302, w_274_1318, w_274_1361, w_274_1374, w_274_1404, w_274_1428, w_274_1480, w_274_1487, w_274_1491, w_274_1512, w_274_1523, w_274_1538, w_274_1576, w_274_1580, w_274_1586, w_274_1597, w_274_1604, w_274_1615, w_274_1618, w_274_1638, w_274_1642, w_274_1644, w_274_1653, w_274_1668, w_274_1669, w_274_1670, w_274_1673, w_274_1698, w_274_1704, w_274_1709, w_274_1714, w_274_1721, w_274_1725, w_274_1737, w_274_1769, w_274_1799, w_274_1802, w_274_1805, w_274_1824, w_274_1863, w_274_1870, w_274_1883, w_274_1884, w_274_1898, w_274_1906, w_274_1910, w_274_1913, w_274_1939, w_274_1957, w_274_1996, w_274_1997, w_274_2005, w_274_2016, w_274_2040, w_274_2056, w_274_2062, w_274_2066, w_274_2084, w_274_2087, w_274_2116, w_274_2119, w_274_2122, w_274_2134, w_274_2140, w_274_2141, w_274_2157, w_274_2196, w_274_2208, w_274_2210, w_274_2214, w_274_2218, w_274_2288, w_274_2292, w_274_2295, w_274_2300, w_274_2306, w_274_2314, w_274_2316, w_274_2329, w_274_2406, w_274_2464, w_274_2504, w_274_2507, w_274_2511, w_274_2532, w_274_2538, w_274_2543, w_274_2560, w_274_2562, w_274_2565, w_274_2578, w_274_2586, w_274_2588, w_274_2602, w_274_2609, w_274_2616, w_274_2620, w_274_2625, w_274_2644, w_274_2646, w_274_2650, w_274_2669, w_274_2708, w_274_2714, w_274_2722, w_274_2731, w_274_2735, w_274_2752, w_274_2767, w_274_2777, w_274_2812, w_274_2820, w_274_2833, w_274_2845, w_274_2848, w_274_2853, w_274_2860, w_274_2881, w_274_2915, w_274_2943, w_274_2950, w_274_2954, w_274_2981, w_274_2982, w_274_2997, w_274_3012, w_274_3015, w_274_3017, w_274_3028, w_274_3040, w_274_3046, w_274_3053, w_274_3064, w_274_3069, w_274_3097, w_274_3167, w_274_3174, w_274_3177, w_274_3210, w_274_3241, w_274_3246, w_274_3295, w_274_3301, w_274_3304, w_274_3317, w_274_3327, w_274_3342, w_274_3358, w_274_3367, w_274_3369, w_274_3385, w_274_3404, w_274_3408, w_274_3418, w_274_3439, w_274_3447, w_274_3450, w_274_3455, w_274_3479, w_274_3507, w_274_3532, w_274_3540, w_274_3567, w_274_3583, w_274_3619, w_274_3628, w_274_3630, w_274_3640, w_274_3642, w_274_3679, w_274_3681, w_274_3691, w_274_3696, w_274_3707, w_274_3710, w_274_3711, w_274_3712, w_274_3713, w_274_3714, w_274_3715, w_274_3716, w_274_3717, w_274_3718, w_274_3719, w_274_3720, w_274_3722;
  wire w_275_000, w_275_001, w_275_002, w_275_003, w_275_005, w_275_007, w_275_012, w_275_015, w_275_020, w_275_022, w_275_023, w_275_026, w_275_028, w_275_038, w_275_047, w_275_048, w_275_050, w_275_054, w_275_057, w_275_058, w_275_060, w_275_064, w_275_065, w_275_066, w_275_067, w_275_069, w_275_071, w_275_082, w_275_087, w_275_093, w_275_096, w_275_101, w_275_103, w_275_107, w_275_120, w_275_124, w_275_132, w_275_133, w_275_134, w_275_146, w_275_163, w_275_167, w_275_170, w_275_181, w_275_183, w_275_185, w_275_186, w_275_192, w_275_193, w_275_198, w_275_202, w_275_203, w_275_208, w_275_214, w_275_217, w_275_218, w_275_220, w_275_221, w_275_236, w_275_239, w_275_240, w_275_241, w_275_247, w_275_251, w_275_260, w_275_276, w_275_279, w_275_283, w_275_287, w_275_290, w_275_293, w_275_295, w_275_297, w_275_299, w_275_305, w_275_308, w_275_310, w_275_312, w_275_323, w_275_326, w_275_327, w_275_343, w_275_349, w_275_353, w_275_357, w_275_360, w_275_361, w_275_368, w_275_369, w_275_371, w_275_378, w_275_388, w_275_399, w_275_400, w_275_410, w_275_411, w_275_413, w_275_418, w_275_419, w_275_424, w_275_433, w_275_445, w_275_446, w_275_451, w_275_458, w_275_466, w_275_467, w_275_473, w_275_475, w_275_479, w_275_489, w_275_496, w_275_499, w_275_505, w_275_513, w_275_518, w_275_523, w_275_524, w_275_526, w_275_527, w_275_529, w_275_532, w_275_533, w_275_539, w_275_541, w_275_544, w_275_546, w_275_550, w_275_553, w_275_556, w_275_561, w_275_572, w_275_573, w_275_574, w_275_591, w_275_593, w_275_600, w_275_605, w_275_608, w_275_610, w_275_622, w_275_624, w_275_635, w_275_641, w_275_642, w_275_653, w_275_656, w_275_658, w_275_660, w_275_662, w_275_665, w_275_666, w_275_671, w_275_681, w_275_683, w_275_686, w_275_687, w_275_688, w_275_691, w_275_714, w_275_717, w_275_719, w_275_721, w_275_723, w_275_728, w_275_732, w_275_733, w_275_738, w_275_741, w_275_743, w_275_744, w_275_757, w_275_758, w_275_766, w_275_767, w_275_769, w_275_774, w_275_778, w_275_789, w_275_798, w_275_804, w_275_811, w_275_813, w_275_817, w_275_820, w_275_843, w_275_845, w_275_848, w_275_850, w_275_862, w_275_870, w_275_872, w_275_873, w_275_880, w_275_889, w_275_900, w_275_901, w_275_902, w_275_906, w_275_916, w_275_931, w_275_940, w_275_954, w_275_962, w_275_964, w_275_965, w_275_970, w_275_971, w_275_973, w_275_985, w_275_987, w_275_1008, w_275_1010, w_275_1019, w_275_1027, w_275_1037, w_275_1052, w_275_1056, w_275_1083, w_275_1089, w_275_1093, w_275_1111, w_275_1117, w_275_1139, w_275_1177, w_275_1181, w_275_1184, w_275_1186, w_275_1195, w_275_1204, w_275_1207, w_275_1213, w_275_1216, w_275_1220, w_275_1226, w_275_1229, w_275_1242, w_275_1244, w_275_1261, w_275_1264, w_275_1274, w_275_1276, w_275_1283, w_275_1286, w_275_1294, w_275_1295, w_275_1302, w_275_1311, w_275_1313, w_275_1315, w_275_1320, w_275_1339, w_275_1340, w_275_1343, w_275_1355, w_275_1359, w_275_1360, w_275_1383, w_275_1388, w_275_1389, w_275_1392, w_275_1397, w_275_1403, w_275_1423, w_275_1433, w_275_1449, w_275_1451, w_275_1461, w_275_1475, w_275_1480, w_275_1487, w_275_1494, w_275_1514, w_275_1519, w_275_1521, w_275_1524, w_275_1530, w_275_1531, w_275_1533, w_275_1542, w_275_1545, w_275_1546, w_275_1551, w_275_1564, w_275_1566, w_275_1581, w_275_1584, w_275_1601, w_275_1604, w_275_1613, w_275_1621, w_275_1625, w_275_1630, w_275_1631, w_275_1634, w_275_1646, w_275_1659, w_275_1675, w_275_1679, w_275_1693, w_275_1702, w_275_1704, w_275_1712, w_275_1715, w_275_1716, w_275_1721, w_275_1727, w_275_1730, w_275_1739, w_275_1748, w_275_1750, w_275_1756, w_275_1762, w_275_1768, w_275_1783, w_275_1792, w_275_1797, w_275_1798, w_275_1807, w_275_1815, w_275_1835, w_275_1883, w_275_1889, w_275_1892, w_275_1899, w_275_1901, w_275_1907, w_275_1914, w_275_1916, w_275_1917, w_275_1934, w_275_1935, w_275_1941, w_275_1945, w_275_1952, w_275_1955, w_275_1966, w_275_1997, w_275_2011, w_275_2027, w_275_2030, w_275_2040, w_275_2050, w_275_2052, w_275_2053, w_275_2055, w_275_2066, w_275_2075, w_275_2076, w_275_2080, w_275_2081, w_275_2095, w_275_2098, w_275_2121, w_275_2124, w_275_2129, w_275_2133, w_275_2141, w_275_2142, w_275_2154, w_275_2159, w_275_2161, w_275_2175, w_275_2176, w_275_2177, w_275_2189, w_275_2192, w_275_2200, w_275_2207, w_275_2211, w_275_2212, w_275_2213, w_275_2229, w_275_2232;
  wire w_276_000, w_276_001, w_276_002, w_276_006, w_276_010, w_276_011, w_276_012, w_276_014, w_276_015, w_276_017, w_276_018, w_276_027, w_276_033, w_276_035, w_276_039, w_276_041, w_276_043, w_276_047, w_276_048, w_276_051, w_276_064, w_276_071, w_276_079, w_276_088, w_276_089, w_276_093, w_276_094, w_276_096, w_276_097, w_276_098, w_276_104, w_276_107, w_276_108, w_276_109, w_276_110, w_276_111, w_276_114, w_276_116, w_276_118, w_276_123, w_276_125, w_276_126, w_276_127, w_276_129, w_276_133, w_276_137, w_276_141, w_276_142, w_276_149, w_276_150, w_276_152, w_276_155, w_276_156, w_276_158, w_276_159, w_276_164, w_276_166, w_276_167, w_276_169, w_276_170, w_276_173, w_276_174, w_276_175, w_276_178, w_276_179, w_276_182, w_276_186, w_276_187, w_276_193, w_276_198, w_276_200, w_276_201, w_276_206, w_276_209, w_276_211, w_276_212, w_276_215, w_276_216, w_276_219, w_276_220, w_276_222, w_276_223, w_276_226, w_276_228, w_276_231, w_276_238, w_276_239, w_276_243, w_276_246, w_276_247, w_276_250, w_276_252, w_276_254, w_276_257, w_276_258, w_276_260, w_276_263, w_276_267, w_276_268, w_276_269, w_276_275, w_276_276, w_276_284, w_276_295, w_276_305, w_276_307, w_276_309, w_276_310, w_276_311, w_276_313, w_276_318, w_276_319, w_276_320, w_276_323, w_276_326, w_276_327, w_276_331, w_276_332, w_276_347, w_276_349, w_276_350, w_276_356, w_276_357, w_276_358, w_276_360, w_276_362, w_276_366, w_276_371, w_276_372, w_276_374, w_276_375, w_276_376, w_276_377, w_276_378, w_276_384, w_276_389, w_276_390, w_276_391, w_276_395, w_276_399, w_276_402, w_276_404, w_276_408, w_276_411, w_276_413, w_276_415, w_276_417, w_276_418, w_276_425, w_276_427, w_276_431, w_276_432, w_276_443, w_276_444, w_276_446, w_276_457, w_276_466, w_276_469, w_276_470, w_276_472, w_276_481, w_276_484, w_276_486, w_276_492, w_276_493, w_276_494, w_276_497, w_276_499, w_276_500, w_276_501, w_276_502, w_276_503, w_276_506, w_276_511, w_276_521, w_276_524, w_276_525, w_276_526, w_276_527, w_276_530, w_276_533, w_276_534, w_276_537, w_276_539, w_276_541, w_276_542, w_276_546, w_276_547, w_276_549, w_276_551, w_276_552, w_276_553, w_276_554, w_276_556, w_276_560, w_276_561, w_276_562, w_276_566, w_276_567, w_276_568, w_276_574, w_276_575, w_276_576, w_276_578, w_276_579, w_276_580, w_276_581, w_276_582, w_276_584, w_276_587, w_276_595, w_276_600, w_276_609, w_276_612, w_276_614, w_276_618, w_276_619, w_276_622, w_276_624, w_276_625, w_276_629, w_276_630, w_276_633, w_276_634, w_276_638, w_276_646, w_276_647, w_276_649, w_276_652, w_276_653, w_276_654, w_276_656, w_276_658, w_276_660, w_276_662, w_276_667, w_276_672, w_276_673, w_276_677, w_276_678, w_276_679, w_276_680, w_276_683, w_276_685, w_276_687, w_276_688, w_276_690, w_276_694, w_276_701, w_276_703, w_276_704, w_276_706, w_276_709, w_276_715, w_276_720, w_276_724, w_276_726, w_276_727, w_276_728, w_276_730, w_276_732, w_276_735, w_276_739, w_276_744, w_276_750, w_276_752, w_276_753, w_276_762, w_276_765, w_276_772, w_276_774, w_276_777, w_276_778, w_276_779, w_276_787, w_276_793, w_276_794, w_276_797, w_276_798, w_276_801, w_276_804, w_276_807, w_276_820, w_276_821, w_276_828, w_276_835, w_276_839, w_276_842, w_276_852, w_276_856, w_276_859, w_276_862, w_276_865, w_276_867, w_276_871, w_276_875, w_276_877, w_276_878, w_276_879, w_276_889, w_276_896, w_276_905, w_276_906, w_276_907, w_276_908, w_276_909, w_276_911, w_276_915, w_276_919, w_276_929, w_276_935, w_276_941, w_276_952, w_276_953, w_276_955, w_276_957, w_276_960, w_276_968, w_276_975, w_276_979, w_276_987, w_276_993, w_276_995, w_276_997, w_276_998, w_276_1005, w_276_1007, w_276_1013, w_276_1014, w_276_1017, w_276_1022, w_276_1030, w_276_1031, w_276_1034, w_276_1037, w_276_1042, w_276_1044, w_276_1064, w_276_1065, w_276_1072, w_276_1077;
  wire w_277_001, w_277_003, w_277_005, w_277_006, w_277_009, w_277_010, w_277_011, w_277_014, w_277_015, w_277_018, w_277_019, w_277_020, w_277_021, w_277_022, w_277_024, w_277_026, w_277_027, w_277_031, w_277_032, w_277_034, w_277_039, w_277_041, w_277_042, w_277_043, w_277_045, w_277_046, w_277_047, w_277_050, w_277_052, w_277_053, w_277_054, w_277_055, w_277_057, w_277_059, w_277_060, w_277_061, w_277_062, w_277_066, w_277_067, w_277_068, w_277_069, w_277_071, w_277_074, w_277_075, w_277_079, w_277_080, w_277_084, w_277_089, w_277_092, w_277_099, w_277_105, w_277_110, w_277_111, w_277_112, w_277_113, w_277_114, w_277_117, w_277_118, w_277_119, w_277_120, w_277_121, w_277_122, w_277_123, w_277_124, w_277_125, w_277_126, w_277_128, w_277_129, w_277_130, w_277_135, w_277_138, w_277_140, w_277_141, w_277_143, w_277_144, w_277_147, w_277_149, w_277_155, w_277_156, w_277_158, w_277_159, w_277_164, w_277_166, w_277_167, w_277_169, w_277_171, w_277_176, w_277_177, w_277_178, w_277_179, w_277_182, w_277_183, w_277_184, w_277_185, w_277_186, w_277_189, w_277_190, w_277_192, w_277_193, w_277_199, w_277_200, w_277_202, w_277_203, w_277_204, w_277_208, w_277_213, w_277_218, w_277_222, w_277_224, w_277_226, w_277_227, w_277_229, w_277_230, w_277_231, w_277_234, w_277_235, w_277_236, w_277_237, w_277_239, w_277_242, w_277_243, w_277_244, w_277_247, w_277_249, w_277_252, w_277_260, w_277_264, w_277_266, w_277_267, w_277_271, w_277_275, w_277_276, w_277_277, w_277_281, w_277_282, w_277_283, w_277_286, w_277_287, w_277_288, w_277_290, w_277_294, w_277_295, w_277_297, w_277_299, w_277_301, w_277_305, w_277_307, w_277_311, w_277_314, w_277_315, w_277_317, w_277_318, w_277_319, w_277_323, w_277_324, w_277_325, w_277_326, w_277_327, w_277_329, w_277_335, w_277_336, w_277_337, w_277_338, w_277_343, w_277_344, w_277_347, w_277_348, w_277_354, w_277_355, w_277_357, w_277_359, w_277_361, w_277_363, w_277_365, w_277_366, w_277_367, w_277_370, w_277_371, w_277_372, w_277_374, w_277_378, w_277_379, w_277_382, w_277_388, w_277_394, w_277_396, w_277_398, w_277_400, w_277_409, w_277_415, w_277_418, w_277_419, w_277_420, w_277_422, w_277_424, w_277_428, w_277_433, w_277_434, w_277_436, w_277_440, w_277_441, w_277_443, w_277_445, w_277_447, w_277_450, w_277_451, w_277_452, w_277_455, w_277_456, w_277_458, w_277_460, w_277_465, w_277_466, w_277_467, w_277_470, w_277_472, w_277_474, w_277_475, w_277_477, w_277_478, w_277_480, w_277_481, w_277_482, w_277_483, w_277_484, w_277_485, w_277_486, w_277_489, w_277_490, w_277_493, w_277_500, w_277_501, w_277_503, w_277_504, w_277_505, w_277_511, w_277_512, w_277_513, w_277_516, w_277_517, w_277_522, w_277_523, w_277_525, w_277_527, w_277_529, w_277_530, w_277_531, w_277_533, w_277_534, w_277_537, w_277_541, w_277_542, w_277_543, w_277_544, w_277_545, w_277_547, w_277_551, w_277_552, w_277_554, w_277_557, w_277_563, w_277_567, w_277_568, w_277_570, w_277_574, w_277_575, w_277_578, w_277_580, w_277_581, w_277_586, w_277_587, w_277_591, w_277_594, w_277_598, w_277_600, w_277_601, w_277_604, w_277_608, w_277_609, w_277_612, w_277_613, w_277_614, w_277_617, w_277_618, w_277_619, w_277_622, w_277_623, w_277_624, w_277_625, w_277_631, w_277_634, w_277_636, w_277_640, w_277_641, w_277_642, w_277_644, w_277_646, w_277_648, w_277_651, w_277_652, w_277_656;
  wire w_278_007, w_278_013, w_278_014, w_278_015, w_278_028, w_278_037, w_278_039, w_278_042, w_278_045, w_278_046, w_278_051, w_278_055, w_278_069, w_278_082, w_278_086, w_278_088, w_278_090, w_278_091, w_278_101, w_278_117, w_278_123, w_278_133, w_278_135, w_278_140, w_278_146, w_278_152, w_278_161, w_278_165, w_278_166, w_278_169, w_278_172, w_278_173, w_278_179, w_278_182, w_278_183, w_278_188, w_278_189, w_278_202, w_278_206, w_278_207, w_278_209, w_278_218, w_278_220, w_278_224, w_278_226, w_278_231, w_278_233, w_278_237, w_278_240, w_278_249, w_278_250, w_278_257, w_278_258, w_278_262, w_278_264, w_278_269, w_278_277, w_278_278, w_278_280, w_278_282, w_278_283, w_278_285, w_278_293, w_278_294, w_278_297, w_278_300, w_278_302, w_278_306, w_278_307, w_278_310, w_278_314, w_278_317, w_278_318, w_278_319, w_278_336, w_278_337, w_278_342, w_278_343, w_278_349, w_278_352, w_278_354, w_278_360, w_278_367, w_278_371, w_278_373, w_278_376, w_278_380, w_278_384, w_278_393, w_278_406, w_278_411, w_278_413, w_278_420, w_278_436, w_278_438, w_278_441, w_278_445, w_278_446, w_278_447, w_278_449, w_278_450, w_278_454, w_278_462, w_278_469, w_278_476, w_278_477, w_278_479, w_278_481, w_278_485, w_278_493, w_278_494, w_278_495, w_278_496, w_278_497, w_278_500, w_278_501, w_278_508, w_278_509, w_278_511, w_278_513, w_278_514, w_278_516, w_278_523, w_278_538, w_278_539, w_278_552, w_278_555, w_278_558, w_278_559, w_278_561, w_278_563, w_278_564, w_278_566, w_278_571, w_278_576, w_278_580, w_278_584, w_278_587, w_278_594, w_278_595, w_278_596, w_278_601, w_278_604, w_278_607, w_278_608, w_278_612, w_278_614, w_278_618, w_278_622, w_278_626, w_278_628, w_278_640, w_278_647, w_278_653, w_278_656, w_278_659, w_278_663, w_278_668, w_278_672, w_278_674, w_278_678, w_278_691, w_278_693, w_278_694, w_278_702, w_278_709, w_278_711, w_278_712, w_278_719, w_278_728, w_278_730, w_278_733, w_278_740, w_278_741, w_278_743, w_278_749, w_278_756, w_278_757, w_278_758, w_278_775, w_278_780, w_278_784, w_278_786, w_278_794, w_278_797, w_278_799, w_278_805, w_278_810, w_278_811, w_278_822, w_278_826, w_278_829, w_278_830, w_278_833, w_278_837, w_278_838, w_278_839, w_278_840, w_278_841, w_278_842, w_278_845, w_278_848, w_278_852, w_278_854, w_278_857, w_278_863, w_278_868, w_278_874, w_278_882, w_278_889, w_278_893, w_278_895, w_278_902, w_278_904, w_278_912, w_278_923, w_278_927, w_278_935, w_278_942, w_278_943, w_278_950, w_278_951, w_278_957, w_278_960, w_278_969, w_278_972, w_278_979, w_278_984, w_278_985, w_278_987, w_278_991, w_278_992, w_278_995, w_278_1009, w_278_1012, w_278_1018, w_278_1020, w_278_1024, w_278_1032, w_278_1033, w_278_1040, w_278_1047, w_278_1055, w_278_1058, w_278_1059, w_278_1065, w_278_1067, w_278_1070, w_278_1075, w_278_1080, w_278_1090, w_278_1097, w_278_1101, w_278_1102, w_278_1104, w_278_1106, w_278_1110, w_278_1113, w_278_1114, w_278_1115, w_278_1119, w_278_1121, w_278_1137, w_278_1138, w_278_1146, w_278_1147, w_278_1168, w_278_1174, w_278_1188, w_278_1196, w_278_1199, w_278_1200, w_278_1205, w_278_1206, w_278_1208, w_278_1211, w_278_1216, w_278_1221, w_278_1225, w_278_1226, w_278_1229, w_278_1232, w_278_1239, w_278_1248, w_278_1251, w_278_1252, w_278_1256, w_278_1259, w_278_1264, w_278_1277, w_278_1280, w_278_1283, w_278_1285, w_278_1286, w_278_1300, w_278_1301, w_278_1305, w_278_1310, w_278_1311, w_278_1312, w_278_1321, w_278_1323, w_278_1338, w_278_1339, w_278_1346, w_278_1347, w_278_1350, w_278_1356, w_278_1368, w_278_1376, w_278_1391, w_278_1399, w_278_1406, w_278_1407, w_278_1408, w_278_1426, w_278_1432, w_278_1435, w_278_1438, w_278_1442, w_278_1454, w_278_1461, w_278_1466, w_278_1468, w_278_1487, w_278_1505, w_278_1509, w_278_1514, w_278_1519, w_278_1520, w_278_1521, w_278_1529, w_278_1535, w_278_1553, w_278_1555, w_278_1558, w_278_1569, w_278_1571, w_278_1585, w_278_1586, w_278_1587, w_278_1595, w_278_1596, w_278_1598, w_278_1605, w_278_1607, w_278_1611, w_278_1624, w_278_1632, w_278_1636, w_278_1642, w_278_1647, w_278_1652, w_278_1656, w_278_1661, w_278_1664, w_278_1668, w_278_1672, w_278_1678, w_278_1680, w_278_1708, w_278_1723, w_278_1724, w_278_1726, w_278_1727, w_278_1730, w_278_1735, w_278_1737, w_278_1740, w_278_1743, w_278_1744, w_278_1752, w_278_1755, w_278_1759, w_278_1768, w_278_1774, w_278_1782, w_278_1786, w_278_1792, w_278_1794, w_278_1803, w_278_1809, w_278_1817, w_278_1818, w_278_1823, w_278_1845, w_278_1846, w_278_1847, w_278_1848, w_278_1849, w_278_1850, w_278_1854, w_278_1855, w_278_1856, w_278_1857, w_278_1859;
  wire w_279_001, w_279_002, w_279_004, w_279_008, w_279_011, w_279_013, w_279_014, w_279_016, w_279_018, w_279_026, w_279_027, w_279_028, w_279_029, w_279_032, w_279_034, w_279_035, w_279_037, w_279_038, w_279_040, w_279_042, w_279_043, w_279_046, w_279_048, w_279_049, w_279_052, w_279_056, w_279_057, w_279_059, w_279_064, w_279_065, w_279_067, w_279_070, w_279_075, w_279_078, w_279_080, w_279_082, w_279_084, w_279_085, w_279_086, w_279_088, w_279_092, w_279_094, w_279_097, w_279_100, w_279_108, w_279_110, w_279_113, w_279_115, w_279_116, w_279_117, w_279_119, w_279_125, w_279_127, w_279_133, w_279_135, w_279_138, w_279_139, w_279_142, w_279_147, w_279_148, w_279_152, w_279_153, w_279_156, w_279_158, w_279_159, w_279_163, w_279_164, w_279_167, w_279_171, w_279_174, w_279_175, w_279_176, w_279_177, w_279_180, w_279_184, w_279_185, w_279_186, w_279_189, w_279_191, w_279_193, w_279_196, w_279_197, w_279_198, w_279_200, w_279_205, w_279_206, w_279_212, w_279_213, w_279_215, w_279_216, w_279_217, w_279_219, w_279_220, w_279_221, w_279_225, w_279_230, w_279_233, w_279_235, w_279_240, w_279_242, w_279_243, w_279_246, w_279_250, w_279_251, w_279_252, w_279_255, w_279_258, w_279_265, w_279_269, w_279_271, w_279_273, w_279_275, w_279_276, w_279_277, w_279_279, w_279_280, w_279_282, w_279_283, w_279_285, w_279_286, w_279_292, w_279_297, w_279_300, w_279_304, w_279_306, w_279_307, w_279_309, w_279_311, w_279_313, w_279_317, w_279_318, w_279_320, w_279_321, w_279_329, w_279_333, w_279_334, w_279_336, w_279_338, w_279_339, w_279_340, w_279_343, w_279_350, w_279_352, w_279_355, w_279_356, w_279_363, w_279_369, w_279_374, w_279_377, w_279_378, w_279_380, w_279_385, w_279_387, w_279_388, w_279_394, w_279_395, w_279_398, w_279_399, w_279_401, w_279_403, w_279_404, w_279_405, w_279_409, w_279_411, w_279_412, w_279_414, w_279_421, w_279_427, w_279_428, w_279_429, w_279_430, w_279_431, w_279_432, w_279_441, w_279_447, w_279_453, w_279_459, w_279_461, w_279_463, w_279_464, w_279_467, w_279_479, w_279_482, w_279_484, w_279_489, w_279_491, w_279_497, w_279_499, w_279_502, w_279_505, w_279_507, w_279_511, w_279_513, w_279_527, w_279_529, w_279_533, w_279_536, w_279_538, w_279_540, w_279_541, w_279_543, w_279_546, w_279_548, w_279_554, w_279_556, w_279_560, w_279_570, w_279_578, w_279_580, w_279_586, w_279_587, w_279_589, w_279_599, w_279_600, w_279_601, w_279_606, w_279_607, w_279_610, w_279_613, w_279_621, w_279_624, w_279_626, w_279_635, w_279_636, w_279_641, w_279_642, w_279_646, w_279_647, w_279_650, w_279_653, w_279_658, w_279_663, w_279_664, w_279_668, w_279_670, w_279_672, w_279_676, w_279_677, w_279_685, w_279_694, w_279_695, w_279_699, w_279_701, w_279_707, w_279_712, w_279_720, w_279_721, w_279_727, w_279_734, w_279_736, w_279_737, w_279_743, w_279_745, w_279_754, w_279_756, w_279_758, w_279_760, w_279_763, w_279_765, w_279_775, w_279_786, w_279_788, w_279_795, w_279_797, w_279_799, w_279_801, w_279_803, w_279_805, w_279_809, w_279_810, w_279_815, w_279_824, w_279_825, w_279_826, w_279_830, w_279_832, w_279_836, w_279_838, w_279_842, w_279_848, w_279_851, w_279_856, w_279_859, w_279_861, w_279_862, w_279_865, w_279_866, w_279_869, w_279_874, w_279_875, w_279_876, w_279_877, w_279_883, w_279_888, w_279_897, w_279_904, w_279_909, w_279_912, w_279_917, w_279_921, w_279_925, w_279_926, w_279_929, w_279_930, w_279_935, w_279_936, w_279_938, w_279_939, w_279_945, w_279_949, w_279_952, w_279_955, w_279_957, w_279_959, w_279_962, w_279_965, w_279_966, w_279_967, w_279_969, w_279_972, w_279_974, w_279_976, w_279_977, w_279_978, w_279_982, w_279_990, w_279_993, w_279_994, w_279_997, w_279_999, w_279_1005, w_279_1007, w_279_1009, w_279_1010, w_279_1012, w_279_1013, w_279_1015, w_279_1020, w_279_1021, w_279_1023, w_279_1026, w_279_1028, w_279_1029, w_279_1033, w_279_1034, w_279_1039, w_279_1044, w_279_1046, w_279_1049, w_279_1055, w_279_1058, w_279_1060, w_279_1073, w_279_1090, w_279_1094, w_279_1096, w_279_1097, w_279_1099, w_279_1102, w_279_1106, w_279_1108, w_279_1109, w_279_1115, w_279_1117, w_279_1119, w_279_1120, w_279_1121, w_279_1124, w_279_1131, w_279_1134, w_279_1149, w_279_1150, w_279_1151, w_279_1152, w_279_1153, w_279_1154, w_279_1155, w_279_1156, w_279_1157, w_279_1158, w_279_1159, w_279_1160, w_279_1164, w_279_1165, w_279_1166, w_279_1167, w_279_1168, w_279_1170;
  wire w_280_003, w_280_005, w_280_006, w_280_012, w_280_026, w_280_037, w_280_038, w_280_041, w_280_043, w_280_054, w_280_066, w_280_068, w_280_077, w_280_079, w_280_082, w_280_085, w_280_091, w_280_105, w_280_111, w_280_113, w_280_115, w_280_119, w_280_128, w_280_138, w_280_143, w_280_148, w_280_149, w_280_152, w_280_158, w_280_170, w_280_180, w_280_181, w_280_183, w_280_185, w_280_192, w_280_193, w_280_194, w_280_201, w_280_204, w_280_208, w_280_209, w_280_218, w_280_220, w_280_222, w_280_225, w_280_229, w_280_232, w_280_236, w_280_240, w_280_243, w_280_246, w_280_252, w_280_253, w_280_257, w_280_267, w_280_271, w_280_273, w_280_275, w_280_284, w_280_292, w_280_307, w_280_308, w_280_318, w_280_321, w_280_336, w_280_338, w_280_344, w_280_358, w_280_361, w_280_385, w_280_394, w_280_399, w_280_400, w_280_402, w_280_404, w_280_430, w_280_432, w_280_434, w_280_438, w_280_454, w_280_455, w_280_464, w_280_471, w_280_472, w_280_487, w_280_501, w_280_502, w_280_505, w_280_506, w_280_509, w_280_512, w_280_516, w_280_519, w_280_521, w_280_539, w_280_540, w_280_544, w_280_549, w_280_553, w_280_554, w_280_556, w_280_558, w_280_563, w_280_564, w_280_581, w_280_583, w_280_591, w_280_596, w_280_604, w_280_609, w_280_610, w_280_623, w_280_624, w_280_626, w_280_642, w_280_645, w_280_648, w_280_650, w_280_651, w_280_652, w_280_655, w_280_658, w_280_659, w_280_660, w_280_665, w_280_668, w_280_674, w_280_675, w_280_693, w_280_696, w_280_700, w_280_726, w_280_744, w_280_775, w_280_776, w_280_778, w_280_781, w_280_782, w_280_786, w_280_789, w_280_790, w_280_793, w_280_801, w_280_806, w_280_814, w_280_816, w_280_825, w_280_829, w_280_840, w_280_847, w_280_866, w_280_873, w_280_882, w_280_893, w_280_897, w_280_909, w_280_923, w_280_926, w_280_929, w_280_940, w_280_959, w_280_963, w_280_967, w_280_970, w_280_994, w_280_998, w_280_999, w_280_1000, w_280_1004, w_280_1006, w_280_1007, w_280_1042, w_280_1046, w_280_1057, w_280_1065, w_280_1070, w_280_1096, w_280_1097, w_280_1102, w_280_1122, w_280_1125, w_280_1126, w_280_1127, w_280_1129, w_280_1131, w_280_1132, w_280_1140, w_280_1148, w_280_1151, w_280_1162, w_280_1163, w_280_1165, w_280_1170, w_280_1188, w_280_1190, w_280_1198, w_280_1205, w_280_1211, w_280_1213, w_280_1215, w_280_1217, w_280_1227, w_280_1244, w_280_1248, w_280_1251, w_280_1253, w_280_1258, w_280_1259, w_280_1265, w_280_1275, w_280_1281, w_280_1326, w_280_1339, w_280_1343, w_280_1344, w_280_1346, w_280_1355, w_280_1381, w_280_1384, w_280_1443, w_280_1445, w_280_1456, w_280_1471, w_280_1473, w_280_1496, w_280_1526, w_280_1539, w_280_1541, w_280_1548, w_280_1566, w_280_1576, w_280_1600, w_280_1619, w_280_1622, w_280_1649, w_280_1680, w_280_1712, w_280_1721, w_280_1730, w_280_1734, w_280_1755, w_280_1766, w_280_1768, w_280_1769, w_280_1797, w_280_1808, w_280_1837, w_280_1852, w_280_1853, w_280_1858, w_280_1865, w_280_1869, w_280_1876, w_280_1888, w_280_1915, w_280_1930, w_280_1933, w_280_1936, w_280_1940, w_280_1949, w_280_1950, w_280_1957, w_280_1969, w_280_2001, w_280_2010, w_280_2029, w_280_2034, w_280_2069, w_280_2072, w_280_2076, w_280_2086, w_280_2101, w_280_2102, w_280_2140, w_280_2152, w_280_2167, w_280_2189, w_280_2194, w_280_2195, w_280_2198, w_280_2205, w_280_2206, w_280_2222, w_280_2225, w_280_2245, w_280_2248, w_280_2252, w_280_2260, w_280_2273, w_280_2277, w_280_2289, w_280_2302, w_280_2327, w_280_2328, w_280_2339, w_280_2350, w_280_2354, w_280_2374, w_280_2378, w_280_2385, w_280_2389, w_280_2413, w_280_2421, w_280_2430, w_280_2431, w_280_2457, w_280_2465, w_280_2513, w_280_2519, w_280_2520, w_280_2526, w_280_2547, w_280_2582, w_280_2591, w_280_2606, w_280_2622, w_280_2624, w_280_2657, w_280_2668, w_280_2669, w_280_2682, w_280_2728, w_280_2743, w_280_2752, w_280_2770, w_280_2771, w_280_2780, w_280_2784, w_280_2786, w_280_2789, w_280_2803, w_280_2812, w_280_2820, w_280_2838, w_280_2839, w_280_2857, w_280_2864, w_280_2883, w_280_2887, w_280_2893, w_280_2916, w_280_2923, w_280_2933, w_280_2939, w_280_2948, w_280_2954, w_280_2968, w_280_3000, w_280_3005, w_280_3009, w_280_3033, w_280_3036, w_280_3040, w_280_3041, w_280_3042, w_280_3048, w_280_3054, w_280_3084, w_280_3097, w_280_3101, w_280_3111, w_280_3120, w_280_3154, w_280_3179, w_280_3187, w_280_3218, w_280_3233, w_280_3243, w_280_3246, w_280_3280, w_280_3300, w_280_3318, w_280_3326, w_280_3345, w_280_3349, w_280_3354, w_280_3376, w_280_3415, w_280_3418, w_280_3421, w_280_3424, w_280_3428, w_280_3453, w_280_3459, w_280_3462, w_280_3473, w_280_3480, w_280_3484, w_280_3498, w_280_3518, w_280_3530, w_280_3532, w_280_3533, w_280_3552, w_280_3556, w_280_3561, w_280_3564, w_280_3565, w_280_3577, w_280_3580, w_280_3616, w_280_3622, w_280_3627, w_280_3635, w_280_3640, w_280_3642, w_280_3653, w_280_3660, w_280_3676, w_280_3678, w_280_3682, w_280_3707;
  wire w_281_008, w_281_010, w_281_015, w_281_017, w_281_023, w_281_033, w_281_044, w_281_045, w_281_052, w_281_060, w_281_062, w_281_064, w_281_068, w_281_084, w_281_085, w_281_089, w_281_100, w_281_103, w_281_108, w_281_120, w_281_123, w_281_124, w_281_136, w_281_143, w_281_150, w_281_157, w_281_168, w_281_181, w_281_189, w_281_191, w_281_192, w_281_193, w_281_200, w_281_215, w_281_223, w_281_227, w_281_238, w_281_248, w_281_249, w_281_250, w_281_257, w_281_258, w_281_260, w_281_266, w_281_267, w_281_269, w_281_277, w_281_289, w_281_304, w_281_314, w_281_322, w_281_333, w_281_348, w_281_358, w_281_396, w_281_406, w_281_413, w_281_415, w_281_427, w_281_428, w_281_433, w_281_447, w_281_472, w_281_476, w_281_491, w_281_539, w_281_544, w_281_545, w_281_548, w_281_550, w_281_552, w_281_554, w_281_557, w_281_576, w_281_581, w_281_604, w_281_614, w_281_624, w_281_634, w_281_652, w_281_656, w_281_659, w_281_706, w_281_716, w_281_737, w_281_740, w_281_753, w_281_763, w_281_773, w_281_776, w_281_777, w_281_793, w_281_816, w_281_818, w_281_839, w_281_854, w_281_857, w_281_877, w_281_887, w_281_919, w_281_940, w_281_941, w_281_944, w_281_981, w_281_996, w_281_999, w_281_1005, w_281_1019, w_281_1027, w_281_1040, w_281_1060, w_281_1065, w_281_1071, w_281_1083, w_281_1089, w_281_1094, w_281_1123, w_281_1127, w_281_1129, w_281_1143, w_281_1163, w_281_1186, w_281_1195, w_281_1247, w_281_1250, w_281_1259, w_281_1269, w_281_1274, w_281_1281, w_281_1314, w_281_1318, w_281_1325, w_281_1329, w_281_1335, w_281_1359, w_281_1365, w_281_1382, w_281_1388, w_281_1406, w_281_1411, w_281_1465, w_281_1470, w_281_1528, w_281_1530, w_281_1550, w_281_1554, w_281_1558, w_281_1559, w_281_1560, w_281_1577, w_281_1593, w_281_1594, w_281_1611, w_281_1647, w_281_1649, w_281_1668, w_281_1688, w_281_1716, w_281_1728, w_281_1729, w_281_1730, w_281_1735, w_281_1740, w_281_1768, w_281_1796, w_281_1807, w_281_1810, w_281_1821, w_281_1824, w_281_1841, w_281_1847, w_281_1857, w_281_1869, w_281_1880, w_281_1927, w_281_1935, w_281_1939, w_281_1946, w_281_1947, w_281_1951, w_281_1986, w_281_2000, w_281_2040, w_281_2047, w_281_2071, w_281_2077, w_281_2079, w_281_2087, w_281_2092, w_281_2100, w_281_2131, w_281_2201, w_281_2217, w_281_2219, w_281_2223, w_281_2227, w_281_2232, w_281_2248, w_281_2249, w_281_2250, w_281_2261, w_281_2264, w_281_2266, w_281_2273, w_281_2296, w_281_2310, w_281_2346, w_281_2348, w_281_2374, w_281_2386, w_281_2406, w_281_2409, w_281_2445, w_281_2465, w_281_2513, w_281_2517, w_281_2518, w_281_2539, w_281_2551, w_281_2563, w_281_2596, w_281_2614, w_281_2630, w_281_2635, w_281_2643, w_281_2650, w_281_2663, w_281_2696, w_281_2702, w_281_2704, w_281_2706, w_281_2717, w_281_2722, w_281_2723, w_281_2759, w_281_2767, w_281_2787, w_281_2798, w_281_2801, w_281_2829, w_281_2853, w_281_2860, w_281_2886, w_281_2892, w_281_2893, w_281_2930, w_281_2931, w_281_2936, w_281_2959, w_281_2989, w_281_2992, w_281_3101, w_281_3146, w_281_3154, w_281_3155, w_281_3159, w_281_3160, w_281_3193, w_281_3194, w_281_3221, w_281_3259, w_281_3272, w_281_3291, w_281_3303, w_281_3327, w_281_3360, w_281_3364, w_281_3383, w_281_3401, w_281_3422, w_281_3445, w_281_3452, w_281_3465, w_281_3480, w_281_3498, w_281_3517, w_281_3539, w_281_3552, w_281_3575, w_281_3583, w_281_3590, w_281_3620, w_281_3669, w_281_3698, w_281_3723, w_281_3737, w_281_3757, w_281_3784, w_281_3823, w_281_3828, w_281_3829, w_281_3834, w_281_3836, w_281_3839, w_281_3853, w_281_3856, w_281_3878, w_281_3881, w_281_3916, w_281_3927, w_281_3928, w_281_3964, w_281_3970, w_281_3983, w_281_3987, w_281_3989, w_281_3994, w_281_3995, w_281_4015, w_281_4042, w_281_4054, w_281_4064, w_281_4080, w_281_4090, w_281_4096, w_281_4105, w_281_4147, w_281_4170, w_281_4172, w_281_4185, w_281_4237, w_281_4238, w_281_4255, w_281_4259, w_281_4261, w_281_4263, w_281_4269, w_281_4282, w_281_4318, w_281_4353, w_281_4360, w_281_4361, w_281_4367, w_281_4373, w_281_4375, w_281_4376, w_281_4394, w_281_4400, w_281_4408, w_281_4419, w_281_4430, w_281_4446, w_281_4455, w_281_4474, w_281_4478, w_281_4487, w_281_4490, w_281_4514, w_281_4515, w_281_4516, w_281_4522, w_281_4542, w_281_4543, w_281_4546, w_281_4547, w_281_4556, w_281_4567, w_281_4571, w_281_4581, w_281_4598, w_281_4599, w_281_4612, w_281_4620, w_281_4627, w_281_4643, w_281_4661, w_281_4666, w_281_4694, w_281_4705, w_281_4706, w_281_4707, w_281_4708, w_281_4709, w_281_4713, w_281_4714, w_281_4715, w_281_4716, w_281_4717, w_281_4718, w_281_4719, w_281_4721;
  wire w_282_007, w_282_012, w_282_014, w_282_016, w_282_020, w_282_021, w_282_023, w_282_028, w_282_033, w_282_034, w_282_038, w_282_039, w_282_041, w_282_042, w_282_043, w_282_047, w_282_049, w_282_050, w_282_069, w_282_073, w_282_074, w_282_076, w_282_077, w_282_080, w_282_084, w_282_086, w_282_087, w_282_094, w_282_096, w_282_097, w_282_100, w_282_101, w_282_102, w_282_107, w_282_108, w_282_109, w_282_110, w_282_116, w_282_118, w_282_119, w_282_123, w_282_126, w_282_128, w_282_130, w_282_133, w_282_136, w_282_144, w_282_152, w_282_153, w_282_157, w_282_160, w_282_165, w_282_169, w_282_173, w_282_176, w_282_177, w_282_178, w_282_185, w_282_187, w_282_197, w_282_201, w_282_205, w_282_206, w_282_207, w_282_208, w_282_209, w_282_212, w_282_220, w_282_223, w_282_224, w_282_227, w_282_231, w_282_232, w_282_237, w_282_239, w_282_243, w_282_246, w_282_256, w_282_261, w_282_262, w_282_264, w_282_270, w_282_271, w_282_272, w_282_274, w_282_275, w_282_278, w_282_284, w_282_286, w_282_294, w_282_295, w_282_296, w_282_297, w_282_303, w_282_306, w_282_307, w_282_310, w_282_311, w_282_312, w_282_318, w_282_328, w_282_330, w_282_333, w_282_335, w_282_339, w_282_342, w_282_345, w_282_348, w_282_350, w_282_351, w_282_352, w_282_355, w_282_359, w_282_361, w_282_362, w_282_365, w_282_366, w_282_371, w_282_373, w_282_374, w_282_376, w_282_378, w_282_381, w_282_385, w_282_386, w_282_393, w_282_394, w_282_395, w_282_399, w_282_402, w_282_403, w_282_404, w_282_406, w_282_412, w_282_415, w_282_418, w_282_423, w_282_424, w_282_425, w_282_427, w_282_428, w_282_430, w_282_443, w_282_450, w_282_454, w_282_455, w_282_456, w_282_459, w_282_461, w_282_463, w_282_464, w_282_468, w_282_471, w_282_472, w_282_476, w_282_477, w_282_479, w_282_480, w_282_487, w_282_488, w_282_492, w_282_499, w_282_501, w_282_505, w_282_506, w_282_508, w_282_521, w_282_523, w_282_524, w_282_525, w_282_533, w_282_535, w_282_536, w_282_538, w_282_540, w_282_542, w_282_544, w_282_545, w_282_547, w_282_549, w_282_550, w_282_553, w_282_561, w_282_562, w_282_566, w_282_570, w_282_584, w_282_590, w_282_591, w_282_592, w_282_607, w_282_608, w_282_614, w_282_619, w_282_624, w_282_635, w_282_636, w_282_642, w_282_644, w_282_646, w_282_649, w_282_650, w_282_660, w_282_662, w_282_663, w_282_667, w_282_671, w_282_674, w_282_676, w_282_679, w_282_681, w_282_685, w_282_688, w_282_691, w_282_692, w_282_694, w_282_696, w_282_699, w_282_702, w_282_706, w_282_716, w_282_717, w_282_720, w_282_728, w_282_735, w_282_740, w_282_747, w_282_759, w_282_764, w_282_766, w_282_773, w_282_777, w_282_781, w_282_782, w_282_784, w_282_785, w_282_788, w_282_789, w_282_790, w_282_792, w_282_793, w_282_802, w_282_803, w_282_805, w_282_809, w_282_813, w_282_817, w_282_821, w_282_823, w_282_824, w_282_825, w_282_827, w_282_831, w_282_832, w_282_836, w_282_837, w_282_839, w_282_842, w_282_843, w_282_846, w_282_848, w_282_852, w_282_854, w_282_855, w_282_860, w_282_862, w_282_866, w_282_867, w_282_871, w_282_874, w_282_876, w_282_877, w_282_883, w_282_885, w_282_889, w_282_891, w_282_892, w_282_901, w_282_909, w_282_910, w_282_912, w_282_913, w_282_914, w_282_915, w_282_917, w_282_918, w_282_922, w_282_941, w_282_944, w_282_946, w_282_947, w_282_949, w_282_959, w_282_960, w_282_963, w_282_964, w_282_972, w_282_976, w_282_977, w_282_981, w_282_985, w_282_989, w_282_990, w_282_997, w_282_998, w_282_1003, w_282_1007, w_282_1011, w_282_1012, w_282_1018, w_282_1021, w_282_1025, w_282_1026, w_282_1029, w_282_1034, w_282_1038, w_282_1041, w_282_1046, w_282_1049, w_282_1050, w_282_1054, w_282_1057, w_282_1060, w_282_1065, w_282_1066, w_282_1071, w_282_1078, w_282_1079, w_282_1082, w_282_1091, w_282_1092, w_282_1093, w_282_1095, w_282_1098, w_282_1105, w_282_1108, w_282_1114, w_282_1115, w_282_1116, w_282_1124;
  wire w_283_003, w_283_004, w_283_005, w_283_009, w_283_011, w_283_013, w_283_016, w_283_017, w_283_020, w_283_022, w_283_026, w_283_029, w_283_038, w_283_040, w_283_042, w_283_046, w_283_049, w_283_054, w_283_071, w_283_079, w_283_082, w_283_088, w_283_092, w_283_108, w_283_120, w_283_122, w_283_126, w_283_136, w_283_143, w_283_154, w_283_163, w_283_166, w_283_176, w_283_181, w_283_185, w_283_193, w_283_196, w_283_197, w_283_198, w_283_201, w_283_204, w_283_236, w_283_243, w_283_245, w_283_246, w_283_248, w_283_252, w_283_254, w_283_256, w_283_269, w_283_274, w_283_279, w_283_280, w_283_284, w_283_287, w_283_288, w_283_292, w_283_295, w_283_301, w_283_307, w_283_320, w_283_329, w_283_330, w_283_333, w_283_335, w_283_341, w_283_347, w_283_349, w_283_351, w_283_352, w_283_360, w_283_361, w_283_375, w_283_376, w_283_382, w_283_384, w_283_385, w_283_386, w_283_391, w_283_395, w_283_396, w_283_401, w_283_405, w_283_414, w_283_422, w_283_425, w_283_426, w_283_435, w_283_442, w_283_449, w_283_451, w_283_454, w_283_470, w_283_474, w_283_480, w_283_484, w_283_500, w_283_510, w_283_513, w_283_515, w_283_521, w_283_522, w_283_524, w_283_529, w_283_533, w_283_549, w_283_560, w_283_566, w_283_569, w_283_582, w_283_594, w_283_599, w_283_603, w_283_606, w_283_612, w_283_616, w_283_626, w_283_633, w_283_634, w_283_638, w_283_640, w_283_649, w_283_650, w_283_652, w_283_654, w_283_662, w_283_664, w_283_665, w_283_666, w_283_669, w_283_675, w_283_676, w_283_678, w_283_683, w_283_686, w_283_688, w_283_692, w_283_694, w_283_703, w_283_707, w_283_709, w_283_712, w_283_723, w_283_731, w_283_735, w_283_751, w_283_759, w_283_761, w_283_771, w_283_774, w_283_776, w_283_781, w_283_786, w_283_788, w_283_790, w_283_792, w_283_795, w_283_799, w_283_809, w_283_813, w_283_817, w_283_818, w_283_820, w_283_824, w_283_827, w_283_831, w_283_834, w_283_838, w_283_841, w_283_844, w_283_852, w_283_857, w_283_859, w_283_875, w_283_884, w_283_890, w_283_894, w_283_898, w_283_899, w_283_902, w_283_904, w_283_908, w_283_909, w_283_912, w_283_914, w_283_915, w_283_920, w_283_924, w_283_927, w_283_933, w_283_935, w_283_937, w_283_939, w_283_946, w_283_947, w_283_960, w_283_962, w_283_965, w_283_966, w_283_969, w_283_971, w_283_976, w_283_979, w_283_980, w_283_985, w_283_986, w_283_991, w_283_994, w_283_997, w_283_1004, w_283_1009, w_283_1014, w_283_1015, w_283_1025, w_283_1032, w_283_1041, w_283_1042, w_283_1044, w_283_1048, w_283_1057, w_283_1069, w_283_1074, w_283_1089, w_283_1090, w_283_1098, w_283_1103, w_283_1104, w_283_1131, w_283_1133, w_283_1145, w_283_1151, w_283_1156, w_283_1164, w_283_1190, w_283_1193, w_283_1194, w_283_1204, w_283_1205, w_283_1211, w_283_1212, w_283_1221, w_283_1226, w_283_1227, w_283_1237, w_283_1239, w_283_1243, w_283_1247, w_283_1251, w_283_1252, w_283_1269, w_283_1292, w_283_1304, w_283_1308, w_283_1313, w_283_1327, w_283_1336, w_283_1339, w_283_1356, w_283_1359, w_283_1361, w_283_1366, w_283_1372, w_283_1381, w_283_1392, w_283_1399, w_283_1405, w_283_1419, w_283_1434, w_283_1441, w_283_1444, w_283_1474, w_283_1480, w_283_1484, w_283_1491, w_283_1493, w_283_1497, w_283_1501, w_283_1503, w_283_1512, w_283_1520, w_283_1524, w_283_1526, w_283_1527, w_283_1529, w_283_1531, w_283_1532, w_283_1533, w_283_1535, w_283_1536, w_283_1539, w_283_1548, w_283_1552, w_283_1557, w_283_1571, w_283_1572, w_283_1583, w_283_1586, w_283_1589, w_283_1591, w_283_1593, w_283_1598, w_283_1601, w_283_1604, w_283_1610, w_283_1615, w_283_1628, w_283_1634, w_283_1637, w_283_1649, w_283_1655, w_283_1664, w_283_1666, w_283_1672, w_283_1679, w_283_1680, w_283_1686, w_283_1687, w_283_1691, w_283_1693, w_283_1694, w_283_1709, w_283_1711, w_283_1724, w_283_1727, w_283_1748, w_283_1763, w_283_1764, w_283_1775, w_283_1778, w_283_1779, w_283_1811, w_283_1821, w_283_1835, w_283_1838, w_283_1840, w_283_1846, w_283_1847, w_283_1853, w_283_1854, w_283_1858, w_283_1859, w_283_1861, w_283_1864, w_283_1880, w_283_1885, w_283_1891, w_283_1892, w_283_1908, w_283_1910, w_283_1916, w_283_1933, w_283_1937, w_283_1943;
  wire w_284_001, w_284_005, w_284_013, w_284_015, w_284_019, w_284_028, w_284_030, w_284_033, w_284_035, w_284_041, w_284_044, w_284_051, w_284_058, w_284_063, w_284_067, w_284_071, w_284_072, w_284_073, w_284_082, w_284_083, w_284_084, w_284_090, w_284_094, w_284_096, w_284_099, w_284_102, w_284_103, w_284_113, w_284_116, w_284_117, w_284_118, w_284_129, w_284_130, w_284_131, w_284_133, w_284_136, w_284_137, w_284_140, w_284_144, w_284_146, w_284_148, w_284_152, w_284_157, w_284_171, w_284_177, w_284_178, w_284_182, w_284_190, w_284_198, w_284_204, w_284_214, w_284_216, w_284_217, w_284_219, w_284_220, w_284_221, w_284_226, w_284_235, w_284_236, w_284_237, w_284_240, w_284_241, w_284_244, w_284_250, w_284_255, w_284_256, w_284_261, w_284_263, w_284_264, w_284_265, w_284_266, w_284_277, w_284_280, w_284_281, w_284_282, w_284_286, w_284_288, w_284_291, w_284_292, w_284_293, w_284_295, w_284_296, w_284_297, w_284_298, w_284_301, w_284_302, w_284_309, w_284_310, w_284_311, w_284_316, w_284_317, w_284_327, w_284_336, w_284_337, w_284_338, w_284_339, w_284_340, w_284_343, w_284_344, w_284_345, w_284_349, w_284_353, w_284_354, w_284_355, w_284_363, w_284_365, w_284_367, w_284_368, w_284_371, w_284_372, w_284_373, w_284_376, w_284_381, w_284_386, w_284_398, w_284_401, w_284_407, w_284_408, w_284_409, w_284_421, w_284_422, w_284_424, w_284_425, w_284_429, w_284_442, w_284_443, w_284_448, w_284_451, w_284_455, w_284_457, w_284_458, w_284_461, w_284_463, w_284_464, w_284_471, w_284_474, w_284_478, w_284_486, w_284_490, w_284_492, w_284_499, w_284_504, w_284_505, w_284_507, w_284_510, w_284_513, w_284_516, w_284_519, w_284_520, w_284_521, w_284_523, w_284_527, w_284_530, w_284_532, w_284_536, w_284_540, w_284_546, w_284_554, w_284_556, w_284_559, w_284_561, w_284_564, w_284_569, w_284_570, w_284_572, w_284_573, w_284_575, w_284_578, w_284_580, w_284_582, w_284_585, w_284_590, w_284_595, w_284_596, w_284_598, w_284_599, w_284_602, w_284_604, w_284_605, w_284_607, w_284_608, w_284_619, w_284_620, w_284_622, w_284_625, w_284_632, w_284_638, w_284_641, w_284_642, w_284_644, w_284_647, w_284_649, w_284_651, w_284_661, w_284_664, w_284_665, w_284_667, w_284_677, w_284_679, w_284_684, w_284_687, w_284_690, w_284_698, w_284_699, w_284_701, w_284_703, w_284_712, w_284_717, w_284_721, w_284_723, w_284_724, w_284_725, w_284_726, w_284_731, w_284_732, w_284_739, w_284_740, w_284_742, w_284_761, w_284_764, w_284_768, w_284_770, w_284_771, w_284_774, w_284_775, w_284_776, w_284_777, w_284_782, w_284_783, w_284_787, w_284_790, w_284_793, w_284_794, w_284_799, w_284_801, w_284_804, w_284_808, w_284_815, w_284_816, w_284_818, w_284_819, w_284_823, w_284_825, w_284_827, w_284_828, w_284_831, w_284_834, w_284_845, w_284_847, w_284_853, w_284_854, w_284_855, w_284_862, w_284_863, w_284_865, w_284_873, w_284_883, w_284_885, w_284_887, w_284_890, w_284_891, w_284_902, w_284_904, w_284_905, w_284_909, w_284_910, w_284_919, w_284_921, w_284_928, w_284_930, w_284_932, w_284_939, w_284_941, w_284_945, w_284_948, w_284_950, w_284_952, w_284_953, w_284_957, w_284_959, w_284_965, w_284_967, w_284_968, w_284_969, w_284_971, w_284_972, w_284_975, w_284_979, w_284_985, w_284_986, w_284_990, w_284_991, w_284_992, w_284_995, w_284_996, w_284_997, w_284_998, w_284_1000, w_284_1013, w_284_1016, w_284_1018, w_284_1035, w_284_1039, w_284_1048, w_284_1049, w_284_1057, w_284_1061, w_284_1066, w_284_1094, w_284_1106, w_284_1111, w_284_1112, w_284_1126, w_284_1127, w_284_1128, w_284_1131, w_284_1138, w_284_1140, w_284_1141, w_284_1148, w_284_1158, w_284_1159, w_284_1167, w_284_1172, w_284_1180, w_284_1181, w_284_1183, w_284_1186, w_284_1190, w_284_1199, w_284_1209, w_284_1214, w_284_1221, w_284_1222, w_284_1223, w_284_1224, w_284_1227, w_284_1229, w_284_1233, w_284_1239, w_284_1240, w_284_1245, w_284_1248, w_284_1264, w_284_1265, w_284_1266, w_284_1271, w_284_1273, w_284_1275, w_284_1276, w_284_1283, w_284_1289, w_284_1307, w_284_1308, w_284_1310, w_284_1311, w_284_1312, w_284_1333, w_284_1334, w_284_1335, w_284_1339, w_284_1340, w_284_1341, w_284_1342, w_284_1343, w_284_1344, w_284_1345, w_284_1347;
  wire w_285_000, w_285_001, w_285_002, w_285_003, w_285_004, w_285_006, w_285_007, w_285_009, w_285_010, w_285_011, w_285_012, w_285_013, w_285_014, w_285_015, w_285_018, w_285_019, w_285_020, w_285_021, w_285_022, w_285_023, w_285_024, w_285_025, w_285_026, w_285_027, w_285_028, w_285_029, w_285_030, w_285_031, w_285_032, w_285_033, w_285_034, w_285_035, w_285_036, w_285_038, w_285_039, w_285_040, w_285_041, w_285_043, w_285_044, w_285_045, w_285_046, w_285_047, w_285_048, w_285_049, w_285_050, w_285_051, w_285_052, w_285_053, w_285_054, w_285_055, w_285_056, w_285_057, w_285_058, w_285_059, w_285_060, w_285_061, w_285_062, w_285_063, w_285_064, w_285_065, w_285_066, w_285_067, w_285_068, w_285_069, w_285_070, w_285_071, w_285_072, w_285_074, w_285_075, w_285_076, w_285_077, w_285_078, w_285_079, w_285_080, w_285_082, w_285_083, w_285_084, w_285_086, w_285_087, w_285_088, w_285_089, w_285_090, w_285_091, w_285_093, w_285_094, w_285_095, w_285_096, w_285_097, w_285_098, w_285_099, w_285_100, w_285_101, w_285_102, w_285_103, w_285_104, w_285_105, w_285_106, w_285_107, w_285_109, w_285_110, w_285_111, w_285_112, w_285_113, w_285_114, w_285_115, w_285_116, w_285_117, w_285_119, w_285_120, w_285_121, w_285_122, w_285_123, w_285_124, w_285_125, w_285_126, w_285_128, w_285_129, w_285_130, w_285_131, w_285_133, w_285_134, w_285_135, w_285_136, w_285_137, w_285_139, w_285_140, w_285_143, w_285_144, w_285_145, w_285_146, w_285_147, w_285_148, w_285_149, w_285_150, w_285_151, w_285_152, w_285_153, w_285_154, w_285_155, w_285_156, w_285_158, w_285_159, w_285_161, w_285_162, w_285_163, w_285_164, w_285_165, w_285_167, w_285_168, w_285_169, w_285_170, w_285_171, w_285_172, w_285_173, w_285_174, w_285_175, w_285_176, w_285_177, w_285_178, w_285_179, w_285_180, w_285_181, w_285_182, w_285_183, w_285_184, w_285_185, w_285_186, w_285_187, w_285_190, w_285_191, w_285_192, w_285_193, w_285_194, w_285_195, w_285_196, w_285_197, w_285_198, w_285_199, w_285_200, w_285_201, w_285_203, w_285_204, w_285_205, w_285_206, w_285_207, w_285_208, w_285_209, w_285_210, w_285_211, w_285_212, w_285_213, w_285_214, w_285_218, w_285_219, w_285_220, w_285_221, w_285_222, w_285_223, w_285_224, w_285_225, w_285_226, w_285_228;
  wire w_286_007, w_286_008, w_286_009, w_286_021, w_286_023, w_286_039, w_286_045, w_286_047, w_286_049, w_286_051, w_286_054, w_286_075, w_286_090, w_286_096, w_286_101, w_286_110, w_286_120, w_286_126, w_286_130, w_286_138, w_286_139, w_286_143, w_286_147, w_286_153, w_286_154, w_286_156, w_286_190, w_286_195, w_286_204, w_286_210, w_286_212, w_286_221, w_286_223, w_286_234, w_286_239, w_286_251, w_286_254, w_286_257, w_286_261, w_286_264, w_286_266, w_286_284, w_286_285, w_286_286, w_286_291, w_286_305, w_286_311, w_286_328, w_286_335, w_286_340, w_286_342, w_286_345, w_286_376, w_286_385, w_286_388, w_286_390, w_286_394, w_286_398, w_286_399, w_286_403, w_286_412, w_286_415, w_286_419, w_286_431, w_286_445, w_286_446, w_286_454, w_286_456, w_286_457, w_286_469, w_286_474, w_286_485, w_286_486, w_286_491, w_286_510, w_286_515, w_286_523, w_286_529, w_286_533, w_286_538, w_286_539, w_286_541, w_286_543, w_286_545, w_286_556, w_286_562, w_286_569, w_286_570, w_286_582, w_286_590, w_286_592, w_286_603, w_286_613, w_286_622, w_286_624, w_286_634, w_286_640, w_286_643, w_286_655, w_286_672, w_286_675, w_286_686, w_286_692, w_286_699, w_286_705, w_286_707, w_286_710, w_286_713, w_286_716, w_286_719, w_286_720, w_286_725, w_286_732, w_286_733, w_286_752, w_286_759, w_286_762, w_286_765, w_286_771, w_286_773, w_286_786, w_286_789, w_286_791, w_286_796, w_286_804, w_286_805, w_286_809, w_286_816, w_286_821, w_286_827, w_286_849, w_286_852, w_286_862, w_286_868, w_286_871, w_286_875, w_286_877, w_286_881, w_286_886, w_286_891, w_286_904, w_286_914, w_286_916, w_286_940, w_286_951, w_286_952, w_286_957, w_286_981, w_286_986, w_286_1010, w_286_1031, w_286_1040, w_286_1056, w_286_1062, w_286_1087, w_286_1114, w_286_1122, w_286_1124, w_286_1128, w_286_1131, w_286_1132, w_286_1173, w_286_1196, w_286_1213, w_286_1218, w_286_1242, w_286_1256, w_286_1259, w_286_1261, w_286_1286, w_286_1309, w_286_1324, w_286_1366, w_286_1410, w_286_1416, w_286_1421, w_286_1425, w_286_1435, w_286_1439, w_286_1457, w_286_1495, w_286_1517, w_286_1519, w_286_1527, w_286_1530, w_286_1535, w_286_1555, w_286_1605, w_286_1606, w_286_1630, w_286_1632, w_286_1644, w_286_1685, w_286_1722, w_286_1739, w_286_1754, w_286_1767, w_286_1814, w_286_1833, w_286_1838, w_286_1839, w_286_1843, w_286_1850, w_286_1863, w_286_1891, w_286_1909, w_286_1911, w_286_1914, w_286_1916, w_286_1925, w_286_1973, w_286_1985, w_286_1992, w_286_2018, w_286_2026, w_286_2027, w_286_2038, w_286_2063, w_286_2068, w_286_2090, w_286_2091, w_286_2106, w_286_2113, w_286_2118, w_286_2128, w_286_2139, w_286_2185, w_286_2200, w_286_2205, w_286_2245, w_286_2256, w_286_2268, w_286_2275, w_286_2284, w_286_2350, w_286_2366, w_286_2369, w_286_2416, w_286_2451, w_286_2452, w_286_2467, w_286_2486, w_286_2518, w_286_2532, w_286_2538, w_286_2569, w_286_2579, w_286_2581, w_286_2601, w_286_2602, w_286_2615, w_286_2626, w_286_2635, w_286_2647, w_286_2673, w_286_2697, w_286_2753, w_286_2754, w_286_2793, w_286_2804, w_286_2818, w_286_2819, w_286_2832, w_286_2843, w_286_2852, w_286_2854, w_286_2855, w_286_2873, w_286_2891, w_286_2892, w_286_2894, w_286_2913, w_286_2915, w_286_2917, w_286_2925, w_286_2931, w_286_2935, w_286_2973, w_286_2982, w_286_2983, w_286_2985, w_286_3005, w_286_3008, w_286_3061, w_286_3072, w_286_3075, w_286_3088, w_286_3095, w_286_3120, w_286_3130, w_286_3142, w_286_3160, w_286_3169, w_286_3173, w_286_3175, w_286_3179, w_286_3194, w_286_3212, w_286_3214, w_286_3220, w_286_3231, w_286_3244, w_286_3255, w_286_3256, w_286_3257, w_286_3258, w_286_3259, w_286_3270, w_286_3280, w_286_3303, w_286_3330, w_286_3356, w_286_3360, w_286_3368, w_286_3384, w_286_3385, w_286_3405, w_286_3431, w_286_3443, w_286_3470, w_286_3481, w_286_3496, w_286_3500, w_286_3501, w_286_3533, w_286_3547, w_286_3566, w_286_3567, w_286_3593, w_286_3612, w_286_3624, w_286_3638, w_286_3648, w_286_3651, w_286_3656, w_286_3663, w_286_3677, w_286_3680, w_286_3696, w_286_3711, w_286_3739, w_286_3759, w_286_3782, w_286_3783, w_286_3786, w_286_3798, w_286_3824, w_286_3845, w_286_3876, w_286_3896, w_286_3965, w_286_3970, w_286_3972, w_286_3985, w_286_4004, w_286_4006, w_286_4007, w_286_4046, w_286_4067, w_286_4087, w_286_4096, w_286_4100, w_286_4105, w_286_4106, w_286_4107, w_286_4108, w_286_4109, w_286_4110, w_286_4111, w_286_4112, w_286_4113, w_286_4114, w_286_4115;
  wire w_287_001, w_287_007, w_287_010, w_287_013, w_287_022, w_287_028, w_287_029, w_287_030, w_287_032, w_287_043, w_287_047, w_287_049, w_287_079, w_287_084, w_287_085, w_287_086, w_287_101, w_287_106, w_287_108, w_287_113, w_287_126, w_287_134, w_287_141, w_287_144, w_287_146, w_287_147, w_287_149, w_287_156, w_287_159, w_287_171, w_287_174, w_287_188, w_287_212, w_287_216, w_287_225, w_287_231, w_287_241, w_287_244, w_287_247, w_287_249, w_287_268, w_287_269, w_287_272, w_287_275, w_287_277, w_287_285, w_287_296, w_287_309, w_287_321, w_287_324, w_287_327, w_287_337, w_287_344, w_287_348, w_287_354, w_287_356, w_287_369, w_287_375, w_287_390, w_287_393, w_287_403, w_287_405, w_287_417, w_287_425, w_287_426, w_287_441, w_287_442, w_287_444, w_287_446, w_287_456, w_287_457, w_287_463, w_287_483, w_287_485, w_287_490, w_287_495, w_287_505, w_287_510, w_287_521, w_287_526, w_287_527, w_287_541, w_287_554, w_287_569, w_287_571, w_287_576, w_287_584, w_287_586, w_287_589, w_287_596, w_287_598, w_287_610, w_287_613, w_287_623, w_287_626, w_287_629, w_287_641, w_287_657, w_287_658, w_287_659, w_287_667, w_287_671, w_287_672, w_287_674, w_287_685, w_287_689, w_287_691, w_287_700, w_287_704, w_287_709, w_287_710, w_287_712, w_287_714, w_287_715, w_287_722, w_287_723, w_287_745, w_287_755, w_287_756, w_287_767, w_287_769, w_287_770, w_287_771, w_287_781, w_287_782, w_287_787, w_287_788, w_287_800, w_287_801, w_287_819, w_287_820, w_287_827, w_287_830, w_287_831, w_287_835, w_287_836, w_287_846, w_287_880, w_287_885, w_287_886, w_287_898, w_287_899, w_287_908, w_287_919, w_287_921, w_287_924, w_287_930, w_287_931, w_287_934, w_287_935, w_287_946, w_287_947, w_287_958, w_287_966, w_287_988, w_287_991, w_287_999, w_287_1000, w_287_1001, w_287_1004, w_287_1032, w_287_1039, w_287_1042, w_287_1050, w_287_1057, w_287_1084, w_287_1093, w_287_1101, w_287_1115, w_287_1119, w_287_1122, w_287_1124, w_287_1128, w_287_1142, w_287_1146, w_287_1153, w_287_1166, w_287_1167, w_287_1178, w_287_1188, w_287_1192, w_287_1203, w_287_1210, w_287_1225, w_287_1234, w_287_1244, w_287_1252, w_287_1255, w_287_1279, w_287_1283, w_287_1307, w_287_1313, w_287_1317, w_287_1329, w_287_1332, w_287_1359, w_287_1372, w_287_1402, w_287_1427, w_287_1457, w_287_1460, w_287_1469, w_287_1475, w_287_1476, w_287_1491, w_287_1493, w_287_1500, w_287_1536, w_287_1540, w_287_1546, w_287_1555, w_287_1561, w_287_1562, w_287_1577, w_287_1585, w_287_1615, w_287_1618, w_287_1645, w_287_1647, w_287_1669, w_287_1721, w_287_1760, w_287_1762, w_287_1814, w_287_1815, w_287_1820, w_287_1839, w_287_1874, w_287_1876, w_287_1885, w_287_1887, w_287_1907, w_287_1915, w_287_1921, w_287_1922, w_287_1975, w_287_1976, w_287_1996, w_287_2008, w_287_2012, w_287_2022, w_287_2026, w_287_2047, w_287_2049, w_287_2053, w_287_2079, w_287_2080, w_287_2084, w_287_2086, w_287_2091, w_287_2109, w_287_2124, w_287_2133, w_287_2143, w_287_2155, w_287_2166, w_287_2187, w_287_2188, w_287_2223, w_287_2250, w_287_2251, w_287_2257, w_287_2259, w_287_2276, w_287_2314, w_287_2330, w_287_2337, w_287_2363, w_287_2386, w_287_2396, w_287_2401, w_287_2407, w_287_2412, w_287_2420, w_287_2438, w_287_2458, w_287_2461, w_287_2466, w_287_2471, w_287_2487, w_287_2503, w_287_2524, w_287_2528, w_287_2541, w_287_2544, w_287_2550, w_287_2552, w_287_2556, w_287_2559, w_287_2561, w_287_2582, w_287_2583, w_287_2589, w_287_2603, w_287_2654, w_287_2671, w_287_2674, w_287_2697, w_287_2724, w_287_2728, w_287_2733, w_287_2747, w_287_2760, w_287_2775, w_287_2788, w_287_2792, w_287_2805, w_287_2810, w_287_2823, w_287_2835, w_287_2844, w_287_2863, w_287_2893, w_287_2904, w_287_2953, w_287_2959, w_287_2977, w_287_2981, w_287_2987, w_287_2992, w_287_2995, w_287_2996, w_287_3017, w_287_3034, w_287_3041, w_287_3046, w_287_3063, w_287_3065, w_287_3081, w_287_3087, w_287_3088, w_287_3106, w_287_3112, w_287_3116, w_287_3118, w_287_3119, w_287_3130, w_287_3152, w_287_3155, w_287_3157, w_287_3172, w_287_3175, w_287_3179, w_287_3194, w_287_3210, w_287_3236, w_287_3262, w_287_3308, w_287_3315, w_287_3333, w_287_3343, w_287_3358, w_287_3359, w_287_3366, w_287_3391, w_287_3400, w_287_3406, w_287_3420, w_287_3424, w_287_3426, w_287_3437, w_287_3444, w_287_3445, w_287_3451, w_287_3476, w_287_3477, w_287_3479, w_287_3503, w_287_3504, w_287_3511, w_287_3517, w_287_3532, w_287_3536, w_287_3550, w_287_3554, w_287_3577, w_287_3591, w_287_3602, w_287_3606, w_287_3618, w_287_3629, w_287_3644, w_287_3667, w_287_3672, w_287_3698, w_287_3702, w_287_3703, w_287_3710, w_287_3726, w_287_3730, w_287_3744, w_287_3756, w_287_3792, w_287_3793, w_287_3802, w_287_3803, w_287_3804, w_287_3805, w_287_3806, w_287_3807, w_287_3811, w_287_3812, w_287_3813, w_287_3814, w_287_3815, w_287_3816, w_287_3817, w_287_3819;
  wire w_288_001, w_288_022, w_288_037, w_288_038, w_288_048, w_288_054, w_288_059, w_288_060, w_288_062, w_288_063, w_288_074, w_288_086, w_288_091, w_288_098, w_288_102, w_288_108, w_288_111, w_288_115, w_288_126, w_288_130, w_288_137, w_288_139, w_288_146, w_288_160, w_288_166, w_288_182, w_288_202, w_288_214, w_288_225, w_288_227, w_288_228, w_288_236, w_288_240, w_288_248, w_288_250, w_288_251, w_288_255, w_288_265, w_288_273, w_288_275, w_288_276, w_288_277, w_288_279, w_288_289, w_288_296, w_288_309, w_288_323, w_288_333, w_288_343, w_288_344, w_288_346, w_288_351, w_288_353, w_288_354, w_288_367, w_288_380, w_288_411, w_288_425, w_288_429, w_288_430, w_288_439, w_288_445, w_288_453, w_288_456, w_288_463, w_288_464, w_288_467, w_288_473, w_288_476, w_288_484, w_288_501, w_288_502, w_288_514, w_288_521, w_288_522, w_288_525, w_288_568, w_288_572, w_288_582, w_288_587, w_288_603, w_288_605, w_288_607, w_288_610, w_288_611, w_288_615, w_288_617, w_288_621, w_288_625, w_288_626, w_288_627, w_288_639, w_288_641, w_288_643, w_288_652, w_288_667, w_288_672, w_288_683, w_288_690, w_288_692, w_288_705, w_288_710, w_288_711, w_288_714, w_288_718, w_288_726, w_288_730, w_288_741, w_288_756, w_288_762, w_288_768, w_288_772, w_288_779, w_288_785, w_288_797, w_288_800, w_288_803, w_288_819, w_288_820, w_288_848, w_288_860, w_288_861, w_288_877, w_288_880, w_288_883, w_288_889, w_288_904, w_288_908, w_288_909, w_288_916, w_288_917, w_288_926, w_288_932, w_288_940, w_288_948, w_288_967, w_288_992, w_288_1004, w_288_1009, w_288_1013, w_288_1015, w_288_1041, w_288_1042, w_288_1044, w_288_1053, w_288_1055, w_288_1062, w_288_1066, w_288_1072, w_288_1074, w_288_1083, w_288_1087, w_288_1113, w_288_1117, w_288_1127, w_288_1133, w_288_1135, w_288_1137, w_288_1139, w_288_1151, w_288_1157, w_288_1159, w_288_1171, w_288_1193, w_288_1200, w_288_1204, w_288_1214, w_288_1218, w_288_1239, w_288_1241, w_288_1257, w_288_1260, w_288_1263, w_288_1270, w_288_1287, w_288_1295, w_288_1308, w_288_1309, w_288_1310, w_288_1316, w_288_1332, w_288_1342, w_288_1344, w_288_1350, w_288_1355, w_288_1364, w_288_1366, w_288_1379, w_288_1381, w_288_1395, w_288_1401, w_288_1402, w_288_1403, w_288_1407, w_288_1411, w_288_1440, w_288_1441, w_288_1468, w_288_1480, w_288_1485, w_288_1489, w_288_1497, w_288_1508, w_288_1511, w_288_1512, w_288_1515, w_288_1530, w_288_1531, w_288_1541, w_288_1543, w_288_1547, w_288_1556, w_288_1562, w_288_1568, w_288_1570, w_288_1573, w_288_1585, w_288_1597, w_288_1602, w_288_1606, w_288_1617, w_288_1624, w_288_1630, w_288_1634, w_288_1637, w_288_1638, w_288_1646, w_288_1655, w_288_1657, w_288_1658, w_288_1664, w_288_1666, w_288_1672, w_288_1674, w_288_1683, w_288_1687, w_288_1688, w_288_1689, w_288_1707, w_288_1710, w_288_1716, w_288_1722, w_288_1726, w_288_1729, w_288_1730, w_288_1735, w_288_1765, w_288_1767, w_288_1770, w_288_1776, w_288_1790, w_288_1791, w_288_1792, w_288_1800, w_288_1843, w_288_1844, w_288_1847, w_288_1859, w_288_1865, w_288_1868, w_288_1873, w_288_1876, w_288_1902, w_288_1906, w_288_1910, w_288_1914, w_288_1921, w_288_1931, w_288_1935, w_288_1939, w_288_1940, w_288_1944, w_288_1949, w_288_1966, w_288_1969, w_288_1980, w_288_2007, w_288_2011, w_288_2012, w_288_2037, w_288_2038, w_288_2041, w_288_2048, w_288_2057, w_288_2062, w_288_2076, w_288_2096, w_288_2097, w_288_2106, w_288_2131, w_288_2149, w_288_2154, w_288_2163, w_288_2250, w_288_2254, w_288_2262, w_288_2273, w_288_2289, w_288_2311, w_288_2319, w_288_2326, w_288_2340, w_288_2358, w_288_2374, w_288_2397, w_288_2408, w_288_2441, w_288_2446, w_288_2447, w_288_2448, w_288_2460, w_288_2467, w_288_2470, w_288_2482, w_288_2503, w_288_2506, w_288_2528, w_288_2556, w_288_2557, w_288_2561, w_288_2565, w_288_2575, w_288_2578, w_288_2582, w_288_2584, w_288_2589, w_288_2612, w_288_2633, w_288_2641, w_288_2642, w_288_2652, w_288_2685, w_288_2696, w_288_2704, w_288_2717, w_288_2739, w_288_2751, w_288_2758, w_288_2774, w_288_2777, w_288_2781, w_288_2785, w_288_2789, w_288_2814, w_288_2818, w_288_2831, w_288_2846, w_288_2852, w_288_2909, w_288_2911, w_288_2931, w_288_2947, w_288_2950, w_288_2965, w_288_2983, w_288_3005, w_288_3007, w_288_3008, w_288_3014, w_288_3038, w_288_3049;
  wire w_289_000, w_289_009, w_289_013, w_289_028, w_289_029, w_289_047, w_289_050, w_289_060, w_289_061, w_289_068, w_289_083, w_289_091, w_289_099, w_289_105, w_289_106, w_289_107, w_289_108, w_289_112, w_289_120, w_289_124, w_289_129, w_289_140, w_289_143, w_289_154, w_289_158, w_289_159, w_289_162, w_289_169, w_289_176, w_289_181, w_289_183, w_289_205, w_289_206, w_289_207, w_289_212, w_289_216, w_289_229, w_289_230, w_289_235, w_289_237, w_289_244, w_289_246, w_289_249, w_289_281, w_289_285, w_289_287, w_289_290, w_289_301, w_289_329, w_289_331, w_289_339, w_289_340, w_289_343, w_289_344, w_289_352, w_289_361, w_289_372, w_289_378, w_289_386, w_289_391, w_289_396, w_289_403, w_289_431, w_289_432, w_289_434, w_289_458, w_289_465, w_289_467, w_289_472, w_289_476, w_289_480, w_289_484, w_289_496, w_289_501, w_289_504, w_289_515, w_289_520, w_289_521, w_289_523, w_289_532, w_289_543, w_289_548, w_289_551, w_289_581, w_289_593, w_289_621, w_289_626, w_289_627, w_289_631, w_289_649, w_289_650, w_289_651, w_289_654, w_289_657, w_289_666, w_289_678, w_289_683, w_289_684, w_289_686, w_289_688, w_289_709, w_289_737, w_289_746, w_289_748, w_289_754, w_289_762, w_289_772, w_289_777, w_289_780, w_289_782, w_289_783, w_289_797, w_289_813, w_289_816, w_289_837, w_289_861, w_289_862, w_289_866, w_289_870, w_289_880, w_289_888, w_289_889, w_289_892, w_289_906, w_289_916, w_289_922, w_289_926, w_289_947, w_289_951, w_289_952, w_289_957, w_289_962, w_289_966, w_289_999, w_289_1000, w_289_1008, w_289_1015, w_289_1020, w_289_1033, w_289_1036, w_289_1038, w_289_1042, w_289_1053, w_289_1059, w_289_1072, w_289_1079, w_289_1084, w_289_1089, w_289_1097, w_289_1103, w_289_1108, w_289_1109, w_289_1110, w_289_1114, w_289_1120, w_289_1121, w_289_1123, w_289_1124, w_289_1126, w_289_1127, w_289_1148, w_289_1150, w_289_1153, w_289_1156, w_289_1160, w_289_1167, w_289_1168, w_289_1173, w_289_1184, w_289_1207, w_289_1220, w_289_1226, w_289_1232, w_289_1243, w_289_1250, w_289_1251, w_289_1255, w_289_1257, w_289_1261, w_289_1267, w_289_1278, w_289_1281, w_289_1292, w_289_1296, w_289_1306, w_289_1308, w_289_1310, w_289_1311, w_289_1328, w_289_1346, w_289_1349, w_289_1354, w_289_1356, w_289_1357, w_289_1359, w_289_1361, w_289_1383, w_289_1384, w_289_1386, w_289_1393, w_289_1425, w_289_1427, w_289_1435, w_289_1455, w_289_1461, w_289_1464, w_289_1466, w_289_1468, w_289_1492, w_289_1495, w_289_1504, w_289_1505, w_289_1506, w_289_1514, w_289_1515, w_289_1516, w_289_1522, w_289_1533, w_289_1537, w_289_1540, w_289_1546, w_289_1555, w_289_1562, w_289_1568, w_289_1572, w_289_1575, w_289_1579, w_289_1605, w_289_1606, w_289_1609, w_289_1612, w_289_1624, w_289_1630, w_289_1631, w_289_1641, w_289_1658, w_289_1661, w_289_1668, w_289_1672, w_289_1673, w_289_1674, w_289_1676, w_289_1681, w_289_1697, w_289_1700, w_289_1702, w_289_1708, w_289_1713, w_289_1714, w_289_1716, w_289_1730, w_289_1740, w_289_1747, w_289_1767, w_289_1773, w_289_1787, w_289_1789, w_289_1800, w_289_1802, w_289_1822, w_289_1829, w_289_1830, w_289_1856, w_289_1858, w_289_1890, w_289_1892, w_289_1897, w_289_1915, w_289_1917, w_289_1924, w_289_1940, w_289_1941, w_289_1945, w_289_1947, w_289_1953, w_289_1961, w_289_1962, w_289_1965, w_289_1975, w_289_1977, w_289_1991, w_289_1996, w_289_2007, w_289_2009, w_289_2010, w_289_2020, w_289_2023, w_289_2036, w_289_2039, w_289_2053, w_289_2059, w_289_2065, w_289_2066, w_289_2073, w_289_2076, w_289_2077, w_289_2081, w_289_2083, w_289_2097, w_289_2113, w_289_2122, w_289_2125, w_289_2130, w_289_2134, w_289_2136, w_289_2143, w_289_2146, w_289_2152, w_289_2153, w_289_2165, w_289_2170, w_289_2171, w_289_2173, w_289_2176, w_289_2190, w_289_2191, w_289_2195, w_289_2197, w_289_2198, w_289_2206, w_289_2216, w_289_2225, w_289_2228, w_289_2229, w_289_2233, w_289_2234, w_289_2237, w_289_2255, w_289_2264, w_289_2266, w_289_2270, w_289_2284, w_289_2292, w_289_2298, w_289_2303, w_289_2311, w_289_2318, w_289_2322, w_289_2323, w_289_2324, w_289_2347, w_289_2354, w_289_2359, w_289_2366, w_289_2379, w_289_2381, w_289_2382, w_289_2383, w_289_2385, w_289_2386, w_289_2391, w_289_2401, w_289_2402, w_289_2408, w_289_2409, w_289_2416, w_289_2420, w_289_2435, w_289_2437, w_289_2462, w_289_2474, w_289_2490, w_289_2494, w_289_2511, w_289_2515, w_289_2527, w_289_2531, w_289_2535, w_289_2538, w_289_2557, w_289_2577, w_289_2591, w_289_2592, w_289_2593, w_289_2594, w_289_2595, w_289_2596, w_289_2597, w_289_2599, w_289_2601, w_289_2602, w_289_2603, w_289_2604, w_289_2605, w_289_2607;
  wire w_290_000, w_290_001, w_290_006, w_290_012, w_290_041, w_290_050, w_290_059, w_290_087, w_290_090, w_290_095, w_290_118, w_290_132, w_290_135, w_290_141, w_290_154, w_290_158, w_290_162, w_290_168, w_290_232, w_290_234, w_290_240, w_290_250, w_290_260, w_290_270, w_290_276, w_290_288, w_290_293, w_290_294, w_290_295, w_290_313, w_290_315, w_290_316, w_290_317, w_290_321, w_290_329, w_290_333, w_290_337, w_290_346, w_290_350, w_290_356, w_290_363, w_290_367, w_290_370, w_290_384, w_290_395, w_290_398, w_290_399, w_290_402, w_290_404, w_290_409, w_290_412, w_290_425, w_290_427, w_290_428, w_290_432, w_290_434, w_290_440, w_290_448, w_290_454, w_290_456, w_290_462, w_290_470, w_290_485, w_290_487, w_290_489, w_290_490, w_290_502, w_290_507, w_290_523, w_290_526, w_290_542, w_290_549, w_290_550, w_290_558, w_290_563, w_290_567, w_290_572, w_290_578, w_290_581, w_290_587, w_290_592, w_290_596, w_290_609, w_290_613, w_290_614, w_290_615, w_290_616, w_290_623, w_290_625, w_290_629, w_290_630, w_290_633, w_290_638, w_290_649, w_290_652, w_290_669, w_290_676, w_290_678, w_290_688, w_290_693, w_290_700, w_290_702, w_290_703, w_290_710, w_290_711, w_290_731, w_290_739, w_290_744, w_290_755, w_290_761, w_290_777, w_290_792, w_290_794, w_290_796, w_290_809, w_290_814, w_290_817, w_290_820, w_290_843, w_290_847, w_290_855, w_290_870, w_290_873, w_290_875, w_290_877, w_290_880, w_290_892, w_290_901, w_290_903, w_290_907, w_290_909, w_290_914, w_290_924, w_290_926, w_290_927, w_290_945, w_290_957, w_290_959, w_290_961, w_290_967, w_290_971, w_290_984, w_290_1003, w_290_1007, w_290_1012, w_290_1017, w_290_1031, w_290_1043, w_290_1047, w_290_1049, w_290_1051, w_290_1053, w_290_1054, w_290_1055, w_290_1058, w_290_1063, w_290_1071, w_290_1075, w_290_1083, w_290_1088, w_290_1089, w_290_1093, w_290_1096, w_290_1102, w_290_1106, w_290_1109, w_290_1110, w_290_1130, w_290_1131, w_290_1141, w_290_1142, w_290_1147, w_290_1159, w_290_1161, w_290_1163, w_290_1180, w_290_1181, w_290_1182, w_290_1191, w_290_1198, w_290_1202, w_290_1212, w_290_1225, w_290_1233, w_290_1242, w_290_1248, w_290_1255, w_290_1261, w_290_1273, w_290_1286, w_290_1291, w_290_1298, w_290_1301, w_290_1308, w_290_1315, w_290_1323, w_290_1329, w_290_1331, w_290_1339, w_290_1344, w_290_1347, w_290_1353, w_290_1355, w_290_1359, w_290_1365, w_290_1368, w_290_1376, w_290_1380, w_290_1386, w_290_1387, w_290_1394, w_290_1410, w_290_1412, w_290_1425, w_290_1428, w_290_1436, w_290_1448, w_290_1456, w_290_1471, w_290_1473, w_290_1484, w_290_1486, w_290_1489, w_290_1491, w_290_1492, w_290_1500, w_290_1508, w_290_1527, w_290_1533, w_290_1538, w_290_1539, w_290_1544, w_290_1551, w_290_1556, w_290_1559, w_290_1568, w_290_1570, w_290_1575, w_290_1579, w_290_1585, w_290_1596, w_290_1620, w_290_1625, w_290_1627, w_290_1631, w_290_1636, w_290_1637, w_290_1638, w_290_1642, w_290_1644, w_290_1654, w_290_1668, w_290_1673, w_290_1682, w_290_1688, w_290_1690, w_290_1693, w_290_1713, w_290_1716, w_290_1717, w_290_1721, w_290_1723, w_290_1736, w_290_1737, w_290_1739, w_290_1766, w_290_1777, w_290_1782, w_290_1783, w_290_1792, w_290_1808, w_290_1824, w_290_1826, w_290_1830, w_290_1831, w_290_1845, w_290_1847, w_290_1852, w_290_1859, w_290_1861, w_290_1875, w_290_1885, w_290_1888, w_290_1896, w_290_1901, w_290_1902, w_290_1909, w_290_1915, w_290_1921, w_290_1935, w_290_1943, w_290_1947, w_290_1950, w_290_1958, w_290_1967, w_290_1968, w_290_1969, w_290_1972, w_290_1973, w_290_1982, w_290_1983, w_290_1987, w_290_1990, w_290_1996, w_290_1998, w_290_2000, w_290_2010, w_290_2022, w_290_2025, w_290_2028, w_290_2029, w_290_2030, w_290_2034, w_290_2041, w_290_2043, w_290_2046, w_290_2059, w_290_2061, w_290_2086, w_290_2089, w_290_2095, w_290_2097, w_290_2104, w_290_2110, w_290_2119, w_290_2126, w_290_2128, w_290_2132, w_290_2161, w_290_2171, w_290_2202, w_290_2216, w_290_2222, w_290_2236, w_290_2253, w_290_2257, w_290_2274, w_290_2277, w_290_2324, w_290_2331, w_290_2372, w_290_2392, w_290_2398, w_290_2400, w_290_2401, w_290_2409, w_290_2425, w_290_2455, w_290_2458, w_290_2468, w_290_2482, w_290_2491, w_290_2492, w_290_2495, w_290_2505, w_290_2506, w_290_2509, w_290_2529, w_290_2535, w_290_2542, w_290_2544, w_290_2552, w_290_2557, w_290_2562, w_290_2576, w_290_2583, w_290_2587, w_290_2595, w_290_2631, w_290_2645, w_290_2646, w_290_2647, w_290_2651, w_290_2659, w_290_2667, w_290_2673, w_290_2715, w_290_2725, w_290_2739, w_290_2742, w_290_2744, w_290_2752, w_290_2757, w_290_2766, w_290_2768, w_290_2771, w_290_2775, w_290_2790, w_290_2795, w_290_2812;
  wire w_291_002, w_291_005, w_291_006, w_291_008, w_291_012, w_291_019, w_291_022, w_291_023, w_291_024, w_291_026, w_291_031, w_291_038, w_291_040, w_291_041, w_291_045, w_291_053, w_291_055, w_291_056, w_291_057, w_291_060, w_291_065, w_291_069, w_291_072, w_291_075, w_291_079, w_291_080, w_291_087, w_291_091, w_291_096, w_291_097, w_291_102, w_291_109, w_291_110, w_291_112, w_291_117, w_291_123, w_291_127, w_291_128, w_291_130, w_291_131, w_291_133, w_291_134, w_291_135, w_291_136, w_291_138, w_291_140, w_291_153, w_291_154, w_291_161, w_291_163, w_291_169, w_291_170, w_291_171, w_291_174, w_291_178, w_291_180, w_291_181, w_291_182, w_291_183, w_291_184, w_291_189, w_291_191, w_291_193, w_291_195, w_291_197, w_291_201, w_291_202, w_291_205, w_291_206, w_291_207, w_291_212, w_291_213, w_291_215, w_291_217, w_291_218, w_291_223, w_291_229, w_291_234, w_291_236, w_291_237, w_291_240, w_291_245, w_291_246, w_291_247, w_291_249, w_291_252, w_291_253, w_291_254, w_291_257, w_291_260, w_291_267, w_291_268, w_291_269, w_291_271, w_291_272, w_291_277, w_291_282, w_291_291, w_291_292, w_291_293, w_291_295, w_291_299, w_291_300, w_291_303, w_291_308, w_291_309, w_291_312, w_291_313, w_291_320, w_291_321, w_291_329, w_291_331, w_291_332, w_291_334, w_291_336, w_291_339, w_291_341, w_291_349, w_291_351, w_291_357, w_291_361, w_291_365, w_291_366, w_291_367, w_291_368, w_291_370, w_291_372, w_291_376, w_291_380, w_291_382, w_291_385, w_291_390, w_291_392, w_291_402, w_291_409, w_291_410, w_291_411, w_291_416, w_291_424, w_291_431, w_291_433, w_291_434, w_291_435, w_291_436, w_291_442, w_291_448, w_291_452, w_291_462, w_291_468, w_291_469, w_291_470, w_291_472, w_291_474, w_291_482, w_291_483, w_291_484, w_291_485, w_291_489, w_291_491, w_291_495, w_291_501, w_291_503, w_291_509, w_291_512, w_291_519, w_291_520, w_291_521, w_291_522, w_291_526, w_291_527, w_291_530, w_291_532, w_291_535, w_291_538, w_291_541, w_291_544, w_291_547, w_291_548, w_291_549, w_291_550, w_291_552, w_291_554, w_291_555, w_291_558, w_291_563, w_291_565, w_291_566, w_291_567, w_291_573, w_291_583, w_291_585, w_291_586, w_291_587, w_291_589, w_291_596, w_291_597, w_291_598, w_291_599, w_291_600, w_291_603, w_291_605, w_291_608, w_291_609, w_291_614, w_291_619, w_291_622, w_291_624, w_291_625, w_291_630, w_291_631, w_291_635, w_291_637, w_291_639, w_291_646, w_291_649, w_291_651, w_291_652, w_291_657, w_291_658, w_291_659, w_291_661, w_291_662, w_291_664, w_291_665, w_291_668, w_291_669, w_291_673, w_291_675, w_291_678, w_291_679, w_291_680, w_291_681, w_291_683, w_291_687, w_291_692, w_291_693, w_291_701, w_291_707, w_291_709, w_291_719, w_291_721, w_291_729, w_291_737, w_291_744, w_291_745, w_291_753, w_291_754, w_291_757, w_291_758, w_291_761, w_291_765, w_291_768, w_291_770, w_291_771, w_291_772, w_291_774, w_291_783, w_291_792, w_291_794, w_291_795, w_291_800, w_291_801, w_291_803, w_291_804, w_291_805, w_291_809, w_291_815, w_291_819, w_291_820, w_291_823, w_291_825, w_291_826, w_291_827, w_291_829, w_291_830, w_291_832, w_291_834, w_291_835, w_291_841, w_291_842, w_291_843, w_291_845, w_291_846, w_291_847, w_291_850, w_291_851, w_291_852, w_291_855, w_291_857, w_291_862, w_291_863, w_291_866, w_291_871, w_291_872, w_291_877, w_291_880, w_291_883, w_291_887, w_291_894, w_291_908, w_291_913, w_291_922, w_291_932, w_291_933, w_291_940, w_291_944, w_291_948, w_291_957, w_291_958, w_291_962, w_291_964, w_291_965, w_291_972, w_291_979, w_291_985, w_291_997, w_291_1000, w_291_1002, w_291_1007, w_291_1008, w_291_1011, w_291_1012, w_291_1022, w_291_1029, w_291_1030, w_291_1031, w_291_1035, w_291_1036, w_291_1037, w_291_1038, w_291_1039, w_291_1040, w_291_1041, w_291_1042, w_291_1044;
  wire w_292_013, w_292_021, w_292_023, w_292_026, w_292_027, w_292_031, w_292_057, w_292_064, w_292_066, w_292_068, w_292_074, w_292_076, w_292_078, w_292_083, w_292_085, w_292_089, w_292_090, w_292_102, w_292_118, w_292_149, w_292_167, w_292_168, w_292_187, w_292_188, w_292_232, w_292_237, w_292_269, w_292_278, w_292_301, w_292_305, w_292_306, w_292_308, w_292_309, w_292_320, w_292_363, w_292_392, w_292_411, w_292_420, w_292_473, w_292_476, w_292_477, w_292_490, w_292_493, w_292_502, w_292_505, w_292_560, w_292_586, w_292_596, w_292_598, w_292_603, w_292_604, w_292_620, w_292_663, w_292_678, w_292_683, w_292_700, w_292_720, w_292_751, w_292_779, w_292_790, w_292_798, w_292_821, w_292_825, w_292_832, w_292_878, w_292_922, w_292_924, w_292_939, w_292_944, w_292_969, w_292_977, w_292_983, w_292_994, w_292_1006, w_292_1062, w_292_1100, w_292_1105, w_292_1109, w_292_1113, w_292_1127, w_292_1151, w_292_1158, w_292_1177, w_292_1189, w_292_1201, w_292_1207, w_292_1220, w_292_1223, w_292_1224, w_292_1230, w_292_1239, w_292_1245, w_292_1249, w_292_1261, w_292_1262, w_292_1279, w_292_1316, w_292_1317, w_292_1366, w_292_1367, w_292_1372, w_292_1385, w_292_1401, w_292_1404, w_292_1406, w_292_1411, w_292_1428, w_292_1436, w_292_1462, w_292_1488, w_292_1529, w_292_1539, w_292_1544, w_292_1546, w_292_1592, w_292_1597, w_292_1602, w_292_1605, w_292_1615, w_292_1621, w_292_1625, w_292_1635, w_292_1651, w_292_1652, w_292_1668, w_292_1681, w_292_1698, w_292_1701, w_292_1703, w_292_1704, w_292_1713, w_292_1725, w_292_1726, w_292_1736, w_292_1756, w_292_1763, w_292_1785, w_292_1789, w_292_1825, w_292_1832, w_292_1861, w_292_1862, w_292_1866, w_292_1867, w_292_1877, w_292_1900, w_292_1915, w_292_1923, w_292_1929, w_292_1932, w_292_1938, w_292_1940, w_292_1942, w_292_1960, w_292_1986, w_292_2002, w_292_2007, w_292_2016, w_292_2077, w_292_2090, w_292_2108, w_292_2114, w_292_2146, w_292_2150, w_292_2185, w_292_2194, w_292_2214, w_292_2229, w_292_2255, w_292_2289, w_292_2291, w_292_2295, w_292_2297, w_292_2301, w_292_2304, w_292_2316, w_292_2368, w_292_2404, w_292_2410, w_292_2433, w_292_2453, w_292_2464, w_292_2471, w_292_2483, w_292_2485, w_292_2500, w_292_2515, w_292_2534, w_292_2541, w_292_2548, w_292_2552, w_292_2588, w_292_2609, w_292_2618, w_292_2629, w_292_2632, w_292_2650, w_292_2654, w_292_2655, w_292_2689, w_292_2690, w_292_2696, w_292_2708, w_292_2735, w_292_2756, w_292_2778, w_292_2783, w_292_2797, w_292_2803, w_292_2808, w_292_2810, w_292_2812, w_292_2840, w_292_2846, w_292_2851, w_292_2876, w_292_2940, w_292_2954, w_292_2962, w_292_2966, w_292_2969, w_292_2975, w_292_2978, w_292_3024, w_292_3032, w_292_3035, w_292_3048, w_292_3070, w_292_3074, w_292_3100, w_292_3101, w_292_3126, w_292_3158, w_292_3181, w_292_3199, w_292_3204, w_292_3206, w_292_3211, w_292_3213, w_292_3217, w_292_3238, w_292_3258, w_292_3278, w_292_3305, w_292_3307, w_292_3313, w_292_3322, w_292_3329, w_292_3332, w_292_3357, w_292_3363, w_292_3370, w_292_3375, w_292_3388, w_292_3401, w_292_3402, w_292_3409, w_292_3412, w_292_3417, w_292_3440, w_292_3455, w_292_3472, w_292_3494, w_292_3551, w_292_3564, w_292_3573, w_292_3575, w_292_3588, w_292_3615, w_292_3628, w_292_3667, w_292_3672, w_292_3674, w_292_3680, w_292_3696, w_292_3732, w_292_3744, w_292_3766, w_292_3772, w_292_3784, w_292_3804, w_292_3846, w_292_3847, w_292_3853, w_292_3859, w_292_3861, w_292_3866, w_292_3871, w_292_3875, w_292_3889, w_292_3892, w_292_3908, w_292_3916, w_292_3917, w_292_3926, w_292_4003, w_292_4005, w_292_4039, w_292_4050, w_292_4055, w_292_4072, w_292_4077, w_292_4082, w_292_4083, w_292_4092, w_292_4100, w_292_4103, w_292_4113, w_292_4128, w_292_4145, w_292_4151, w_292_4155, w_292_4173, w_292_4177, w_292_4180, w_292_4193, w_292_4222, w_292_4228, w_292_4234, w_292_4235, w_292_4248, w_292_4261, w_292_4266, w_292_4280, w_292_4284, w_292_4285, w_292_4298, w_292_4310, w_292_4319, w_292_4328, w_292_4329, w_292_4335, w_292_4338, w_292_4350, w_292_4351, w_292_4355, w_292_4357, w_292_4367, w_292_4371, w_292_4378, w_292_4399, w_292_4414, w_292_4419, w_292_4422, w_292_4423, w_292_4424, w_292_4457, w_292_4469, w_292_4484, w_292_4486, w_292_4492, w_292_4503, w_292_4543, w_292_4592, w_292_4611, w_292_4620, w_292_4634, w_292_4654, w_292_4659, w_292_4670, w_292_4699, w_292_4710, w_292_4711, w_292_4726, w_292_4735, w_292_4738, w_292_4747, w_292_4761, w_292_4771, w_292_4782, w_292_4803, w_292_4807, w_292_4819, w_292_4825, w_292_4828, w_292_4830, w_292_4837, w_292_4844, w_292_4861, w_292_4887, w_292_4892;
  wire w_293_001, w_293_002, w_293_010, w_293_018, w_293_022, w_293_026, w_293_033, w_293_036, w_293_041, w_293_046, w_293_049, w_293_051, w_293_053, w_293_057, w_293_059, w_293_061, w_293_065, w_293_068, w_293_075, w_293_081, w_293_083, w_293_085, w_293_091, w_293_097, w_293_100, w_293_104, w_293_105, w_293_107, w_293_111, w_293_112, w_293_115, w_293_124, w_293_128, w_293_133, w_293_134, w_293_136, w_293_139, w_293_141, w_293_143, w_293_146, w_293_148, w_293_151, w_293_154, w_293_157, w_293_158, w_293_159, w_293_168, w_293_170, w_293_186, w_293_187, w_293_201, w_293_207, w_293_208, w_293_217, w_293_234, w_293_235, w_293_236, w_293_241, w_293_243, w_293_250, w_293_256, w_293_257, w_293_265, w_293_269, w_293_281, w_293_282, w_293_285, w_293_286, w_293_299, w_293_301, w_293_302, w_293_307, w_293_313, w_293_315, w_293_317, w_293_318, w_293_322, w_293_325, w_293_326, w_293_330, w_293_331, w_293_334, w_293_335, w_293_336, w_293_337, w_293_338, w_293_348, w_293_357, w_293_358, w_293_361, w_293_365, w_293_366, w_293_367, w_293_373, w_293_376, w_293_391, w_293_392, w_293_393, w_293_399, w_293_402, w_293_407, w_293_410, w_293_413, w_293_414, w_293_415, w_293_416, w_293_418, w_293_419, w_293_425, w_293_428, w_293_431, w_293_436, w_293_438, w_293_439, w_293_442, w_293_443, w_293_449, w_293_451, w_293_453, w_293_454, w_293_457, w_293_462, w_293_463, w_293_464, w_293_468, w_293_472, w_293_477, w_293_479, w_293_480, w_293_484, w_293_485, w_293_491, w_293_492, w_293_495, w_293_504, w_293_508, w_293_509, w_293_512, w_293_518, w_293_520, w_293_530, w_293_533, w_293_536, w_293_537, w_293_539, w_293_550, w_293_553, w_293_555, w_293_561, w_293_563, w_293_569, w_293_571, w_293_572, w_293_576, w_293_578, w_293_584, w_293_586, w_293_588, w_293_590, w_293_604, w_293_613, w_293_623, w_293_626, w_293_628, w_293_640, w_293_642, w_293_644, w_293_649, w_293_660, w_293_665, w_293_675, w_293_676, w_293_678, w_293_680, w_293_685, w_293_687, w_293_689, w_293_690, w_293_691, w_293_696, w_293_703, w_293_709, w_293_712, w_293_715, w_293_717, w_293_720, w_293_722, w_293_727, w_293_729, w_293_735, w_293_736, w_293_746, w_293_749, w_293_750, w_293_757, w_293_767, w_293_777, w_293_778, w_293_780, w_293_784, w_293_789, w_293_791, w_293_797, w_293_801, w_293_802, w_293_807, w_293_808, w_293_810, w_293_812, w_293_814, w_293_822, w_293_828, w_293_831, w_293_835, w_293_839, w_293_840, w_293_850, w_293_852, w_293_854, w_293_858, w_293_859, w_293_865, w_293_867, w_293_871, w_293_872, w_293_873, w_293_875, w_293_876, w_293_883, w_293_885, w_293_888, w_293_892, w_293_896, w_293_897, w_293_900, w_293_918, w_293_923, w_293_937, w_293_944, w_293_947, w_293_962, w_293_973, w_293_975, w_293_978, w_293_992, w_293_1005, w_293_1008, w_293_1009, w_293_1014, w_293_1019, w_293_1021, w_293_1022, w_293_1026, w_293_1028, w_293_1031, w_293_1034, w_293_1035, w_293_1041, w_293_1059, w_293_1063, w_293_1064, w_293_1069, w_293_1070, w_293_1078, w_293_1083, w_293_1086, w_293_1087, w_293_1089, w_293_1099, w_293_1108, w_293_1114, w_293_1126, w_293_1131, w_293_1132, w_293_1134, w_293_1136, w_293_1137, w_293_1139, w_293_1157, w_293_1161, w_293_1175, w_293_1186, w_293_1197, w_293_1207, w_293_1215, w_293_1227, w_293_1229, w_293_1232, w_293_1233, w_293_1234, w_293_1237, w_293_1239, w_293_1240, w_293_1244, w_293_1245, w_293_1251, w_293_1258, w_293_1271, w_293_1275, w_293_1279, w_293_1281, w_293_1297, w_293_1299, w_293_1302, w_293_1303, w_293_1305, w_293_1309, w_293_1311, w_293_1315, w_293_1321, w_293_1325, w_293_1335, w_293_1341, w_293_1344, w_293_1356, w_293_1357, w_293_1360, w_293_1368, w_293_1369, w_293_1370, w_293_1372;
  wire w_294_000, w_294_006, w_294_010, w_294_012, w_294_018, w_294_019, w_294_045, w_294_048, w_294_050, w_294_063, w_294_071, w_294_104, w_294_108, w_294_110, w_294_126, w_294_134, w_294_139, w_294_156, w_294_171, w_294_180, w_294_215, w_294_217, w_294_220, w_294_222, w_294_223, w_294_225, w_294_236, w_294_240, w_294_248, w_294_258, w_294_279, w_294_290, w_294_294, w_294_300, w_294_309, w_294_316, w_294_319, w_294_323, w_294_324, w_294_334, w_294_339, w_294_352, w_294_353, w_294_361, w_294_364, w_294_365, w_294_375, w_294_381, w_294_387, w_294_388, w_294_392, w_294_398, w_294_403, w_294_423, w_294_443, w_294_447, w_294_454, w_294_468, w_294_478, w_294_492, w_294_502, w_294_506, w_294_513, w_294_522, w_294_527, w_294_533, w_294_563, w_294_576, w_294_582, w_294_586, w_294_589, w_294_590, w_294_595, w_294_601, w_294_615, w_294_617, w_294_623, w_294_630, w_294_635, w_294_649, w_294_655, w_294_660, w_294_662, w_294_669, w_294_681, w_294_692, w_294_694, w_294_699, w_294_701, w_294_712, w_294_721, w_294_729, w_294_738, w_294_739, w_294_740, w_294_742, w_294_750, w_294_756, w_294_770, w_294_779, w_294_788, w_294_798, w_294_803, w_294_846, w_294_847, w_294_853, w_294_856, w_294_858, w_294_874, w_294_901, w_294_902, w_294_916, w_294_919, w_294_931, w_294_942, w_294_947, w_294_950, w_294_955, w_294_957, w_294_965, w_294_971, w_294_972, w_294_977, w_294_982, w_294_991, w_294_996, w_294_1020, w_294_1035, w_294_1036, w_294_1038, w_294_1071, w_294_1072, w_294_1077, w_294_1083, w_294_1099, w_294_1100, w_294_1104, w_294_1106, w_294_1129, w_294_1132, w_294_1134, w_294_1135, w_294_1138, w_294_1155, w_294_1179, w_294_1184, w_294_1194, w_294_1200, w_294_1209, w_294_1223, w_294_1229, w_294_1241, w_294_1244, w_294_1259, w_294_1275, w_294_1292, w_294_1303, w_294_1326, w_294_1342, w_294_1365, w_294_1396, w_294_1402, w_294_1424, w_294_1439, w_294_1454, w_294_1467, w_294_1469, w_294_1495, w_294_1499, w_294_1506, w_294_1562, w_294_1573, w_294_1580, w_294_1589, w_294_1594, w_294_1603, w_294_1609, w_294_1619, w_294_1654, w_294_1658, w_294_1668, w_294_1673, w_294_1676, w_294_1696, w_294_1738, w_294_1747, w_294_1800, w_294_1834, w_294_1841, w_294_1856, w_294_1858, w_294_1863, w_294_1873, w_294_1892, w_294_1900, w_294_1909, w_294_1935, w_294_1945, w_294_1955, w_294_1960, w_294_1996, w_294_2011, w_294_2029, w_294_2038, w_294_2057, w_294_2061, w_294_2068, w_294_2096, w_294_2105, w_294_2112, w_294_2122, w_294_2126, w_294_2131, w_294_2140, w_294_2141, w_294_2151, w_294_2160, w_294_2193, w_294_2204, w_294_2266, w_294_2285, w_294_2287, w_294_2297, w_294_2334, w_294_2336, w_294_2341, w_294_2350, w_294_2357, w_294_2362, w_294_2417, w_294_2421, w_294_2445, w_294_2448, w_294_2493, w_294_2506, w_294_2511, w_294_2526, w_294_2539, w_294_2542, w_294_2545, w_294_2548, w_294_2562, w_294_2563, w_294_2595, w_294_2600, w_294_2631, w_294_2647, w_294_2675, w_294_2709, w_294_2721, w_294_2723, w_294_2729, w_294_2753, w_294_2756, w_294_2759, w_294_2764, w_294_2791, w_294_2793, w_294_2796, w_294_2803, w_294_2804, w_294_2832, w_294_2837, w_294_2845, w_294_2874, w_294_2880, w_294_2897, w_294_2917, w_294_2946, w_294_2964, w_294_2969, w_294_2972, w_294_3019, w_294_3035, w_294_3048, w_294_3075, w_294_3079, w_294_3111, w_294_3121, w_294_3131, w_294_3135, w_294_3141, w_294_3160, w_294_3164, w_294_3168, w_294_3171, w_294_3190, w_294_3211, w_294_3247, w_294_3259, w_294_3270, w_294_3293, w_294_3294, w_294_3300, w_294_3311, w_294_3322, w_294_3337, w_294_3348, w_294_3363, w_294_3380, w_294_3381, w_294_3386, w_294_3392, w_294_3397, w_294_3399, w_294_3416, w_294_3422, w_294_3428, w_294_3444, w_294_3447, w_294_3454, w_294_3461, w_294_3476, w_294_3537, w_294_3543, w_294_3553, w_294_3561, w_294_3596, w_294_3601, w_294_3608, w_294_3616, w_294_3707, w_294_3714, w_294_3725, w_294_3731, w_294_3737, w_294_3766, w_294_3777, w_294_3778, w_294_3780, w_294_3795, w_294_3806, w_294_3809, w_294_3810, w_294_3812, w_294_3819, w_294_3845, w_294_3875, w_294_3882, w_294_3889, w_294_3894, w_294_3896, w_294_3897, w_294_3916, w_294_3924, w_294_3961, w_294_3982, w_294_3996, w_294_3998, w_294_4024, w_294_4025, w_294_4028, w_294_4033, w_294_4043, w_294_4058, w_294_4061, w_294_4062, w_294_4063, w_294_4064;
  wire w_295_000, w_295_009, w_295_010, w_295_011, w_295_012, w_295_014, w_295_017, w_295_022, w_295_025, w_295_029, w_295_034, w_295_039, w_295_043, w_295_044, w_295_045, w_295_047, w_295_050, w_295_051, w_295_053, w_295_059, w_295_060, w_295_062, w_295_063, w_295_065, w_295_068, w_295_070, w_295_071, w_295_073, w_295_074, w_295_075, w_295_076, w_295_078, w_295_080, w_295_084, w_295_089, w_295_090, w_295_091, w_295_093, w_295_094, w_295_097, w_295_100, w_295_102, w_295_112, w_295_114, w_295_117, w_295_118, w_295_120, w_295_121, w_295_125, w_295_127, w_295_131, w_295_136, w_295_137, w_295_138, w_295_140, w_295_144, w_295_147, w_295_148, w_295_149, w_295_158, w_295_160, w_295_162, w_295_165, w_295_176, w_295_178, w_295_182, w_295_187, w_295_192, w_295_199, w_295_201, w_295_202, w_295_203, w_295_205, w_295_226, w_295_228, w_295_230, w_295_231, w_295_234, w_295_236, w_295_240, w_295_243, w_295_246, w_295_248, w_295_249, w_295_251, w_295_257, w_295_263, w_295_266, w_295_268, w_295_272, w_295_273, w_295_276, w_295_278, w_295_280, w_295_281, w_295_284, w_295_285, w_295_292, w_295_300, w_295_301, w_295_307, w_295_310, w_295_311, w_295_312, w_295_314, w_295_315, w_295_320, w_295_324, w_295_347, w_295_348, w_295_349, w_295_352, w_295_353, w_295_354, w_295_356, w_295_357, w_295_359, w_295_365, w_295_366, w_295_368, w_295_371, w_295_375, w_295_379, w_295_381, w_295_384, w_295_385, w_295_386, w_295_389, w_295_390, w_295_395, w_295_397, w_295_403, w_295_406, w_295_407, w_295_417, w_295_418, w_295_421, w_295_422, w_295_425, w_295_426, w_295_433, w_295_435, w_295_437, w_295_445, w_295_447, w_295_454, w_295_455, w_295_457, w_295_459, w_295_462, w_295_465, w_295_466, w_295_472, w_295_480, w_295_482, w_295_483, w_295_493, w_295_494, w_295_505, w_295_508, w_295_509, w_295_512, w_295_514, w_295_518, w_295_520, w_295_521, w_295_525, w_295_526, w_295_533, w_295_534, w_295_535, w_295_539, w_295_540, w_295_548, w_295_551, w_295_552, w_295_554, w_295_555, w_295_557, w_295_558, w_295_559, w_295_562, w_295_567, w_295_574, w_295_583, w_295_584, w_295_591, w_295_594, w_295_595, w_295_598, w_295_602, w_295_603, w_295_604, w_295_606, w_295_608, w_295_610, w_295_611, w_295_613, w_295_618, w_295_619, w_295_620, w_295_621, w_295_625, w_295_627, w_295_628, w_295_629, w_295_634, w_295_636, w_295_640, w_295_648, w_295_650, w_295_651, w_295_652, w_295_654, w_295_655, w_295_658, w_295_661, w_295_663, w_295_666, w_295_672, w_295_673, w_295_674, w_295_675, w_295_677, w_295_681, w_295_682, w_295_691, w_295_692, w_295_695, w_295_696, w_295_698, w_295_701, w_295_702, w_295_705, w_295_707, w_295_709, w_295_710, w_295_711, w_295_712, w_295_714, w_295_716, w_295_726, w_295_727, w_295_732, w_295_734, w_295_736, w_295_739, w_295_740, w_295_741, w_295_749, w_295_753, w_295_754, w_295_764, w_295_765, w_295_766, w_295_768, w_295_771, w_295_772, w_295_773, w_295_775, w_295_778, w_295_779, w_295_781, w_295_783, w_295_784, w_295_786, w_295_790, w_295_791, w_295_792, w_295_793, w_295_794, w_295_796, w_295_800, w_295_802, w_295_803, w_295_806, w_295_807, w_295_811, w_295_814, w_295_820, w_295_823, w_295_827, w_295_835, w_295_838, w_295_840, w_295_845, w_295_846, w_295_849, w_295_856, w_295_857, w_295_858, w_295_871, w_295_876, w_295_882, w_295_893, w_295_894, w_295_898, w_295_899, w_295_904, w_295_908, w_295_910, w_295_913, w_295_914, w_295_916, w_295_919, w_295_921, w_295_929, w_295_937, w_295_951, w_295_954, w_295_956, w_295_965, w_295_970, w_295_973, w_295_979, w_295_989, w_295_992, w_295_996, w_295_997, w_295_1004, w_295_1005, w_295_1008, w_295_1009, w_295_1011, w_295_1015, w_295_1016, w_295_1020, w_295_1021, w_295_1031, w_295_1032, w_295_1033, w_295_1038, w_295_1040, w_295_1041, w_295_1048;
  wire w_296_012, w_296_024, w_296_025, w_296_033, w_296_042, w_296_062, w_296_069, w_296_085, w_296_088, w_296_103, w_296_104, w_296_110, w_296_113, w_296_119, w_296_120, w_296_136, w_296_145, w_296_149, w_296_150, w_296_157, w_296_170, w_296_173, w_296_175, w_296_176, w_296_179, w_296_182, w_296_205, w_296_206, w_296_207, w_296_209, w_296_217, w_296_220, w_296_244, w_296_245, w_296_251, w_296_254, w_296_258, w_296_264, w_296_280, w_296_283, w_296_286, w_296_291, w_296_292, w_296_293, w_296_320, w_296_327, w_296_329, w_296_330, w_296_345, w_296_350, w_296_352, w_296_355, w_296_369, w_296_371, w_296_372, w_296_376, w_296_383, w_296_387, w_296_398, w_296_412, w_296_429, w_296_437, w_296_441, w_296_442, w_296_446, w_296_458, w_296_460, w_296_479, w_296_483, w_296_489, w_296_501, w_296_505, w_296_526, w_296_532, w_296_537, w_296_542, w_296_543, w_296_545, w_296_558, w_296_563, w_296_577, w_296_578, w_296_602, w_296_605, w_296_609, w_296_611, w_296_619, w_296_623, w_296_631, w_296_635, w_296_645, w_296_648, w_296_661, w_296_666, w_296_672, w_296_673, w_296_684, w_296_701, w_296_729, w_296_732, w_296_750, w_296_763, w_296_768, w_296_779, w_296_780, w_296_799, w_296_811, w_296_812, w_296_815, w_296_824, w_296_828, w_296_830, w_296_839, w_296_849, w_296_851, w_296_858, w_296_873, w_296_875, w_296_881, w_296_892, w_296_897, w_296_925, w_296_959, w_296_961, w_296_997, w_296_1002, w_296_1003, w_296_1016, w_296_1023, w_296_1032, w_296_1034, w_296_1044, w_296_1056, w_296_1059, w_296_1060, w_296_1061, w_296_1062, w_296_1068, w_296_1082, w_296_1083, w_296_1087, w_296_1095, w_296_1104, w_296_1110, w_296_1122, w_296_1124, w_296_1146, w_296_1149, w_296_1159, w_296_1185, w_296_1187, w_296_1189, w_296_1199, w_296_1200, w_296_1210, w_296_1227, w_296_1246, w_296_1248, w_296_1256, w_296_1258, w_296_1270, w_296_1272, w_296_1273, w_296_1279, w_296_1285, w_296_1287, w_296_1289, w_296_1294, w_296_1303, w_296_1304, w_296_1307, w_296_1311, w_296_1315, w_296_1321, w_296_1327, w_296_1348, w_296_1349, w_296_1351, w_296_1357, w_296_1360, w_296_1362, w_296_1367, w_296_1375, w_296_1396, w_296_1397, w_296_1401, w_296_1405, w_296_1410, w_296_1414, w_296_1416, w_296_1417, w_296_1420, w_296_1422, w_296_1435, w_296_1439, w_296_1457, w_296_1464, w_296_1467, w_296_1468, w_296_1469, w_296_1476, w_296_1489, w_296_1491, w_296_1492, w_296_1508, w_296_1522, w_296_1532, w_296_1533, w_296_1538, w_296_1544, w_296_1546, w_296_1561, w_296_1565, w_296_1567, w_296_1572, w_296_1576, w_296_1588, w_296_1595, w_296_1597, w_296_1617, w_296_1633, w_296_1647, w_296_1650, w_296_1663, w_296_1673, w_296_1705, w_296_1710, w_296_1714, w_296_1718, w_296_1724, w_296_1729, w_296_1732, w_296_1733, w_296_1735, w_296_1739, w_296_1759, w_296_1769, w_296_1775, w_296_1789, w_296_1790, w_296_1793, w_296_1796, w_296_1800, w_296_1807, w_296_1822, w_296_1823, w_296_1827, w_296_1842, w_296_1848, w_296_1853, w_296_1860, w_296_1867, w_296_1871, w_296_1892, w_296_1894, w_296_1905, w_296_1908, w_296_1918, w_296_1921, w_296_1928, w_296_1931, w_296_1935, w_296_1942, w_296_1950, w_296_1952, w_296_1953, w_296_1960, w_296_1961, w_296_1968, w_296_1969, w_296_1971, w_296_1977, w_296_1982, w_296_1984, w_296_1988, w_296_1994, w_296_2000, w_296_2001, w_296_2004, w_296_2010, w_296_2013, w_296_2018, w_296_2021, w_296_2022, w_296_2033, w_296_2035, w_296_2044, w_296_2046, w_296_2047, w_296_2052, w_296_2055, w_296_2070, w_296_2076, w_296_2077, w_296_2091, w_296_2095, w_296_2104, w_296_2108, w_296_2117, w_296_2127, w_296_2128, w_296_2131, w_296_2139, w_296_2148, w_296_2160, w_296_2162, w_296_2164, w_296_2172, w_296_2180, w_296_2274, w_296_2300, w_296_2305, w_296_2356, w_296_2380, w_296_2403, w_296_2404, w_296_2407, w_296_2413, w_296_2427, w_296_2433, w_296_2438, w_296_2444, w_296_2446, w_296_2447, w_296_2468, w_296_2490, w_296_2519, w_296_2532, w_296_2572, w_296_2580, w_296_2585, w_296_2591, w_296_2593, w_296_2594, w_296_2638, w_296_2657, w_296_2702, w_296_2703, w_296_2708, w_296_2718, w_296_2746, w_296_2827, w_296_2843, w_296_2845;
  wire w_297_002, w_297_004, w_297_010, w_297_011, w_297_012, w_297_014, w_297_016, w_297_020, w_297_024, w_297_031, w_297_037, w_297_043, w_297_048, w_297_055, w_297_057, w_297_059, w_297_072, w_297_076, w_297_081, w_297_082, w_297_083, w_297_087, w_297_088, w_297_089, w_297_093, w_297_099, w_297_104, w_297_105, w_297_110, w_297_114, w_297_116, w_297_123, w_297_127, w_297_138, w_297_141, w_297_144, w_297_149, w_297_150, w_297_157, w_297_160, w_297_163, w_297_166, w_297_176, w_297_177, w_297_184, w_297_185, w_297_189, w_297_193, w_297_199, w_297_203, w_297_213, w_297_221, w_297_224, w_297_230, w_297_236, w_297_239, w_297_242, w_297_248, w_297_251, w_297_253, w_297_257, w_297_258, w_297_259, w_297_261, w_297_269, w_297_277, w_297_279, w_297_289, w_297_293, w_297_297, w_297_307, w_297_330, w_297_336, w_297_342, w_297_345, w_297_354, w_297_360, w_297_363, w_297_367, w_297_369, w_297_377, w_297_383, w_297_389, w_297_392, w_297_398, w_297_401, w_297_416, w_297_419, w_297_421, w_297_433, w_297_439, w_297_440, w_297_442, w_297_445, w_297_450, w_297_458, w_297_462, w_297_464, w_297_470, w_297_477, w_297_483, w_297_490, w_297_493, w_297_496, w_297_507, w_297_511, w_297_520, w_297_524, w_297_534, w_297_536, w_297_540, w_297_543, w_297_545, w_297_553, w_297_560, w_297_566, w_297_580, w_297_585, w_297_586, w_297_588, w_297_600, w_297_603, w_297_614, w_297_617, w_297_618, w_297_619, w_297_626, w_297_633, w_297_638, w_297_640, w_297_641, w_297_646, w_297_647, w_297_649, w_297_661, w_297_662, w_297_665, w_297_668, w_297_670, w_297_674, w_297_677, w_297_681, w_297_685, w_297_688, w_297_689, w_297_691, w_297_710, w_297_711, w_297_712, w_297_715, w_297_726, w_297_728, w_297_731, w_297_732, w_297_734, w_297_737, w_297_743, w_297_744, w_297_763, w_297_766, w_297_774, w_297_777, w_297_785, w_297_808, w_297_821, w_297_829, w_297_838, w_297_841, w_297_842, w_297_854, w_297_856, w_297_860, w_297_861, w_297_864, w_297_867, w_297_869, w_297_870, w_297_873, w_297_874, w_297_881, w_297_891, w_297_893, w_297_904, w_297_907, w_297_920, w_297_929, w_297_941, w_297_942, w_297_946, w_297_947, w_297_962, w_297_970, w_297_977, w_297_999, w_297_1008, w_297_1009, w_297_1016, w_297_1017, w_297_1022, w_297_1036, w_297_1037, w_297_1041, w_297_1044, w_297_1051, w_297_1054, w_297_1055, w_297_1066, w_297_1081, w_297_1087, w_297_1088, w_297_1093, w_297_1095, w_297_1097, w_297_1103, w_297_1113, w_297_1121, w_297_1129, w_297_1131, w_297_1139, w_297_1146, w_297_1157, w_297_1163, w_297_1170, w_297_1172, w_297_1176, w_297_1182, w_297_1186, w_297_1195, w_297_1197, w_297_1208, w_297_1209, w_297_1215, w_297_1217, w_297_1219, w_297_1222, w_297_1225, w_297_1226, w_297_1236, w_297_1237, w_297_1242, w_297_1264, w_297_1274, w_297_1279, w_297_1282, w_297_1284, w_297_1292, w_297_1296, w_297_1301, w_297_1307, w_297_1310, w_297_1329, w_297_1336, w_297_1339, w_297_1347, w_297_1350, w_297_1356, w_297_1363, w_297_1370, w_297_1391, w_297_1400, w_297_1401, w_297_1409, w_297_1422, w_297_1431, w_297_1435, w_297_1443, w_297_1454, w_297_1462, w_297_1467, w_297_1475, w_297_1477, w_297_1479, w_297_1486, w_297_1487, w_297_1491, w_297_1496, w_297_1501, w_297_1507, w_297_1513, w_297_1540, w_297_1544, w_297_1545, w_297_1549, w_297_1560, w_297_1566, w_297_1571, w_297_1573, w_297_1574, w_297_1576, w_297_1577, w_297_1579, w_297_1608, w_297_1618, w_297_1620, w_297_1624, w_297_1629, w_297_1630, w_297_1639, w_297_1643, w_297_1644, w_297_1647, w_297_1670, w_297_1671, w_297_1682, w_297_1686, w_297_1688, w_297_1698, w_297_1699, w_297_1701, w_297_1708, w_297_1728, w_297_1731, w_297_1737, w_297_1748, w_297_1751, w_297_1753, w_297_1774, w_297_1775, w_297_1776, w_297_1787, w_297_1814, w_297_1817, w_297_1821, w_297_1826, w_297_1833, w_297_1835, w_297_1837, w_297_1845, w_297_1855, w_297_1858, w_297_1870, w_297_1873, w_297_1880, w_297_1881, w_297_1901, w_297_1905, w_297_1909, w_297_1917, w_297_1938, w_297_1943, w_297_1949, w_297_1954, w_297_1965, w_297_1968, w_297_1984, w_297_1992, w_297_1997, w_297_2002, w_297_2005, w_297_2009, w_297_2017, w_297_2024, w_297_2025, w_297_2035, w_297_2037, w_297_2038, w_297_2039, w_297_2040, w_297_2041, w_297_2042, w_297_2043, w_297_2044, w_297_2045, w_297_2047, w_297_2049, w_297_2050, w_297_2051, w_297_2055, w_297_2056, w_297_2057, w_297_2058, w_297_2059, w_297_2060, w_297_2062;
  wire w_298_001, w_298_009, w_298_015, w_298_020, w_298_024, w_298_031, w_298_036, w_298_040, w_298_055, w_298_073, w_298_083, w_298_099, w_298_103, w_298_120, w_298_128, w_298_133, w_298_140, w_298_144, w_298_171, w_298_172, w_298_174, w_298_193, w_298_195, w_298_197, w_298_206, w_298_209, w_298_218, w_298_226, w_298_254, w_298_262, w_298_267, w_298_268, w_298_274, w_298_281, w_298_282, w_298_285, w_298_287, w_298_298, w_298_315, w_298_318, w_298_319, w_298_322, w_298_325, w_298_345, w_298_387, w_298_388, w_298_391, w_298_394, w_298_399, w_298_403, w_298_404, w_298_427, w_298_429, w_298_439, w_298_444, w_298_445, w_298_447, w_298_448, w_298_449, w_298_463, w_298_469, w_298_474, w_298_485, w_298_504, w_298_508, w_298_511, w_298_512, w_298_518, w_298_523, w_298_530, w_298_542, w_298_553, w_298_582, w_298_583, w_298_600, w_298_611, w_298_638, w_298_644, w_298_652, w_298_656, w_298_658, w_298_659, w_298_661, w_298_671, w_298_672, w_298_680, w_298_686, w_298_696, w_298_698, w_298_715, w_298_716, w_298_745, w_298_750, w_298_778, w_298_781, w_298_784, w_298_791, w_298_813, w_298_827, w_298_830, w_298_842, w_298_849, w_298_855, w_298_870, w_298_882, w_298_884, w_298_885, w_298_886, w_298_888, w_298_890, w_298_891, w_298_892, w_298_900, w_298_909, w_298_917, w_298_942, w_298_943, w_298_947, w_298_953, w_298_963, w_298_966, w_298_980, w_298_981, w_298_982, w_298_984, w_298_985, w_298_987, w_298_989, w_298_1001, w_298_1006, w_298_1024, w_298_1030, w_298_1032, w_298_1048, w_298_1050, w_298_1055, w_298_1062, w_298_1071, w_298_1078, w_298_1080, w_298_1082, w_298_1083, w_298_1090, w_298_1092, w_298_1094, w_298_1098, w_298_1102, w_298_1105, w_298_1108, w_298_1125, w_298_1128, w_298_1131, w_298_1144, w_298_1149, w_298_1152, w_298_1155, w_298_1171, w_298_1177, w_298_1188, w_298_1198, w_298_1203, w_298_1204, w_298_1205, w_298_1226, w_298_1244, w_298_1247, w_298_1249, w_298_1254, w_298_1258, w_298_1260, w_298_1264, w_298_1265, w_298_1277, w_298_1283, w_298_1288, w_298_1302, w_298_1311, w_298_1325, w_298_1340, w_298_1341, w_298_1344, w_298_1355, w_298_1356, w_298_1362, w_298_1364, w_298_1365, w_298_1381, w_298_1387, w_298_1398, w_298_1406, w_298_1416, w_298_1417, w_298_1444, w_298_1447, w_298_1455, w_298_1456, w_298_1466, w_298_1487, w_298_1492, w_298_1500, w_298_1503, w_298_1505, w_298_1514, w_298_1516, w_298_1517, w_298_1520, w_298_1523, w_298_1526, w_298_1528, w_298_1533, w_298_1536, w_298_1540, w_298_1546, w_298_1565, w_298_1571, w_298_1582, w_298_1587, w_298_1590, w_298_1597, w_298_1618, w_298_1631, w_298_1645, w_298_1656, w_298_1671, w_298_1686, w_298_1688, w_298_1693, w_298_1704, w_298_1708, w_298_1714, w_298_1731, w_298_1735, w_298_1739, w_298_1743, w_298_1747, w_298_1748, w_298_1754, w_298_1759, w_298_1762, w_298_1779, w_298_1786, w_298_1791, w_298_1795, w_298_1811, w_298_1817, w_298_1824, w_298_1827, w_298_1828, w_298_1843, w_298_1846, w_298_1847, w_298_1854, w_298_1862, w_298_1865, w_298_1876, w_298_1883, w_298_1884, w_298_1891, w_298_1894, w_298_1931, w_298_1933, w_298_1938, w_298_1943, w_298_1952, w_298_1959, w_298_1960, w_298_1976, w_298_1978, w_298_1981, w_298_2005, w_298_2012, w_298_2016, w_298_2042, w_298_2053, w_298_2055, w_298_2068, w_298_2076, w_298_2086, w_298_2106, w_298_2122, w_298_2130, w_298_2140, w_298_2150, w_298_2152, w_298_2162, w_298_2177, w_298_2179, w_298_2227, w_298_2238, w_298_2246, w_298_2250, w_298_2252, w_298_2300, w_298_2320, w_298_2337, w_298_2350, w_298_2352, w_298_2355, w_298_2369, w_298_2373, w_298_2383, w_298_2386, w_298_2412, w_298_2417, w_298_2432, w_298_2433, w_298_2444, w_298_2473, w_298_2490, w_298_2504, w_298_2516, w_298_2528, w_298_2535, w_298_2559, w_298_2561, w_298_2564, w_298_2567, w_298_2568, w_298_2580, w_298_2582, w_298_2583, w_298_2599, w_298_2612, w_298_2625, w_298_2643, w_298_2644, w_298_2660, w_298_2667, w_298_2675, w_298_2700, w_298_2723, w_298_2732, w_298_2737, w_298_2741, w_298_2758, w_298_2765, w_298_2790, w_298_2793, w_298_2794, w_298_2810, w_298_2821, w_298_2832, w_298_2833, w_298_2843, w_298_2865, w_298_2904, w_298_2941, w_298_2966, w_298_2967, w_298_2974, w_298_2975, w_298_2976, w_298_2977, w_298_2978, w_298_2979;
  wire w_299_001, w_299_002, w_299_006, w_299_008, w_299_016, w_299_032, w_299_034, w_299_036, w_299_041, w_299_046, w_299_053, w_299_059, w_299_060, w_299_063, w_299_064, w_299_065, w_299_068, w_299_072, w_299_074, w_299_076, w_299_079, w_299_088, w_299_092, w_299_098, w_299_099, w_299_101, w_299_109, w_299_114, w_299_119, w_299_126, w_299_153, w_299_169, w_299_170, w_299_172, w_299_176, w_299_184, w_299_191, w_299_196, w_299_219, w_299_226, w_299_230, w_299_236, w_299_237, w_299_238, w_299_242, w_299_249, w_299_251, w_299_257, w_299_277, w_299_278, w_299_279, w_299_293, w_299_294, w_299_311, w_299_313, w_299_316, w_299_324, w_299_333, w_299_334, w_299_335, w_299_339, w_299_340, w_299_346, w_299_375, w_299_377, w_299_383, w_299_397, w_299_401, w_299_404, w_299_418, w_299_422, w_299_423, w_299_437, w_299_445, w_299_446, w_299_449, w_299_460, w_299_469, w_299_470, w_299_475, w_299_477, w_299_485, w_299_486, w_299_494, w_299_495, w_299_517, w_299_535, w_299_585, w_299_588, w_299_590, w_299_591, w_299_680, w_299_687, w_299_690, w_299_701, w_299_714, w_299_742, w_299_746, w_299_778, w_299_786, w_299_795, w_299_812, w_299_826, w_299_831, w_299_837, w_299_843, w_299_863, w_299_887, w_299_888, w_299_893, w_299_922, w_299_924, w_299_928, w_299_959, w_299_962, w_299_1022, w_299_1083, w_299_1099, w_299_1100, w_299_1105, w_299_1115, w_299_1148, w_299_1188, w_299_1211, w_299_1213, w_299_1239, w_299_1243, w_299_1247, w_299_1273, w_299_1308, w_299_1312, w_299_1321, w_299_1326, w_299_1343, w_299_1352, w_299_1357, w_299_1367, w_299_1408, w_299_1412, w_299_1415, w_299_1442, w_299_1453, w_299_1475, w_299_1492, w_299_1494, w_299_1624, w_299_1650, w_299_1675, w_299_1693, w_299_1717, w_299_1719, w_299_1724, w_299_1728, w_299_1749, w_299_1753, w_299_1761, w_299_1767, w_299_1769, w_299_1778, w_299_1779, w_299_1810, w_299_1816, w_299_1821, w_299_1826, w_299_1842, w_299_1845, w_299_1881, w_299_1890, w_299_1894, w_299_1918, w_299_1928, w_299_1934, w_299_1971, w_299_1989, w_299_2031, w_299_2037, w_299_2041, w_299_2070, w_299_2121, w_299_2123, w_299_2138, w_299_2143, w_299_2166, w_299_2169, w_299_2171, w_299_2174, w_299_2177, w_299_2181, w_299_2190, w_299_2196, w_299_2197, w_299_2207, w_299_2217, w_299_2231, w_299_2284, w_299_2287, w_299_2298, w_299_2317, w_299_2319, w_299_2326, w_299_2364, w_299_2400, w_299_2406, w_299_2429, w_299_2452, w_299_2475, w_299_2516, w_299_2552, w_299_2557, w_299_2560, w_299_2571, w_299_2574, w_299_2580, w_299_2602, w_299_2606, w_299_2614, w_299_2656, w_299_2661, w_299_2669, w_299_2695, w_299_2699, w_299_2704, w_299_2710, w_299_2721, w_299_2725, w_299_2739, w_299_2746, w_299_2752, w_299_2754, w_299_2761, w_299_2767, w_299_2786, w_299_2824, w_299_2828, w_299_2835, w_299_2874, w_299_2887, w_299_2893, w_299_2894, w_299_2906, w_299_2907, w_299_2921, w_299_2927, w_299_2934, w_299_2972, w_299_2988, w_299_2995, w_299_3014, w_299_3015, w_299_3037, w_299_3038, w_299_3041, w_299_3049, w_299_3079, w_299_3088, w_299_3098, w_299_3121, w_299_3125, w_299_3143, w_299_3154, w_299_3158, w_299_3167, w_299_3192, w_299_3209, w_299_3230, w_299_3251, w_299_3253, w_299_3270, w_299_3273, w_299_3280, w_299_3282, w_299_3291, w_299_3304, w_299_3359, w_299_3366, w_299_3373, w_299_3379, w_299_3419, w_299_3422, w_299_3449, w_299_3452, w_299_3454, w_299_3460, w_299_3463, w_299_3467, w_299_3469, w_299_3494, w_299_3496, w_299_3512, w_299_3529, w_299_3531, w_299_3534, w_299_3546, w_299_3547, w_299_3568, w_299_3608, w_299_3617, w_299_3619, w_299_3655, w_299_3705, w_299_3741, w_299_3747, w_299_3750, w_299_3753, w_299_3761, w_299_3762, w_299_3770, w_299_3773, w_299_3791, w_299_3803, w_299_3804, w_299_3819, w_299_3824, w_299_3832, w_299_3839, w_299_3850, w_299_3878, w_299_3906, w_299_3908, w_299_3916, w_299_3929, w_299_3944, w_299_3961, w_299_3967, w_299_3989, w_299_4000, w_299_4001, w_299_4003, w_299_4017, w_299_4026, w_299_4040, w_299_4063, w_299_4083, w_299_4088, w_299_4117, w_299_4122, w_299_4139, w_299_4156, w_299_4158, w_299_4174, w_299_4177, w_299_4231, w_299_4243, w_299_4258, w_299_4265, w_299_4280, w_299_4298, w_299_4299, w_299_4328, w_299_4332, w_299_4362, w_299_4364, w_299_4390, w_299_4400, w_299_4405, w_299_4411, w_299_4418, w_299_4423, w_299_4436, w_299_4452, w_299_4453, w_299_4460, w_299_4485, w_299_4520;
  wire w_300_002, w_300_006, w_300_010, w_300_012, w_300_014, w_300_016, w_300_017, w_300_022, w_300_025, w_300_027, w_300_029, w_300_032, w_300_037, w_300_039, w_300_040, w_300_046, w_300_050, w_300_070, w_300_075, w_300_078, w_300_079, w_300_083, w_300_092, w_300_099, w_300_102, w_300_106, w_300_110, w_300_114, w_300_115, w_300_123, w_300_134, w_300_143, w_300_147, w_300_151, w_300_155, w_300_156, w_300_158, w_300_162, w_300_163, w_300_171, w_300_172, w_300_173, w_300_180, w_300_184, w_300_190, w_300_191, w_300_194, w_300_202, w_300_203, w_300_217, w_300_221, w_300_225, w_300_226, w_300_229, w_300_237, w_300_244, w_300_254, w_300_256, w_300_275, w_300_277, w_300_285, w_300_302, w_300_304, w_300_308, w_300_310, w_300_311, w_300_335, w_300_339, w_300_350, w_300_351, w_300_356, w_300_358, w_300_368, w_300_372, w_300_375, w_300_378, w_300_382, w_300_386, w_300_388, w_300_393, w_300_397, w_300_412, w_300_413, w_300_423, w_300_425, w_300_426, w_300_431, w_300_438, w_300_439, w_300_446, w_300_449, w_300_454, w_300_466, w_300_471, w_300_472, w_300_474, w_300_479, w_300_490, w_300_494, w_300_495, w_300_498, w_300_526, w_300_530, w_300_534, w_300_543, w_300_546, w_300_547, w_300_548, w_300_553, w_300_560, w_300_562, w_300_564, w_300_580, w_300_591, w_300_594, w_300_613, w_300_618, w_300_628, w_300_633, w_300_640, w_300_646, w_300_655, w_300_656, w_300_657, w_300_659, w_300_663, w_300_667, w_300_669, w_300_670, w_300_671, w_300_676, w_300_677, w_300_690, w_300_692, w_300_707, w_300_708, w_300_711, w_300_716, w_300_723, w_300_728, w_300_749, w_300_761, w_300_765, w_300_767, w_300_768, w_300_769, w_300_770, w_300_772, w_300_773, w_300_779, w_300_796, w_300_802, w_300_804, w_300_805, w_300_808, w_300_813, w_300_814, w_300_815, w_300_825, w_300_829, w_300_833, w_300_844, w_300_845, w_300_848, w_300_851, w_300_859, w_300_865, w_300_877, w_300_881, w_300_884, w_300_886, w_300_887, w_300_894, w_300_898, w_300_899, w_300_902, w_300_908, w_300_909, w_300_910, w_300_914, w_300_916, w_300_918, w_300_922, w_300_923, w_300_929, w_300_935, w_300_939, w_300_954, w_300_955, w_300_965, w_300_985, w_300_988, w_300_1000, w_300_1001, w_300_1006, w_300_1007, w_300_1017, w_300_1019, w_300_1020, w_300_1021, w_300_1027, w_300_1034, w_300_1041, w_300_1044, w_300_1046, w_300_1053, w_300_1055, w_300_1056, w_300_1063, w_300_1072, w_300_1078, w_300_1081, w_300_1086, w_300_1090, w_300_1109, w_300_1112, w_300_1116, w_300_1117, w_300_1119, w_300_1125, w_300_1129, w_300_1133, w_300_1150, w_300_1152, w_300_1154, w_300_1161, w_300_1164, w_300_1165, w_300_1166, w_300_1167, w_300_1168, w_300_1175, w_300_1177, w_300_1182, w_300_1188, w_300_1198, w_300_1208, w_300_1215, w_300_1224, w_300_1230, w_300_1232, w_300_1236, w_300_1237, w_300_1239, w_300_1240, w_300_1242, w_300_1259, w_300_1260, w_300_1266, w_300_1274, w_300_1276, w_300_1285, w_300_1297, w_300_1298, w_300_1299, w_300_1304, w_300_1306, w_300_1309, w_300_1311, w_300_1323, w_300_1324, w_300_1327, w_300_1339, w_300_1342, w_300_1343, w_300_1349, w_300_1355, w_300_1359, w_300_1360, w_300_1363, w_300_1365, w_300_1366, w_300_1378, w_300_1386, w_300_1389, w_300_1391, w_300_1402, w_300_1404, w_300_1407, w_300_1410, w_300_1416, w_300_1419, w_300_1422, w_300_1425, w_300_1426, w_300_1428, w_300_1430, w_300_1438, w_300_1454, w_300_1457, w_300_1461, w_300_1463, w_300_1472, w_300_1474, w_300_1475, w_300_1483, w_300_1484, w_300_1497, w_300_1498, w_300_1503, w_300_1506, w_300_1509, w_300_1511, w_300_1513, w_300_1514, w_300_1529, w_300_1530, w_300_1533, w_300_1539, w_300_1547, w_300_1551, w_300_1552, w_300_1554, w_300_1556, w_300_1562, w_300_1565, w_300_1566, w_300_1574, w_300_1581, w_300_1582, w_300_1588, w_300_1593, w_300_1594, w_300_1597, w_300_1601, w_300_1609, w_300_1622, w_300_1624, w_300_1625;
  wire w_301_000, w_301_001, w_301_002, w_301_003, w_301_004, w_301_005, w_301_006, w_301_007, w_301_008, w_301_009, w_301_010, w_301_011, w_301_012, w_301_013, w_301_018, w_301_019, w_301_020, w_301_021, w_301_022, w_301_023, w_301_026, w_301_027, w_301_028, w_301_029, w_301_030, w_301_031, w_301_032, w_301_033, w_301_034, w_301_035, w_301_037, w_301_038, w_301_039, w_301_040, w_301_041, w_301_042, w_301_043, w_301_044, w_301_045, w_301_046, w_301_047, w_301_048, w_301_050, w_301_051, w_301_052, w_301_053, w_301_054, w_301_055, w_301_056, w_301_057, w_301_058, w_301_059, w_301_060, w_301_061, w_301_063, w_301_065, w_301_066, w_301_067, w_301_068, w_301_071, w_301_075, w_301_077, w_301_078, w_301_079, w_301_080, w_301_081, w_301_082, w_301_084, w_301_085, w_301_086, w_301_087, w_301_088, w_301_091, w_301_092, w_301_093, w_301_094, w_301_095, w_301_096, w_301_097, w_301_099, w_301_101, w_301_102, w_301_103, w_301_104, w_301_105, w_301_106, w_301_107, w_301_108, w_301_109, w_301_110, w_301_112, w_301_113, w_301_114, w_301_115, w_301_116, w_301_117, w_301_118, w_301_119, w_301_120, w_301_122, w_301_123, w_301_124, w_301_125, w_301_126, w_301_127, w_301_129, w_301_130, w_301_131, w_301_132, w_301_133, w_301_137, w_301_139, w_301_140, w_301_141, w_301_142, w_301_143, w_301_144, w_301_145, w_301_146, w_301_148, w_301_149, w_301_150, w_301_151, w_301_152, w_301_154, w_301_155, w_301_157, w_301_159, w_301_162, w_301_164, w_301_165, w_301_167, w_301_168, w_301_169, w_301_171, w_301_172, w_301_173, w_301_174, w_301_175, w_301_176, w_301_177, w_301_178, w_301_179, w_301_180, w_301_181, w_301_182, w_301_183, w_301_184, w_301_185, w_301_186, w_301_187, w_301_188, w_301_189, w_301_190, w_301_191, w_301_193, w_301_194, w_301_195, w_301_196, w_301_197, w_301_198, w_301_199, w_301_200, w_301_202, w_301_203, w_301_204, w_301_205, w_301_207, w_301_208, w_301_209, w_301_212, w_301_213, w_301_214, w_301_215, w_301_216, w_301_217, w_301_218, w_301_219, w_301_221, w_301_222;
  wire w_302_000, w_302_001, w_302_002, w_302_003, w_302_004, w_302_005, w_302_006, w_302_007, w_302_008, w_302_009, w_302_010, w_302_011, w_302_012, w_302_013, w_302_014, w_302_015, w_302_016, w_302_018, w_302_019, w_302_020, w_302_021, w_302_022, w_302_023, w_302_024, w_302_025, w_302_026, w_302_027, w_302_028, w_302_029;
  wire w_303_003, w_303_013, w_303_014, w_303_018, w_303_025, w_303_028, w_303_035, w_303_036, w_303_037, w_303_039, w_303_044, w_303_046, w_303_050, w_303_056, w_303_067, w_303_068, w_303_071, w_303_078, w_303_079, w_303_089, w_303_090, w_303_092, w_303_099, w_303_100, w_303_107, w_303_108, w_303_122, w_303_124, w_303_127, w_303_128, w_303_131, w_303_133, w_303_134, w_303_139, w_303_141, w_303_144, w_303_159, w_303_160, w_303_161, w_303_163, w_303_167, w_303_172, w_303_174, w_303_179, w_303_180, w_303_185, w_303_191, w_303_193, w_303_194, w_303_195, w_303_198, w_303_200, w_303_201, w_303_204, w_303_214, w_303_217, w_303_219, w_303_220, w_303_222, w_303_228, w_303_230, w_303_234, w_303_237, w_303_240, w_303_241, w_303_242, w_303_253, w_303_256, w_303_260, w_303_269, w_303_271, w_303_272, w_303_276, w_303_284, w_303_294, w_303_296, w_303_297, w_303_299, w_303_301, w_303_307, w_303_313, w_303_314, w_303_316, w_303_322, w_303_324, w_303_326, w_303_332, w_303_333, w_303_337, w_303_338, w_303_339, w_303_341, w_303_361, w_303_369, w_303_373, w_303_374, w_303_379, w_303_383, w_303_384, w_303_389, w_303_391, w_303_398, w_303_403, w_303_405, w_303_408, w_303_412, w_303_414, w_303_418, w_303_421, w_303_424, w_303_425, w_303_436, w_303_438, w_303_441, w_303_442, w_303_451, w_303_453, w_303_455, w_303_457, w_303_458, w_303_461, w_303_462, w_303_463, w_303_471, w_303_473, w_303_475, w_303_476, w_303_482, w_303_487, w_303_493, w_303_495, w_303_502, w_303_504, w_303_506, w_303_517, w_303_524, w_303_525, w_303_527, w_303_530, w_303_533, w_303_537, w_303_540, w_303_547, w_303_549, w_303_550, w_303_551, w_303_554, w_303_555, w_303_558, w_303_564, w_303_571, w_303_582, w_303_583, w_303_584, w_303_587, w_303_589, w_303_597, w_303_598, w_303_603, w_303_604, w_303_616, w_303_623, w_303_625, w_303_626, w_303_632, w_303_635, w_303_636, w_303_643, w_303_647, w_303_652, w_303_654, w_303_664, w_303_665, w_303_670, w_303_675, w_303_680, w_303_683, w_303_686, w_303_687, w_303_693, w_303_703, w_303_704, w_303_706, w_303_712, w_303_714, w_303_718, w_303_719, w_303_728, w_303_730, w_303_732, w_303_733, w_303_735, w_303_740, w_303_743, w_303_747, w_303_753, w_303_761, w_303_768, w_303_784, w_303_787, w_303_792, w_303_794, w_303_799, w_303_803, w_303_804, w_303_807, w_303_808, w_303_815, w_303_830, w_303_841, w_303_844, w_303_855, w_303_856, w_303_860, w_303_862, w_303_863, w_303_868, w_303_870, w_303_872, w_303_879, w_303_880, w_303_887, w_303_889, w_303_891, w_303_904, w_303_910, w_303_911, w_303_922, w_303_923, w_303_925, w_303_930, w_303_940, w_303_943, w_303_945, w_303_954, w_303_958, w_303_969, w_303_976, w_303_980, w_303_988, w_303_992, w_303_994, w_303_995, w_303_996, w_303_997, w_303_1000, w_303_1023, w_303_1025, w_303_1029, w_303_1030, w_303_1032, w_303_1033, w_303_1048, w_303_1052, w_303_1058, w_303_1060, w_303_1067, w_303_1068, w_303_1071, w_303_1072, w_303_1075, w_303_1077, w_303_1078, w_303_1082, w_303_1089, w_303_1100, w_303_1101, w_303_1103, w_303_1110, w_303_1114, w_303_1116, w_303_1117, w_303_1125, w_303_1128, w_303_1133, w_303_1135, w_303_1140, w_303_1142, w_303_1153, w_303_1156, w_303_1157, w_303_1161, w_303_1163, w_303_1168, w_303_1173, w_303_1178, w_303_1180, w_303_1189, w_303_1205, w_303_1208, w_303_1210, w_303_1211, w_303_1215, w_303_1221, w_303_1229, w_303_1240, w_303_1241, w_303_1247, w_303_1249, w_303_1253, w_303_1256, w_303_1264, w_303_1266, w_303_1270, w_303_1271, w_303_1274, w_303_1275, w_303_1278, w_303_1285, w_303_1289, w_303_1296, w_303_1308, w_303_1314, w_303_1324, w_303_1347, w_303_1351, w_303_1352, w_303_1354, w_303_1356, w_303_1357, w_303_1360, w_303_1367, w_303_1369, w_303_1371, w_303_1376, w_303_1381, w_303_1386, w_303_1395, w_303_1400, w_303_1401, w_303_1402, w_303_1404, w_303_1438, w_303_1439, w_303_1440, w_303_1442, w_303_1445, w_303_1448, w_303_1450, w_303_1453, w_303_1456, w_303_1462, w_303_1464, w_303_1466, w_303_1468;
  wire w_304_003, w_304_004, w_304_006, w_304_007, w_304_008, w_304_009, w_304_013, w_304_018, w_304_020, w_304_023, w_304_025, w_304_032, w_304_041, w_304_043, w_304_044, w_304_046, w_304_048, w_304_049, w_304_051, w_304_057, w_304_059, w_304_060, w_304_061, w_304_067, w_304_068, w_304_070, w_304_074, w_304_078, w_304_080, w_304_097, w_304_099, w_304_101, w_304_102, w_304_103, w_304_114, w_304_126, w_304_130, w_304_143, w_304_145, w_304_147, w_304_148, w_304_159, w_304_160, w_304_161, w_304_167, w_304_169, w_304_170, w_304_171, w_304_173, w_304_174, w_304_180, w_304_185, w_304_188, w_304_190, w_304_191, w_304_192, w_304_195, w_304_199, w_304_203, w_304_204, w_304_205, w_304_210, w_304_211, w_304_214, w_304_215, w_304_216, w_304_218, w_304_222, w_304_227, w_304_229, w_304_232, w_304_235, w_304_237, w_304_238, w_304_239, w_304_241, w_304_247, w_304_257, w_304_264, w_304_265, w_304_266, w_304_270, w_304_277, w_304_279, w_304_284, w_304_285, w_304_286, w_304_287, w_304_288, w_304_290, w_304_292, w_304_295, w_304_296, w_304_302, w_304_303, w_304_306, w_304_314, w_304_318, w_304_320, w_304_323, w_304_324, w_304_328, w_304_329, w_304_331, w_304_332, w_304_336, w_304_341, w_304_345, w_304_353, w_304_354, w_304_377, w_304_383, w_304_388, w_304_390, w_304_408, w_304_409, w_304_413, w_304_417, w_304_420, w_304_423, w_304_425, w_304_428, w_304_439, w_304_441, w_304_444, w_304_446, w_304_447, w_304_449, w_304_453, w_304_460, w_304_463, w_304_467, w_304_476, w_304_483, w_304_487, w_304_494, w_304_496, w_304_505, w_304_517, w_304_525, w_304_527, w_304_540, w_304_541, w_304_549, w_304_552, w_304_555, w_304_556, w_304_558, w_304_560, w_304_570, w_304_571, w_304_574, w_304_576, w_304_577, w_304_580, w_304_586, w_304_597, w_304_602, w_304_614, w_304_618, w_304_619, w_304_634, w_304_637, w_304_641, w_304_643, w_304_648, w_304_651, w_304_654, w_304_655, w_304_658, w_304_663, w_304_665, w_304_669, w_304_675, w_304_682, w_304_692, w_304_696, w_304_697, w_304_709, w_304_712, w_304_713, w_304_714, w_304_716, w_304_717, w_304_721, w_304_726, w_304_729, w_304_731, w_304_736, w_304_741, w_304_748, w_304_750, w_304_751, w_304_754, w_304_756, w_304_764, w_304_769, w_304_770, w_304_772, w_304_777, w_304_778, w_304_782, w_304_788, w_304_790, w_304_795, w_304_797, w_304_804, w_304_810, w_304_812, w_304_818, w_304_822, w_304_823, w_304_828, w_304_833, w_304_841, w_304_843, w_304_844, w_304_850, w_304_852, w_304_862, w_304_864, w_304_869, w_304_877, w_304_878, w_304_881, w_304_884, w_304_888, w_304_892, w_304_903, w_304_904, w_304_911, w_304_915, w_304_916, w_304_926, w_304_941, w_304_950, w_304_956, w_304_957, w_304_958, w_304_963, w_304_972, w_304_975, w_304_981, w_304_984, w_304_991, w_304_995, w_304_1005, w_304_1006, w_304_1009, w_304_1014, w_304_1024, w_304_1027, w_304_1028, w_304_1030, w_304_1036, w_304_1037, w_304_1038, w_304_1040, w_304_1041, w_304_1042, w_304_1045, w_304_1062, w_304_1064, w_304_1066, w_304_1071, w_304_1079, w_304_1080, w_304_1085, w_304_1087, w_304_1091, w_304_1096, w_304_1110, w_304_1113, w_304_1118, w_304_1119, w_304_1126, w_304_1127, w_304_1136, w_304_1150, w_304_1158, w_304_1169, w_304_1170, w_304_1171, w_304_1172, w_304_1174, w_304_1175, w_304_1176, w_304_1177, w_304_1178, w_304_1179, w_304_1181, w_304_1182, w_304_1191, w_304_1194, w_304_1196, w_304_1200, w_304_1205, w_304_1214, w_304_1216, w_304_1221, w_304_1222, w_304_1224, w_304_1225, w_304_1227, w_304_1232, w_304_1243, w_304_1247, w_304_1251, w_304_1258, w_304_1260, w_304_1261, w_304_1262, w_304_1278, w_304_1281, w_304_1282, w_304_1283, w_304_1287, w_304_1288, w_304_1292, w_304_1294, w_304_1300, w_304_1302, w_304_1306, w_304_1316, w_304_1317, w_304_1318, w_304_1320, w_304_1328, w_304_1339, w_304_1345, w_304_1349, w_304_1350, w_304_1353, w_304_1359, w_304_1362, w_304_1372, w_304_1374, w_304_1375, w_304_1381, w_304_1394, w_304_1399, w_304_1401, w_304_1402;
  wire w_305_007, w_305_013, w_305_021, w_305_023, w_305_033, w_305_046, w_305_049, w_305_052, w_305_059, w_305_071, w_305_072, w_305_075, w_305_083, w_305_086, w_305_090, w_305_095, w_305_099, w_305_100, w_305_114, w_305_115, w_305_131, w_305_144, w_305_149, w_305_159, w_305_161, w_305_163, w_305_164, w_305_190, w_305_192, w_305_197, w_305_198, w_305_202, w_305_207, w_305_238, w_305_253, w_305_263, w_305_272, w_305_292, w_305_302, w_305_307, w_305_324, w_305_330, w_305_358, w_305_376, w_305_380, w_305_384, w_305_387, w_305_394, w_305_420, w_305_426, w_305_427, w_305_461, w_305_478, w_305_485, w_305_488, w_305_518, w_305_537, w_305_538, w_305_543, w_305_551, w_305_606, w_305_619, w_305_625, w_305_628, w_305_638, w_305_652, w_305_658, w_305_665, w_305_670, w_305_681, w_305_713, w_305_728, w_305_756, w_305_760, w_305_780, w_305_826, w_305_829, w_305_830, w_305_845, w_305_855, w_305_857, w_305_870, w_305_886, w_305_900, w_305_905, w_305_907, w_305_925, w_305_933, w_305_939, w_305_944, w_305_945, w_305_948, w_305_951, w_305_960, w_305_983, w_305_989, w_305_996, w_305_1000, w_305_1009, w_305_1043, w_305_1053, w_305_1055, w_305_1077, w_305_1089, w_305_1105, w_305_1109, w_305_1150, w_305_1157, w_305_1188, w_305_1212, w_305_1234, w_305_1243, w_305_1255, w_305_1343, w_305_1353, w_305_1358, w_305_1365, w_305_1380, w_305_1407, w_305_1418, w_305_1429, w_305_1434, w_305_1438, w_305_1463, w_305_1466, w_305_1472, w_305_1489, w_305_1497, w_305_1504, w_305_1514, w_305_1522, w_305_1539, w_305_1542, w_305_1569, w_305_1576, w_305_1584, w_305_1597, w_305_1602, w_305_1619, w_305_1645, w_305_1667, w_305_1672, w_305_1679, w_305_1683, w_305_1719, w_305_1725, w_305_1764, w_305_1766, w_305_1787, w_305_1789, w_305_1794, w_305_1801, w_305_1834, w_305_1853, w_305_1881, w_305_1892, w_305_1893, w_305_1911, w_305_1915, w_305_1917, w_305_1918, w_305_1958, w_305_1963, w_305_1966, w_305_1967, w_305_1979, w_305_1984, w_305_1990, w_305_2001, w_305_2002, w_305_2003, w_305_2011, w_305_2025, w_305_2050, w_305_2055, w_305_2086, w_305_2090, w_305_2094, w_305_2108, w_305_2109, w_305_2128, w_305_2140, w_305_2169, w_305_2184, w_305_2208, w_305_2216, w_305_2229, w_305_2292, w_305_2308, w_305_2317, w_305_2318, w_305_2322, w_305_2351, w_305_2372, w_305_2386, w_305_2403, w_305_2406, w_305_2419, w_305_2443, w_305_2446, w_305_2466, w_305_2471, w_305_2473, w_305_2474, w_305_2482, w_305_2489, w_305_2509, w_305_2512, w_305_2567, w_305_2569, w_305_2576, w_305_2579, w_305_2594, w_305_2595, w_305_2607, w_305_2626, w_305_2630, w_305_2634, w_305_2635, w_305_2655, w_305_2664, w_305_2688, w_305_2714, w_305_2716, w_305_2718, w_305_2721, w_305_2722, w_305_2742, w_305_2753, w_305_2786, w_305_2789, w_305_2799, w_305_2805, w_305_2819, w_305_2877, w_305_2880, w_305_2884, w_305_2919, w_305_2922, w_305_2943, w_305_2970, w_305_2971, w_305_3006, w_305_3016, w_305_3054, w_305_3084, w_305_3104, w_305_3113, w_305_3117, w_305_3139, w_305_3155, w_305_3165, w_305_3184, w_305_3196, w_305_3203, w_305_3216, w_305_3219, w_305_3221, w_305_3223, w_305_3262, w_305_3265, w_305_3266, w_305_3289, w_305_3298, w_305_3330, w_305_3339, w_305_3348, w_305_3358, w_305_3363, w_305_3369, w_305_3377, w_305_3394, w_305_3397, w_305_3412, w_305_3445, w_305_3468, w_305_3471, w_305_3481, w_305_3484, w_305_3485, w_305_3510, w_305_3517, w_305_3530, w_305_3545, w_305_3547, w_305_3567, w_305_3570, w_305_3571, w_305_3599, w_305_3603, w_305_3616, w_305_3636, w_305_3640, w_305_3641, w_305_3643, w_305_3644, w_305_3658, w_305_3695, w_305_3699, w_305_3700, w_305_3710, w_305_3714, w_305_3738, w_305_3741, w_305_3754, w_305_3761, w_305_3766, w_305_3795, w_305_3799, w_305_3801, w_305_3805, w_305_3815, w_305_3821, w_305_3827, w_305_3842, w_305_3865, w_305_3873, w_305_3876, w_305_3879, w_305_3904, w_305_3938, w_305_3942, w_305_3990, w_305_4027, w_305_4083, w_305_4084, w_305_4090, w_305_4092, w_305_4097, w_305_4101, w_305_4109, w_305_4111, w_305_4112, w_305_4114, w_305_4120, w_305_4132, w_305_4140, w_305_4185, w_305_4195, w_305_4224, w_305_4227, w_305_4234, w_305_4251, w_305_4262, w_305_4263, w_305_4287, w_305_4289, w_305_4298, w_305_4319, w_305_4329, w_305_4342, w_305_4365, w_305_4369, w_305_4391, w_305_4394, w_305_4401, w_305_4424, w_305_4452, w_305_4462, w_305_4464, w_305_4494, w_305_4534, w_305_4538, w_305_4576, w_305_4582, w_305_4583, w_305_4587, w_305_4596, w_305_4612, w_305_4623, w_305_4626, w_305_4647, w_305_4650, w_305_4682, w_305_4706, w_305_4716, w_305_4753, w_305_4758, w_305_4769;
  wire w_306_001, w_306_004, w_306_005, w_306_014, w_306_018, w_306_024, w_306_033, w_306_036, w_306_044, w_306_045, w_306_046, w_306_050, w_306_052, w_306_056, w_306_061, w_306_064, w_306_065, w_306_067, w_306_071, w_306_073, w_306_075, w_306_082, w_306_086, w_306_097, w_306_099, w_306_119, w_306_121, w_306_123, w_306_130, w_306_141, w_306_142, w_306_146, w_306_157, w_306_159, w_306_160, w_306_163, w_306_166, w_306_167, w_306_170, w_306_171, w_306_181, w_306_190, w_306_194, w_306_195, w_306_196, w_306_199, w_306_202, w_306_208, w_306_213, w_306_216, w_306_219, w_306_222, w_306_223, w_306_226, w_306_231, w_306_232, w_306_238, w_306_247, w_306_253, w_306_255, w_306_262, w_306_264, w_306_267, w_306_268, w_306_274, w_306_275, w_306_282, w_306_287, w_306_289, w_306_305, w_306_308, w_306_311, w_306_315, w_306_316, w_306_323, w_306_324, w_306_329, w_306_332, w_306_334, w_306_339, w_306_340, w_306_347, w_306_350, w_306_352, w_306_359, w_306_371, w_306_393, w_306_395, w_306_401, w_306_402, w_306_403, w_306_407, w_306_410, w_306_412, w_306_416, w_306_425, w_306_431, w_306_433, w_306_441, w_306_445, w_306_452, w_306_459, w_306_477, w_306_490, w_306_492, w_306_494, w_306_497, w_306_502, w_306_504, w_306_506, w_306_511, w_306_513, w_306_514, w_306_515, w_306_521, w_306_533, w_306_537, w_306_538, w_306_542, w_306_543, w_306_545, w_306_561, w_306_571, w_306_577, w_306_581, w_306_583, w_306_584, w_306_596, w_306_599, w_306_612, w_306_614, w_306_616, w_306_617, w_306_618, w_306_620, w_306_625, w_306_639, w_306_651, w_306_653, w_306_658, w_306_673, w_306_680, w_306_683, w_306_685, w_306_687, w_306_690, w_306_704, w_306_706, w_306_712, w_306_715, w_306_717, w_306_720, w_306_721, w_306_733, w_306_744, w_306_745, w_306_763, w_306_766, w_306_771, w_306_782, w_306_784, w_306_794, w_306_796, w_306_799, w_306_804, w_306_807, w_306_818, w_306_823, w_306_825, w_306_826, w_306_827, w_306_829, w_306_830, w_306_834, w_306_837, w_306_847, w_306_850, w_306_851, w_306_855, w_306_857, w_306_862, w_306_870, w_306_874, w_306_879, w_306_881, w_306_883, w_306_885, w_306_891, w_306_894, w_306_896, w_306_898, w_306_901, w_306_903, w_306_906, w_306_913, w_306_933, w_306_936, w_306_939, w_306_944, w_306_951, w_306_978, w_306_984, w_306_990, w_306_993, w_306_995, w_306_1000, w_306_1002, w_306_1003, w_306_1005, w_306_1014, w_306_1017, w_306_1023, w_306_1027, w_306_1030, w_306_1033, w_306_1037, w_306_1042, w_306_1045, w_306_1048, w_306_1053, w_306_1066, w_306_1069, w_306_1072, w_306_1073, w_306_1074, w_306_1087, w_306_1094, w_306_1095, w_306_1097, w_306_1101, w_306_1103, w_306_1106, w_306_1107, w_306_1112, w_306_1116, w_306_1120, w_306_1137, w_306_1138, w_306_1139, w_306_1140, w_306_1141, w_306_1144, w_306_1145, w_306_1150, w_306_1156, w_306_1181, w_306_1185, w_306_1190, w_306_1192, w_306_1199, w_306_1202, w_306_1204, w_306_1206, w_306_1209, w_306_1215, w_306_1218, w_306_1220, w_306_1222, w_306_1225, w_306_1226, w_306_1233, w_306_1234, w_306_1237, w_306_1243, w_306_1244, w_306_1245, w_306_1248, w_306_1249, w_306_1250, w_306_1252, w_306_1253, w_306_1257, w_306_1261, w_306_1265, w_306_1282, w_306_1285, w_306_1293, w_306_1309, w_306_1316, w_306_1328, w_306_1329, w_306_1344, w_306_1363, w_306_1370, w_306_1377, w_306_1385, w_306_1390, w_306_1391, w_306_1392, w_306_1410, w_306_1417, w_306_1430, w_306_1433, w_306_1440, w_306_1443, w_306_1446, w_306_1451, w_306_1470, w_306_1479, w_306_1480, w_306_1498, w_306_1514, w_306_1517, w_306_1520, w_306_1521, w_306_1532, w_306_1539, w_306_1542, w_306_1547, w_306_1548, w_306_1561, w_306_1564, w_306_1585, w_306_1588, w_306_1593, w_306_1605, w_306_1607, w_306_1617, w_306_1624, w_306_1642, w_306_1647, w_306_1651, w_306_1657, w_306_1669, w_306_1674, w_306_1679, w_306_1685, w_306_1688, w_306_1694, w_306_1699, w_306_1704, w_306_1726, w_306_1734, w_306_1737, w_306_1741, w_306_1751, w_306_1770, w_306_1776, w_306_1785, w_306_1787, w_306_1790, w_306_1799;
  wire w_307_003, w_307_004, w_307_011, w_307_024, w_307_034, w_307_051, w_307_054, w_307_058, w_307_059, w_307_080, w_307_084, w_307_088, w_307_089, w_307_097, w_307_100, w_307_102, w_307_115, w_307_123, w_307_127, w_307_133, w_307_137, w_307_146, w_307_153, w_307_156, w_307_162, w_307_188, w_307_194, w_307_197, w_307_201, w_307_213, w_307_217, w_307_226, w_307_233, w_307_235, w_307_243, w_307_252, w_307_254, w_307_256, w_307_286, w_307_291, w_307_307, w_307_308, w_307_311, w_307_313, w_307_326, w_307_337, w_307_341, w_307_344, w_307_349, w_307_350, w_307_353, w_307_359, w_307_365, w_307_369, w_307_373, w_307_391, w_307_418, w_307_432, w_307_440, w_307_445, w_307_454, w_307_460, w_307_462, w_307_463, w_307_493, w_307_494, w_307_497, w_307_507, w_307_516, w_307_519, w_307_521, w_307_527, w_307_540, w_307_542, w_307_543, w_307_553, w_307_574, w_307_579, w_307_582, w_307_592, w_307_618, w_307_625, w_307_637, w_307_670, w_307_678, w_307_679, w_307_687, w_307_690, w_307_702, w_307_709, w_307_717, w_307_725, w_307_729, w_307_732, w_307_747, w_307_752, w_307_755, w_307_763, w_307_766, w_307_772, w_307_773, w_307_777, w_307_783, w_307_787, w_307_791, w_307_793, w_307_795, w_307_805, w_307_820, w_307_827, w_307_837, w_307_838, w_307_850, w_307_872, w_307_874, w_307_882, w_307_894, w_307_902, w_307_909, w_307_916, w_307_932, w_307_933, w_307_941, w_307_948, w_307_955, w_307_961, w_307_974, w_307_981, w_307_986, w_307_988, w_307_1001, w_307_1009, w_307_1013, w_307_1016, w_307_1020, w_307_1026, w_307_1036, w_307_1039, w_307_1044, w_307_1066, w_307_1071, w_307_1076, w_307_1079, w_307_1086, w_307_1087, w_307_1097, w_307_1098, w_307_1099, w_307_1108, w_307_1120, w_307_1121, w_307_1122, w_307_1138, w_307_1139, w_307_1142, w_307_1145, w_307_1148, w_307_1151, w_307_1168, w_307_1169, w_307_1194, w_307_1212, w_307_1213, w_307_1217, w_307_1220, w_307_1227, w_307_1229, w_307_1230, w_307_1244, w_307_1246, w_307_1249, w_307_1252, w_307_1255, w_307_1257, w_307_1260, w_307_1264, w_307_1280, w_307_1281, w_307_1291, w_307_1313, w_307_1320, w_307_1324, w_307_1331, w_307_1332, w_307_1334, w_307_1335, w_307_1339, w_307_1344, w_307_1348, w_307_1353, w_307_1363, w_307_1370, w_307_1379, w_307_1387, w_307_1424, w_307_1436, w_307_1470, w_307_1496, w_307_1524, w_307_1537, w_307_1541, w_307_1546, w_307_1548, w_307_1552, w_307_1586, w_307_1587, w_307_1594, w_307_1614, w_307_1618, w_307_1625, w_307_1626, w_307_1630, w_307_1693, w_307_1695, w_307_1712, w_307_1717, w_307_1718, w_307_1724, w_307_1733, w_307_1779, w_307_1804, w_307_1810, w_307_1817, w_307_1829, w_307_1838, w_307_1847, w_307_1886, w_307_1898, w_307_1910, w_307_1911, w_307_1939, w_307_1945, w_307_1951, w_307_1985, w_307_1997, w_307_2002, w_307_2012, w_307_2022, w_307_2023, w_307_2037, w_307_2054, w_307_2058, w_307_2064, w_307_2065, w_307_2082, w_307_2105, w_307_2125, w_307_2143, w_307_2182, w_307_2188, w_307_2195, w_307_2201, w_307_2215, w_307_2222, w_307_2234, w_307_2236, w_307_2259, w_307_2261, w_307_2274, w_307_2278, w_307_2279, w_307_2284, w_307_2299, w_307_2302, w_307_2311, w_307_2316, w_307_2325, w_307_2333, w_307_2337, w_307_2348, w_307_2351, w_307_2363, w_307_2369, w_307_2400, w_307_2410, w_307_2417, w_307_2453, w_307_2461, w_307_2469, w_307_2482, w_307_2488, w_307_2490, w_307_2500, w_307_2505, w_307_2513, w_307_2522, w_307_2527, w_307_2541, w_307_2559, w_307_2562, w_307_2565, w_307_2569, w_307_2572, w_307_2580, w_307_2602, w_307_2609, w_307_2612, w_307_2615, w_307_2617, w_307_2650, w_307_2683, w_307_2688, w_307_2689, w_307_2697, w_307_2722, w_307_2728, w_307_2729, w_307_2746, w_307_2772, w_307_2775, w_307_2780, w_307_2809, w_307_2830, w_307_2835, w_307_2870, w_307_2913, w_307_2917, w_307_2922, w_307_2946, w_307_2972, w_307_2991, w_307_3023, w_307_3048, w_307_3059, w_307_3066, w_307_3076, w_307_3093, w_307_3100, w_307_3135, w_307_3179, w_307_3207, w_307_3217, w_307_3221, w_307_3229, w_307_3231, w_307_3250, w_307_3254, w_307_3286, w_307_3291, w_307_3294, w_307_3319, w_307_3322, w_307_3350, w_307_3365, w_307_3370, w_307_3371, w_307_3375, w_307_3384, w_307_3391, w_307_3392, w_307_3413, w_307_3415, w_307_3433, w_307_3462, w_307_3474, w_307_3476, w_307_3494, w_307_3527, w_307_3551, w_307_3554, w_307_3564, w_307_3572, w_307_3584, w_307_3587, w_307_3599, w_307_3606;
  wire w_308_000, w_308_002, w_308_008, w_308_010, w_308_011, w_308_013, w_308_016, w_308_017, w_308_020, w_308_021, w_308_022, w_308_031, w_308_034, w_308_047, w_308_050, w_308_052, w_308_053, w_308_054, w_308_056, w_308_058, w_308_060, w_308_068, w_308_084, w_308_086, w_308_090, w_308_091, w_308_105, w_308_110, w_308_111, w_308_122, w_308_128, w_308_132, w_308_134, w_308_136, w_308_139, w_308_142, w_308_146, w_308_150, w_308_152, w_308_158, w_308_167, w_308_171, w_308_179, w_308_182, w_308_184, w_308_191, w_308_193, w_308_197, w_308_199, w_308_210, w_308_212, w_308_214, w_308_215, w_308_228, w_308_230, w_308_232, w_308_235, w_308_249, w_308_254, w_308_258, w_308_261, w_308_263, w_308_267, w_308_275, w_308_277, w_308_279, w_308_290, w_308_298, w_308_300, w_308_301, w_308_306, w_308_312, w_308_313, w_308_321, w_308_322, w_308_327, w_308_332, w_308_333, w_308_336, w_308_337, w_308_344, w_308_350, w_308_356, w_308_358, w_308_359, w_308_361, w_308_365, w_308_376, w_308_381, w_308_385, w_308_388, w_308_393, w_308_394, w_308_400, w_308_402, w_308_419, w_308_428, w_308_432, w_308_434, w_308_435, w_308_438, w_308_440, w_308_441, w_308_442, w_308_448, w_308_449, w_308_458, w_308_460, w_308_463, w_308_467, w_308_468, w_308_469, w_308_472, w_308_475, w_308_478, w_308_482, w_308_484, w_308_485, w_308_488, w_308_500, w_308_502, w_308_507, w_308_508, w_308_511, w_308_515, w_308_517, w_308_518, w_308_523, w_308_524, w_308_526, w_308_529, w_308_536, w_308_537, w_308_539, w_308_542, w_308_543, w_308_544, w_308_546, w_308_547, w_308_548, w_308_558, w_308_559, w_308_565, w_308_572, w_308_573, w_308_575, w_308_583, w_308_587, w_308_596, w_308_597, w_308_608, w_308_610, w_308_619, w_308_620, w_308_623, w_308_626, w_308_634, w_308_636, w_308_640, w_308_641, w_308_646, w_308_654, w_308_656, w_308_659, w_308_660, w_308_661, w_308_667, w_308_676, w_308_678, w_308_680, w_308_688, w_308_689, w_308_694, w_308_696, w_308_697, w_308_709, w_308_712, w_308_721, w_308_723, w_308_730, w_308_731, w_308_737, w_308_740, w_308_742, w_308_743, w_308_748, w_308_754, w_308_758, w_308_762, w_308_764, w_308_766, w_308_767, w_308_769, w_308_773, w_308_775, w_308_780, w_308_782, w_308_784, w_308_793, w_308_798, w_308_801, w_308_805, w_308_806, w_308_816, w_308_824, w_308_827, w_308_829, w_308_832, w_308_833, w_308_834, w_308_839, w_308_842, w_308_846, w_308_847, w_308_849, w_308_852, w_308_855, w_308_864, w_308_865, w_308_868, w_308_873, w_308_878, w_308_881, w_308_889, w_308_897, w_308_907, w_308_908, w_308_912, w_308_913, w_308_915, w_308_916, w_308_918, w_308_920, w_308_930, w_308_931, w_308_936, w_308_937, w_308_943, w_308_944, w_308_957, w_308_959, w_308_961, w_308_962, w_308_968, w_308_979, w_308_980, w_308_982, w_308_984, w_308_986, w_308_988, w_308_989, w_308_993, w_308_994, w_308_995, w_308_1000, w_308_1001, w_308_1008, w_308_1013, w_308_1017, w_308_1018, w_308_1019, w_308_1022, w_308_1023, w_308_1024, w_308_1027, w_308_1031, w_308_1032, w_308_1035, w_308_1043, w_308_1047, w_308_1062, w_308_1065, w_308_1067, w_308_1068, w_308_1069, w_308_1070, w_308_1072, w_308_1078, w_308_1082, w_308_1088, w_308_1094, w_308_1096, w_308_1098, w_308_1099, w_308_1100, w_308_1101, w_308_1105, w_308_1106, w_308_1110, w_308_1111, w_308_1117, w_308_1118, w_308_1126, w_308_1127, w_308_1128, w_308_1143, w_308_1167, w_308_1172, w_308_1173, w_308_1176, w_308_1178, w_308_1180, w_308_1184, w_308_1186, w_308_1195, w_308_1196, w_308_1201, w_308_1203, w_308_1204, w_308_1208, w_308_1222, w_308_1223, w_308_1226, w_308_1231, w_308_1233, w_308_1236, w_308_1241, w_308_1249, w_308_1254, w_308_1258, w_308_1275, w_308_1280, w_308_1286;
  wire w_309_001, w_309_004, w_309_011, w_309_013, w_309_016, w_309_024, w_309_028, w_309_029, w_309_031, w_309_033, w_309_043, w_309_044, w_309_064, w_309_078, w_309_079, w_309_080, w_309_081, w_309_086, w_309_088, w_309_107, w_309_114, w_309_115, w_309_129, w_309_130, w_309_134, w_309_136, w_309_138, w_309_139, w_309_142, w_309_149, w_309_156, w_309_157, w_309_165, w_309_166, w_309_168, w_309_171, w_309_180, w_309_182, w_309_186, w_309_189, w_309_190, w_309_192, w_309_194, w_309_205, w_309_207, w_309_223, w_309_232, w_309_233, w_309_234, w_309_238, w_309_249, w_309_250, w_309_252, w_309_256, w_309_257, w_309_261, w_309_266, w_309_267, w_309_272, w_309_274, w_309_275, w_309_288, w_309_292, w_309_294, w_309_296, w_309_300, w_309_305, w_309_311, w_309_314, w_309_315, w_309_317, w_309_319, w_309_326, w_309_339, w_309_343, w_309_346, w_309_347, w_309_363, w_309_364, w_309_366, w_309_367, w_309_368, w_309_369, w_309_372, w_309_373, w_309_383, w_309_386, w_309_395, w_309_407, w_309_413, w_309_419, w_309_427, w_309_429, w_309_435, w_309_452, w_309_460, w_309_461, w_309_465, w_309_478, w_309_480, w_309_484, w_309_485, w_309_497, w_309_503, w_309_509, w_309_510, w_309_527, w_309_531, w_309_550, w_309_553, w_309_555, w_309_556, w_309_568, w_309_586, w_309_593, w_309_598, w_309_599, w_309_603, w_309_619, w_309_628, w_309_645, w_309_647, w_309_655, w_309_664, w_309_665, w_309_667, w_309_669, w_309_678, w_309_684, w_309_698, w_309_703, w_309_710, w_309_711, w_309_712, w_309_718, w_309_720, w_309_728, w_309_730, w_309_731, w_309_734, w_309_744, w_309_750, w_309_756, w_309_760, w_309_762, w_309_763, w_309_776, w_309_788, w_309_791, w_309_793, w_309_794, w_309_800, w_309_801, w_309_806, w_309_823, w_309_832, w_309_837, w_309_839, w_309_845, w_309_848, w_309_853, w_309_858, w_309_863, w_309_865, w_309_867, w_309_883, w_309_890, w_309_891, w_309_897, w_309_900, w_309_904, w_309_913, w_309_931, w_309_939, w_309_957, w_309_959, w_309_960, w_309_963, w_309_964, w_309_969, w_309_970, w_309_971, w_309_972, w_309_977, w_309_981, w_309_982, w_309_983, w_309_987, w_309_991, w_309_992, w_309_993, w_309_998, w_309_999, w_309_1004, w_309_1012, w_309_1013, w_309_1015, w_309_1017, w_309_1018, w_309_1025, w_309_1029, w_309_1031, w_309_1034, w_309_1036, w_309_1045, w_309_1050, w_309_1058, w_309_1060, w_309_1067, w_309_1068, w_309_1069, w_309_1072, w_309_1074, w_309_1076, w_309_1077, w_309_1080, w_309_1092, w_309_1094, w_309_1096, w_309_1100, w_309_1101, w_309_1113, w_309_1114, w_309_1120, w_309_1127, w_309_1130, w_309_1131, w_309_1137, w_309_1150, w_309_1162, w_309_1166, w_309_1172, w_309_1173, w_309_1188, w_309_1192, w_309_1197, w_309_1199, w_309_1200, w_309_1201, w_309_1212, w_309_1223, w_309_1224, w_309_1231, w_309_1238, w_309_1249, w_309_1252, w_309_1253, w_309_1256, w_309_1258, w_309_1264, w_309_1268, w_309_1276, w_309_1279, w_309_1280, w_309_1281, w_309_1286, w_309_1299, w_309_1314, w_309_1319, w_309_1323, w_309_1326, w_309_1337, w_309_1353, w_309_1354, w_309_1358, w_309_1360, w_309_1367, w_309_1374, w_309_1376, w_309_1380, w_309_1385, w_309_1388, w_309_1390, w_309_1392, w_309_1398, w_309_1403, w_309_1409, w_309_1410, w_309_1413, w_309_1419, w_309_1437, w_309_1440, w_309_1441, w_309_1445, w_309_1449, w_309_1460, w_309_1463, w_309_1502, w_309_1521, w_309_1523, w_309_1528, w_309_1529, w_309_1530, w_309_1556, w_309_1560, w_309_1575, w_309_1578, w_309_1579, w_309_1583, w_309_1606, w_309_1612, w_309_1625, w_309_1639, w_309_1672, w_309_1689, w_309_1699, w_309_1715, w_309_1730, w_309_1751, w_309_1753, w_309_1757, w_309_1777, w_309_1784, w_309_1785, w_309_1796, w_309_1800, w_309_1806, w_309_1812, w_309_1819, w_309_1824, w_309_1840, w_309_1841, w_309_1849, w_309_1858, w_309_1865, w_309_1872, w_309_1888, w_309_1896, w_309_1910, w_309_1911, w_309_1914, w_309_1920, w_309_1921, w_309_1928, w_309_1936, w_309_1941, w_309_1949;
  wire w_310_001, w_310_004, w_310_005, w_310_008, w_310_009, w_310_010, w_310_011, w_310_012, w_310_013, w_310_014, w_310_015, w_310_016, w_310_017, w_310_018, w_310_019, w_310_020, w_310_021, w_310_022, w_310_023, w_310_024, w_310_025, w_310_026, w_310_027, w_310_028, w_310_032, w_310_033, w_310_037, w_310_040, w_310_041, w_310_044, w_310_045, w_310_046, w_310_047, w_310_048, w_310_049, w_310_051, w_310_053, w_310_054, w_310_055, w_310_056, w_310_057, w_310_059, w_310_061, w_310_062, w_310_063, w_310_064, w_310_065, w_310_066, w_310_067, w_310_068, w_310_070, w_310_071, w_310_072, w_310_074, w_310_075, w_310_076, w_310_077, w_310_079, w_310_080, w_310_082, w_310_083, w_310_084, w_310_085, w_310_088, w_310_089, w_310_093, w_310_094, w_310_095, w_310_098, w_310_099, w_310_100, w_310_101, w_310_102, w_310_103, w_310_104, w_310_105, w_310_106, w_310_108, w_310_109, w_310_110, w_310_111, w_310_112, w_310_114, w_310_115, w_310_116, w_310_117, w_310_119, w_310_120, w_310_121, w_310_122, w_310_123, w_310_124, w_310_126, w_310_127, w_310_129, w_310_130, w_310_132, w_310_133, w_310_134, w_310_136, w_310_137, w_310_138, w_310_139, w_310_140, w_310_141, w_310_143, w_310_144, w_310_146, w_310_147, w_310_148, w_310_150, w_310_153, w_310_154, w_310_155, w_310_156, w_310_157, w_310_158, w_310_160, w_310_161, w_310_162, w_310_163, w_310_164, w_310_165, w_310_170, w_310_171, w_310_174, w_310_175, w_310_176, w_310_178, w_310_179, w_310_180, w_310_181, w_310_182, w_310_183, w_310_184, w_310_186, w_310_187, w_310_188, w_310_191, w_310_192, w_310_193, w_310_194, w_310_198, w_310_199, w_310_200, w_310_201, w_310_202, w_310_203, w_310_205, w_310_206, w_310_207, w_310_208, w_310_209, w_310_210, w_310_211, w_310_212, w_310_213, w_310_214, w_310_215, w_310_216, w_310_217, w_310_218, w_310_219, w_310_220, w_310_221, w_310_222, w_310_223, w_310_225, w_310_226, w_310_228, w_310_229, w_310_230, w_310_231, w_310_232, w_310_233, w_310_234, w_310_235, w_310_236, w_310_237, w_310_239, w_310_241, w_310_242, w_310_243, w_310_244, w_310_245, w_310_246, w_310_247, w_310_248, w_310_250, w_310_251;
  wire w_311_005, w_311_008, w_311_009, w_311_011, w_311_021, w_311_036, w_311_041, w_311_055, w_311_061, w_311_073, w_311_079, w_311_094, w_311_114, w_311_117, w_311_121, w_311_129, w_311_144, w_311_153, w_311_159, w_311_165, w_311_180, w_311_192, w_311_195, w_311_196, w_311_200, w_311_203, w_311_220, w_311_236, w_311_239, w_311_243, w_311_248, w_311_254, w_311_257, w_311_271, w_311_276, w_311_278, w_311_281, w_311_285, w_311_288, w_311_304, w_311_312, w_311_317, w_311_328, w_311_329, w_311_336, w_311_337, w_311_344, w_311_345, w_311_349, w_311_361, w_311_364, w_311_372, w_311_373, w_311_383, w_311_384, w_311_403, w_311_406, w_311_419, w_311_420, w_311_425, w_311_426, w_311_430, w_311_433, w_311_447, w_311_455, w_311_458, w_311_470, w_311_474, w_311_483, w_311_487, w_311_507, w_311_527, w_311_530, w_311_533, w_311_538, w_311_549, w_311_550, w_311_554, w_311_575, w_311_576, w_311_578, w_311_583, w_311_588, w_311_599, w_311_603, w_311_604, w_311_606, w_311_612, w_311_613, w_311_628, w_311_632, w_311_634, w_311_644, w_311_654, w_311_660, w_311_681, w_311_690, w_311_691, w_311_701, w_311_707, w_311_710, w_311_738, w_311_766, w_311_775, w_311_776, w_311_794, w_311_799, w_311_803, w_311_807, w_311_813, w_311_825, w_311_826, w_311_827, w_311_832, w_311_834, w_311_842, w_311_846, w_311_850, w_311_857, w_311_874, w_311_882, w_311_897, w_311_926, w_311_939, w_311_942, w_311_965, w_311_984, w_311_985, w_311_994, w_311_1000, w_311_1020, w_311_1022, w_311_1032, w_311_1049, w_311_1062, w_311_1066, w_311_1072, w_311_1082, w_311_1085, w_311_1103, w_311_1107, w_311_1118, w_311_1131, w_311_1136, w_311_1139, w_311_1149, w_311_1150, w_311_1152, w_311_1164, w_311_1194, w_311_1201, w_311_1205, w_311_1208, w_311_1211, w_311_1218, w_311_1236, w_311_1274, w_311_1280, w_311_1282, w_311_1295, w_311_1324, w_311_1348, w_311_1415, w_311_1441, w_311_1444, w_311_1489, w_311_1497, w_311_1500, w_311_1501, w_311_1525, w_311_1536, w_311_1544, w_311_1573, w_311_1576, w_311_1589, w_311_1596, w_311_1606, w_311_1610, w_311_1618, w_311_1627, w_311_1630, w_311_1636, w_311_1654, w_311_1673, w_311_1731, w_311_1735, w_311_1737, w_311_1741, w_311_1760, w_311_1782, w_311_1790, w_311_1791, w_311_1798, w_311_1801, w_311_1855, w_311_1865, w_311_1879, w_311_1927, w_311_1954, w_311_1972, w_311_1974, w_311_1994, w_311_1998, w_311_2023, w_311_2033, w_311_2037, w_311_2056, w_311_2065, w_311_2075, w_311_2078, w_311_2104, w_311_2128, w_311_2137, w_311_2138, w_311_2156, w_311_2162, w_311_2184, w_311_2214, w_311_2216, w_311_2229, w_311_2257, w_311_2286, w_311_2298, w_311_2326, w_311_2330, w_311_2348, w_311_2360, w_311_2365, w_311_2392, w_311_2401, w_311_2424, w_311_2438, w_311_2456, w_311_2463, w_311_2482, w_311_2504, w_311_2508, w_311_2510, w_311_2535, w_311_2542, w_311_2546, w_311_2560, w_311_2588, w_311_2635, w_311_2674, w_311_2680, w_311_2681, w_311_2696, w_311_2717, w_311_2718, w_311_2722, w_311_2731, w_311_2760, w_311_2774, w_311_2804, w_311_2825, w_311_2830, w_311_2843, w_311_2856, w_311_2864, w_311_2870, w_311_2885, w_311_2910, w_311_2921, w_311_2929, w_311_2947, w_311_2969, w_311_3020, w_311_3030, w_311_3032, w_311_3046, w_311_3080, w_311_3108, w_311_3122, w_311_3126, w_311_3131, w_311_3142, w_311_3157, w_311_3167, w_311_3174, w_311_3190, w_311_3192, w_311_3214, w_311_3218, w_311_3237, w_311_3257, w_311_3283, w_311_3320, w_311_3340, w_311_3342, w_311_3355, w_311_3359, w_311_3383, w_311_3390, w_311_3403, w_311_3420, w_311_3423, w_311_3454, w_311_3462, w_311_3474, w_311_3476, w_311_3480, w_311_3514, w_311_3534, w_311_3545, w_311_3560, w_311_3562, w_311_3583, w_311_3600, w_311_3657, w_311_3668, w_311_3669, w_311_3690, w_311_3714, w_311_3723, w_311_3725, w_311_3737, w_311_3754, w_311_3773, w_311_3803, w_311_3811, w_311_3819, w_311_3821, w_311_3830, w_311_3831;
  wire w_312_001, w_312_007, w_312_009, w_312_012, w_312_015, w_312_016, w_312_017, w_312_020, w_312_021, w_312_024, w_312_028, w_312_030, w_312_032, w_312_041, w_312_047, w_312_051, w_312_052, w_312_053, w_312_056, w_312_060, w_312_062, w_312_071, w_312_081, w_312_082, w_312_084, w_312_085, w_312_087, w_312_104, w_312_105, w_312_107, w_312_108, w_312_116, w_312_120, w_312_121, w_312_127, w_312_128, w_312_134, w_312_141, w_312_142, w_312_151, w_312_154, w_312_156, w_312_160, w_312_164, w_312_170, w_312_176, w_312_180, w_312_186, w_312_188, w_312_189, w_312_191, w_312_192, w_312_198, w_312_199, w_312_204, w_312_207, w_312_214, w_312_227, w_312_242, w_312_246, w_312_256, w_312_257, w_312_260, w_312_263, w_312_264, w_312_269, w_312_278, w_312_283, w_312_301, w_312_308, w_312_316, w_312_317, w_312_322, w_312_325, w_312_339, w_312_344, w_312_345, w_312_352, w_312_357, w_312_370, w_312_371, w_312_378, w_312_382, w_312_384, w_312_386, w_312_393, w_312_394, w_312_395, w_312_400, w_312_401, w_312_405, w_312_422, w_312_427, w_312_433, w_312_435, w_312_437, w_312_441, w_312_443, w_312_449, w_312_450, w_312_457, w_312_463, w_312_466, w_312_467, w_312_468, w_312_471, w_312_477, w_312_485, w_312_488, w_312_496, w_312_498, w_312_505, w_312_506, w_312_507, w_312_518, w_312_521, w_312_527, w_312_535, w_312_543, w_312_547, w_312_550, w_312_552, w_312_555, w_312_556, w_312_562, w_312_564, w_312_568, w_312_570, w_312_586, w_312_591, w_312_596, w_312_610, w_312_614, w_312_617, w_312_624, w_312_626, w_312_633, w_312_634, w_312_635, w_312_640, w_312_642, w_312_646, w_312_647, w_312_653, w_312_667, w_312_668, w_312_669, w_312_674, w_312_685, w_312_686, w_312_739, w_312_746, w_312_753, w_312_756, w_312_758, w_312_764, w_312_768, w_312_783, w_312_785, w_312_796, w_312_798, w_312_806, w_312_825, w_312_827, w_312_829, w_312_839, w_312_840, w_312_842, w_312_845, w_312_848, w_312_849, w_312_852, w_312_855, w_312_856, w_312_857, w_312_861, w_312_874, w_312_882, w_312_886, w_312_887, w_312_891, w_312_896, w_312_904, w_312_907, w_312_909, w_312_912, w_312_916, w_312_941, w_312_942, w_312_946, w_312_947, w_312_950, w_312_962, w_312_963, w_312_969, w_312_970, w_312_984, w_312_989, w_312_993, w_312_994, w_312_1001, w_312_1010, w_312_1013, w_312_1017, w_312_1018, w_312_1024, w_312_1027, w_312_1034, w_312_1043, w_312_1049, w_312_1054, w_312_1064, w_312_1069, w_312_1079, w_312_1090, w_312_1092, w_312_1094, w_312_1097, w_312_1101, w_312_1102, w_312_1112, w_312_1118, w_312_1121, w_312_1124, w_312_1126, w_312_1130, w_312_1141, w_312_1153, w_312_1157, w_312_1159, w_312_1160, w_312_1164, w_312_1167, w_312_1168, w_312_1171, w_312_1180, w_312_1183, w_312_1187, w_312_1189, w_312_1190, w_312_1196, w_312_1197, w_312_1202, w_312_1203, w_312_1211, w_312_1213, w_312_1216, w_312_1218, w_312_1228, w_312_1230, w_312_1232, w_312_1233, w_312_1247, w_312_1251, w_312_1258, w_312_1267, w_312_1270, w_312_1272, w_312_1276, w_312_1277, w_312_1282, w_312_1286, w_312_1288, w_312_1289, w_312_1291, w_312_1304, w_312_1312, w_312_1313, w_312_1315, w_312_1322, w_312_1324, w_312_1325, w_312_1326, w_312_1339, w_312_1343, w_312_1345, w_312_1347, w_312_1352, w_312_1357, w_312_1367, w_312_1368, w_312_1374, w_312_1375, w_312_1379, w_312_1380, w_312_1389, w_312_1390, w_312_1391, w_312_1395, w_312_1396, w_312_1402, w_312_1407, w_312_1413, w_312_1419, w_312_1420, w_312_1424, w_312_1426, w_312_1428, w_312_1433, w_312_1434, w_312_1455, w_312_1458, w_312_1465, w_312_1489, w_312_1490, w_312_1494, w_312_1499, w_312_1502, w_312_1503, w_312_1507, w_312_1509, w_312_1516, w_312_1517, w_312_1518, w_312_1533, w_312_1539, w_312_1540, w_312_1561, w_312_1562, w_312_1564, w_312_1581, w_312_1595, w_312_1600, w_312_1603, w_312_1607, w_312_1609;
  wire w_313_001, w_313_005, w_313_007, w_313_016, w_313_028, w_313_030, w_313_047, w_313_048, w_313_092, w_313_093, w_313_100, w_313_142, w_313_157, w_313_158, w_313_160, w_313_165, w_313_171, w_313_173, w_313_175, w_313_183, w_313_185, w_313_195, w_313_201, w_313_203, w_313_218, w_313_221, w_313_241, w_313_245, w_313_249, w_313_252, w_313_256, w_313_260, w_313_268, w_313_269, w_313_289, w_313_297, w_313_310, w_313_322, w_313_328, w_313_329, w_313_330, w_313_331, w_313_332, w_313_335, w_313_343, w_313_349, w_313_353, w_313_357, w_313_371, w_313_380, w_313_392, w_313_404, w_313_411, w_313_417, w_313_422, w_313_424, w_313_434, w_313_470, w_313_475, w_313_486, w_313_501, w_313_504, w_313_505, w_313_519, w_313_525, w_313_527, w_313_550, w_313_563, w_313_564, w_313_570, w_313_591, w_313_595, w_313_611, w_313_620, w_313_622, w_313_628, w_313_653, w_313_681, w_313_702, w_313_723, w_313_726, w_313_754, w_313_765, w_313_784, w_313_819, w_313_826, w_313_835, w_313_840, w_313_861, w_313_883, w_313_890, w_313_894, w_313_914, w_313_920, w_313_931, w_313_950, w_313_959, w_313_989, w_313_990, w_313_993, w_313_994, w_313_1004, w_313_1005, w_313_1013, w_313_1016, w_313_1028, w_313_1031, w_313_1035, w_313_1053, w_313_1084, w_313_1093, w_313_1151, w_313_1167, w_313_1198, w_313_1225, w_313_1264, w_313_1275, w_313_1280, w_313_1284, w_313_1329, w_313_1355, w_313_1413, w_313_1441, w_313_1469, w_313_1479, w_313_1480, w_313_1484, w_313_1502, w_313_1503, w_313_1530, w_313_1577, w_313_1599, w_313_1610, w_313_1611, w_313_1613, w_313_1641, w_313_1663, w_313_1668, w_313_1669, w_313_1670, w_313_1673, w_313_1739, w_313_1760, w_313_1790, w_313_1798, w_313_1808, w_313_1832, w_313_1837, w_313_1847, w_313_1864, w_313_1873, w_313_1902, w_313_1904, w_313_1931, w_313_1933, w_313_1952, w_313_1962, w_313_1968, w_313_2006, w_313_2007, w_313_2044, w_313_2048, w_313_2062, w_313_2107, w_313_2109, w_313_2117, w_313_2122, w_313_2130, w_313_2143, w_313_2151, w_313_2166, w_313_2195, w_313_2197, w_313_2228, w_313_2267, w_313_2277, w_313_2293, w_313_2316, w_313_2347, w_313_2352, w_313_2355, w_313_2359, w_313_2376, w_313_2383, w_313_2393, w_313_2399, w_313_2425, w_313_2433, w_313_2438, w_313_2483, w_313_2492, w_313_2508, w_313_2526, w_313_2536, w_313_2537, w_313_2553, w_313_2569, w_313_2575, w_313_2582, w_313_2584, w_313_2651, w_313_2665, w_313_2669, w_313_2681, w_313_2684, w_313_2687, w_313_2699, w_313_2712, w_313_2718, w_313_2722, w_313_2733, w_313_2782, w_313_2787, w_313_2796, w_313_2797, w_313_2813, w_313_2827, w_313_2828, w_313_2845, w_313_2851, w_313_2858, w_313_2901, w_313_2910, w_313_2922, w_313_2926, w_313_2927, w_313_2955, w_313_3028, w_313_3045, w_313_3051, w_313_3074, w_313_3079, w_313_3093, w_313_3098, w_313_3118, w_313_3144, w_313_3148, w_313_3180, w_313_3211, w_313_3227, w_313_3238, w_313_3241, w_313_3246, w_313_3247, w_313_3257, w_313_3264, w_313_3300, w_313_3325, w_313_3354, w_313_3368, w_313_3384, w_313_3406, w_313_3462, w_313_3471, w_313_3493, w_313_3494, w_313_3545, w_313_3553, w_313_3569, w_313_3576, w_313_3580, w_313_3598, w_313_3601, w_313_3634, w_313_3637, w_313_3638, w_313_3642, w_313_3647, w_313_3730, w_313_3731, w_313_3765, w_313_3788, w_313_3790, w_313_3797, w_313_3802, w_313_3804, w_313_3808, w_313_3814, w_313_3840, w_313_3867, w_313_3886, w_313_3889, w_313_3898, w_313_3926, w_313_3952, w_313_3958, w_313_3967, w_313_3975, w_313_3976, w_313_3997, w_313_4017, w_313_4050, w_313_4063, w_313_4066, w_313_4069, w_313_4087, w_313_4091, w_313_4095, w_313_4098, w_313_4099, w_313_4100, w_313_4102, w_313_4108, w_313_4123, w_313_4126, w_313_4135, w_313_4144, w_313_4148, w_313_4211, w_313_4251, w_313_4252, w_313_4263, w_313_4265, w_313_4295, w_313_4297, w_313_4320, w_313_4322, w_313_4324, w_313_4329, w_313_4375;
  wire w_314_002, w_314_003, w_314_008, w_314_015, w_314_026, w_314_036, w_314_039, w_314_049, w_314_076, w_314_079, w_314_081, w_314_082, w_314_083, w_314_091, w_314_098, w_314_100, w_314_111, w_314_124, w_314_132, w_314_143, w_314_149, w_314_158, w_314_160, w_314_162, w_314_171, w_314_172, w_314_174, w_314_175, w_314_178, w_314_186, w_314_188, w_314_200, w_314_211, w_314_219, w_314_225, w_314_230, w_314_231, w_314_242, w_314_245, w_314_256, w_314_271, w_314_275, w_314_278, w_314_281, w_314_294, w_314_311, w_314_315, w_314_334, w_314_341, w_314_350, w_314_355, w_314_358, w_314_360, w_314_363, w_314_368, w_314_377, w_314_387, w_314_398, w_314_407, w_314_419, w_314_421, w_314_423, w_314_428, w_314_444, w_314_447, w_314_451, w_314_453, w_314_457, w_314_461, w_314_472, w_314_477, w_314_482, w_314_485, w_314_487, w_314_500, w_314_504, w_314_507, w_314_508, w_314_510, w_314_517, w_314_553, w_314_554, w_314_561, w_314_562, w_314_563, w_314_566, w_314_572, w_314_593, w_314_599, w_314_600, w_314_611, w_314_614, w_314_619, w_314_623, w_314_631, w_314_648, w_314_654, w_314_655, w_314_667, w_314_669, w_314_680, w_314_693, w_314_694, w_314_751, w_314_769, w_314_782, w_314_783, w_314_809, w_314_814, w_314_823, w_314_825, w_314_826, w_314_827, w_314_855, w_314_858, w_314_875, w_314_878, w_314_881, w_314_892, w_314_893, w_314_901, w_314_902, w_314_909, w_314_916, w_314_921, w_314_922, w_314_931, w_314_932, w_314_934, w_314_941, w_314_958, w_314_963, w_314_964, w_314_973, w_314_976, w_314_980, w_314_981, w_314_985, w_314_993, w_314_1007, w_314_1029, w_314_1035, w_314_1036, w_314_1046, w_314_1059, w_314_1067, w_314_1068, w_314_1078, w_314_1098, w_314_1109, w_314_1120, w_314_1139, w_314_1154, w_314_1155, w_314_1176, w_314_1178, w_314_1186, w_314_1243, w_314_1249, w_314_1254, w_314_1260, w_314_1261, w_314_1265, w_314_1269, w_314_1271, w_314_1284, w_314_1288, w_314_1298, w_314_1302, w_314_1308, w_314_1319, w_314_1332, w_314_1341, w_314_1342, w_314_1345, w_314_1346, w_314_1371, w_314_1373, w_314_1389, w_314_1390, w_314_1394, w_314_1397, w_314_1407, w_314_1411, w_314_1414, w_314_1416, w_314_1417, w_314_1434, w_314_1451, w_314_1454, w_314_1456, w_314_1457, w_314_1461, w_314_1468, w_314_1476, w_314_1477, w_314_1479, w_314_1480, w_314_1489, w_314_1491, w_314_1501, w_314_1510, w_314_1525, w_314_1534, w_314_1538, w_314_1571, w_314_1623, w_314_1634, w_314_1668, w_314_1692, w_314_1694, w_314_1722, w_314_1745, w_314_1753, w_314_1765, w_314_1768, w_314_1784, w_314_1796, w_314_1835, w_314_1845, w_314_1850, w_314_1858, w_314_1861, w_314_1866, w_314_1867, w_314_1874, w_314_1902, w_314_1914, w_314_1930, w_314_1945, w_314_1958, w_314_1969, w_314_1982, w_314_1996, w_314_2001, w_314_2009, w_314_2064, w_314_2089, w_314_2093, w_314_2113, w_314_2125, w_314_2128, w_314_2133, w_314_2194, w_314_2197, w_314_2214, w_314_2235, w_314_2243, w_314_2270, w_314_2310, w_314_2342, w_314_2361, w_314_2368, w_314_2372, w_314_2374, w_314_2386, w_314_2393, w_314_2428, w_314_2442, w_314_2445, w_314_2475, w_314_2486, w_314_2492, w_314_2497, w_314_2537, w_314_2541, w_314_2544, w_314_2548, w_314_2561, w_314_2562, w_314_2564, w_314_2566, w_314_2570, w_314_2581, w_314_2592, w_314_2594, w_314_2605, w_314_2633, w_314_2657, w_314_2670, w_314_2672, w_314_2677, w_314_2680, w_314_2684, w_314_2700, w_314_2713, w_314_2733, w_314_2736, w_314_2739, w_314_2756, w_314_2758, w_314_2762, w_314_2765, w_314_2777, w_314_2782, w_314_2804, w_314_2857, w_314_2860, w_314_2869, w_314_2891, w_314_2909, w_314_2919, w_314_2940, w_314_2941, w_314_2951, w_314_3011, w_314_3014, w_314_3039, w_314_3048, w_314_3053, w_314_3058, w_314_3061, w_314_3077, w_314_3085, w_314_3115, w_314_3125, w_314_3135, w_314_3168, w_314_3169, w_314_3223, w_314_3257, w_314_3260, w_314_3275, w_314_3289, w_314_3295, w_314_3317, w_314_3331, w_314_3339, w_314_3340, w_314_3377, w_314_3381, w_314_3406, w_314_3420, w_314_3439;
  wire w_315_007, w_315_010, w_315_025, w_315_029, w_315_034, w_315_039, w_315_041, w_315_044, w_315_063, w_315_075, w_315_083, w_315_085, w_315_096, w_315_103, w_315_111, w_315_115, w_315_137, w_315_154, w_315_155, w_315_164, w_315_190, w_315_193, w_315_198, w_315_206, w_315_211, w_315_215, w_315_216, w_315_219, w_315_226, w_315_233, w_315_258, w_315_260, w_315_285, w_315_292, w_315_297, w_315_303, w_315_306, w_315_312, w_315_324, w_315_330, w_315_338, w_315_343, w_315_392, w_315_394, w_315_399, w_315_412, w_315_417, w_315_425, w_315_441, w_315_496, w_315_498, w_315_541, w_315_549, w_315_574, w_315_575, w_315_577, w_315_591, w_315_618, w_315_654, w_315_669, w_315_729, w_315_739, w_315_745, w_315_762, w_315_781, w_315_783, w_315_811, w_315_815, w_315_818, w_315_862, w_315_867, w_315_868, w_315_871, w_315_875, w_315_880, w_315_881, w_315_907, w_315_915, w_315_927, w_315_940, w_315_955, w_315_973, w_315_1004, w_315_1010, w_315_1015, w_315_1027, w_315_1039, w_315_1053, w_315_1082, w_315_1110, w_315_1123, w_315_1124, w_315_1135, w_315_1147, w_315_1150, w_315_1182, w_315_1188, w_315_1205, w_315_1214, w_315_1243, w_315_1289, w_315_1304, w_315_1317, w_315_1327, w_315_1333, w_315_1349, w_315_1363, w_315_1387, w_315_1388, w_315_1389, w_315_1446, w_315_1456, w_315_1476, w_315_1480, w_315_1490, w_315_1505, w_315_1531, w_315_1540, w_315_1566, w_315_1589, w_315_1627, w_315_1651, w_315_1710, w_315_1730, w_315_1737, w_315_1754, w_315_1759, w_315_1806, w_315_1827, w_315_1831, w_315_1856, w_315_1885, w_315_1897, w_315_1924, w_315_1936, w_315_1949, w_315_1991, w_315_2007, w_315_2018, w_315_2028, w_315_2062, w_315_2077, w_315_2108, w_315_2112, w_315_2114, w_315_2124, w_315_2131, w_315_2179, w_315_2207, w_315_2211, w_315_2222, w_315_2234, w_315_2246, w_315_2260, w_315_2316, w_315_2327, w_315_2331, w_315_2362, w_315_2367, w_315_2385, w_315_2394, w_315_2399, w_315_2415, w_315_2430, w_315_2461, w_315_2467, w_315_2481, w_315_2484, w_315_2497, w_315_2498, w_315_2502, w_315_2515, w_315_2550, w_315_2552, w_315_2561, w_315_2562, w_315_2569, w_315_2587, w_315_2590, w_315_2624, w_315_2639, w_315_2653, w_315_2661, w_315_2718, w_315_2727, w_315_2730, w_315_2756, w_315_2778, w_315_2815, w_315_2827, w_315_2836, w_315_2865, w_315_2886, w_315_2889, w_315_2935, w_315_2939, w_315_2950, w_315_2956, w_315_3000, w_315_3001, w_315_3015, w_315_3030, w_315_3040, w_315_3048, w_315_3059, w_315_3066, w_315_3069, w_315_3114, w_315_3124, w_315_3141, w_315_3146, w_315_3149, w_315_3158, w_315_3189, w_315_3247, w_315_3286, w_315_3295, w_315_3366, w_315_3445, w_315_3455, w_315_3461, w_315_3489, w_315_3530, w_315_3533, w_315_3546, w_315_3568, w_315_3575, w_315_3579, w_315_3580, w_315_3611, w_315_3618, w_315_3629, w_315_3631, w_315_3632, w_315_3644, w_315_3666, w_315_3714, w_315_3718, w_315_3719, w_315_3730, w_315_3769, w_315_3773, w_315_3777, w_315_3778, w_315_3785, w_315_3790, w_315_3853, w_315_3855, w_315_3874, w_315_3908, w_315_3940, w_315_3949, w_315_3954, w_315_3994, w_315_4004, w_315_4018, w_315_4036, w_315_4047, w_315_4070, w_315_4116, w_315_4126, w_315_4162, w_315_4163, w_315_4166, w_315_4171, w_315_4176, w_315_4178, w_315_4193, w_315_4197, w_315_4198, w_315_4213, w_315_4237, w_315_4272, w_315_4274, w_315_4295, w_315_4296, w_315_4338, w_315_4369, w_315_4377, w_315_4384, w_315_4387, w_315_4405, w_315_4446, w_315_4450, w_315_4475, w_315_4547, w_315_4555, w_315_4557, w_315_4580, w_315_4624;
  wire w_316_003, w_316_007, w_316_009, w_316_010, w_316_011, w_316_013, w_316_014, w_316_016, w_316_017, w_316_021, w_316_024, w_316_025, w_316_027, w_316_028, w_316_036, w_316_037, w_316_041, w_316_044, w_316_045, w_316_051, w_316_052, w_316_053, w_316_055, w_316_056, w_316_057, w_316_058, w_316_059, w_316_061, w_316_063, w_316_064, w_316_066, w_316_067, w_316_075, w_316_079, w_316_082, w_316_083, w_316_089, w_316_091, w_316_093, w_316_097, w_316_098, w_316_099, w_316_100, w_316_103, w_316_105, w_316_112, w_316_116, w_316_120, w_316_124, w_316_127, w_316_129, w_316_131, w_316_132, w_316_133, w_316_136, w_316_138, w_316_139, w_316_141, w_316_143, w_316_144, w_316_153, w_316_155, w_316_157, w_316_160, w_316_162, w_316_163, w_316_167, w_316_169, w_316_171, w_316_175, w_316_180, w_316_182, w_316_183, w_316_186, w_316_187, w_316_188, w_316_193, w_316_194, w_316_196, w_316_198, w_316_200, w_316_204, w_316_206, w_316_209, w_316_211, w_316_213, w_316_214, w_316_223, w_316_226, w_316_230, w_316_234, w_316_235, w_316_236, w_316_237, w_316_239, w_316_241, w_316_243, w_316_249, w_316_250, w_316_251, w_316_255, w_316_256, w_316_257, w_316_259, w_316_261, w_316_264, w_316_265, w_316_274, w_316_278, w_316_286, w_316_288, w_316_289, w_316_290, w_316_291, w_316_292, w_316_293, w_316_297, w_316_299, w_316_304, w_316_309, w_316_310, w_316_311, w_316_312, w_316_315, w_316_318, w_316_323, w_316_324, w_316_327, w_316_331, w_316_343, w_316_344, w_316_352, w_316_353, w_316_355, w_316_356, w_316_359, w_316_365, w_316_368, w_316_369, w_316_371, w_316_377, w_316_380, w_316_381, w_316_382, w_316_385, w_316_388, w_316_389, w_316_390, w_316_391, w_316_393, w_316_394, w_316_396, w_316_400, w_316_403, w_316_406, w_316_409, w_316_417, w_316_419, w_316_423, w_316_426, w_316_430, w_316_432, w_316_433, w_316_434, w_316_441, w_316_446, w_316_447, w_316_449, w_316_452, w_316_456, w_316_462, w_316_463, w_316_464, w_316_465, w_316_471, w_316_472, w_316_474, w_316_476, w_316_480, w_316_482, w_316_484, w_316_486, w_316_489, w_316_491, w_316_495, w_316_496, w_316_498, w_316_499, w_316_503, w_316_505, w_316_509, w_316_510, w_316_514, w_316_517, w_316_518, w_316_526, w_316_528, w_316_530, w_316_535, w_316_536, w_316_538, w_316_543, w_316_547, w_316_549, w_316_550, w_316_551, w_316_554, w_316_555, w_316_558, w_316_561, w_316_567, w_316_572, w_316_580, w_316_581, w_316_583, w_316_584, w_316_586, w_316_587, w_316_590, w_316_591, w_316_592, w_316_593, w_316_595, w_316_596, w_316_597, w_316_600, w_316_601, w_316_602, w_316_603, w_316_604, w_316_605, w_316_607, w_316_609, w_316_612, w_316_613, w_316_616, w_316_617, w_316_618, w_316_622, w_316_623, w_316_624, w_316_625, w_316_631, w_316_632, w_316_633, w_316_641, w_316_642, w_316_645, w_316_647, w_316_652, w_316_655, w_316_656, w_316_658, w_316_663, w_316_671, w_316_673, w_316_681, w_316_682, w_316_684, w_316_685, w_316_689, w_316_691, w_316_692, w_316_693, w_316_694, w_316_700, w_316_701, w_316_709, w_316_712, w_316_713, w_316_716, w_316_717, w_316_718;
  wire w_317_010, w_317_019, w_317_024, w_317_029, w_317_031, w_317_034, w_317_038, w_317_039, w_317_061, w_317_066, w_317_088, w_317_109, w_317_121, w_317_122, w_317_124, w_317_128, w_317_131, w_317_134, w_317_135, w_317_139, w_317_142, w_317_155, w_317_157, w_317_166, w_317_167, w_317_169, w_317_171, w_317_183, w_317_189, w_317_193, w_317_208, w_317_217, w_317_223, w_317_224, w_317_230, w_317_232, w_317_235, w_317_236, w_317_244, w_317_246, w_317_254, w_317_256, w_317_258, w_317_259, w_317_263, w_317_264, w_317_269, w_317_271, w_317_273, w_317_280, w_317_287, w_317_295, w_317_318, w_317_326, w_317_329, w_317_334, w_317_336, w_317_337, w_317_340, w_317_345, w_317_360, w_317_362, w_317_369, w_317_373, w_317_374, w_317_384, w_317_396, w_317_403, w_317_404, w_317_410, w_317_420, w_317_422, w_317_426, w_317_432, w_317_434, w_317_446, w_317_449, w_317_452, w_317_455, w_317_460, w_317_462, w_317_467, w_317_469, w_317_470, w_317_476, w_317_485, w_317_488, w_317_492, w_317_500, w_317_508, w_317_509, w_317_514, w_317_520, w_317_521, w_317_524, w_317_535, w_317_539, w_317_543, w_317_552, w_317_555, w_317_560, w_317_565, w_317_570, w_317_571, w_317_583, w_317_599, w_317_608, w_317_609, w_317_616, w_317_621, w_317_622, w_317_623, w_317_633, w_317_635, w_317_636, w_317_648, w_317_651, w_317_654, w_317_655, w_317_668, w_317_669, w_317_672, w_317_675, w_317_681, w_317_690, w_317_701, w_317_702, w_317_705, w_317_710, w_317_719, w_317_723, w_317_724, w_317_731, w_317_734, w_317_735, w_317_739, w_317_743, w_317_744, w_317_745, w_317_748, w_317_749, w_317_750, w_317_754, w_317_755, w_317_756, w_317_759, w_317_767, w_317_771, w_317_789, w_317_791, w_317_807, w_317_808, w_317_814, w_317_815, w_317_817, w_317_831, w_317_838, w_317_840, w_317_841, w_317_842, w_317_848, w_317_850, w_317_851, w_317_861, w_317_864, w_317_867, w_317_872, w_317_873, w_317_881, w_317_883, w_317_887, w_317_891, w_317_898, w_317_903, w_317_909, w_317_919, w_317_922, w_317_925, w_317_937, w_317_943, w_317_944, w_317_946, w_317_948, w_317_957, w_317_961, w_317_967, w_317_972, w_317_977, w_317_980, w_317_981, w_317_986, w_317_992, w_317_1007, w_317_1011, w_317_1012, w_317_1036, w_317_1038, w_317_1039, w_317_1040, w_317_1048, w_317_1051, w_317_1056, w_317_1071, w_317_1075, w_317_1084, w_317_1085, w_317_1086, w_317_1087, w_317_1094, w_317_1103, w_317_1105, w_317_1129, w_317_1130, w_317_1131, w_317_1136, w_317_1137, w_317_1138, w_317_1140, w_317_1143, w_317_1144, w_317_1149, w_317_1157, w_317_1158, w_317_1161, w_317_1165, w_317_1172, w_317_1184, w_317_1185, w_317_1197, w_317_1212, w_317_1214, w_317_1220, w_317_1227, w_317_1231, w_317_1234, w_317_1239, w_317_1256, w_317_1260, w_317_1263, w_317_1265, w_317_1266, w_317_1275, w_317_1277, w_317_1281, w_317_1290, w_317_1292, w_317_1293, w_317_1309, w_317_1313, w_317_1318, w_317_1330, w_317_1345, w_317_1346, w_317_1358, w_317_1376, w_317_1379, w_317_1388, w_317_1389, w_317_1401, w_317_1402, w_317_1407, w_317_1426, w_317_1430, w_317_1431, w_317_1460, w_317_1462, w_317_1468, w_317_1479, w_317_1486, w_317_1493, w_317_1511, w_317_1517, w_317_1521, w_317_1523, w_317_1524, w_317_1527, w_317_1535, w_317_1552, w_317_1566, w_317_1568, w_317_1571, w_317_1577, w_317_1579, w_317_1583, w_317_1586, w_317_1596, w_317_1599, w_317_1600, w_317_1608, w_317_1615, w_317_1617, w_317_1626, w_317_1631, w_317_1640, w_317_1645, w_317_1664, w_317_1668, w_317_1673, w_317_1674, w_317_1685, w_317_1686, w_317_1696, w_317_1700, w_317_1706, w_317_1709, w_317_1721, w_317_1725, w_317_1728, w_317_1730, w_317_1733, w_317_1742, w_317_1748, w_317_1761, w_317_1787, w_317_1796, w_317_1803, w_317_1804, w_317_1828, w_317_1829, w_317_1833, w_317_1835, w_317_1837, w_317_1862, w_317_1863, w_317_1889, w_317_1891, w_317_1893, w_317_1903, w_317_1912, w_317_1917, w_317_1934, w_317_1957, w_317_1958, w_317_1959, w_317_1968, w_317_1972, w_317_1988, w_317_1990, w_317_1991, w_317_1992;
  wire w_318_002, w_318_007, w_318_008, w_318_009, w_318_010, w_318_013, w_318_015, w_318_018, w_318_019, w_318_022, w_318_033, w_318_039, w_318_043, w_318_044, w_318_045, w_318_046, w_318_049, w_318_050, w_318_055, w_318_057, w_318_065, w_318_066, w_318_067, w_318_068, w_318_072, w_318_074, w_318_080, w_318_082, w_318_085, w_318_086, w_318_088, w_318_094, w_318_096, w_318_102, w_318_103, w_318_104, w_318_109, w_318_112, w_318_115, w_318_116, w_318_118, w_318_119, w_318_121, w_318_122, w_318_124, w_318_127, w_318_132, w_318_134, w_318_137, w_318_138, w_318_140, w_318_142, w_318_149, w_318_154, w_318_158, w_318_163, w_318_165, w_318_167, w_318_171, w_318_172, w_318_174, w_318_178, w_318_185, w_318_186, w_318_189, w_318_193, w_318_196, w_318_197, w_318_198, w_318_201, w_318_202, w_318_203, w_318_205, w_318_208, w_318_210, w_318_222, w_318_234, w_318_236, w_318_238, w_318_244, w_318_246, w_318_249, w_318_251, w_318_260, w_318_261, w_318_265, w_318_266, w_318_271, w_318_279, w_318_281, w_318_282, w_318_300, w_318_306, w_318_308, w_318_311, w_318_312, w_318_315, w_318_316, w_318_321, w_318_322, w_318_324, w_318_326, w_318_331, w_318_332, w_318_333, w_318_341, w_318_344, w_318_345, w_318_359, w_318_361, w_318_364, w_318_366, w_318_367, w_318_369, w_318_371, w_318_372, w_318_381, w_318_391, w_318_396, w_318_401, w_318_407, w_318_413, w_318_416, w_318_418, w_318_422, w_318_425, w_318_436, w_318_442, w_318_448, w_318_449, w_318_460, w_318_467, w_318_468, w_318_472, w_318_474, w_318_475, w_318_482, w_318_492, w_318_499, w_318_508, w_318_512, w_318_515, w_318_520, w_318_527, w_318_533, w_318_534, w_318_535, w_318_540, w_318_541, w_318_544, w_318_555, w_318_558, w_318_564, w_318_569, w_318_571, w_318_572, w_318_576, w_318_584, w_318_588, w_318_593, w_318_596, w_318_597, w_318_608, w_318_609, w_318_613, w_318_619, w_318_628, w_318_632, w_318_637, w_318_640, w_318_644, w_318_650, w_318_651, w_318_654, w_318_659, w_318_661, w_318_662, w_318_664, w_318_666, w_318_667, w_318_674, w_318_677, w_318_678, w_318_682, w_318_685, w_318_695, w_318_708, w_318_713, w_318_722, w_318_728, w_318_738, w_318_739, w_318_740, w_318_742, w_318_745, w_318_750, w_318_754, w_318_755, w_318_756, w_318_759, w_318_760, w_318_762, w_318_765, w_318_769, w_318_775, w_318_776, w_318_785, w_318_786, w_318_787, w_318_791, w_318_794, w_318_796, w_318_797, w_318_800, w_318_802, w_318_805, w_318_809, w_318_813, w_318_814, w_318_823, w_318_825, w_318_828, w_318_830, w_318_839, w_318_842, w_318_844, w_318_846, w_318_850, w_318_852, w_318_857, w_318_865, w_318_868, w_318_869, w_318_871, w_318_872, w_318_873, w_318_874, w_318_877, w_318_881, w_318_888, w_318_889, w_318_894, w_318_899, w_318_901, w_318_903, w_318_904, w_318_905, w_318_919, w_318_925, w_318_932, w_318_934, w_318_940, w_318_945, w_318_947, w_318_952, w_318_957, w_318_961, w_318_962, w_318_963, w_318_964, w_318_965, w_318_969, w_318_973, w_318_978, w_318_981, w_318_985, w_318_993, w_318_1000, w_318_1001, w_318_1008, w_318_1010, w_318_1014, w_318_1021, w_318_1024, w_318_1027, w_318_1035, w_318_1040, w_318_1050, w_318_1063, w_318_1064, w_318_1066, w_318_1068, w_318_1074, w_318_1081, w_318_1082, w_318_1090, w_318_1091, w_318_1092, w_318_1096, w_318_1098, w_318_1114, w_318_1115, w_318_1120, w_318_1123, w_318_1124, w_318_1136, w_318_1139, w_318_1141, w_318_1155, w_318_1172, w_318_1182, w_318_1183, w_318_1184, w_318_1187;
  wire w_319_000, w_319_002, w_319_008, w_319_019, w_319_023, w_319_025, w_319_032, w_319_039, w_319_042, w_319_047, w_319_055, w_319_056, w_319_057, w_319_058, w_319_059, w_319_060, w_319_061, w_319_063, w_319_068, w_319_069, w_319_073, w_319_078, w_319_080, w_319_087, w_319_092, w_319_104, w_319_132, w_319_135, w_319_136, w_319_147, w_319_148, w_319_150, w_319_159, w_319_164, w_319_165, w_319_166, w_319_172, w_319_177, w_319_183, w_319_184, w_319_190, w_319_194, w_319_205, w_319_209, w_319_215, w_319_223, w_319_225, w_319_226, w_319_227, w_319_229, w_319_231, w_319_232, w_319_234, w_319_235, w_319_236, w_319_240, w_319_241, w_319_245, w_319_246, w_319_251, w_319_255, w_319_256, w_319_263, w_319_264, w_319_266, w_319_269, w_319_272, w_319_287, w_319_290, w_319_296, w_319_302, w_319_306, w_319_309, w_319_320, w_319_326, w_319_328, w_319_330, w_319_338, w_319_340, w_319_354, w_319_356, w_319_360, w_319_362, w_319_365, w_319_366, w_319_379, w_319_386, w_319_395, w_319_402, w_319_409, w_319_412, w_319_413, w_319_414, w_319_415, w_319_419, w_319_422, w_319_424, w_319_425, w_319_429, w_319_438, w_319_444, w_319_447, w_319_456, w_319_465, w_319_468, w_319_469, w_319_472, w_319_476, w_319_479, w_319_488, w_319_508, w_319_518, w_319_521, w_319_523, w_319_528, w_319_534, w_319_536, w_319_547, w_319_550, w_319_552, w_319_553, w_319_557, w_319_559, w_319_561, w_319_564, w_319_571, w_319_578, w_319_584, w_319_589, w_319_590, w_319_591, w_319_593, w_319_611, w_319_619, w_319_621, w_319_625, w_319_629, w_319_632, w_319_634, w_319_639, w_319_641, w_319_650, w_319_655, w_319_658, w_319_669, w_319_677, w_319_682, w_319_687, w_319_689, w_319_690, w_319_709, w_319_710, w_319_720, w_319_725, w_319_727, w_319_730, w_319_732, w_319_733, w_319_738, w_319_743, w_319_758, w_319_760, w_319_764, w_319_769, w_319_771, w_319_775, w_319_780, w_319_787, w_319_788, w_319_791, w_319_796, w_319_799, w_319_804, w_319_806, w_319_821, w_319_823, w_319_825, w_319_829, w_319_835, w_319_836, w_319_839, w_319_848, w_319_851, w_319_852, w_319_858, w_319_862, w_319_875, w_319_880, w_319_885, w_319_889, w_319_897, w_319_902, w_319_923, w_319_933, w_319_936, w_319_938, w_319_939, w_319_940, w_319_942, w_319_948, w_319_949, w_319_957, w_319_960, w_319_962, w_319_964, w_319_969, w_319_979, w_319_989, w_319_992, w_319_996, w_319_998, w_319_1001, w_319_1009, w_319_1017, w_319_1026, w_319_1028, w_319_1037, w_319_1038, w_319_1040, w_319_1042, w_319_1043, w_319_1047, w_319_1051, w_319_1056, w_319_1065, w_319_1069, w_319_1071, w_319_1089, w_319_1101, w_319_1117, w_319_1122, w_319_1124, w_319_1125, w_319_1129, w_319_1135, w_319_1144, w_319_1148, w_319_1150, w_319_1152, w_319_1154, w_319_1159, w_319_1162, w_319_1169, w_319_1171, w_319_1177, w_319_1187, w_319_1193, w_319_1207, w_319_1212, w_319_1216, w_319_1222, w_319_1240, w_319_1242, w_319_1261, w_319_1264, w_319_1270, w_319_1276, w_319_1282, w_319_1283, w_319_1284, w_319_1285, w_319_1299, w_319_1303, w_319_1304, w_319_1307, w_319_1312, w_319_1314, w_319_1315, w_319_1318, w_319_1320, w_319_1321, w_319_1324, w_319_1326, w_319_1329, w_319_1332, w_319_1336, w_319_1345, w_319_1347, w_319_1353, w_319_1355, w_319_1356, w_319_1369, w_319_1382, w_319_1397, w_319_1405, w_319_1410, w_319_1412, w_319_1413, w_319_1415, w_319_1418, w_319_1423, w_319_1424, w_319_1426, w_319_1427, w_319_1428, w_319_1429, w_319_1433, w_319_1434, w_319_1442, w_319_1443, w_319_1455, w_319_1461, w_319_1463, w_319_1465, w_319_1471, w_319_1472, w_319_1473, w_319_1475, w_319_1481, w_319_1483, w_319_1486, w_319_1492, w_319_1499, w_319_1525, w_319_1526, w_319_1535, w_319_1543, w_319_1548, w_319_1553, w_319_1567, w_319_1572, w_319_1574, w_319_1576;
  wire w_320_001, w_320_005, w_320_008, w_320_013, w_320_016, w_320_018, w_320_025, w_320_033, w_320_038, w_320_039, w_320_050, w_320_053, w_320_063, w_320_070, w_320_078, w_320_096, w_320_098, w_320_107, w_320_119, w_320_120, w_320_122, w_320_128, w_320_132, w_320_142, w_320_144, w_320_147, w_320_149, w_320_152, w_320_153, w_320_166, w_320_175, w_320_187, w_320_188, w_320_195, w_320_197, w_320_228, w_320_230, w_320_236, w_320_237, w_320_238, w_320_239, w_320_242, w_320_245, w_320_255, w_320_257, w_320_258, w_320_260, w_320_262, w_320_268, w_320_273, w_320_276, w_320_278, w_320_289, w_320_290, w_320_292, w_320_309, w_320_314, w_320_324, w_320_327, w_320_336, w_320_338, w_320_340, w_320_348, w_320_367, w_320_376, w_320_382, w_320_388, w_320_392, w_320_398, w_320_399, w_320_404, w_320_414, w_320_415, w_320_418, w_320_421, w_320_429, w_320_430, w_320_440, w_320_444, w_320_473, w_320_475, w_320_476, w_320_477, w_320_478, w_320_484, w_320_489, w_320_494, w_320_496, w_320_505, w_320_517, w_320_520, w_320_522, w_320_529, w_320_544, w_320_565, w_320_585, w_320_586, w_320_587, w_320_595, w_320_615, w_320_627, w_320_649, w_320_653, w_320_670, w_320_673, w_320_686, w_320_694, w_320_695, w_320_702, w_320_713, w_320_714, w_320_716, w_320_717, w_320_721, w_320_748, w_320_749, w_320_751, w_320_757, w_320_760, w_320_761, w_320_767, w_320_769, w_320_778, w_320_781, w_320_791, w_320_796, w_320_798, w_320_801, w_320_814, w_320_817, w_320_834, w_320_836, w_320_840, w_320_845, w_320_848, w_320_852, w_320_855, w_320_861, w_320_868, w_320_869, w_320_871, w_320_877, w_320_906, w_320_907, w_320_911, w_320_913, w_320_917, w_320_925, w_320_928, w_320_935, w_320_937, w_320_955, w_320_961, w_320_964, w_320_983, w_320_998, w_320_1010, w_320_1024, w_320_1035, w_320_1036, w_320_1039, w_320_1052, w_320_1062, w_320_1069, w_320_1079, w_320_1091, w_320_1094, w_320_1112, w_320_1115, w_320_1122, w_320_1123, w_320_1149, w_320_1157, w_320_1158, w_320_1162, w_320_1168, w_320_1169, w_320_1190, w_320_1192, w_320_1196, w_320_1208, w_320_1214, w_320_1234, w_320_1238, w_320_1239, w_320_1240, w_320_1247, w_320_1248, w_320_1255, w_320_1257, w_320_1263, w_320_1266, w_320_1270, w_320_1273, w_320_1275, w_320_1277, w_320_1299, w_320_1300, w_320_1303, w_320_1337, w_320_1346, w_320_1356, w_320_1360, w_320_1364, w_320_1372, w_320_1387, w_320_1388, w_320_1392, w_320_1399, w_320_1408, w_320_1410, w_320_1439, w_320_1451, w_320_1466, w_320_1467, w_320_1470, w_320_1471, w_320_1472, w_320_1496, w_320_1500, w_320_1506, w_320_1508, w_320_1516, w_320_1520, w_320_1541, w_320_1581, w_320_1582, w_320_1589, w_320_1591, w_320_1599, w_320_1602, w_320_1615, w_320_1617, w_320_1623, w_320_1630, w_320_1632, w_320_1633, w_320_1634, w_320_1637, w_320_1639, w_320_1641, w_320_1645, w_320_1650, w_320_1654, w_320_1667, w_320_1680, w_320_1683, w_320_1687, w_320_1692, w_320_1696, w_320_1710, w_320_1711, w_320_1719, w_320_1723, w_320_1737, w_320_1741, w_320_1749, w_320_1763, w_320_1765, w_320_1769, w_320_1788, w_320_1791, w_320_1792, w_320_1799, w_320_1816, w_320_1836, w_320_1842, w_320_1843, w_320_1845, w_320_1848, w_320_1857, w_320_1859, w_320_1866, w_320_1875, w_320_1885, w_320_1890, w_320_1911, w_320_1913, w_320_1917, w_320_1918, w_320_1928, w_320_1931, w_320_1934, w_320_1939, w_320_1942, w_320_1949, w_320_1953, w_320_1958, w_320_1965, w_320_1980, w_320_1988, w_320_1989, w_320_2005, w_320_2010, w_320_2031, w_320_2032, w_320_2033, w_320_2034, w_320_2035, w_320_2036, w_320_2037, w_320_2038, w_320_2039, w_320_2040, w_320_2041, w_320_2043;
  wire w_321_002, w_321_010, w_321_012, w_321_014, w_321_022, w_321_023, w_321_024, w_321_028, w_321_032, w_321_033, w_321_047, w_321_051, w_321_054, w_321_056, w_321_064, w_321_070, w_321_073, w_321_074, w_321_075, w_321_078, w_321_080, w_321_087, w_321_089, w_321_090, w_321_096, w_321_097, w_321_102, w_321_103, w_321_106, w_321_114, w_321_115, w_321_116, w_321_121, w_321_128, w_321_131, w_321_132, w_321_133, w_321_134, w_321_135, w_321_138, w_321_139, w_321_142, w_321_144, w_321_147, w_321_154, w_321_155, w_321_160, w_321_161, w_321_164, w_321_167, w_321_169, w_321_170, w_321_173, w_321_177, w_321_179, w_321_182, w_321_186, w_321_187, w_321_188, w_321_192, w_321_195, w_321_197, w_321_201, w_321_202, w_321_204, w_321_207, w_321_214, w_321_216, w_321_220, w_321_224, w_321_225, w_321_231, w_321_236, w_321_246, w_321_248, w_321_256, w_321_258, w_321_259, w_321_260, w_321_262, w_321_264, w_321_265, w_321_267, w_321_270, w_321_273, w_321_275, w_321_279, w_321_280, w_321_282, w_321_284, w_321_288, w_321_293, w_321_298, w_321_299, w_321_302, w_321_308, w_321_314, w_321_315, w_321_316, w_321_317, w_321_318, w_321_320, w_321_321, w_321_331, w_321_336, w_321_345, w_321_348, w_321_355, w_321_360, w_321_363, w_321_367, w_321_369, w_321_370, w_321_375, w_321_379, w_321_388, w_321_393, w_321_394, w_321_396, w_321_398, w_321_405, w_321_406, w_321_407, w_321_411, w_321_413, w_321_420, w_321_421, w_321_425, w_321_431, w_321_432, w_321_438, w_321_440, w_321_447, w_321_448, w_321_458, w_321_460, w_321_462, w_321_463, w_321_467, w_321_469, w_321_470, w_321_471, w_321_474, w_321_482, w_321_488, w_321_492, w_321_493, w_321_495, w_321_497, w_321_499, w_321_501, w_321_503, w_321_506, w_321_509, w_321_513, w_321_514, w_321_522, w_321_524, w_321_530, w_321_531, w_321_537, w_321_538, w_321_540, w_321_544, w_321_545, w_321_547, w_321_548, w_321_553, w_321_554, w_321_555, w_321_557, w_321_558, w_321_559, w_321_560, w_321_565, w_321_567, w_321_569, w_321_571, w_321_576, w_321_580, w_321_585, w_321_586, w_321_587, w_321_589, w_321_591, w_321_592, w_321_606, w_321_619, w_321_621, w_321_622, w_321_623, w_321_626, w_321_633, w_321_635, w_321_636, w_321_640, w_321_641, w_321_643, w_321_651, w_321_654, w_321_657, w_321_659, w_321_669, w_321_670, w_321_671, w_321_678, w_321_681, w_321_683, w_321_684, w_321_689, w_321_692, w_321_693, w_321_696, w_321_699, w_321_700, w_321_702, w_321_710, w_321_712, w_321_715, w_321_719, w_321_720, w_321_724, w_321_725, w_321_726, w_321_730, w_321_731, w_321_733, w_321_736, w_321_741, w_321_754, w_321_757, w_321_772, w_321_774, w_321_781, w_321_787, w_321_790, w_321_797, w_321_799, w_321_800, w_321_801, w_321_803, w_321_809, w_321_812, w_321_814, w_321_817, w_321_825, w_321_826, w_321_829, w_321_831, w_321_833, w_321_840, w_321_843, w_321_845, w_321_847, w_321_848, w_321_851, w_321_854, w_321_857, w_321_866, w_321_867, w_321_868, w_321_875, w_321_878, w_321_889, w_321_890, w_321_895, w_321_901, w_321_903, w_321_908, w_321_910, w_321_911, w_321_912, w_321_915, w_321_920, w_321_921, w_321_922, w_321_923, w_321_925, w_321_926, w_321_935, w_321_943, w_321_944, w_321_946, w_321_953, w_321_954, w_321_955, w_321_967, w_321_974, w_321_977, w_321_978, w_321_981, w_321_983, w_321_985, w_321_986, w_321_997, w_321_1001, w_321_1004, w_321_1010, w_321_1011, w_321_1026, w_321_1027;
  wire w_322_000, w_322_005, w_322_020, w_322_021, w_322_025, w_322_029, w_322_046, w_322_050, w_322_051, w_322_056, w_322_058, w_322_061, w_322_064, w_322_069, w_322_071, w_322_075, w_322_079, w_322_088, w_322_095, w_322_101, w_322_111, w_322_112, w_322_115, w_322_126, w_322_129, w_322_135, w_322_138, w_322_142, w_322_145, w_322_150, w_322_153, w_322_156, w_322_159, w_322_164, w_322_166, w_322_169, w_322_172, w_322_179, w_322_182, w_322_191, w_322_199, w_322_201, w_322_204, w_322_208, w_322_214, w_322_221, w_322_225, w_322_226, w_322_228, w_322_239, w_322_247, w_322_248, w_322_250, w_322_251, w_322_263, w_322_264, w_322_266, w_322_268, w_322_274, w_322_280, w_322_287, w_322_303, w_322_305, w_322_307, w_322_309, w_322_310, w_322_318, w_322_328, w_322_329, w_322_330, w_322_336, w_322_338, w_322_348, w_322_350, w_322_357, w_322_359, w_322_365, w_322_366, w_322_373, w_322_377, w_322_381, w_322_386, w_322_388, w_322_393, w_322_411, w_322_412, w_322_413, w_322_419, w_322_421, w_322_424, w_322_428, w_322_436, w_322_437, w_322_441, w_322_457, w_322_461, w_322_463, w_322_478, w_322_488, w_322_497, w_322_499, w_322_502, w_322_507, w_322_510, w_322_516, w_322_519, w_322_520, w_322_521, w_322_523, w_322_527, w_322_533, w_322_542, w_322_556, w_322_562, w_322_572, w_322_573, w_322_577, w_322_583, w_322_588, w_322_589, w_322_595, w_322_596, w_322_598, w_322_603, w_322_620, w_322_630, w_322_633, w_322_635, w_322_644, w_322_645, w_322_648, w_322_649, w_322_656, w_322_658, w_322_659, w_322_666, w_322_674, w_322_677, w_322_679, w_322_682, w_322_689, w_322_690, w_322_698, w_322_700, w_322_702, w_322_718, w_322_720, w_322_726, w_322_732, w_322_739, w_322_746, w_322_749, w_322_751, w_322_752, w_322_755, w_322_757, w_322_763, w_322_765, w_322_766, w_322_773, w_322_776, w_322_777, w_322_779, w_322_788, w_322_789, w_322_790, w_322_811, w_322_816, w_322_821, w_322_825, w_322_841, w_322_843, w_322_845, w_322_848, w_322_856, w_322_859, w_322_864, w_322_865, w_322_887, w_322_892, w_322_893, w_322_901, w_322_921, w_322_928, w_322_936, w_322_942, w_322_943, w_322_946, w_322_956, w_322_957, w_322_959, w_322_960, w_322_969, w_322_972, w_322_975, w_322_976, w_322_988, w_322_989, w_322_1008, w_322_1011, w_322_1012, w_322_1016, w_322_1021, w_322_1029, w_322_1030, w_322_1035, w_322_1036, w_322_1038, w_322_1040, w_322_1045, w_322_1052, w_322_1053, w_322_1055, w_322_1067, w_322_1071, w_322_1076, w_322_1078, w_322_1094, w_322_1095, w_322_1098, w_322_1110, w_322_1113, w_322_1115, w_322_1116, w_322_1123, w_322_1127, w_322_1134, w_322_1142, w_322_1152, w_322_1154, w_322_1156, w_322_1159, w_322_1161, w_322_1168, w_322_1181, w_322_1186, w_322_1189, w_322_1191, w_322_1192, w_322_1202, w_322_1215, w_322_1220, w_322_1222, w_322_1225, w_322_1226, w_322_1227, w_322_1228, w_322_1235, w_322_1243, w_322_1250, w_322_1258, w_322_1263, w_322_1269, w_322_1274, w_322_1283, w_322_1284, w_322_1302, w_322_1316, w_322_1323, w_322_1325, w_322_1332, w_322_1335, w_322_1340, w_322_1346, w_322_1351, w_322_1354, w_322_1365, w_322_1374, w_322_1379, w_322_1382, w_322_1388, w_322_1394, w_322_1395, w_322_1405, w_322_1414, w_322_1419, w_322_1427, w_322_1437, w_322_1445, w_322_1478, w_322_1495, w_322_1498, w_322_1506, w_322_1513, w_322_1514, w_322_1536, w_322_1547, w_322_1562, w_322_1566, w_322_1575, w_322_1580, w_322_1584, w_322_1594, w_322_1604, w_322_1607, w_322_1612, w_322_1613, w_322_1639, w_322_1641, w_322_1643, w_322_1644, w_322_1648, w_322_1664, w_322_1667, w_322_1670, w_322_1689, w_322_1692, w_322_1709, w_322_1745, w_322_1751, w_322_1765, w_322_1781, w_322_1782, w_322_1783, w_322_1790, w_322_1794, w_322_1812, w_322_1814, w_322_1828, w_322_1830, w_322_1831, w_322_1854, w_322_1855, w_322_1857;
  wire w_323_000, w_323_004, w_323_021, w_323_026, w_323_027, w_323_037, w_323_044, w_323_046, w_323_053, w_323_055, w_323_067, w_323_077, w_323_083, w_323_095, w_323_106, w_323_132, w_323_166, w_323_168, w_323_171, w_323_177, w_323_185, w_323_199, w_323_203, w_323_204, w_323_205, w_323_224, w_323_230, w_323_232, w_323_238, w_323_239, w_323_261, w_323_262, w_323_265, w_323_277, w_323_295, w_323_296, w_323_300, w_323_324, w_323_329, w_323_334, w_323_344, w_323_349, w_323_350, w_323_356, w_323_361, w_323_362, w_323_379, w_323_391, w_323_412, w_323_417, w_323_429, w_323_450, w_323_458, w_323_467, w_323_479, w_323_500, w_323_521, w_323_534, w_323_535, w_323_545, w_323_550, w_323_556, w_323_574, w_323_589, w_323_597, w_323_600, w_323_607, w_323_611, w_323_619, w_323_621, w_323_622, w_323_631, w_323_633, w_323_643, w_323_649, w_323_654, w_323_665, w_323_674, w_323_689, w_323_691, w_323_701, w_323_710, w_323_729, w_323_738, w_323_742, w_323_747, w_323_757, w_323_759, w_323_777, w_323_785, w_323_795, w_323_805, w_323_812, w_323_830, w_323_853, w_323_858, w_323_862, w_323_879, w_323_888, w_323_896, w_323_903, w_323_907, w_323_914, w_323_926, w_323_930, w_323_937, w_323_947, w_323_961, w_323_963, w_323_971, w_323_1014, w_323_1017, w_323_1024, w_323_1025, w_323_1045, w_323_1046, w_323_1048, w_323_1052, w_323_1053, w_323_1062, w_323_1065, w_323_1068, w_323_1077, w_323_1084, w_323_1085, w_323_1098, w_323_1116, w_323_1121, w_323_1142, w_323_1152, w_323_1154, w_323_1158, w_323_1165, w_323_1171, w_323_1183, w_323_1201, w_323_1204, w_323_1208, w_323_1209, w_323_1210, w_323_1215, w_323_1218, w_323_1219, w_323_1221, w_323_1229, w_323_1254, w_323_1282, w_323_1289, w_323_1298, w_323_1316, w_323_1326, w_323_1329, w_323_1351, w_323_1359, w_323_1364, w_323_1367, w_323_1379, w_323_1381, w_323_1383, w_323_1386, w_323_1387, w_323_1394, w_323_1396, w_323_1409, w_323_1425, w_323_1449, w_323_1454, w_323_1467, w_323_1469, w_323_1492, w_323_1497, w_323_1500, w_323_1511, w_323_1516, w_323_1518, w_323_1520, w_323_1528, w_323_1538, w_323_1554, w_323_1557, w_323_1558, w_323_1572, w_323_1576, w_323_1579, w_323_1584, w_323_1594, w_323_1602, w_323_1629, w_323_1632, w_323_1644, w_323_1650, w_323_1651, w_323_1653, w_323_1665, w_323_1666, w_323_1673, w_323_1693, w_323_1698, w_323_1702, w_323_1705, w_323_1706, w_323_1708, w_323_1729, w_323_1742, w_323_1747, w_323_1765, w_323_1794, w_323_1796, w_323_1807, w_323_1832, w_323_1833, w_323_1850, w_323_1854, w_323_1857, w_323_1866, w_323_1870, w_323_1881, w_323_1886, w_323_1892, w_323_1901, w_323_1909, w_323_1923, w_323_1930, w_323_1931, w_323_1934, w_323_1941, w_323_1953, w_323_1957, w_323_1969, w_323_1978, w_323_1983, w_323_1989, w_323_2024, w_323_2042, w_323_2043, w_323_2060, w_323_2095, w_323_2122, w_323_2130, w_323_2170, w_323_2192, w_323_2193, w_323_2205, w_323_2208, w_323_2210, w_323_2266, w_323_2279, w_323_2290, w_323_2294, w_323_2314, w_323_2320, w_323_2354, w_323_2356, w_323_2397, w_323_2403, w_323_2409, w_323_2465, w_323_2467, w_323_2474, w_323_2477, w_323_2489, w_323_2505, w_323_2507, w_323_2533, w_323_2539, w_323_2541, w_323_2564, w_323_2591, w_323_2598, w_323_2599, w_323_2606, w_323_2610, w_323_2613, w_323_2654, w_323_2655, w_323_2660, w_323_2695, w_323_2714, w_323_2733, w_323_2739, w_323_2744, w_323_2758, w_323_2769, w_323_2771, w_323_2837, w_323_2842, w_323_2864, w_323_2885, w_323_2890, w_323_2908, w_323_2912, w_323_2918, w_323_2919, w_323_2925, w_323_2961, w_323_2986, w_323_3006, w_323_3012, w_323_3021, w_323_3022, w_323_3023, w_323_3024;
  wire w_324_018, w_324_028, w_324_030, w_324_038, w_324_053, w_324_055, w_324_081, w_324_082, w_324_092, w_324_093, w_324_101, w_324_104, w_324_108, w_324_111, w_324_116, w_324_125, w_324_136, w_324_138, w_324_139, w_324_143, w_324_162, w_324_165, w_324_170, w_324_172, w_324_187, w_324_202, w_324_208, w_324_215, w_324_224, w_324_226, w_324_242, w_324_258, w_324_262, w_324_277, w_324_294, w_324_306, w_324_310, w_324_328, w_324_330, w_324_343, w_324_344, w_324_353, w_324_354, w_324_358, w_324_359, w_324_369, w_324_372, w_324_379, w_324_388, w_324_392, w_324_394, w_324_399, w_324_406, w_324_412, w_324_431, w_324_435, w_324_438, w_324_446, w_324_451, w_324_453, w_324_459, w_324_462, w_324_465, w_324_468, w_324_475, w_324_478, w_324_490, w_324_493, w_324_496, w_324_497, w_324_498, w_324_502, w_324_505, w_324_507, w_324_514, w_324_523, w_324_528, w_324_530, w_324_536, w_324_537, w_324_540, w_324_542, w_324_547, w_324_552, w_324_555, w_324_570, w_324_575, w_324_584, w_324_585, w_324_592, w_324_594, w_324_598, w_324_606, w_324_645, w_324_647, w_324_650, w_324_655, w_324_656, w_324_671, w_324_674, w_324_678, w_324_679, w_324_683, w_324_688, w_324_690, w_324_692, w_324_697, w_324_712, w_324_725, w_324_728, w_324_734, w_324_737, w_324_739, w_324_744, w_324_753, w_324_756, w_324_758, w_324_759, w_324_762, w_324_770, w_324_773, w_324_776, w_324_783, w_324_786, w_324_795, w_324_797, w_324_803, w_324_812, w_324_813, w_324_816, w_324_817, w_324_827, w_324_828, w_324_840, w_324_841, w_324_844, w_324_857, w_324_862, w_324_870, w_324_878, w_324_888, w_324_890, w_324_891, w_324_910, w_324_924, w_324_927, w_324_934, w_324_936, w_324_951, w_324_957, w_324_958, w_324_969, w_324_977, w_324_980, w_324_990, w_324_991, w_324_997, w_324_1006, w_324_1017, w_324_1019, w_324_1021, w_324_1031, w_324_1045, w_324_1049, w_324_1091, w_324_1098, w_324_1128, w_324_1132, w_324_1134, w_324_1137, w_324_1140, w_324_1153, w_324_1163, w_324_1172, w_324_1177, w_324_1188, w_324_1189, w_324_1210, w_324_1215, w_324_1223, w_324_1225, w_324_1245, w_324_1254, w_324_1261, w_324_1268, w_324_1271, w_324_1273, w_324_1281, w_324_1284, w_324_1293, w_324_1298, w_324_1308, w_324_1312, w_324_1323, w_324_1336, w_324_1365, w_324_1374, w_324_1396, w_324_1420, w_324_1422, w_324_1431, w_324_1432, w_324_1439, w_324_1441, w_324_1445, w_324_1452, w_324_1458, w_324_1462, w_324_1497, w_324_1498, w_324_1504, w_324_1507, w_324_1519, w_324_1520, w_324_1530, w_324_1541, w_324_1544, w_324_1577, w_324_1579, w_324_1589, w_324_1592, w_324_1594, w_324_1602, w_324_1614, w_324_1616, w_324_1620, w_324_1621, w_324_1622, w_324_1623, w_324_1628, w_324_1637, w_324_1642, w_324_1650, w_324_1665, w_324_1667, w_324_1671, w_324_1686, w_324_1693, w_324_1715, w_324_1718, w_324_1741, w_324_1743, w_324_1756, w_324_1770, w_324_1771, w_324_1772, w_324_1775, w_324_1801, w_324_1802, w_324_1803, w_324_1806, w_324_1808, w_324_1811, w_324_1812, w_324_1839, w_324_1840, w_324_1846, w_324_1850, w_324_1858, w_324_1899, w_324_1900, w_324_1909, w_324_1911, w_324_1922, w_324_1923, w_324_1929, w_324_1935, w_324_1936, w_324_1942, w_324_1945, w_324_1946, w_324_1947, w_324_1980, w_324_1983, w_324_1988, w_324_1996, w_324_1998, w_324_2016, w_324_2042, w_324_2064, w_324_2071, w_324_2091, w_324_2112, w_324_2119, w_324_2126, w_324_2131, w_324_2156, w_324_2252, w_324_2253, w_324_2311, w_324_2350, w_324_2366, w_324_2368, w_324_2386, w_324_2388, w_324_2401, w_324_2402, w_324_2432, w_324_2442, w_324_2455, w_324_2467, w_324_2476, w_324_2491, w_324_2492, w_324_2503, w_324_2504, w_324_2513, w_324_2527, w_324_2542, w_324_2545, w_324_2555, w_324_2558, w_324_2562, w_324_2593, w_324_2603, w_324_2604, w_324_2608, w_324_2622, w_324_2624, w_324_2650, w_324_2663, w_324_2676, w_324_2686, w_324_2688, w_324_2720, w_324_2722, w_324_2734, w_324_2738, w_324_2748, w_324_2751, w_324_2757, w_324_2772, w_324_2774, w_324_2783, w_324_2788, w_324_2791, w_324_2799, w_324_2830, w_324_2839, w_324_2916, w_324_2936, w_324_2940, w_324_2950, w_324_2971, w_324_2974, w_324_2987, w_324_2988, w_324_2989, w_324_2990;
  wire w_325_008, w_325_011, w_325_012, w_325_019, w_325_028, w_325_029, w_325_037, w_325_050, w_325_057, w_325_064, w_325_067, w_325_086, w_325_090, w_325_091, w_325_092, w_325_097, w_325_105, w_325_111, w_325_113, w_325_115, w_325_126, w_325_150, w_325_152, w_325_155, w_325_157, w_325_162, w_325_168, w_325_169, w_325_172, w_325_174, w_325_175, w_325_178, w_325_184, w_325_186, w_325_191, w_325_203, w_325_212, w_325_213, w_325_220, w_325_225, w_325_232, w_325_233, w_325_239, w_325_246, w_325_256, w_325_278, w_325_280, w_325_306, w_325_336, w_325_338, w_325_349, w_325_352, w_325_366, w_325_386, w_325_406, w_325_413, w_325_418, w_325_432, w_325_437, w_325_441, w_325_444, w_325_456, w_325_461, w_325_462, w_325_477, w_325_481, w_325_485, w_325_500, w_325_502, w_325_504, w_325_505, w_325_507, w_325_508, w_325_517, w_325_522, w_325_536, w_325_537, w_325_546, w_325_552, w_325_561, w_325_569, w_325_588, w_325_589, w_325_615, w_325_618, w_325_621, w_325_629, w_325_657, w_325_658, w_325_661, w_325_688, w_325_697, w_325_712, w_325_717, w_325_729, w_325_730, w_325_731, w_325_744, w_325_748, w_325_762, w_325_772, w_325_783, w_325_789, w_325_792, w_325_806, w_325_809, w_325_815, w_325_826, w_325_845, w_325_851, w_325_853, w_325_858, w_325_869, w_325_875, w_325_876, w_325_882, w_325_886, w_325_897, w_325_899, w_325_903, w_325_907, w_325_932, w_325_945, w_325_958, w_325_965, w_325_1000, w_325_1020, w_325_1038, w_325_1042, w_325_1059, w_325_1068, w_325_1080, w_325_1089, w_325_1095, w_325_1104, w_325_1124, w_325_1132, w_325_1174, w_325_1226, w_325_1238, w_325_1244, w_325_1251, w_325_1272, w_325_1281, w_325_1312, w_325_1323, w_325_1332, w_325_1387, w_325_1402, w_325_1408, w_325_1414, w_325_1464, w_325_1480, w_325_1504, w_325_1518, w_325_1521, w_325_1524, w_325_1561, w_325_1565, w_325_1570, w_325_1587, w_325_1601, w_325_1614, w_325_1617, w_325_1660, w_325_1671, w_325_1702, w_325_1724, w_325_1739, w_325_1763, w_325_1771, w_325_1791, w_325_1805, w_325_1809, w_325_1828, w_325_1832, w_325_1842, w_325_1874, w_325_1880, w_325_1901, w_325_1903, w_325_1928, w_325_1932, w_325_1949, w_325_1983, w_325_1985, w_325_2019, w_325_2032, w_325_2082, w_325_2100, w_325_2102, w_325_2110, w_325_2115, w_325_2119, w_325_2121, w_325_2127, w_325_2165, w_325_2176, w_325_2190, w_325_2255, w_325_2315, w_325_2338, w_325_2356, w_325_2363, w_325_2413, w_325_2428, w_325_2431, w_325_2435, w_325_2445, w_325_2450, w_325_2472, w_325_2475, w_325_2497, w_325_2509, w_325_2527, w_325_2537, w_325_2546, w_325_2551, w_325_2570, w_325_2584, w_325_2598, w_325_2609, w_325_2612, w_325_2670, w_325_2673, w_325_2675, w_325_2714, w_325_2717, w_325_2757, w_325_2782, w_325_2788, w_325_2814, w_325_2817, w_325_2818, w_325_2819, w_325_2829, w_325_2846, w_325_2859, w_325_2906, w_325_2953, w_325_2970, w_325_3013, w_325_3014, w_325_3029, w_325_3040, w_325_3088, w_325_3089, w_325_3104, w_325_3105, w_325_3123, w_325_3125, w_325_3127, w_325_3134, w_325_3139, w_325_3140, w_325_3146, w_325_3178, w_325_3186, w_325_3191, w_325_3228, w_325_3250, w_325_3268, w_325_3277, w_325_3284, w_325_3285, w_325_3288, w_325_3309, w_325_3319, w_325_3331, w_325_3345, w_325_3350, w_325_3359, w_325_3360, w_325_3379, w_325_3383, w_325_3388, w_325_3393, w_325_3430, w_325_3442, w_325_3444, w_325_3448, w_325_3497, w_325_3518, w_325_3522, w_325_3531, w_325_3537, w_325_3544, w_325_3591, w_325_3619, w_325_3719, w_325_3747, w_325_3753, w_325_3813, w_325_3858, w_325_3860, w_325_3882, w_325_3895, w_325_3927, w_325_3932, w_325_3943, w_325_3977, w_325_4022, w_325_4024, w_325_4052, w_325_4089, w_325_4104, w_325_4112, w_325_4113, w_325_4114, w_325_4115, w_325_4116, w_325_4117, w_325_4118, w_325_4119, w_325_4120, w_325_4121, w_325_4122, w_325_4123, w_325_4127, w_325_4128, w_325_4129, w_325_4130, w_325_4132;
  wire w_326_001, w_326_005, w_326_018, w_326_020, w_326_034, w_326_036, w_326_041, w_326_044, w_326_045, w_326_048, w_326_054, w_326_057, w_326_067, w_326_068, w_326_072, w_326_078, w_326_081, w_326_088, w_326_089, w_326_104, w_326_109, w_326_111, w_326_113, w_326_116, w_326_117, w_326_118, w_326_124, w_326_131, w_326_135, w_326_141, w_326_145, w_326_147, w_326_151, w_326_152, w_326_154, w_326_166, w_326_170, w_326_173, w_326_186, w_326_187, w_326_188, w_326_192, w_326_193, w_326_194, w_326_195, w_326_197, w_326_205, w_326_215, w_326_216, w_326_221, w_326_227, w_326_235, w_326_246, w_326_256, w_326_258, w_326_259, w_326_262, w_326_266, w_326_271, w_326_305, w_326_320, w_326_326, w_326_332, w_326_350, w_326_357, w_326_378, w_326_385, w_326_386, w_326_391, w_326_392, w_326_395, w_326_397, w_326_411, w_326_413, w_326_425, w_326_429, w_326_433, w_326_438, w_326_445, w_326_455, w_326_464, w_326_480, w_326_485, w_326_487, w_326_499, w_326_508, w_326_511, w_326_524, w_326_526, w_326_528, w_326_537, w_326_539, w_326_540, w_326_541, w_326_551, w_326_565, w_326_573, w_326_576, w_326_582, w_326_584, w_326_585, w_326_587, w_326_591, w_326_598, w_326_606, w_326_613, w_326_616, w_326_627, w_326_633, w_326_637, w_326_644, w_326_646, w_326_649, w_326_651, w_326_661, w_326_675, w_326_680, w_326_682, w_326_684, w_326_686, w_326_689, w_326_690, w_326_693, w_326_701, w_326_704, w_326_713, w_326_714, w_326_717, w_326_719, w_326_724, w_326_726, w_326_727, w_326_733, w_326_738, w_326_740, w_326_752, w_326_755, w_326_758, w_326_759, w_326_763, w_326_780, w_326_787, w_326_790, w_326_793, w_326_796, w_326_797, w_326_799, w_326_804, w_326_821, w_326_825, w_326_833, w_326_835, w_326_836, w_326_847, w_326_850, w_326_851, w_326_852, w_326_860, w_326_862, w_326_863, w_326_868, w_326_875, w_326_878, w_326_879, w_326_903, w_326_904, w_326_907, w_326_926, w_326_944, w_326_947, w_326_950, w_326_961, w_326_962, w_326_969, w_326_978, w_326_986, w_326_990, w_326_996, w_326_998, w_326_1002, w_326_1012, w_326_1013, w_326_1016, w_326_1018, w_326_1020, w_326_1023, w_326_1028, w_326_1033, w_326_1045, w_326_1049, w_326_1051, w_326_1056, w_326_1057, w_326_1065, w_326_1071, w_326_1073, w_326_1077, w_326_1078, w_326_1081, w_326_1083, w_326_1089, w_326_1095, w_326_1097, w_326_1101, w_326_1105, w_326_1108, w_326_1118, w_326_1139, w_326_1140, w_326_1143, w_326_1146, w_326_1148, w_326_1156, w_326_1162, w_326_1173, w_326_1183, w_326_1185, w_326_1191, w_326_1194, w_326_1200, w_326_1206, w_326_1214, w_326_1217, w_326_1223, w_326_1224, w_326_1227, w_326_1235, w_326_1239, w_326_1241, w_326_1243, w_326_1244, w_326_1249, w_326_1253, w_326_1254, w_326_1260, w_326_1262, w_326_1265, w_326_1266, w_326_1280, w_326_1296, w_326_1301, w_326_1307, w_326_1318, w_326_1323, w_326_1331, w_326_1333, w_326_1337, w_326_1339, w_326_1347, w_326_1357, w_326_1364, w_326_1374, w_326_1380, w_326_1385, w_326_1386, w_326_1389, w_326_1393, w_326_1394, w_326_1398, w_326_1417, w_326_1420, w_326_1425, w_326_1434, w_326_1440, w_326_1441, w_326_1443, w_326_1454, w_326_1456, w_326_1465, w_326_1467, w_326_1474, w_326_1476, w_326_1477, w_326_1485, w_326_1487, w_326_1488, w_326_1490, w_326_1511, w_326_1512, w_326_1517, w_326_1520, w_326_1522, w_326_1533, w_326_1546, w_326_1552, w_326_1557, w_326_1562, w_326_1566, w_326_1567, w_326_1579, w_326_1584, w_326_1585, w_326_1586, w_326_1587, w_326_1604, w_326_1613, w_326_1624, w_326_1630;
  wire w_327_007, w_327_019, w_327_022, w_327_023, w_327_024, w_327_034, w_327_041, w_327_050, w_327_053, w_327_055, w_327_058, w_327_059, w_327_064, w_327_069, w_327_098, w_327_107, w_327_126, w_327_128, w_327_135, w_327_151, w_327_170, w_327_178, w_327_191, w_327_196, w_327_197, w_327_212, w_327_213, w_327_220, w_327_228, w_327_248, w_327_252, w_327_253, w_327_257, w_327_275, w_327_302, w_327_315, w_327_321, w_327_327, w_327_336, w_327_351, w_327_354, w_327_364, w_327_380, w_327_383, w_327_387, w_327_391, w_327_399, w_327_403, w_327_411, w_327_414, w_327_416, w_327_417, w_327_420, w_327_439, w_327_454, w_327_483, w_327_504, w_327_514, w_327_526, w_327_527, w_327_528, w_327_530, w_327_533, w_327_556, w_327_557, w_327_562, w_327_568, w_327_585, w_327_607, w_327_623, w_327_628, w_327_647, w_327_660, w_327_664, w_327_665, w_327_675, w_327_698, w_327_718, w_327_720, w_327_728, w_327_729, w_327_737, w_327_744, w_327_746, w_327_747, w_327_754, w_327_755, w_327_770, w_327_792, w_327_819, w_327_828, w_327_833, w_327_835, w_327_853, w_327_872, w_327_874, w_327_877, w_327_880, w_327_897, w_327_923, w_327_926, w_327_928, w_327_941, w_327_947, w_327_948, w_327_951, w_327_953, w_327_956, w_327_963, w_327_972, w_327_1004, w_327_1005, w_327_1008, w_327_1023, w_327_1028, w_327_1043, w_327_1060, w_327_1061, w_327_1071, w_327_1080, w_327_1081, w_327_1093, w_327_1108, w_327_1118, w_327_1136, w_327_1144, w_327_1148, w_327_1150, w_327_1168, w_327_1183, w_327_1186, w_327_1189, w_327_1190, w_327_1205, w_327_1209, w_327_1226, w_327_1250, w_327_1256, w_327_1260, w_327_1269, w_327_1279, w_327_1284, w_327_1285, w_327_1286, w_327_1312, w_327_1316, w_327_1324, w_327_1326, w_327_1332, w_327_1333, w_327_1334, w_327_1372, w_327_1377, w_327_1379, w_327_1392, w_327_1414, w_327_1420, w_327_1436, w_327_1442, w_327_1446, w_327_1451, w_327_1454, w_327_1460, w_327_1464, w_327_1493, w_327_1497, w_327_1502, w_327_1503, w_327_1517, w_327_1531, w_327_1533, w_327_1534, w_327_1538, w_327_1551, w_327_1558, w_327_1566, w_327_1568, w_327_1572, w_327_1604, w_327_1615, w_327_1617, w_327_1618, w_327_1647, w_327_1653, w_327_1659, w_327_1677, w_327_1684, w_327_1686, w_327_1689, w_327_1718, w_327_1725, w_327_1736, w_327_1741, w_327_1742, w_327_1753, w_327_1761, w_327_1764, w_327_1772, w_327_1776, w_327_1779, w_327_1796, w_327_1803, w_327_1832, w_327_1870, w_327_1881, w_327_1889, w_327_1910, w_327_1914, w_327_1924, w_327_1959, w_327_2015, w_327_2046, w_327_2055, w_327_2061, w_327_2068, w_327_2097, w_327_2118, w_327_2130, w_327_2132, w_327_2172, w_327_2181, w_327_2204, w_327_2236, w_327_2264, w_327_2283, w_327_2318, w_327_2362, w_327_2381, w_327_2404, w_327_2406, w_327_2462, w_327_2478, w_327_2491, w_327_2501, w_327_2524, w_327_2539, w_327_2553, w_327_2574, w_327_2575, w_327_2582, w_327_2628, w_327_2639, w_327_2640, w_327_2652, w_327_2655, w_327_2665, w_327_2670, w_327_2672, w_327_2688, w_327_2702, w_327_2707, w_327_2738, w_327_2741, w_327_2747, w_327_2751, w_327_2790, w_327_2798, w_327_2823, w_327_2824, w_327_2827, w_327_2886, w_327_2918, w_327_2919, w_327_2971, w_327_2994, w_327_3016, w_327_3029, w_327_3037, w_327_3080, w_327_3115, w_327_3125, w_327_3164, w_327_3197, w_327_3225, w_327_3234, w_327_3242, w_327_3252, w_327_3253, w_327_3270, w_327_3284, w_327_3285, w_327_3288, w_327_3297, w_327_3303, w_327_3310, w_327_3311, w_327_3312, w_327_3313, w_327_3314, w_327_3315, w_327_3316, w_327_3317, w_327_3318, w_327_3319, w_327_3320, w_327_3321;
  wire w_328_000, w_328_003, w_328_009, w_328_012, w_328_014, w_328_021, w_328_025, w_328_032, w_328_044, w_328_048, w_328_049, w_328_052, w_328_053, w_328_061, w_328_062, w_328_064, w_328_066, w_328_071, w_328_073, w_328_074, w_328_083, w_328_093, w_328_098, w_328_099, w_328_109, w_328_117, w_328_123, w_328_128, w_328_139, w_328_142, w_328_144, w_328_147, w_328_148, w_328_153, w_328_164, w_328_171, w_328_175, w_328_177, w_328_184, w_328_188, w_328_189, w_328_192, w_328_193, w_328_202, w_328_204, w_328_206, w_328_214, w_328_217, w_328_222, w_328_227, w_328_235, w_328_245, w_328_256, w_328_279, w_328_287, w_328_295, w_328_297, w_328_305, w_328_309, w_328_316, w_328_320, w_328_329, w_328_332, w_328_348, w_328_359, w_328_362, w_328_365, w_328_368, w_328_386, w_328_389, w_328_393, w_328_397, w_328_405, w_328_406, w_328_407, w_328_410, w_328_411, w_328_413, w_328_417, w_328_418, w_328_425, w_328_428, w_328_437, w_328_440, w_328_445, w_328_446, w_328_447, w_328_454, w_328_461, w_328_463, w_328_472, w_328_477, w_328_480, w_328_486, w_328_488, w_328_492, w_328_494, w_328_498, w_328_503, w_328_507, w_328_509, w_328_512, w_328_514, w_328_516, w_328_530, w_328_531, w_328_546, w_328_562, w_328_579, w_328_582, w_328_585, w_328_590, w_328_596, w_328_615, w_328_617, w_328_624, w_328_628, w_328_629, w_328_630, w_328_634, w_328_659, w_328_663, w_328_665, w_328_673, w_328_675, w_328_676, w_328_682, w_328_686, w_328_689, w_328_690, w_328_694, w_328_695, w_328_697, w_328_712, w_328_713, w_328_714, w_328_733, w_328_739, w_328_747, w_328_752, w_328_755, w_328_764, w_328_772, w_328_774, w_328_777, w_328_796, w_328_802, w_328_807, w_328_822, w_328_824, w_328_840, w_328_849, w_328_852, w_328_853, w_328_870, w_328_885, w_328_889, w_328_896, w_328_899, w_328_903, w_328_921, w_328_922, w_328_924, w_328_943, w_328_966, w_328_975, w_328_983, w_328_985, w_328_986, w_328_992, w_328_996, w_328_1015, w_328_1025, w_328_1043, w_328_1045, w_328_1049, w_328_1050, w_328_1061, w_328_1066, w_328_1069, w_328_1080, w_328_1089, w_328_1110, w_328_1116, w_328_1122, w_328_1129, w_328_1138, w_328_1160, w_328_1171, w_328_1175, w_328_1182, w_328_1183, w_328_1184, w_328_1187, w_328_1188, w_328_1203, w_328_1208, w_328_1221, w_328_1225, w_328_1227, w_328_1230, w_328_1233, w_328_1245, w_328_1252, w_328_1256, w_328_1261, w_328_1265, w_328_1271, w_328_1277, w_328_1281, w_328_1290, w_328_1291, w_328_1293, w_328_1296, w_328_1311, w_328_1312, w_328_1314, w_328_1317, w_328_1319, w_328_1324, w_328_1333, w_328_1336, w_328_1345, w_328_1353, w_328_1359, w_328_1366, w_328_1393, w_328_1414, w_328_1419, w_328_1428, w_328_1444, w_328_1450, w_328_1454, w_328_1457, w_328_1476, w_328_1493, w_328_1503, w_328_1505, w_328_1510, w_328_1515, w_328_1526, w_328_1539, w_328_1559, w_328_1561, w_328_1567, w_328_1572, w_328_1577, w_328_1580, w_328_1592, w_328_1597, w_328_1604, w_328_1613, w_328_1624, w_328_1627, w_328_1631, w_328_1642, w_328_1650, w_328_1663, w_328_1673, w_328_1676, w_328_1681, w_328_1688, w_328_1696, w_328_1709, w_328_1726, w_328_1728, w_328_1764, w_328_1772, w_328_1775, w_328_1783, w_328_1787, w_328_1793, w_328_1794, w_328_1822, w_328_1824, w_328_1830, w_328_1839, w_328_1849, w_328_1855, w_328_1874, w_328_1876, w_328_1879, w_328_1902, w_328_1917, w_328_1920, w_328_1925, w_328_1927, w_328_1933, w_328_1936, w_328_1938, w_328_1939, w_328_1950, w_328_1959, w_328_1966, w_328_1977, w_328_1978, w_328_1985, w_328_1990, w_328_2010, w_328_2015, w_328_2018, w_328_2019, w_328_2037, w_328_2039, w_328_2043, w_328_2051, w_328_2052, w_328_2054, w_328_2071, w_328_2087, w_328_2090, w_328_2098, w_328_2100, w_328_2101, w_328_2108, w_328_2119, w_328_2140, w_328_2144, w_328_2162, w_328_2172, w_328_2187, w_328_2194, w_328_2201, w_328_2202, w_328_2203, w_328_2204, w_328_2205, w_328_2206, w_328_2207, w_328_2209, w_328_2211, w_328_2212, w_328_2213, w_328_2214, w_328_2215, w_328_2216, w_328_2217, w_328_2218, w_328_2219, w_328_2220, w_328_2222;
  wire w_329_022, w_329_040, w_329_045, w_329_049, w_329_053, w_329_057, w_329_058, w_329_062, w_329_064, w_329_082, w_329_085, w_329_086, w_329_088, w_329_091, w_329_104, w_329_116, w_329_123, w_329_127, w_329_139, w_329_141, w_329_142, w_329_144, w_329_160, w_329_167, w_329_188, w_329_190, w_329_191, w_329_193, w_329_227, w_329_234, w_329_238, w_329_245, w_329_257, w_329_258, w_329_259, w_329_269, w_329_276, w_329_279, w_329_300, w_329_304, w_329_309, w_329_323, w_329_332, w_329_339, w_329_340, w_329_346, w_329_360, w_329_374, w_329_388, w_329_393, w_329_396, w_329_420, w_329_430, w_329_448, w_329_458, w_329_467, w_329_490, w_329_503, w_329_543, w_329_561, w_329_562, w_329_565, w_329_578, w_329_581, w_329_583, w_329_586, w_329_597, w_329_607, w_329_613, w_329_614, w_329_617, w_329_663, w_329_664, w_329_670, w_329_671, w_329_677, w_329_685, w_329_695, w_329_719, w_329_728, w_329_734, w_329_737, w_329_742, w_329_757, w_329_765, w_329_777, w_329_789, w_329_790, w_329_795, w_329_797, w_329_829, w_329_843, w_329_850, w_329_853, w_329_879, w_329_885, w_329_889, w_329_895, w_329_937, w_329_959, w_329_982, w_329_990, w_329_1003, w_329_1013, w_329_1019, w_329_1053, w_329_1068, w_329_1071, w_329_1089, w_329_1091, w_329_1095, w_329_1148, w_329_1158, w_329_1185, w_329_1188, w_329_1197, w_329_1235, w_329_1241, w_329_1242, w_329_1253, w_329_1257, w_329_1271, w_329_1281, w_329_1289, w_329_1297, w_329_1323, w_329_1337, w_329_1354, w_329_1367, w_329_1377, w_329_1388, w_329_1395, w_329_1416, w_329_1432, w_329_1461, w_329_1470, w_329_1495, w_329_1517, w_329_1520, w_329_1581, w_329_1589, w_329_1591, w_329_1639, w_329_1643, w_329_1644, w_329_1653, w_329_1663, w_329_1665, w_329_1680, w_329_1690, w_329_1705, w_329_1710, w_329_1715, w_329_1716, w_329_1719, w_329_1723, w_329_1750, w_329_1782, w_329_1785, w_329_1802, w_329_1811, w_329_1822, w_329_1827, w_329_1829, w_329_1838, w_329_1839, w_329_1863, w_329_1875, w_329_1889, w_329_1914, w_329_1932, w_329_1939, w_329_1959, w_329_1960, w_329_1968, w_329_1973, w_329_1994, w_329_2026, w_329_2049, w_329_2057, w_329_2064, w_329_2076, w_329_2090, w_329_2092, w_329_2097, w_329_2164, w_329_2167, w_329_2170, w_329_2189, w_329_2198, w_329_2202, w_329_2212, w_329_2239, w_329_2254, w_329_2262, w_329_2279, w_329_2298, w_329_2330, w_329_2351, w_329_2357, w_329_2391, w_329_2414, w_329_2417, w_329_2436, w_329_2446, w_329_2463, w_329_2468, w_329_2475, w_329_2486, w_329_2493, w_329_2499, w_329_2502, w_329_2505, w_329_2517, w_329_2544, w_329_2564, w_329_2566, w_329_2569, w_329_2570, w_329_2576, w_329_2593, w_329_2596, w_329_2622, w_329_2628, w_329_2629, w_329_2630, w_329_2644, w_329_2653, w_329_2662, w_329_2679, w_329_2681, w_329_2693, w_329_2713, w_329_2722, w_329_2729, w_329_2730, w_329_2736, w_329_2755, w_329_2783, w_329_2813, w_329_2821, w_329_2841, w_329_2857, w_329_2862, w_329_2984, w_329_2990, w_329_3004, w_329_3018, w_329_3020, w_329_3021, w_329_3037, w_329_3039, w_329_3042, w_329_3043, w_329_3050, w_329_3066, w_329_3073, w_329_3075, w_329_3083, w_329_3091, w_329_3103, w_329_3132, w_329_3136, w_329_3178, w_329_3189, w_329_3192, w_329_3201, w_329_3230, w_329_3271, w_329_3275, w_329_3288, w_329_3298, w_329_3304, w_329_3332, w_329_3351, w_329_3356, w_329_3364, w_329_3426, w_329_3430, w_329_3470, w_329_3481, w_329_3488, w_329_3503, w_329_3538, w_329_3595, w_329_3601, w_329_3620, w_329_3633, w_329_3654, w_329_3711, w_329_3714, w_329_3722, w_329_3726, w_329_3750, w_329_3770, w_329_3771, w_329_3781, w_329_3789, w_329_3790, w_329_3809, w_329_3814, w_329_3840, w_329_3854, w_329_3917, w_329_3926, w_329_3939, w_329_3942, w_329_3970, w_329_4006, w_329_4050;
  wire w_330_004, w_330_014, w_330_018, w_330_027, w_330_030, w_330_031, w_330_036, w_330_037, w_330_042, w_330_046, w_330_057, w_330_060, w_330_065, w_330_066, w_330_070, w_330_071, w_330_074, w_330_078, w_330_083, w_330_107, w_330_111, w_330_127, w_330_133, w_330_136, w_330_139, w_330_145, w_330_149, w_330_160, w_330_164, w_330_165, w_330_167, w_330_171, w_330_174, w_330_175, w_330_183, w_330_189, w_330_198, w_330_220, w_330_222, w_330_228, w_330_237, w_330_238, w_330_257, w_330_258, w_330_265, w_330_266, w_330_271, w_330_289, w_330_298, w_330_299, w_330_309, w_330_312, w_330_314, w_330_316, w_330_321, w_330_323, w_330_327, w_330_332, w_330_335, w_330_338, w_330_340, w_330_342, w_330_345, w_330_346, w_330_354, w_330_358, w_330_360, w_330_373, w_330_377, w_330_384, w_330_386, w_330_396, w_330_407, w_330_411, w_330_423, w_330_426, w_330_428, w_330_429, w_330_437, w_330_439, w_330_440, w_330_442, w_330_443, w_330_450, w_330_451, w_330_452, w_330_453, w_330_457, w_330_466, w_330_477, w_330_481, w_330_482, w_330_487, w_330_491, w_330_500, w_330_512, w_330_519, w_330_520, w_330_524, w_330_531, w_330_532, w_330_535, w_330_539, w_330_540, w_330_541, w_330_549, w_330_553, w_330_558, w_330_561, w_330_562, w_330_566, w_330_570, w_330_586, w_330_587, w_330_596, w_330_620, w_330_638, w_330_641, w_330_646, w_330_653, w_330_655, w_330_656, w_330_661, w_330_666, w_330_676, w_330_684, w_330_687, w_330_694, w_330_699, w_330_717, w_330_732, w_330_739, w_330_750, w_330_770, w_330_771, w_330_773, w_330_780, w_330_796, w_330_799, w_330_802, w_330_836, w_330_850, w_330_852, w_330_862, w_330_866, w_330_868, w_330_870, w_330_873, w_330_878, w_330_883, w_330_887, w_330_898, w_330_916, w_330_931, w_330_937, w_330_951, w_330_956, w_330_962, w_330_987, w_330_995, w_330_1027, w_330_1030, w_330_1032, w_330_1037, w_330_1053, w_330_1056, w_330_1057, w_330_1090, w_330_1105, w_330_1107, w_330_1109, w_330_1117, w_330_1121, w_330_1127, w_330_1128, w_330_1134, w_330_1144, w_330_1147, w_330_1153, w_330_1158, w_330_1163, w_330_1174, w_330_1191, w_330_1207, w_330_1208, w_330_1209, w_330_1219, w_330_1222, w_330_1224, w_330_1247, w_330_1260, w_330_1271, w_330_1273, w_330_1279, w_330_1289, w_330_1290, w_330_1292, w_330_1322, w_330_1328, w_330_1342, w_330_1364, w_330_1368, w_330_1370, w_330_1376, w_330_1397, w_330_1399, w_330_1406, w_330_1417, w_330_1425, w_330_1432, w_330_1433, w_330_1443, w_330_1445, w_330_1451, w_330_1457, w_330_1462, w_330_1471, w_330_1496, w_330_1513, w_330_1529, w_330_1547, w_330_1556, w_330_1566, w_330_1571, w_330_1582, w_330_1588, w_330_1595, w_330_1609, w_330_1612, w_330_1619, w_330_1624, w_330_1626, w_330_1630, w_330_1631, w_330_1637, w_330_1643, w_330_1650, w_330_1654, w_330_1655, w_330_1666, w_330_1667, w_330_1671, w_330_1676, w_330_1677, w_330_1683, w_330_1685, w_330_1692, w_330_1698, w_330_1717, w_330_1718, w_330_1737, w_330_1740, w_330_1750, w_330_1759, w_330_1760, w_330_1761, w_330_1772, w_330_1795, w_330_1806, w_330_1825, w_330_1844, w_330_1859, w_330_1872, w_330_1873, w_330_1880, w_330_1884, w_330_1887, w_330_1888, w_330_1904, w_330_1907, w_330_1928, w_330_1930, w_330_1932, w_330_1939, w_330_1947, w_330_1952, w_330_1960, w_330_1961, w_330_1969, w_330_1971, w_330_1981, w_330_1992, w_330_1999, w_330_2008, w_330_2015, w_330_2020, w_330_2032, w_330_2033, w_330_2034, w_330_2049, w_330_2051, w_330_2056, w_330_2058, w_330_2060, w_330_2075, w_330_2084, w_330_2114, w_330_2120, w_330_2135, w_330_2191, w_330_2194, w_330_2209, w_330_2211, w_330_2214, w_330_2233, w_330_2234, w_330_2235, w_330_2236, w_330_2237, w_330_2238, w_330_2239, w_330_2240, w_330_2241, w_330_2242, w_330_2246, w_330_2247, w_330_2248, w_330_2249, w_330_2250, w_330_2251, w_330_2252;
  wire w_331_003, w_331_006, w_331_023, w_331_030, w_331_039, w_331_069, w_331_070, w_331_074, w_331_075, w_331_077, w_331_086, w_331_088, w_331_093, w_331_100, w_331_103, w_331_105, w_331_113, w_331_117, w_331_125, w_331_130, w_331_164, w_331_187, w_331_189, w_331_191, w_331_192, w_331_201, w_331_206, w_331_214, w_331_230, w_331_241, w_331_247, w_331_260, w_331_271, w_331_272, w_331_281, w_331_286, w_331_300, w_331_313, w_331_329, w_331_344, w_331_355, w_331_365, w_331_369, w_331_376, w_331_377, w_331_379, w_331_392, w_331_406, w_331_415, w_331_416, w_331_419, w_331_420, w_331_430, w_331_439, w_331_442, w_331_443, w_331_446, w_331_482, w_331_487, w_331_491, w_331_498, w_331_502, w_331_507, w_331_516, w_331_519, w_331_529, w_331_549, w_331_550, w_331_557, w_331_562, w_331_565, w_331_575, w_331_578, w_331_588, w_331_595, w_331_613, w_331_631, w_331_646, w_331_659, w_331_661, w_331_667, w_331_686, w_331_708, w_331_719, w_331_721, w_331_722, w_331_726, w_331_727, w_331_733, w_331_735, w_331_753, w_331_762, w_331_773, w_331_776, w_331_788, w_331_794, w_331_813, w_331_816, w_331_824, w_331_829, w_331_839, w_331_844, w_331_846, w_331_849, w_331_865, w_331_867, w_331_871, w_331_876, w_331_882, w_331_883, w_331_892, w_331_909, w_331_914, w_331_945, w_331_947, w_331_974, w_331_977, w_331_978, w_331_982, w_331_994, w_331_999, w_331_1026, w_331_1027, w_331_1034, w_331_1042, w_331_1043, w_331_1054, w_331_1056, w_331_1067, w_331_1073, w_331_1093, w_331_1105, w_331_1106, w_331_1113, w_331_1116, w_331_1122, w_331_1125, w_331_1131, w_331_1136, w_331_1151, w_331_1158, w_331_1159, w_331_1174, w_331_1201, w_331_1202, w_331_1203, w_331_1216, w_331_1218, w_331_1227, w_331_1235, w_331_1254, w_331_1257, w_331_1272, w_331_1273, w_331_1298, w_331_1319, w_331_1324, w_331_1330, w_331_1333, w_331_1340, w_331_1354, w_331_1361, w_331_1364, w_331_1366, w_331_1379, w_331_1387, w_331_1394, w_331_1420, w_331_1422, w_331_1426, w_331_1428, w_331_1429, w_331_1430, w_331_1434, w_331_1439, w_331_1446, w_331_1460, w_331_1477, w_331_1479, w_331_1489, w_331_1490, w_331_1495, w_331_1500, w_331_1513, w_331_1528, w_331_1532, w_331_1537, w_331_1540, w_331_1547, w_331_1549, w_331_1552, w_331_1565, w_331_1586, w_331_1593, w_331_1597, w_331_1612, w_331_1619, w_331_1625, w_331_1626, w_331_1641, w_331_1658, w_331_1672, w_331_1690, w_331_1693, w_331_1703, w_331_1704, w_331_1705, w_331_1706, w_331_1709, w_331_1720, w_331_1727, w_331_1741, w_331_1747, w_331_1750, w_331_1759, w_331_1771, w_331_1773, w_331_1780, w_331_1845, w_331_1861, w_331_1868, w_331_1879, w_331_1899, w_331_1902, w_331_1917, w_331_1960, w_331_1997, w_331_2001, w_331_2002, w_331_2003, w_331_2034, w_331_2036, w_331_2039, w_331_2050, w_331_2082, w_331_2086, w_331_2089, w_331_2106, w_331_2108, w_331_2138, w_331_2169, w_331_2198, w_331_2201, w_331_2219, w_331_2223, w_331_2237, w_331_2238, w_331_2245, w_331_2246, w_331_2255, w_331_2278, w_331_2279, w_331_2301, w_331_2310, w_331_2333, w_331_2350, w_331_2361, w_331_2368, w_331_2387, w_331_2406, w_331_2420, w_331_2426, w_331_2447, w_331_2453, w_331_2484, w_331_2497, w_331_2501, w_331_2510, w_331_2511, w_331_2517, w_331_2527, w_331_2533, w_331_2540, w_331_2570, w_331_2611, w_331_2612, w_331_2617, w_331_2624, w_331_2639, w_331_2656, w_331_2660, w_331_2671, w_331_2674, w_331_2683, w_331_2691, w_331_2726, w_331_2756, w_331_2795, w_331_2863, w_331_2877, w_331_2883, w_331_2923, w_331_2929, w_331_2952, w_331_2961, w_331_2982, w_331_2990, w_331_2994, w_331_3010, w_331_3013, w_331_3024, w_331_3041, w_331_3054, w_331_3068, w_331_3086, w_331_3097, w_331_3104, w_331_3109, w_331_3110, w_331_3118, w_331_3149, w_331_3184, w_331_3192, w_331_3228, w_331_3232;
  wire w_332_004, w_332_007, w_332_033, w_332_044, w_332_048, w_332_060, w_332_063, w_332_082, w_332_091, w_332_099, w_332_100, w_332_106, w_332_107, w_332_114, w_332_125, w_332_127, w_332_132, w_332_133, w_332_144, w_332_149, w_332_150, w_332_152, w_332_154, w_332_157, w_332_167, w_332_175, w_332_188, w_332_191, w_332_197, w_332_202, w_332_210, w_332_216, w_332_223, w_332_241, w_332_245, w_332_256, w_332_267, w_332_292, w_332_296, w_332_307, w_332_311, w_332_328, w_332_335, w_332_356, w_332_359, w_332_382, w_332_388, w_332_395, w_332_398, w_332_412, w_332_420, w_332_425, w_332_437, w_332_448, w_332_478, w_332_480, w_332_482, w_332_496, w_332_514, w_332_520, w_332_522, w_332_523, w_332_544, w_332_547, w_332_548, w_332_567, w_332_614, w_332_619, w_332_621, w_332_635, w_332_643, w_332_647, w_332_648, w_332_649, w_332_663, w_332_669, w_332_706, w_332_747, w_332_752, w_332_773, w_332_774, w_332_775, w_332_790, w_332_797, w_332_800, w_332_816, w_332_820, w_332_842, w_332_927, w_332_928, w_332_949, w_332_976, w_332_985, w_332_986, w_332_1003, w_332_1017, w_332_1029, w_332_1034, w_332_1038, w_332_1042, w_332_1054, w_332_1058, w_332_1061, w_332_1062, w_332_1063, w_332_1099, w_332_1123, w_332_1143, w_332_1155, w_332_1162, w_332_1189, w_332_1236, w_332_1240, w_332_1305, w_332_1306, w_332_1316, w_332_1338, w_332_1369, w_332_1377, w_332_1389, w_332_1404, w_332_1407, w_332_1418, w_332_1419, w_332_1422, w_332_1448, w_332_1459, w_332_1465, w_332_1483, w_332_1497, w_332_1531, w_332_1566, w_332_1608, w_332_1613, w_332_1630, w_332_1644, w_332_1649, w_332_1667, w_332_1669, w_332_1683, w_332_1687, w_332_1695, w_332_1701, w_332_1712, w_332_1719, w_332_1720, w_332_1794, w_